��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���o�*��]�1�Z=����y���<��(�����R���D���qcUT�'桴*�xO��nck��+���/Y뷇�Ė���
:p�=��7��Iw�|��9r��G��i@�A26~kǻJ_�/�iĬ� ��Y~ *��jN���Kdp�[�<G{�Ml�zn,�춣���u�[��kbJ�^�\]{3�6U�qq�g�|b�5�+��yc��@��T��U��h�Ϟ(r�@B"|�Pn�7u��>������&�U~d�w2f+$��=���y2��g���A�v�����n�B����w�vҦ�:�[y�_Ť��7�Z�0�9ʹ�Y�xkQ�7�単ؐy)�е�� �C�1(JD
N�yb�5J��ItpAz�֤���������o������Cc��
�㎧-�+�^6bQ�誩K~~� ~�A�l�z�[(C��ބ��u��n�R��e��q��hkY	��ul�dqߟ">���vf?��p}�f�&�/��ei�<�gۖVá{�َ��e�;6�d_���U���fA(veV��6n���{V�-9���z)e�o=>Y[�`�Z���vUw���W��k9G�i�H�
<�z�lE1&���K�KA{�,����Q�?g�_�o�[1/1q���3x���5���q`{� ����3�A}JM�6g���XD����3����8(����fiT��Icᖬ�޹�7��$�bYa����
/"3L$��=�1���qDՕ2�&�ïF���LP���X
��rC�Y�8�G�xj��h�I΢��Ի��ˀ!�43�K��DK��1��7��X\}���Z�:3�����ߺE�a�r8���
��E�v�ݞL���w������������s�ng�*8(Y�&J�}ط�֐M�g��9����Ԃ��rB�@�zz�:P�	j��=B�����f0�z��lO�@w���[=p ���x[L�cJ�������FҞ��t�u���Ȏ�\%�����<0���PWK��PNm)�l�h�&0,EQ�wÈ圗�rV����<cN�V6	�����[ֹ?�@���p����v$�b�S���
1���
�+��������<���߷]��2h{h�aCk�GQ%'��J����&����F=�_o>;�M\�5O����2�?E�۰�F�n-=A���̦�+h�c�I�
N��';�����ʼ���Ss�i�tl!���MH�(ƵvDt����R�?���k�!�%�v������d� m� ið�
r�+(Ǧ~����!��A����f�q>�>���<9�6��N��$:�x����Xn��N��vni��I�UT+�_�N�E�5eΆ��:~]�k�?b>�k��&<�u>vؤ��N�S"O@�'$5
���d���zW7�������7�� �B1�N4��Ω�V�}6�e��MA��mO�4����<�[�7�L�/�s�sg�b��dɮ<1�m�aV�	M!�����o���m��).�w�9�t
(l��dﵿ�W�D4��&����"e���3���
�)����7%t��e�?���J�,ϓ|x�k=��Ov-B��hАܗw���a��zf���1�8o�T����=^��O�BG�[Oq0���j��z\������<�ډ"���?��11�?�%D����o +q�ĩ������D)�1�E��t*I�6�3�a28��]�$M�F�&@�ֿ�h�Z�ЂR���J�!����\r-�#�R�������@�_���{���݄�����'�~�n�XUa��d't>�|A�!Τ�w?�̽��0檅���+
՗k������`��Aىl�������,"]�����ӟXF�nj2�x�G/5�
�P���2Ǣ?��Q֝���v
�mH�%���V��L�$��_����Whe#N�2Di�:ޠy5@�Q8@lL��l��T�l(O�㗭�|��nMw~	X�eZA�]G��6`)ғ�8&�=l��σ�h-?�l-}��쉩�VGB�q��ߙ�����4j�2�Ԧ�'6�t�4��U�k)�`CH-OL�]̹�>}B���u�L"��n��c���3���2��e�p�cQ7���8��P�){���\��	^Lt������2�_2�{�V�}לc���,	�࣏���fAn����/����̐w
���F
"Pg#�r� �/��Ư��=+<�yu�M���6�[�Td�M��w�TR:G<��v�X�􉴈*��Ze^��O����ir!�+�P{�?O�-��b�B!���@ud��cg	E��{\���|l'^7��йٸS1N�4B(���-U��>�Y�����E4z�PY�S8$��]ތ^ �?�FA�s��{� �n���ϒ����{PVW ,����J0\�C$2r�ИJ؜�f�.Q��~���0GD�s�6�����k��9;6���W��` �n�*�R�I�����lg���0�,��p��p��{���9�C����tX݆�b;)K'�Ǡg�:����SǜK����e�_ �t�Xp�h�hH=��r�c��s����.w��m<W'Ŕ��8���}�z+#��%������
��V�I�И�>U���ta2�ȘrH6`C���L3e�Pêۓo���3hS�B�dF���o�?��F1��qV>"$�.͊%e����幥�����X�yu@_�Y1��擄>+������Y��*�*�6};�@��x���([���YYF�"�4�۸�E��~��$X�%C���re�;�B��@���E��7�A����H<����n䝛s��F����<�O�Ǉ�|���ˬ�aa?����F���L���!��"���K�%�>{��_�W>�6�$��#���Ud�
���	ҏo�����@�uQR�����7T�:�l�h�����gI�������H