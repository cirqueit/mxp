`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
PYOXaMtUZ4kZi/idKooYt3ON7rxKonYg00Pgy+xMJTa78IwvFpR4M5na+asuRCtxNxWHTEJmx6dD
qnDjGl81Zf8lWjSCKKEWC4lvlisfJwnq6uGkcEjjM7yvHaMOEtXFuoJHyRrpIs6/FaxEKg18U6Z4
MOPo8x/JDTiK5P9rFtWhN4sDAJWVVN6Ws+mohywi7Fk/KDtdlwRosr3Q+NDFrX0cuHV9ypd4oqAJ
spyCqga8aCMtq67EG7Rk10cr06dZ87B/PrtGF/0AuyHOo4GqnPC+exV4QKnHey48hq88Pdl3HnQn
LCEEFArPpxo4+jL8+7WY53eY6iUcziBGN1UZs9hN7KQjHlxqSZWCeHly8ywSSGOVjtfOH24t8TYg
xfJK8bmpfOrkQT8sFmWQhNMSLD+5hUaac05RV0jHkwmEoY+2GmwnOZqfuY+btyr20u98eb66Y/vX
toQh89w0Yisfp0e1Ibaz70nCNBi32Y9JkAGyrRCMm3RK/2BcbJ9jy2TdS7u2lTwH2S0PiaASfRjP
3nWWeMfBTwzlberIsIKthnqtLxZ919JMdYcz5Nu3PGrqJb/X9b5FSmVrEmacIS0pPDqfMwbWBXcy
Y13PRfm0ovPKg3g4LT3lzEXBLDb3GxX5CYsIkCKqsM383z2wYNtgfN7YTKCDWluzAo5H+yeHSgLs
teroOmOZybO2Rs+GT087C6pLfUywR4y4V/7NroBybHiGmwbL+/qDaQRPGO4coOp/asDNsxhPZs1r
BG6+7l+mobpc0JB96pHTCH/8lmdjh6pFn4yxL4W+ujwAxsCHSBZ9UQ9E/6eN0Sn6XH/FYHCONZhS
qTp5sdgAfSPmZTrBP75KcKL2Iank8FTObhRj4PzLYWNJbMPhXWyQzxFxA2uBdVYu8T5Ccs30bmPo
Ynz8vhVq78BKkA8WUqwN8j2nIuU0BaCDF2mq+Nnxfg/I8fvIBRke9tjsagzle2KI7nlKLbAcFQHo
J3pEG2mCRFCXyUU4daCd5JnC/NYlVRtsUl8iANn1ux8guS9BjOG9W5hMDFDfZiMAVFRZB2CbejWT
1UCamYvVSZ425xnjElgcATE5SZttv9tJvC/DSEdx+GWM8yTZrXeftIw/dvXfjBp71tJ6kK9amN1f
1ad9Z2A3dey/ay4r57KRt5RnpVElz0OzP8HEaUSBqu6kD1OG277DdGXnyUEOBFevX/wOrICPR88t
3sB0KZNY6HK/7tTdeBnoQwMFun1DkI1QRjahjXrgKK/m79uNx4A2B8pJ6sgaQIZ7H8uOMQNhe3lv
SvyRnLAaZa2ymjQAcLPhg6z/OjqNX4HWG+48iGvdlxDywZTNcPDbt5vPnlLw7kP0DVfebl7HLzv8
FOSQUJKF/zdQ48abINB1dfZP9Vikj7nmMe/umSfrwNocfwxWTdc7oBkA6pUITkKm34IUrj//Ndlm
04RcGZdZ/1xoOvQjBPz6Ax7/5lTF87Y+N47BuHDycwvMBs73CpndHdwK6YflBLCiTpFzREJLw46g
pA1aOghcIUMJ+87/zTCJzHveMVRT2SskNbqPpHISqj+SSPw0GMy/SPzRlTXP7qDcLVXJD5oe3NA6
nBYPXUbM66TVkA5SD7uYrDL0HIvogidEWdtj5paNjQA4VILpsQJm3y5xuNEzSkv4TwevxvUXgSZQ
UztBfiD4D+6ks6I85xqIe3fjBUU8GB52hCbhZGquvTQE9bCNSlqDuo+YmWq7YjiMaOHGuCPFv2PZ
3cuG8O5yLG6TNO3v3Xp2mOMqWPaUF/SemjZ3g41B59VVH4Tf0vj3x7g4Tm0EfgeK3zBYPQnTNi2l
3tzqhOa+vLdiQhXKI69IBbMhiSsvFNaW5R88gOVThlaGCwECPnNgc1JpRIFBpgZQ6TCmb0qt3w2N
qPzSdAUsq43Y79ItcmvO1/I6MLLBSV0iogmr+OqBU66amdb/M2siaJD+mHrA2lagOrtobMdDJSvh
I9sjHCAD5s5Qia2BD+P15gcNEULYq6Z72gLgQmuyR4RftbqcQZW7JmMXGXzb4zRG+iGjb8MLxuLw
9gA0pa2vtQfFtYfKqEwyQGx8Fp1sC61AxXnSqi5OhN+wt1U7t7PfPE+2WmH0HjDQtLBiSaAINwFI
TrmY5pOkj0VzX8srMzEqIlJrN5ebkeTMIZEUDAxlHx/wwqYawcto7G3RgJotntCQueATgmZRMjFF
cfSv6jsMRNoHQctRSwgUOJS6FXkzmEz9HjsaH7tvw6zJL4fez3h79sqoFsDhrTSCSYx5AvJQAJYi
aNuluGl7lL6e1DoQlGihzmp0YLORO5kuhFmxiW5j2KTbBSWTjL4HKL5o0fOURZ3kjXRTGfmANii4
Q15o+2vnsn/0F879+6y9Y/xXqXiLk2uGdF21xuCSwJFIVj2ph5ROfvQ9USYHmF/gOJkXYVUl6vNJ
Zjh4vn+cLWDA1+Uefrb6Bs0OBMrCelF3S6Y8ZxPbUfczEkRUBQIz+LZ7GrCUDfqpiZsQJfuSTusI
lQfzic4O/ZzNECrKstzT5GgBX4XWT2+qBtt9G+DXQSouzN9v8nKapLn0L+e/WdM6ltfpkiEzjXwi
g24EWXcvQuon5dcAXJG8z+328twrV9+rT6JhxqSlXUdICxkSe0kNOpswcqKB9OKfPmvKyY1KwMUQ
f7yQrhOF50ReOFP0qDEIF1/1yAFKHTyVfGgxc+y5AXnhQL9bZMFLjjEPFAlfp3atFfMg7umAT09/
PlXLq+2EF8gj6XKRYoPQqwrnznz+/d/XWkJT/4Ez45n/MgVjbcxPdSZ9UdrsneKIcGfuakfoMUnc
x86RpO+CKILZY+JyBCuYc7eF5cMuvI483ahASRBr4NfEnkjlXOszpBspvCBVrycZv9VqudUq2r5W
ysd0/Z5dcr0mu6kBh+o0re2FrXRMz52RB3aXuT0zWsKHJWrY+mFbr7zem1GO+GC5Jn63qnf7q83P
ey0nyt/jJMO0egH7o4WezbQP8+5de3p2U36/FE8lhWBg95kkfHyNh+gna9o0hgTKBeyZcj3FIZsL
tZynOxzfCmvMevs+gPPqL2he8YGuiy7FtKZ0VAqWjiH4HhQB4q4n3vZJBtJEnTj47O3J7KMjLnQf
7rUi5PX3gsqHfK7aysT+u+E9rpn6Rd7ZJegxh8qxbWud2zLEGxabxv3eJ165kxjt2vXoQ7WqzM2Z
QPzlfpfCegVUWEo3flvuc6TgwIQ3GG+b6MRZRbN8IJ4NUMhTFjhJ1rOo56MxJz45aY+0F9UUmtf9
MnpdC8pR6A0Vb54Nsv6lyJVMWiwVoI9sGPW0FeUdavGi81DAIdq7KaKPfQ+32v3zcTEq6T27jF2c
XZnWfoJ2mE3Qxg4JYneRP/YM+MSTKGM6eXh6CQgzVHssXueZlKMNtCwplGG6jZdGadty5f5o0jPr
WwHCqsPZodkOMkonuak48EcZKIHkXqPUDwHmIOrUEhADSvpOO82sRSJgunhofdGVTevBx096rXRy
eXEqWlPbzTd8OJF9bucjibg9HcFnCtfzrroX0eK1jPJo/FEmAfmX82DJTHAwCFIreXWDySvy5eMh
7KBaMiWFw5l6DmpH7uB1+WjdzkYI/wbGE4fxXFz5zBdRxB9HgH+sbai/WfoYqp2zMrP3NQWDYr5E
GyTCHyFc++DftbT0puk2PUfZjfuM+dIt16c+6WAxDE5SCL/wjrM4mmpQIJiH7qH2NWkMJWahRXA6
ym0T9uw+wB10oPG8+e/+EM/u1h8psySbEo0EpGzBGIb7OQEFUQqqMV6G4OK0t1AWHcrcc/Ofz6Qc
/BTxMcTmBqYqrfZqiexLAfzJethN2+TBGjn7sVYUSZ+FCEY24ydEVeDCz+kgpaoPk1MawlhfELCN
nZMP85SVzvyXo71u3MwdJfjm2kKHqNCNpObgSxL+xdPVgS3V/hJX57v9h8BFT1ZaWHc/37wx7qsh
Fzx5lk2u+KD3LIusGRwrGp0Zl8r1CmxxOeipwdazfwRo0jwboze6t25tQ8oSZ9WYyEbKIyxxpPO7
pNmU/nnEAZeQoK1X6ryULpBbx8g8H4leDaly8XZ8H7CxwEH4Tx4NOtrN6C64vPt6UG1p0UUXeekp
gCkO9Kx5SdJyXeLGi1GWRrdq1TAxPaXfbvUV4ANe4hSbwoB6g+8Pgeplw3U1Ymgz2HQk5JtF3ZrE
YzjeWVtbsqnK+pEhUOByZ9SldOFZb8tYiN4g88oM2lusJIjgGJezTI+9v1BAm1phALlTrKqTXe1U
FSc+UGj3EQhabprQYYFtRjqBZcCHn6qO0eJ7T01TZAtE/o9arIwAWc1GRGwP4Ndu6LHH7bYD+h0f
aD5Dlfw+f3UicUk5cNZ3ZOvXIW9M8z8GbSFf7/S3PVvA3dalLYZrwleOycPqbslwq0xsA8QG1RCv
+jZvsVV+Mj32z2DD31H6EqhUac5xdx5zr7Ul9Xg8lrvjY3+slir02IJFJ1JE0k+doL4J3GX33hin
yAYOizHq+nzp8/P76MC6IYNwwHepdeVWuyJY/dVtm13RnJhZ55x2zGy+KCFdD/2kbanWhLNG3725
4tTw98nUYlov2T5kqXdjQgvbJTuxm6YE1E387h4wj4JZJPliOe4PtsPhK6M4oNgQFeSLMYXUKbE0
2oMNJSRpI36ERCep3nFB8euLAulcEp+ELeRHQcbxbXTskJAv1Tf+3tpkUzQHYGFLbhiUPkPJP+AX
ELxPtI0lxp6k9zHUAY0wbw7U7mZOvO5ydqMNz6OKToG8Mi0IM/wTn/b6TvMjU8Kl01afAlSqCsQc
ejn3x2Ml5AD0lLoUmMMvCG7g8DodsrpFr6gTtIIvcRGMY1wJ/pAE679zo6Oo0/np5osQt9xZcwDj
rNQiKqn/eOClDVs6L7f+3xY5xBmfLJLUOJeuX3h2E4/HwcruxHoQXyAbakA/7THVzCH2KOJRiqXP
2CYnEOsXRfmpFD4NQtHDlSDxGgE+KjO4LVF83lJ/m6RsAGNmmhj94ZcRhD1O7STYzmnU5tHLBhyl
of1M1XA9udu8o1zNgEfH32SfBwSnbEEacbiMhps18NVeKZ5jwCa31GVHp5wJL77M+PIowfuQxvnw
WvPFLnr1jPWzb7BZdUMm3SdFrrIJEWBphxV0iFXnnz71H7AoyyEzcPvs5LrT4A3UWyd0TEAQOiSN
6tLED+n3ukkW3r7eCtPFtaFwBxEXAVPcYlPuDj2W7e0uR297yXeisguKUb2EDmk+soRcS73pfvYa
AERvyXKufT147DHj026GLRrNhSqoDOaRT1Snr1ZcdJlb2JKrhvyuVR2XmOKmztwS25NMeMte+2UB
AZQxbQKEjDGzA0TzOnl+pRCc2wV9uO6899XUXCW6rcRcHZdg6sli9SlpUsLA054anf4ovwrdSj4t
Y5U1Y65/bXoLdfBF64ZELYba9x7f70MIHQIYMjH4xxSXt7/feT4JLGw/wtuFcf0pwQjOXcj+BfKB
tXpuYKJQWmBbqEzzXx7t7X+h+DusJS+FCAgBFbcvmCBOCY/oEj7wWndsbPI2Z6pR71TevqDq/6XP
Cdo/389kjSJNuHw0hfiXjizWD9KunGG7HhQbMDOI2JkfhnMUQyBd0wZU18bsUgnivuJmMUv8i3AF
VjmUtxOlewD93VTjipXKdHgmCUV4DY05E2yeoAdN6LHYM3a0VWp+UaAODSI79gGYnWV+sXmrMieU
5Y8ihvZOgLbXdRF0jZu/dxinpU6n3DMBA2Ir1YAGbBP7q1okC/+JbvTAwqAi+CVhLWJCFBrYGz0+
T9xzLGobwXul7Oe/6zyCinFCOBu8M3vyuX95ygSVndwc5aEYb6y49KQxWUshMLaAoNHq/rVzHmkd
Ry6yfwwU9m/BFppvz7KZgCQaZ7iiPCzPeMr51jJxvXW/WODQkj4oT2UgKPynTqVeKi0fhc1DN/5P
zVem1H+w1gL6/4B5zfW1Tis7L/Lla2IAWhPfWrm0gNnYtdyzxXDqpK1mCaRpUpvrVn1na8SIImin
Ow/x5FqQvAW/A/wLw0X17RZ/v5L+WpiQRqLtxghvut2YCDm7Ww94/egOxrgcyldXk0bi1P7iSiev
0jF0YMjpwRvadPhD/yO2v1YzzZt7S2Vhtxgciu7avOBlWAvSTxCx9+eP/zasFbN3w6P5ngKSQqeR
/oB4dmiquWCmfh+r3L+Ago+WrRBUBtA7scxAm8F/lXP+e8fnlr/qQcAOM17quEnTxo+drqMYOrcL
F6kcdNrkpvQ7WBTbiElp+OvaGeLmtKDo9acYjb8qcnLeHn2SAZd7ruIpwxiIcIr2KjpLvC1fvLAv
TGcv+w2QucghK+EJh41PlZQNOZ69t6h0/+WRguMeAASpqPdYkJbeKsrcI4YzLGntvNtqQ47XXCNc
IhapsmNCouzAS4lBfb/Q01GWHcsh7I8fBQnStuKDxNVcluLjo1vCiicBEbfC3lucC0kracR75RD2
Kp1a9JqSbDFOAq1PO1ZJ7WMRQfWsbP1OHaKl8gKFyGHGsX+ppGuHbn34IhyBuvVDjOkQRsBLYc37
eorxEZEh/y+mkvxkd5jm1CcbEwduWLWsNSQ5NtYX0kgDNZQivFGg5/NscxIyb2r8bJpL48uwAqZ3
2BMDhFXsiM71Qy1gXzG2CYquD2UhozLNXU564zblLZNIXHbOcQu5KegjBLxRuXoA7XJQzkVGc9zr
6rI7OopUwW1Q9ou2Hx3Ry4L8gnDOcWVJfnhjhN0NBtlcTYNJbcqVhlx0krhuMUN/WgRN9DzrKxOy
3UO0azvu6ccQ+Dpc/B4tQ268Fwi0PbSVQmw1J6iAzEkueftDYWS0rUOvTcg0MMqp7S/lol7z/BZM
oJrhB8d673/8bWTQ0iDSQT37VqGoHPRbafq73hcC2aDmNPRG4fSpKGM9RHuJHqmFEA4xHKm+glDt
Hp0jU2GZMhCRifhW5HQIyZ21gPL/khAvJGD+mII7xFv/Qt+IlMuGlzSCPe1UiHoNFS47x6Ekmoh/
tC0sNmkd8iUZQ0kpYlPKcUe20sfQh6Ns6wEUScbWe5KjfbTnoU3jV9AzaNOiTDkLJ5hhAUDzu4r/
GOGSHqoK1O+ON/JYiuzZBPMGXKDEBhHqD1rALot2ubFNsi3pit7aVcBDKEM8kl1MB+dsueYr/pXD
Amsl6PkgAvvr9OhlBOfi3r+cif0YAxkfyzCfkllj/LgkR9Bx6X4/OZvEknZF1u5CB2Ea4PSFWf9g
lT8kj+mYqAiyaJdEnGOvwVprk9JIP1cnDjbOtR+D73T3ZDb4rYgpLnXD+QwoxZGPxB6l4NZBjolA
3TuR1tZo6t1nbCzYKheH8PiI+SKKTWuVzwMhrUTC2l5yczFSLOPrlDENssEkEZNJRbR8vaBPBawb
088CS42/dtIYUpD9b5/KIa5PjeKCRTgGWcNvKSXXDT/+0pxFIcieW8wTTMtTsOoSwhr/1IGnn2i6
pSYkrmZrpkbbQODjRPT+SvvSui4puk6/kD3lhvt/yNLZAg3GWQ8vpmhT8io+9TYacMwAOnFQaQo3
D9fVIHBB5TRMTdxP9Knsd4CN0flQwy2k3bHAz7K1MGkucKW/Seq7/3gSghzLC1KoY6gDJAqMhnY8
gD8FgjODD9vJioRaaMvhhCpWzSgwA2t+//ZAK5tCTqql7dJ2HJot3g4v9jTQsWBsGg5vp6TVW7dS
+8vXcRkCT7b0i+c9ylJXHfuWbERWYrdEA7YBZrDYkPT9gyUC32RAFpszb7K+V04IuDEyrN1+mI0/
FHviAVKtERtAzaX171VAQDt2y23rrsJTSN9+lbkMOtEb45eidl3O28OXK4aDVphgx4MxBu5GXpWP
NKQoPELUUipFL26MMlblUkSVnj7Q+uiq7bmXMOEdirGVC+sqTrkrZrsxhBRKeZkGnHspmV6KAKGh
GxCVw8XAdHZMJqU8ujUMCJix8GZlArMDUoNtymUF93Pn+0RRLnGzHPlzR6A1w/5eeZRQKrB0w62O
4aP+VWaJDQI9WBvYzyz+oS/JoNMioEMU9U9uQ74fGFVph34+YzxuTmJR4Bksmu4p6cC9x25xxW/g
8pghToY5GRDQp1viYnSplzVClkyqFcR+k23nUEbE7NEGMxAfS7GonCfI5bHDGfyv471aaXWs9U2Z
Lro1YE8B0hO9tcngnY+FGjuOnLYW//GHTSX7WRFjJUMq0FFcoKo3S0WTDl4iYa59xp/xPK+iaSEn
Ya0+CpjWC2QoiGtXsPypXRBiGahejs2XGPTNZegdppHZf4O7xVuSmySgnHtWRNNMaytrkYDiOzA/
6HYMduFfBCD1lG/skA+hM3QxubzTG4HiXri387AyBLtyHIAAlcOHn647q0yD8L5Q8f+D3hh+y0Or
zw5wzU1L1XOiLVpNvJT/Ep32xa+OqeTSJpQS/iXj+XnvSgBQaVvvLVm08K1/+yHVxVWwpSK+3WcV
w29lAwUC90bTQEgPWBIEE9DnBoxyFFe/jeH6/zjW86PSkm/t+RiRSxl8WcBwKEqyifBP3RPtbToB
YKvb0+Xp9BMvGc1I89LpqXHjLubMcDedXaElQ+i8OeV0LtLDzHJ0RwiRgWAzRbIkrTa9B8J5jDbK
qMkmB2+N7aJDB6K1iigXmUr7G+PgeSxUyxvV4OkH0YKhEzA7SPhv+okd3JzxrAXC3UkhZjC7aeQr
BwuF6hWT+JaRCBN/kMmiuJtC58C+qAOaXhW6Gs0X1YH5yC9F8kAAVcHHY5qKO/PC9VtaZAlMMllk
jc9fuC3e3LD6YB7yfqz6MQwZWjfdcFQVliMTvLwGnEWy+bR3V3+DEabFOMepjRo8GjiAUCKys/dd
8/61OLmjJKWk/ivozWR5tpdIIE8jBp89e/4LlA7Rd1g0Rqwk8xyoNo3orU1U4U7TplxdzA2nmjTX
LbcjhHIeBuZ7NHLIIrS6UnqwETeQlEmnOUU2YlyMSkvOZ8FchrsSoJ2CFuSxtDOXHMImzE2PC48r
PhsAW7JKFmJd7/xeom8wJDmdWtw6scSDWj+ZS7rOH0isxpWSHaHrsLZ686mNvfVTsps/wNCpWsZc
Up40nHlS1E/kiWwnb7mqmSy+BAzxpffJmWKC7vZHU8rQSxo89zBMmuKRj3WgncPJBHrvZLHTey4A
VYtv9jw/OBdFmDChI1GYQHfAlS2IYdJrYELFHYe7/UuZPI8Fkm+z6YPkZZtAF/oy4dCpeD5tbGjS
eBx20v6o4L6g0S5y9AdaBzXTd4VdsyY6+5euw8MTz1ZbiaobGW4p6zzQM7MhMZktcJStT9hrJkws
m+3wZm1uwQkY4WpzsZz6p6vO04neU+uxh1C+y5vVUiKUm6IJk2JWcC/pw7D0/aAq8vN2kuhnO9oJ
h6zHlHRVo7zJjiBp7/Y6WRsQFKhqhNiAVevN0j+Z8qDOCRxdY0q7wf16HsXDDf4nBHz5rjp+3tAZ
H4UPSqevxB4RWhD3pBPVbUptyA7TW8YgWPQUCqQryD5m7T/y4s084ue3EoRxljok0F3O4hlQk5VP
zSC8ccAyl3NOsTY38tsFg/sooZXOiis9KR5O3xd0uXDkmwreX+beoeuyAmh7EN5rHVuUzOmhlgy0
k3puiKmWZVH1vwbGf6eK4xjnC9MVuTRcmv+Pvf8EkesB+yF5WXxitXgaBwFDGPkgIJDi+9yq2+wd
JUbvUmUdHswzT+GgpjQU71W4sZdEVP2TzCLWq4Ikqj9tipoPVSHiJk5WclF5o5qoUVaiclddqeyc
ZOgUMHCaY0nlmp+4lALk6ssYoeZK/vajDZzpaj+boo4MlgXRMQIo/cv9NqqeMj700r3CBux+FV50
b+qmHw1NFRet2sxuzbx7hHLtZD+yxZCkcA2TFDH0kD+ho0etulT6D4p/CPtffxzyqRZBsAea/j0I
fCF58o0VOZkmKAQ5GB7FnJc0q+TqV75QtuvMIuG1ow+KKceKhxkTC7qck2SpgaQac0mtcsSdZKF+
y2VRY13Ym0fcxm6mfEfCS37DyzPnCNMDx+kLEoMyu1TbwR++2fWQVr66tuX9QKeUP/ROceKeGLxg
/Plu97rmW4RVPBdgFzKWyLCL7s2qHdJmBU+oMd/nhuCWj2QEHIfFm82kwRxi9vX6tWTiMqH1427h
srdegA8rM/Ura1yAy11hES+r7tDm8dXPGIHZUK4VAM8nMIQRyqTZiBHoH9sgbhlb5CQInxeLOeQj
pw9y+me9Uil3SRG6ObVOLEs7v59Y0TNjAeF4yxpzuGlbtnlGQgKHKUdADuRm7bokglhTO9/DWw/e
LE0hKRz5TuMlTfW5BLL5Rk76MGALo4ywhrnfP37d7Jl1j4LdVa24HmM29KzO80gnNLNvm+zijopX
8nXaTDAIF9QkqBdNkOzi6+B3b2ZlK9XkuQRoD3w3xvRB814qj8sJSFclO/ZTKgEVJGmph7xRTmz0
Bd4T8ASlXUEwo7UHlvb/+tEUuKWu3J7EhBQ01bbL9W0X+loMhVWPli+hzwBMfo4RmzgHbW0KkYdL
yeziWYIQ3TRfpUF7lI0Nhban988irrGSAuSOcVPQpmYkZH091Fk9g0gjhKYtrVIxIYZf6Lp7q7cg
RC/57V2CbeJXgO6kvsSdsij5bJdgmjBn/JTjqLfCLf+uhhohSU1aiLs4tDB6oB/0mKeistKlgOtz
UlWwlbyTEC8u3tN0IfX8otKgrGA/Ei5ioxUU3BELcAjjZxh1vrFsuvmw8ugRjN9/fz9RKuj0LWJa
KNtN4YhX/vCFbevBiFS+R9QAV5p7Ee5orgUqb9pijS70BkwYFhC3bMl16xYy4dsx1ouNq3Vzzi5q
O9g2SjrRB5AoW1u2d4pPBUnWJwN5H0g4YrvaAelvwu624KCC+BgUHmL7zLB43Q2mgiHRI3Q0r1pG
rhnHMBWiT/+pHKlToTrYj3GKvjQvM2MSVPC4CYi+FYjMsP8n6yPUkWxEXEVd4ExpA36tueWjZu/Z
xZuYgmGIPcQ8mWpHVYxvXR+4/Kl76bWKZcRp+MDjpkCpeDBnHnQ0GVD3037MQ4UB7mebA01di1KH
zMWkXqm/zh+ph5lZZJyVOrXGaKR13NYm2Y89w8qqJHPkFFlRPYZ841G6Yxsc+HS0QPOBg4NB1qx4
m5wE128S9stRyYjUwI/Gr5GSWM7CgcKfFbjfhLRxJSooM88EB092Ox9pOlahymgJ4n8rThfFOAgG
urTu+C2CcrtCD3pivK2WVlHg5DastxaASEO4hG/Qpj5qOtP7I+IiXDpnNmRBKH6iAQ1hXHgzKhEe
zxYmePfcAiX+pOW9/x53j39XMrxPQ/uT5Tces1A8YQg4U3rc936rRURwU0b2XpzJNcrXmknkKNPN
6tRKyHoid7tzkB47aaZK3+pOzyfWwnc6LKKUR+k2SB4Hwe75ZeY4Xk6JXQPH9BdgsYvTEWpSuDX1
KVr8DpXPwtJMSWHW46drz/0ttueBj0Ab3uWZlDsO0rBaQXZjzRSJ/t1b5zROnOl70W+WHcGq215t
9fGijmvyJeaWt5s2b8GY1sIaCSLe+1CTCz3cMKrPWNua0aNPoDEaPsLkNodlyf4d9D+ecMyFb7ur
IBaqPZzn0Y/jtodmiJd4GQIxA4xTuVf2nuE1dS7+wifkS4YD2Az8lnhnLB3yVicBblBQigJMbWAd
Y0/16GejSTu5ihj/qIMswloUys8Y1nEpOebXVevJFjEc3iNOoaxzEch5D8aXGDsPKeADP42gmNSR
xAhd0LUBS0yY4cH0i0+stM54VTLKMb7wSbUknmriktxvNyHa/q2ndCquu0lXh6wiuXiWDHG5sw+c
Qs6zzdDrFHvTLA/DEcYFbm9Oyx4C1cZQGSc9ZpABx97UI4hxr+3nix1/mSVRwts8ulifMG6z8Pas
u07zP30HFUOzDcf4pKCkdYew6Ly0c+NV6ew5WriAmpdz30NzDcogOFxKlQpI485EKvf8J5/AYqrU
k315PZDljtggbQLJnoV2pSBcxfuTfpe+bkgCIVprge/pKpPzUFXyOMSeXqpxsQg38rPMk12Q4M9F
A7NosVDaioj3sc2ZgBb0jvb8rKcby87tUwSqX9RHrS9eFIjaDBl+rR+8apvXbSd9pfHPfBwrUz+u
6fgCp4kbaEOCGjWvzVH4ztyf6DQwGdMYC1ddRTRXtd1SUQ1M3+20aU2q13lwuW0sGdRYaSyYJw4A
AaATc/WtA/IEgrsPxLhrvIoroU+/cNvEsBql/Q2sjSPJjCdUnWM1P7AuHo24Q+xsZhdH7FVJrRgY
dJhUBetDHk2xRWnTCFXJkgxOJHThipfcnCg4yYzm9zool0VXSicBZZTp5dmcsiOduju+AdqWV59p
jHkO+pm8/HCV6+PLjLO9uGO6g8QqlmSLppimbiTxo3tWwiGDKzy+Tv+M4/NU+qsWHS1b9ZAVAa9L
RcCjQqTtDzvaFmMatMlUSAh3ObxA5deKHB2gPXgc+rDotEOurI4qOTht/oP1NgLgrt47l8xFt6qx
o37lpLDS7DsN0C0sULvCWQ/H0f19SCkWFyQEnnAfde13JtZKsajoSpKzFFTetQlS6d8KYftHa0Mk
ewmwiFTMTaj0e4Se9N2eVz4v2VJcLFLaSo5GnHonIXLLBzP9PsIgsyoC9NqZnKmiK1r38bM7AH5Q
9RmtF1HyhjLpwz8u/rF/XEw7KtceRLnhNdl3MFGvxcclzgWs1tccRjTFq3SLgwK237hlhodq5TMR
WGtFjsur+nYEPWI+3HS9l9iCavELPyJRRlhznTocGfv61uE2kRv9EfICw9hUNjptj/bP2ipjLhw3
cJ35lx4y7/uKHjsUtsXk6BQdz1j8MJZtt66VAhUM3AGA3AoJdMbTNp9MySES9DzHAD3awpHAPv3J
nsCCdluN02KZFDiUce1jflspszYYrH9DqOTBqaHqp9/FqgKGfwBo3Qbc1IajVGWZMXEor0NuQII4
cZX7d8h2ahItVJR7RjYsBZvk6VzpI9Sp/hSCtShy/KixPulsAAB+DRA/HX6mRUJFlbm98+DkoFRI
PVmY+VsnalApE6Rm/VnFGJrZwp2qaWGPRJCPsJ3YakhNiDkDNFtZ46eSAdEUR51vOxweqwX2r5Tk
OZtXSxF9FpxcvjsLOa81RLeKU7vJqAvzXMJS3SK2diO219QZJnObWJGHqeidviatvRfadoF9jdOy
C2A06O61pSk9LIBWad2/Ybkc6zRjv8eEBugiZdqjqzpuQS8WnZLl2MLWhVIbiaAGhl9MZLl0lH8r
/THJQDpd1MLCYAcg/Stk3U0ebFkQn4eVycG/ird95k/2JnZmeMZ6z2HVnnOQKCvHZ8kpzfR7pT0b
mg4buF5FbhDmeWAvFwDhFwlqT0JaV7FXcWDowNnAzuFd7afBN++ofk19efQo6tuJeAryrSxyJTqR
V+hU/k2OTR6NxvqYPAtpQyJvnqMq0da4pNJcNXiIDI4uxlyZQdsOx6r38YOIGHR52dE1jHaOQX+b
d2VhYjCyDBfK5INIukl8hum2CzHjKdRufyOAMoCdHJ1Po3i8sRJrgsYd4UbYKPz0SkejvzFklc9i
g5w7i3ymc0EJQZJxd6tv2c9KMDCg71Us8dGv4mYviwsu2NTiiZjNLWLv5AETtUBwIx2MVb7b/b3q
LI21qUrDKXZ3Anur0CBV06mtdXsPa6d3otnlzYCbs7SD3Tb1oz8FtGpEY7ntFtZVWoQZahdhdiFP
4EGjPS0SyBPYM43ugIgG5mFz3wE2zfIFyXU0aF1slPp4JXAb47bdEE1Kq4UDHT14/TOV2eUn0k/1
FLopatagQo/Z1WaM21yEmMoMa/5cYjyHmwb+2xDFZg5WbPRqGxQ8Eu1ZuXJs1KmtwwewCHliUAKu
wdvf+/m8Wj0vtP+i9GfUJJ5sdl/eD/5OPpNVRdelWrjTMoiBowRtPrQE0Z5fqQmFo8OHaRML6Ero
3hNKjqJ/W47rDll4mpRsPmwAtQaHebZ9SG0MjVbI7lCk5GAPHAC8Ogh30GKpFianvFpz6YTZaX2w
iBCZsadDIvb6C8VU0l7BtwuOGBL8rcAfEjOxOYGVgHyIFyyySw6GgcI8c0gKRrTZT4zSQEWui6qL
5Ym/IilE+2hk6OLLTQedmfNHUg5A3PVTiQNUVTz5k+xc1Yrl1bWFag+Nxy8ny202LMXyDoO85M9p
NlREG8nm9fAQcyMyhw1Ssnf4vmHtDPfoYNAgoZY4KkJoU3wxtPc=
`protect end_protected
