XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���kl�HKT�;˺p���5�zB�$kբ�`�z!��?� a� ��+4��f��=�f3�BH0�a���ԦHs<"�k�����me�u����2�>���/�Z�>��+�5Jd�ն5��8�u�m���I�PE��y��k-�{��\:��@�o�s�CF" ����e�2��!6o�?ˀ�L��vY}K���Z׵�9�iNX�Z%��jn���6��f�<�(�F3Pvp��ijW�:�L�+T;�^��y:[���Ma��v���,�Q�	<UK�ˍ~ڮv�2��~�]�|�#������_��Ī��'H��}є�lk߫2�|��Q*��T���%b���)�B�h゘ ��]ߎȠP��*
���[�p;V�碭�+���i8q�C}�;J�b�L�f���l#"j����M�N [���gI�"1��[�$䨦T��y�V�B���E�
mG����}�,� ���A�+�J�ٽV�_Ԉ#����A�^��}c�c�����3�ak3��]�D� ۘJQ���W��q��E�9���xT��I'^�+c��C�IZ�Ǆ���>�g���-on|s���;1���D��K�+�Jo�H��{d0.�� ��фLD���G���枯#|� ��zw_~Fj��� ��	egi�kHM9kO��*@n~�3_�w��&s)Z*�~pdt��6�p��:&Ǌ&�}g98�B��䗼�T�f���}
��u�ׂ2��v2�0�FXlxVHYEB     400     190� �>Y(�Q��v�v����w���C��s�!,���h�''�H�8���?#����p�?��j+�e�X��:kFQ�~��%�F`^B<|L褝�����B�&Uo0̻Ͳ� �������HC�1�r�.�qɧ
'���,˛�)���R�xe\�K��Y%�#.�ry.B���,��2�����%�Ů�D��q�=v�q��X,�-����a�< �`S��w*��̋ը��l��,(���1K���gŧ������č��\�-�(�l&�bV��V�u��ц7�	�2��Tq�eV@�\�+ʵs�7+̍I{�g��C�K{�˧�j�A9�;�������o-Gzp��K�_.�L��Z��h%�z�:��HKX�xm&��924VXlxVHYEB     400     1f0�t3U3#�8;�� <A��i�欹[�2ʦ���"�@��?;{S󀬍���y{%���B� �q�k����sT��D�_���y���s3W2�����ā�k>����~1���m���"yw�5v��TǪ~*q}n�����he�|N���Xː9���2r����ϊwu�\�}]KE�.��nw�+�ꈮ���N�m�OW�������q�)=8�o�1�)�m��@���jf�ܾ��?�� ��:��P�:X��.�r����3V��gh�J�kv��Ҩ#��	1��?��W�ja̢�v��A�أ#c�����qk�1��W#r]��[�'���D��������n/��j��(��Wh�@PZ����e>�/_��r�3d�����ځ��[�}-l�Qlk7+v�mĸ7���	O���l�����/5�����` *�e��Z��f]+	�*���'�
��V�I�B��H�
�7�������XlxVHYEB     400     200�S��=�,oB1a���{9��>HM�m�,E抹m���ĕE3u����o�e���*�
���5�
4���ǯFq�p�����'sA9R,��lK������H*��ߎdg�^���AUՃ����l0�&WR>,Y:�NH�1v�OHߨ5C�]�aZg���B"gr�	�'��n����,qq#��L���.���$��(�o�����ImK�P�!�Usk�y0r���\iR!�0;���k���98�[�Ѻ]W^ճCh���v���/�G�
��n*F	��&T�[�\.�A�	�gӗ�����T��x\P�������`K}PN�IQ�w��d UX�h��&O�Z� �0d��%z��
�l�sx.j��[7���ccO�!��@���K�qԹ�?��SJ
I�W\����*����8�2pS��K��Į�4F2IqJ�s�H����<��93�KHܢ-�s�j 6���,>���=�Fu�H�xew�T�JѮz��<ϕB7��<���XlxVHYEB     197      f0q�C(�V~��*��3T�����rw��[�q��=8*M2��k|;���K�o��l�'� Q�7��d��n�at��,���_`��JD�6��(Kr�.؝�wE�
��z>LW��p�s88^�j��Iw�`�5��[=j�.�:Ԝ�w�Z �BUױG_�]����g�L[2�ȧ]ٷ.��}w�/�>������POt,m�b�@Ś15W�;"Ӽ�mKWr=��