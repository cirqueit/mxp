XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���BQ@��S�P�� ��Ӭ���Ș�Ii�[��nz��U��|x.\�zV�͝������q�;M;�����~��h%��h�&(V������$�3"_�$�~aD��0����"o]�Ya�tѐ�W�z٢0�a�/��f�o"jG\Q�K�:&*��u�0��d��h�p{�5dc*�6�a�C;��k�,�0(�I;�~�U��-����*��(��z_#[^�2�c� �}��[P,wZP!#���X�?�K��$���s0@�����I�l��E g�>�S\C9�d�a�?7��d)�Mq�]�&޸��̰E��s��}rD�R[�#���5M���)�G Ww6j�n �	F�H���"��;�pW_�����[�CӐ��T9����O�l�P���[#;��~�eA��?����Fa�w��l�Ev��v��`f��M�8(�Z�)H(0�u�,�����Vb� ud;{8��С��r�5��z��ct�`;�erw8=��>�%A�D9���*
t2v>ŷMhl���h� �����BQ栉���A\��Q��B�� ��gӟ��n�@�v��7�F�P1�#��Ғ��N�2��y�p�Z�¿-�$��'��l�΅��#��[��QG0E(�P�lQI�mΠ�����}l�5Z�y�z������j�hV1!-_(n���Ď\2�'�Eؚ>�D0�B���X?r��U$Y��G3C���Q��̯*�'Y�9LT{1ll��c��;�&��_�MȉXlxVHYEB     400     1f0�5��g�2?6tHpҏ�
s��ԫ�qs��V����FD�p���/����o�n��W�׮����;szNۧU��+�crGA��8���~U��wAm���$l&�� ��ZO��g�4?�ګ�
s����M�C�2l[�e4"�6(�F�&? +��Va��c���Sϱ;`�!u&�u��ᰦ�!Z{w����\4�^�ň�o��q
�a��ʧ�k��Rl}����� �w����=[ �dp�µv�x�cnJ�^�icD{�B��
��"Ûk��.���C��]-�?b����~k��,�n�	�>c�Ϙ����30v�E>6��rN��AR:��sq���}�Zy��%|(�ɘ�������B�خ�f�b��Hp�
�#7E�����nՙ���s{ԻO���矄�1��.ޯ��W�Gm���`�A��<�?�x?{w�ن5$��P˔I�_��ĸs!PH z>zyt/XlxVHYEB     400     130�ů�
>�a��}Hwi���8C��&Ku�eA>8Aܘ֗�D�p�3���QJ*�x��^�t,Z7�d#�_媴�( _��o���41�H���7K�G����o�� �|�=؈�����a!��7�+��zܶ
�x���6@Ю�6�$�f���_l8VtVB�0���7��pA�(L��%���5P)��~�/��-F�-Yn��]{�%Dj�����yE>�K.L�D�2s�f�]f��Ru���2�M&.�\uS���]�8gP�Ȏi�A%���5�X��w�N�/;G��&�-��sXXlxVHYEB     400     120­vY�E"�Z�g:��s�R�x�`��t�E��<��e�n=�������|��ۻ?Ь��y�[�������P�T����@oC��>�Hh~dgx����̶TX�Сq%���\(�Ww�u�L�6�[�v�:���x��;^�;zl�W���(Q�I<�̜�ahF.��� ���>c� ͤu��m�����E><��I�^��9�RwĞ��XH	�\�7 ��d\5�����Rr�X�	%�pg�{�!2���)�֧!��.�`��*�7��C��|8�OXlxVHYEB     400     130�(`�o׷�H�T��x�нːϹ�t�=
+5?d��f��g���-��%x�cF"mu������&ѧ�	��w��w	Ş�ұpn�6��z���G�(��"�&��4 UM}������;Qh�}l������0�/K��%��g"SChu}���o�*Pv=O�9�!��!4r�a�I3B��ʖ~Yof��x�����N(�R,��
dR�L'�<�˥"7�eNL
N�g���}&xp��"G1XB�s��S^����bD�\Пe�	=8e���cOZ���X �[>yN2��&�����>�rn��XlxVHYEB     400     140��:�dy/X*ـ�T���p.@E�*h5��ع���]p�p���V��=��t��
�,0�O��A�;��e�s[���Q���a?���h���:�~7����vE���g�J�� !���$�"��h4x�Cl�����ӿ����q�Ӹ�$���D�wzQ��-���:t��JU�x�ų�=0��C��3�ZA{�¸b�w�ܟ�ĜoC-���;~zw8�]��\@��T/b���=�Uu��'	�t�ݲs"$?w$��pqAEW�<��N��E� E%z=Y�iO�`p#�{=�����B�txaL�\���<�»XlxVHYEB     400     180Y7��g�?�����g�1�Y ��+N��1��/੄�n��Ed�T�����	d�ᆜ3��4W�#�t}��p��7����~����������5��E�jEWt���JE�S0C�6�&<i�<|�<�<U֥C������s��Kf�棋���U��b�%��TOsI�9�m����4'�̖6����!�"*y����x;�� 3u�-�	z*��%J�|�G���n�t,��g��|~Btv��1�_�����X+�w�bD���?��L�����p��x�W�K���t �tb�.��A��e�L1�G�N��8��pY_�
<����?�����ﾟ(��=���f��8�u������{E�|$k�XlxVHYEB     400      f0��#�G��j ����֔�Cv��W[}JG��S�d�D�'������/��' .x�+#�QRk-a���'p5ה��b�Hb����7�����u�x� ��K�|�z���w��D��-�`��ܡ{���ʺ1�d��K��⁵m��)�lz�D����m�����jk� 3�ۦ. ��3�W�Z�\!7�M�c|�0]����h/u����G�I7�*�8��o��XlxVHYEB     400     150K��/�a#O�FYL�A��u0w�G�WL�I䖸/؃�:\~'eI��q`K�P���K'��%t���+�EJ�2�ԦQ2y^�r�A��r�j�-O��������2qX��z�W�<�>D��]�Is��s_'�4�@,��Z{hWSՊ��5o��q��M��ś���d�o2�� �
6Uv.�+$�z�662��`��4B�+�-��8qep�M��=�v�7X�H$��a�ǘJ�uq��҅�`Tm���LU����Sĥ�A�z)zj�R�k�W[�eD�������e�*�pM��	��QĨ���S�b��W�!Q�ޞi�X�x�`�X�XlxVHYEB      b5      70��ҟ�3@7��&��pf���ē�@�����7�z]���,��-���4a�M�;$����7��@��Dm*;��ɫ�>'B8T_;�X��R�q�X����H@��н�