XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_�$[B�xq��,=�t�W��S!�BZw�ҧ�d	��rERs��B��0��!-�s������ᦦ�(�R���JrH1�d����'�j|�*���� ��}�v#��=��cqjz�)�}Q��
1�Q6�Czp����gT���NyxW��:��%���$�@GD�S��>�ƫ���b#dFw�b�yD���{m�^�z؟��&�_�E9����C:��6���x�����WO½b&ׇr�lë�_0�;���`���9c�	j�� ��,Z�VK�%]�}��U8�x����@_�=��4UC��bt�ʇY��H�3��*K�\���m�
@�7T �B�I����D���c����G��e��,*���Ay��B@�K?�Y�;�U��}I7��d��ֳr"�S���i���9{��������`@�1�� �*Q-˯z�_}ڜ?�� �yd�*��2�{�F��yea=e��e���$��_@>�E��M�<�S*�P=����ыIؙΒ�Lz��{�g��Y�5�Z�)PMRc+��z��$��L8��Q{z~-A��9���h��;�� �O[�^"B��A#k���g7�VVQ �}.}/��O˜c�\���^Q�L�N25t�����^��U��(�P�Of�|�KlX�wN�_��=������E�Ic�R����Y�"�s��Y�U��2��Jg�dat�q����Z^��U�ĝ��D��'��~򤵖�1q��RתaE�@����]��XlxVHYEB     400     1d0͠ր0��S=���*� ���,�p@Mp0O�����/[�'߁��Y�10��D�9��C�Hm>E��u*��>��4Ɉyж g
Aʅ�E�ˢX޻'i���)ϸR��10i'��#hgJ��e�e�ˏ!du�Z�0��x�k������:%�V~:v,�w�X0KET��]m��̯)y�<����Y$~ዌ��(-n�I��9�-���hr�/*��`�<�=���X���DEM� \�:�vm$N=�U���;Ƨ~18[��R��j67xK�����Ҁ���OD��-�M`��c(��Q�\dw��T�J+�ce�d/�j�rZ�I;U��Nq|�ى�T��á�#D����2�����N��)�R�z��T����"Ɓ�Tb ��c��~_#Rs��=0Wp��!����w��T�mU��0�ng���rgܿ��؂i�@���JJ*�E���XlxVHYEB     400     180h��?�'�qs)�1���9�� ��k~ ��<Ӑ��Ii������tO0����+^���d���H+5Z��{��k�<��4��!�����tU�l�3�d��F��me��ǃ\�(� ꐛ1�o�~�$�}�e��f)�7q?�x���t~#�%y4���z���l��
��[6^����~�%��+!��2[��<��^}ޕ�~�޼o"b7�w��i��E��צSA�h���r,��<s�1loHρ���z�7۷Nd�k�A�Ui��'k���i�@��½�v�a�L
��ņ�K��  1��m~��q���h�h'e���d�o.Yq��;Q�Ȗ��޼-�-�g���'�x}wLL� Ӟu����+N
 όb��p�XlxVHYEB     400     140��͊�C��_�/�'�?n:���z�/�3Ko@GFuZ�C�Ք|��H���@�r"-BK�� �����O�B��Kbz�Yݪ��b&���N�����\���)�8�FuQ<hΎ����:l�8Y�VI�Fd��_͂����j4�Z����/�[m��t6�B�B�Qh�;	�3��]@*���|AKW�9��4Xǹ"y/?��[�LѶ.�e��c;J��We1r�N��;}�ڂ��(X�|�S�/��v�`Dw��>�f������ K90�v�0"&�����L���.�l����k'�=�Q�G�S��XlxVHYEB     400     110��[ͽ(��j���h�H&`d�Ş�Y��?�ۇ�k��w��%���Gged%0r�qP���+��N8=f���Z�cNA�W��+�&d����l��v�V���
��s[���?y�J��;�p��vP��J��y��vr�z�Z?L��/.��q��T����0����L%L8���v9BGn
</�tAj��w<�#J�-e^���,Jy'E������'���f�D�w��Cjb��5��h�*y�t��,e��P�eݱx�/��2
O_��(�XlxVHYEB     400     130���)�W���`uk�J����!��n�Gԉ
���Aٶd�G�ԡ|���@��<����#��
��nm�ډ��m��$����|�.��ǹSg_.��4�p�":���MmR���I���~	"��{�D��d ]͟>�
[����%��:��-���2\����� �,����qь��"��F�����{�dBD�wXb� ���-�W LUsh�����"�6z�{<Y���Q�n��4A����Ϗ�{X�V
��@��֬��h��v4�6��_�)Ѽ���F�Lt�Cb_XlxVHYEB     400     150�[,�:!F��a�X0I�|������w��xØTM,���ĸԇx����(�AH�:��~f�Վ_J `du��1=q�Be�Z��d���4����vH	�IRS�Cc$�(�x��Iyp���">��D�I��"K���{[�_���B�`��Q;�<�Y�U?UE�`�o�OrT�� �Y\�Rs����h�c��ؐe���Z+�-1|@�vh�E6[�W�Tu�� ��T�������W8��~�n��߈�`K1�E�i�-@K���2<����SN�?P��U�l��T��2�~�w���B�_o���Ĵ �=q4��c߅MU�XlxVHYEB     400     110�ZI1��Ы�@M#����i6sfO���#�ҫVO�	�{!\QkfO/�Ac���O���Sql	�a�BC��Ih�v�4GK}PZ,)5'YZX7��b�/M+�9���Cf9�,�-���=�����P��S��E��St�8�����^1��A��cS�G؞�œ��0�	;��U����)-�(������/u�g�t0������x�sS���}h�g��pW��'5TI���صVl�� ���qԪ,s��h�J| %!(XlxVHYEB     400     1c0")fǈ��2���!���x2����A�Q��lr}iHl�Z��@kYgz��F\�D,�t!�0������dDz�N\�(]'��}/����{`��$`1� |�L� �~��3�G;b�6�B���{��n�$��y�9�A,�N)�jKط�Xȥ\�W�N!Fɱ��|8_g[Oz
B�n�vqx&mz�f,Ȉ�z:К� 8R��('���QEbV�	kY�����0!8�R�ܧPP�?[�{;i,'C;�_�d�v%@�� ��E����ck��p��$(|g���o�V��rF�&6�!�Cu�ٌ Nlߛ�C9��(��'����J��-��d9�����Uq��7З��c>�D� rCoS��_~�|� ���.R�_�u�%ԅ]�X��J3��n�*�`��8�[�
E+!ڜj+=
����8�0���Vw��PZj�P�Kv`ZqXlxVHYEB     400     150�.�3�(9/�����%���G��������1$��;�Y̘ca���e���ᡲQ���;#�>{5���{����Ckﾑ�4��Uf ��I�c�!���/u����v���fY�����T��m>9	r	A�:���_ �]�ϖ�GU�(N�%�i��gE�Pt��ܨ��8#J�t��p�a�5��mr��
���
��a+E�2���i��w!�ʌƔy�Pv��*�+H�_�Fl"iʏ{k��}���v�7�eDV �>�Z���o���oYJb�+(</���@;��os�r��+���u��LVc�j�w���XlxVHYEB     400     170����R.,Wŵ�D�"d���6;��Շ��`y������s���U��[�3��C��A/�p�#����Ϡ�'ݓ���
2��I(��@��J����Ёi�H>^@c�Ȱw�
���oib��*�k���a�M���U
&��i���\�9L/
s_����韚�_X�f:ˮ���y8s������D�����\d}$�߱X���v�^�Kz��v9�d!,*��k��9D�$�L@C5؈���{}#ɳZY��^��ׅ��*��dזTv!7o#2��w��;��M�qR3�D�a�(��D_jM��̘��E��'AUG�i���1�m�n�'8���E9جDH�	�{��%����XlxVHYEB     400     170�>�8`%D��v�~V��e*ȅś���7¿]
���a|>"�%��1���uи�O��S~c�~�ڃ���6BP�M�,��e���+#W��{k`�O���&�@L�[��X �f�~����V&DՆ߉�d{Q��Fa?-�K�.�#Y�w*b����wr*O�kTjh��Ou��x2(����CS2�$P/{bw� '�
R*WT�~����WVJ�~VHp�@���#ٱ���ktg���]å�钭Y?� ���,�|J��M�6����Td�8$��N�	�����nb^�_�%7���g�=Zdah��;I}��fT���'qI�o�F��xP��]��R�:�����f��GXlxVHYEB     400     1f0�=n֕t�mA	�r	���/B���Ҽ�g=���s���l��.iҏω��e��Ch��q(a��x��rmG�|Yڏjjb��S��$�n��(���?�>0.um���ˎ	�S�^`�j��o�4��+����VM7�#�ߖ3b�z�\<�q;�EeG�Z��	y���K�6g�?��(
s�|-��G(B ��d�W b�X��dF�R=.�!\��Reer.Tpl��u��I-�,!��6@L �:�{(�����(���6�����۷�3֗�i���n�\!>
lԩ-2i ~8- �xX�Mxq�U��D��.�f�<h*��sG�S�����k���+?PUl��媬�!���ޕW�?�}Zyh�ͼ/l�i��kDY�"�&�U�1�(l�95��-�G&�m��qؾC~k��W��T�]q��U��3�1f�B��a����,w5��L\�x���:Y'�鿂��K=[��To�!h��3٘��~�XlxVHYEB     400     170��x��\�u��L�����r;o��J�X]�k�S�8Yf���I����B�D�h�4�w`-�����ۥ������7g���!m��}s\�F*Q�F%�(�/ �e�&���Ź�I�@���C�⧊��/Kn���\-gi�Nl�K;baYY�SO���p�.��])*�0k����px�\Z���Ë^2�H�z�*����;'tD�/��q8��&�W6I��؁��	����ޟ쌏.^�6�����Z����>j�zw�/6�N1!ß��J��$��nR��+ii9�(�D#����=�i�.%�}O�3�"���kô{R��cB�Rb�������;�Vf��V�J�?P��XlxVHYEB     400     190	������Xe�<��"�O����cAC� �*��q/�F�M���9�#%� ��q��:W:�9��
3L@����D���B��	H[^]3�1����{0�}'�ʑG6�GE>�CFWm=��(*q3��f�e����abw�`�| r(/tlWݪH�B��N"Ki�v5ל�b����-k)҆�do��c>! ��c��#s�4��oO?����'/y���'Y+<�� �Ƚ�=�x
E�Az`��WJ��g���bū$~�ڊ��Ւ�I0dS�n��a�z��ɢ�D�t��ˍ@��ii/�jn5��8F������t�����=s��9&l���Dȿ&҄���cf�Sq.�Ƒdi�REӭaX��$k�n�C0��f�TG�",�x�ĐD"��XlxVHYEB     21f      e0��9��Wr��^�J�����Wk�	��kS������p��B���	���Y��}� ����k��'��@ܼ����q�l�O��Y�[��nћ��\i��T��� �J�G��{09pL��^2�-�Q���������nV2�r���(ǐɒ2*_����K��0j����p�&|�na��g��$]���i���
�7���*���}������mZ�l��