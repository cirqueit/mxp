`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53104)
`protect data_block
3m78KoNT7Bsz2RciJrRxQ09gxIQSprPc5Vm0RpXV1b8v84VmmLahGM8aVxl2Q9pF5+1hvPOz6mV7
+6z8Um0qim8qSfrHUHmo08NUIVilvKJZZlVh+THUxHjtZwiThohgLQcJwPR+VP1QAGtoBqKAuqXf
5QkVj6QuVDLr88R1BHmYnbs/bx9TG8ebKmIC6zojvwwKbABGNOGtr0M2ASw9QVky2sQSy+pCxHr6
wbyfYb5U3OJcPYs0GkW7V+u555oDKc+46kRPmHB63I8zlctoVxHuoy6r+2ENiwfiHcoZxevQqNxu
U9bocsnwcdG50tODNorRG1pThQxjUj4CzEwLDZIhc1eJulWPQMfAzue6QR14Gnjg5eU41s5trMmg
4mzNkEbXkH9ym+rIs6OhCuiDyKH+H3RAe/dnncP/XzqK4PUovmEAuQk0UlyjXK6GHWWbRS8fUAbD
ds5CGlvlTXo9shoBgSCw8DslISTyu/p3t804IzKSbfcWddvRmq7Yw6iQ4Gk47L3+xgyj2+vFN0LF
PbVzPtkUBMBZvuCTDO5RTmmdhiI6b/xylhZvBgEKboxijqLhMz2cBDzKYVCX0oDSpXTpCrLfsuh6
TRrDSI41audKa5/wRyQZbHBHIw8b1Po9JgwuGk3GQo4JzmtGcs34aLaJxodyKL8ban0Br7nGbQFr
YihNnAureJgqUmJwgdUxVrBcs4CeUsEfTRyOXgQB0V/1TUJTLeik7AHvNWXWkPx2xOgbcB9oXFRC
uEoxJ9Nw53bIWxOJGBflMEYjx5SYbpVsnWP1+uki/cQAqstOwnsmpqNSqwgEJkd4XYvn5kvC/C0c
imNr6wWnudfOcc/j2YctamtE+GBOIIKBAzn6Vlf7V8M/D/kK5UjiF/pvve6WJ2itKjKFD6rRNV90
rA7T2mCeuiM3k3u8ibT5HQsYJLYhucwm8b7nnreEoU+q7D0Yscozen5F2QpLDmnwoIE/yDb5OdAA
DlkFrpF8mUYeDsW0i52UDDuEZ4EQ7i6/gLYheow70Ciynfp116rZoIwT1d/BisymoK1E/7A91eoP
YN8qY92+jkDaoDk6TMgsRE80Okug5HAb9FEIFqmfcbvPq3OLdo6BcTKO3Z9OM5cmAYgK3V+wzDtk
tbUeh6uORKN3wp2H7qLzFzJ6oqB2oD83gcV4Zu45kiFyMFEne0w6UIOoBOWI9Q5ww7eFz7aRtL9P
PzMoyRcDI/5HAFqbqxXQQoBthMr5jeMbq0K/uOL1lUcSV3EkwBUwFFmANBjga++4MDD+2kj+8CVo
aGJ+NWK9/7SFRCjYxLUCSn8DWgz9K3l+Ttj4Z9yXs+FDcuTUcPSjjXalCdxVzqbZVyB4082Jf5Mi
JGXOaEL673IyzVM4J0iKDkXp/wO0Xz2jRrXm9wmd9dbyIG5BVg2mFQSjpqBgBQooSW33irNS87RS
MVw7q0y4rFWGWGMvVz0iRMsVhy8oXj/l7jJas5bAod7BvyTCRTKgjxRGY+Gu4j/NZQhq5FZN7fXb
g38nA31cXg+5U+eJRS2MhiWoqcyAyFqO5r9Taig1kKcBv6hC0rBFZmErD4W54ZJJJZ1oCxLTpECs
mawHxEJ++LDkm1CkQHHkQvlAGQFOYiz3hT0qTwhR5IOWKsbe0ix69W6GMidD4M5Gsqw/xuMYN0Dp
oU0Rps5825J065YQk04I1/XjFva1eQAbykAeUGeABOPbCd0+naOyLxLNJpGsYkVOtaZ5zKirk/av
mVdBf2YuhnbQUonWeg261Bok/MqXPVaD3CIRnKk5rTdpGd9KI5RwFMXP3fRm8lBhu2oCBUJIzuOn
CbTwyd5frdDPUd5hA5ks+5RALuUpm7lrZP22yuBsVycZ2rw737nzXDFh2UrDUx50yhg3v8Imtqwv
L6K4rA4ceM52HS9nhh7d2UYnuUllq4hj3T/X4zcEne3pScXB5DABTBB0EdAvFigKCVjoV/sKGu8o
nCCljY1s2LvZ8ke6NzWPPXVjx7jiNzgZeUSxLSRk5vVZF3hRlWDVxAoQZzccgORBeZ+X98iTCmIB
WPvovQ+lpP0c/Lnej9ooMe7I/K4/DuKtZWSXg3zao27sb/8qCISgxjlhn9f7+dwXV363hmJi204i
JIY2IyreSIFGKM57ajZ3F0sQjQChvLhKcG4JwBJi8KzFptXTIKitQ0b7ezKlsu8xgDTpnlwTdhCA
s8BqLySpi3aC2IFwxpwk122u8TKF1pAAOaMqebYNMKvC47PO3+7y3IF0J8+A/ZwTkYavd0Jrwm6M
vP1wp52GNJnvz5vhdFmTReMLv2ZxWl1VMB+0nrxo+faA0w/38h4TmabesKqpgYwC+vqzixBKWzLx
YymrGY96DpTxgL8rthGbuG6C4/6R4n4kYziagIwVYIHlOl8rgqZJhmsYsNc+H4vjyqzEyr18ovTY
bx3O3SaKF24QeSShyB8lVsdWnirgucfaz8eNguohVzQ/o0PVJ5394FuNWIHe3mWOK75qEINOSQKt
UCXjhPCbMrOyPSpT51qMbzauAyHIR0xuOIYBfObkWOiXcVgHfXVTmWJT2RJpawd+WCs4LlCPf3c6
Oi6Sv+SnMtVrHtGS0kWESZk/TuLWaL18JfSfpe1qRYC6mrq/aysaBX1Pvd0F7mrYvbMlaLAl/aME
qIX1QVjeeDEJQTAMcZS+GR4zhYaKjlx09V26ZNy8it1RMNI/70fSKe8iw3kBWFWM5SlYh7JqBsoT
WTu/1wlnBUOuj0DuuPVXRCPfMqWwuetmFM+jJ/4BmOkBwASamQcVqERH2i3RYb8VeM+RQWPckAUQ
AuIBhh8S5vVjoUxCmRbc5nFteF8kDpqAQOvqcFsNO3Ft2AHBih+9jpGED2VzF+Acgh4yrfeY+63a
EHLVNmhF67Lic8jEnMaX1jrvA/vz+fPd6IoalLnTiNls0a1ZuT3LJtcZIbtShGtpa9gmJRzwiG0f
EM4hvUT/5E2RyQHoFCpkl+akRPGel683ASuLma0jbZZ59oNCS775O+HdornOgZVh57Zcck2420rK
pyZOvk1R0rdl44UUn5F/qnV2Iolx6nD0wO2Q+ZBQtIlbwBSffq+ZlWC74La9U0x29wK+vM7/RNAj
S2XlxXlm9h7Olssw3D/s5GX2MBO8QTieXPqd5z2fW+skQCSMhTnhl0UbkVT2Y96iTAobJj0wdEZV
VVm6kgkyqLivS5INaNI5hO+hDF8P+M8iTiZVL2iHkmthxPC4mb82l3GzZeTXE+eVjJ2Ou+m+Z67Z
gd1Pyg4xAuMik5oQT6Zu0Ya+Zer408+qztVAb3kAs0JKG47IO+Z+eGnGeEqUsnBRodTE0iO3h6of
ha5UeOg+pOv7syHWJ83U3MHQrVu5PFOWKWiAljaR7uMQb7NmoWoaZV0iJxi6G+s81iE8hLlWNSAw
6KpzsnLlmm5YJ/G+CWE/R61Evo0iePuoEMov9ZbJZoOaK+SawSmavNpnmJlZqMPu0gO6LYyVQwAW
O5md3NhXDOMFjBOlH18nUrahH7gVLxxcHn/b/7TutRRkM8kZE3BP+TT25fGi5f1PIuoj5E+nIJci
ZALhZw3sLndYrYTMUA2OGiFlLI1NxWY/Jqqj2q4ZE4URdZ78ysgUTxtZBifEj+ywYOTtiRgHAlEg
13wcAzYbZDcRzK7gvjTvgAMwgxHYijIXktN7NpGJcbpHadqXWEn4epGF30sHqkJQfgzZqD6m1iig
FW6Phpav53KwKaSoqojLPWWThILLSsddU3YNH4beiAgz7vGv4AIKAjptTb/myVwOQMc8ir/IZbzp
uSrUsd0rbsd10JAntqZE7VpUsWqvprbEJa/DVGvNwKKzNA6khktr3aZHmtfLDTZpbB9HiyB63zQf
PHzsOeRnPpHoMPfnLd6x7hCg9BcIwAQzyrlqTf6CUCuF6mhCTeYhfeozdK3zwSxwH3XefC1MHjjv
6XcT0pQISkSBT0AqR4xq+5zkIA48OhA+64fCYh5D+EFmuae24J7/O930ToOrsv1g9XNvZw0l6KL9
65ST9T247GzAUqOjWXulWs+8xiq9Mf7eFMn5ay7p10TcrVM8gsdQ36FWPYQSvgXHuf/5lvUKpaUC
yZVWesuE19UFkdIFKHpQ0buAlx99BsTX82WmlJtUDTlWJ0R/du0Mrbb5zINwxvWNTvs+q6qpOU3y
/HBpCv9yNoqits02pLMRgqsKccfVrhvoLmVAMLhtDs1AcdKF3qBuzQcfJvwZkvvxv/iH0e1WwyAi
4SQ4B96485NcsZdgggFdk9SEZRj49whOTptolOAKKzaYTHR3u0gpvKQxJwZzKVruZn7Urplj8AWy
ZLNifcRoqP62ZL1OAItSHEVRN9UwvDWy1N3dNO/GqHcFBmS4QSWex738IgrRgN8lfG0pP0O7178q
HmBmX91R9wLZTce3Fp++L9AjkVGxhII4eOHFcrp96ICdrAKDvSGOH9OFQMxJsj9/gL/lddK+KtwS
J+U11OfhFoRao88g/FHZzIO27Z+T5pSF13SDpoXbupdZcGYuoR6wHxSS7y1IHKcqladaiwtUloV/
24Y3dmJEVkTEAPZ+m5V2UR5wdGQ1IZAXEyaINn+6u/sw9nBkuOnBqcKYByCI8lJLnZ4tE5wNF3/M
tCTFU4XrhlJhyB9h9jDL/PYKTLdIS5H6YOwXZYg0abSW4ie1lacuBH1zpgsZ2nZunwOjREcnZ7/8
Q8SZ6qQvfm1gm4A61XNP64ZvgQy4iyDCFDnt3C12n8D4LmTSHEjM5Q5Evq59+wvsQVuxGsC8snUr
O061wuFH3JIQ+9OgD/X9SfAFKJjxJlgxguAP5Y+9B/pb/TdGsjby4MnuCD9mEHnKr52iWo/Xt2d4
O92C5thAh3pbnK5bAXYQCPSPUpdF+OzX3mFvaCnfhEEMvY5sgjeGVeb3YOUISEgfzk/C+uGxfYhW
h/HfSuvET1J7ZgJwpyGrii8sKtUIpFCnu7+Xft3GJm/D5Z9aK6Y0vRk4grRsQMtA6Sfp5v0V7aoc
OjMp3B5OUTDXAZu4sAZx+DiGosxjPAIhapV7CLiP84MgwKgl9FXzM8LO+DnjpPHzAZ6gYJVuNK+w
pVAKEkW/GCmkVhQjtNw/yzlXpaqntTsYMbOmwOHbYEvGUX3IWdkyd1wEVbPL+NvFmn7304GLHnos
WtNKB972vRNi330JcbE7lzfLquJnGELlakl46jYq6jUICdUUrxD5rcv0OCXuChgj95pb7w/XQVo3
sTVu5WRYfz3io5xsCHrk38ja95+PkmPCLVV6MszUGk6UlCnIaBoPO8mFB+XTdJqmyB+3xbgofoa7
1bSMkJ9t3BdwaS2Xj61TBPjXVyeAOTYzlIYyAc22cp8AIN4y247wYhJorsUg5WCsZH2mCuUUcFYC
Awp4PBJ/zqSol2GB4lpmu6ES3nYlpNfG3h4fYfEjhmH0XDVPw5Igue2/xgeFuswA2My6CIg2+dNI
06KqqEgzMBztLx1uNHQYsWC9KdwOcgZmEEhmM99uemmHN0uxtRgrqCgXXAGgediyootGvibGX2Dv
P64CJeII28Nva+NyoKOlhNGnEpSOKD8f20WSxQtwhOXWIcJwk4V92OXjAAKvjaBDLYiNDPnEmhVr
UnbzJCar2H2988B6v6R3/ItjgkEeQLoJdMqKLToE1CjR03TcmmUNxGfXJG3a/AHvJyo3KvYSKaEx
sPveAayUkMNRQY3JoKBB6RqAyEnYLSMx6SJnwLg2Mlen2esQ4BO5qpyKMxMsfjzfYyF5rVmofiiy
XR36ZuGARvw9mlX7uBXDbomQ305TeeXvA9NC0P40bdzAdJX7r4uj7jh6uvLWmMqDjLDkpmgM7HI/
uoJQrXrG3zdgYWJmQ2cnCgMF9WsDGowUz7sTItKHGbqklauJ+X85r++Y8DBmGH+UuZnAPMwp+G5X
Ffwy6dmShw3mp8F/xwo3/eeUa40VPmjnw8vTBM6oviG1+rZuCzeRtjrp7w+WJM6wheOhlEY6lM0d
HjJMzV7Uryh8gW9vfLuWc7u+vCwzSkk7dZ84qM8FqxN96Rg9+1iqcdPqmi7I2yAdbgX9bSd9si7l
LmzI7x+eXMZRkD3g728zVLDvnW0OCuWS5s7uEmxeV6bJejd4hD75KByXxbpAbMXjOFBZ7OSr6NLi
zTWcKFylEk72vMqYwDrhPPGZQ0sSaS0irLHuz3svOHS7vY81DLlYTPROH3VbOBzPWhscRro5TDeZ
cGwRlr1XHyxU9s5Znqcy0HnwXuuEimJUBbLW6acpH28divFny5pUOF/s8x1bYFWp4dIxB2Wgb+4f
q9Knq600sTMygHY9OCijAP02h8npsFxbBRCJyYoLO81akeodtWP2oXfcnEe8asOUCZueXVIAWTGb
knx3Roj8XsF/6zqnZydQKJqBGu0OcRuCndbNG/5vwoqh0DJl+odooPDRZSIStUh7ekhV4m2+sbrn
iDQpE3TIXODHlx46fpq4gx22ByBez1FKt+TkyOJ+HZ/wIxLa/6hEXcZew6UCOTbQ1thomcKVciWN
Ly8/3Gl1OPsRUPNXzZKkbIGokRCpTGItYpGbWymF60skxl1ZDVuhj6r5nTOB5igQY51bD/9MCygW
OvO2wVUEPR+5XkNEUhkhrLoFZhoKuk2efyfOsLz/85UadaPVTZGWCq0P2xTZog2//hSly9hA/rNw
YDw193VMgMTAjhtbNq0wLd4/aHlKDBsqKq1RXx3tSlZ2z5Et/FZL96x5pmsQDnh4rTpfIBirnBcc
kLV6fX6ASO5V+YiwoFT7nQdEYcqTGa23rlXWmuwlwEiN4cE5MZm4pts2+qlqRpW5Wj2fa4M69KPt
Y0jYpNmXoQIZHgSVcVLISlZo2EXrRumrASOPd5QLvghRI+M7oSNExdrP8wMXggiX8slxsbU0GOkn
uWjnsTXhIM9s5P8iZSUB50C+xgMN4MQ3SVkdL5hcA2yHQ0BBq42Aq95IpuKfhQNPy5kTu3r/fQp4
JMmVQRI2HdXm1WqHDsG53cY6ebyIDWQQZpIDzwXdb8DOpf1zT3WzEy906OyfUUL4reJg/+8UegaJ
Qok9hJPKsozi3Ro6gP2t4yErJqMZKLaQGjKnYdjEugmpnUvH2flv/dbc08pHO8Nhj1BjMRRzYPdW
bev1/gAUyx7ILb1VAHRJwN+7Sd3UkzyKp0/fe3JdcT1q23v/u2EIwBRNa5KmQ92F4IK1/UICnOMW
ujgLzaw7PAu0NfHRf7TlW9eyAQ9t5c2wf14Sb5hRJ6SD4ZkHclf7+YsTjAH2EhA3+CSipK6JJYp+
M/K9HTCzPwGuazdAugoLnws5pTlbet8Ja5oQBkXLFw/edTe9Dw2I+kjMZfjfgT0DqpAwQN9ZXLvF
LtG8Bdt901YrDrWIWHgUHEWcWxfq2FerXw/JNbRUf7xyQeC5f0p37+tfnb2a4iYB5yvy0CFyHieW
sDvKTqht7GbhyFsbAaR9Uq2+pPgiQkdIuYoYfL0K8q3GJSRIX0j+QEIs2xTnbW6pixgGb4P8sVWp
tlW2RV68JqrMeTqsS+hgAJRktGNlb4sU4CYF33VNYSC1j7RM79WN6SOQZjlJ8dt7YXzAoSEYPhuD
gr+8j2+PO83nig1wIrTa2VcNIf0493OMwocj3M+g4PUImtDan56PGD98g2BNKWOCv33VH2koy9zk
2ANIFIcaQ3uTZbWL/WY7AzVw8XCezwcKof+Cv5lzy88h/QGQLlDWfg7MrWxMVko5rvi4Tnr7PWII
SsGoq0SgOPFynUkjsDb35qxXfQpkjTzmbDp6BI+UzUjSgqdInNa/bTjwCA1M4iWJ072OONQsOmeM
6MSHj3vjrbqpriVEgwUlIFrWJvcnjiUmPneOdKC28HByXUBkoI3/zMt2SRgHq0OawQzy8SjYAja3
F1r6v3xl65dVw64V9PG1naFeR+D2CYQbazYJ2G9g9Vj3kF89lvcuFfQpxJy1PJntsKZ07FXKDslR
3Zp59MdcBouddBnX0V1+ecw3NSuP4M7hEMDcJS2g5AjAweGBH/6kZc06jXPG8TJibIca5bdabulY
3sajSJmIL56pYsrH4+dTbVVJ43pR22UOq5CiH7LAjggQj7gWnWoFTCM5p6RP6OFhKVd5EDE9oOY0
U/ODETDYNCfsKPZID6PpkweH9KkB+ub4I4hhCjRNCQxmviEWGlRik0KCf3jYHueih17+c79D+E23
phmAMeGFrRg9DrBG7WLPLzINz8H/FySure4Ny5Dj79sbba1gmnicBtrKQ8T30gWjV1am5vh4COmG
O1lfCIF1jS5aSV5bYhRYDKRDx52V3hbVW/2t+TES3bkK+a4YJu32a0FcOsyV78APfqNKpMQFg0Gm
SOq84LB3RYVldyICOwz07Jc74kA4DlIxvU1f4TpcTqRHrS8EyqiSBt5j+Rlry6qeB10vqP7lOLfx
a3rQ24hScHWlCPT0fw657fAQLSW58TJNyUIS0MA+5reEZp5dKUIMX59boCZSZuiPUUeefhz2KpK2
xbluYCBT4LIpG0+fExSWfUNEfu9VxirckJVVHsHHnomorNDd6cBFA/wRTEzx3S6YzADMgA4Tydy2
eWL/YANY1DDfl2JhYFwlLLlutR/eD7rlri5S31R9UHYIQ7/iIcPAMy4vWBlhfpOJc4JVIGpl7MYw
OKube1VbBXf26m6WLXggaKRnSKNVTR+qwu5WuZbLxenmcuuk8LjF04GcVMcRXUTL6B4pZiKfCQfP
Ul60tHhb2RLYl7Q45KCjna7zy5OQYzzLNQcOpRaofEzT9i6BFgg9wEC7jcrRkClY0yX9m6qW/rN6
mXhuu0rYD58ha/9w14J2rF8iIqj7rdqDitGXbwgTQBKi7XY6sNts6PigY9/qsFJcAPv4DhkHUovN
9cxbTPMjRtQ/B3pj1MLpkJOmqKGQ+KgZRmGUPGOwe9mn/i6Zkbv4Q3xe8YVNIc6LfGVZ6GVQfkAQ
A0uV0ECYgJRxQcRBQLOXnhuAk+FWaWg4Lep2IEm8p8CQ1etAEAIF6LTBgQxVNheRD+M8joOqY5Fq
xmexpF8N2fhTaltsbeYEg6jgmOvk9KMlLNmuqyUT4NLhWsmIH6njjfuVOgMs0SJMUYmh4JF7FB7i
RdPe2mGEwJtYyB95nnt/NSzg0e3RuapMYrxmw3oHtjL/BGkuoGDvA8auIVMAiYCLznBGt/v+k5K9
Ho9uW96UxKvoDh4t/tECOmUh61V8wLSMEyIPdtDmIJdS9SRuSxnpWcCQ5s7VhZ86JnyBa4A6yqjA
4P1fzrWraytPVfS4MAStwE+fvnEn3MHXK4AUsb4vFilhQfKKW+aVeqJQ5XkneZ9ryq0YFvSOEBGT
QVDMCOaTSWWsH15ibGI6NlQ3SvGh2T7PeRd9CKTwi0tPsSQyb4APbGv8JbY1iEolEpP3H6VLXj4f
ExJSt4Bh+VmpNOSUc7WEWSadpQ2J3tOW8zfCzhYd0m1I6yiKLyJGRLKvWx4qOeDyyMF6lSb4r5uu
peRZ/e7L6KuwsOUmesUw0emmqohQwZ8bOkoxbwYittykWy//J4pMxbx3M5ztav+1D6YFXYatnxTV
l2QAZtgIK2HUiYB3+zRkCxGVTkCwYAeFrQBEX7vUMjyBAba9JVkUiGW180QcQ1waSfVKacWm7cdR
KQ/e3j6S74Nq7LTJM47/A3o4BASerXYui1lPx3I+GOfq0RkddSR1VadU8UAaNyNUIFzSHm8Ai09F
V7PKEXjw78eVH8mtDw9W2CIL5qtKXOYZ5EzCmJNvh1tPXT/c+BheYDXroWqzYeu75OpOyz5tX4ZT
xD94WghYxATuW7jum6GO5Np5Shall5XCnVb2ga6dDexf7/56GQf6qAjS46V0WKzXwDso20mvp9Q+
RG2aVULSEHFHt4nwkF93JjB2yWhmNHj6nZlcxnIIcK9gdf/5NYErNS43S3jDnI4sTQA945zvumud
uOU5BPm7ucAEWoc7hjH+8VZr+tzUHjOsTMb42OvPUHzU0a0/zUylk2ce0t+PE6i36SiUrQ+nqIoF
SeuFjsuQScouaEDV0x0+T4kKnnvZ4MHL8zKP6ooYyq/1qGoUwUq8ioueKEhmKL2nlph9rqs1YW5B
NjaBSFeI41IczZEQgaQRJD3OOvHWnZIRFqlOL+qm6nTd+kA1uCc1ICKQxkx73T2VIdBn/gXb7zyK
D1S0Eecolz7XEL1EQ/9aMhglyUws0jzM75fmLLQSjMpJK7h+g5PdFIG9KRx30mGWw+a3hqvZQvuz
aOJrg9tYi4MEwRkPrcgJDBi0c93TTE6l5Px9RiLQcI0WeE/SdGrMxDP31JO75bUrxokiH4lK3Kgq
+kx+H/iEnes12wUTZeZrUxMLbvN9V3L6tUzEAUw1BBPD3PNwWkt/PIVSvHvIP3EZA8yr+QgN6AlN
/ZyrdMT0tdUAUn8yGC9m3XtuPGcna/dFCeS0X9xTMnEseld+Ghqq0Drk0BP/l2B/xEBFg3WIwOmW
upxpin+84hEbgF59d9vptGZ6l8uQsN4bCg5I6ocDcICeR3bLUS6BgpbHbmQnqkeuy7ZDH4merBBF
B+2NkTsKI+WaF8ELMhUDEW2PM7MrkQrp8s+UGJklYpcp4F4lUCnBGqeMEb2Px5pTz1pAjJpUnKxU
/kvKC6GYZzyFycx1SJRJLybkeKbX8X7sjiG2dZz/RVjSJw40i6lNlJaJk2a5WqOBjp/Ckfru/xsN
sMlvks5TA994nlzAvfjbeh3G2tAlcLd7saXZwMiIurtHh9zE9EuK06Ov8dMO59tOfaNkDUMlnU6Q
60dim6hrreZyeEvFDvaMPZZwhp5RcSUU5syFHhLiGB6mUHgdppbvwrH29bJn8MZZu1neao8lDch2
yWP/ViYm9/CINwEqWBK/AqjTrC+DI6J5mVwMIIAjDJaseSutzMWdekb2oSkMDATYB08lGu6D6FgM
7EPtzC/1tBBU4WBYo6RK/edN+IHvS6nre3pnPKF34YZr7yoxYXj1BKYBXASjEy/CIUuY46uoqY0P
DxUNjH2M+5128klWrIpiGHL1Kzl76oMZXuaWBpJALC47hiDpgPL3JQEzJEZz4oVWPhIPnVmCBJ3D
xgu2q29gORCHe2MQEzoo2D6Ms8ZUfFFJnKba8OazapW3D1zq7rc3BM5uM92YGoqikgfrldy38+Dl
1g687GvkiKBaAdKsXSrWzIOPbhs7OISz2mtOSUd4HFKuJuy/Np84UlCau4uBndE8GeNgwQBtJH3N
nljouQf3/Ukp7dswb2LoQJorKLofPhuceJdhE9m/7cE2ifjFBL6f3auGQBMZLEYebcnygSFQIOKW
fQNPV2osx8qKVDcXQF08dIAoXwMjZXOzMQNn2ZzD5eDJnUPfXmSVWrsgB7xyj99S9a7/SgHd1V6x
YJjD7R3Lw8OB0Tq+PbvXUitYX96hXcEQoz5wkrdUNJVI4tVhT2zwFkIpDHxeNre029D5+Hcpulqd
8x4vWafXOfbSri6APR5B5n/6xPiwh2YktFl/7cPkmz+Az/ILKk+PBJfa3WvWfq/AqydD+Kzxf/Dv
vPylY1OI53LNkj2dhnuMpXkjlFgcYe5HcrpjsgIYnq/3zaRFwNW+i+D/o5O6D9YYHxpBRgpBTQKP
ZXZXPYgICYH5z7ez3I61zsirngHNUmLDg25BttPQxZ2jWsbOAC4yKxcnqrCPcoYiAv9SGuXcFnAW
1ThvDBhlFcXFF1AovFmrTQY0Rsd+/Q7YrpaILec0UDOThaUPWWJym9QEKlQy0OjTEqhmBK28F309
uU8LHUQNY6Ss3xuA/OLe0YmsuzxRg9Ke8Klb2p7K52D5e/Ol7qun/RO3sgM8z0B1Uc03K6IOuSjq
uV6I8fSENhtObru+pZFo5Be3QvpueG4+mRbwFBZOjh9w+fMNF2CQVcfkMwvCp7OPR+QbMB3o5J+7
8uWM6bGb7S8wP8Ao4BCK1T7dcjBwmGfzHpvfpE/RjgVOWo/W0/pOg1GFPPHnQeVzngr4UWsDogrf
l0FWKf2rKkAxTM8OgsZGz8WfyJLG2xSk2rexJ/zQXH1MEcROe/GKIVlqaIYgVhKg6Qcd0np29+OS
/aKkZZbSlH4chfBCciZ7nSvwC+B6GvBkrO9EZhYPGDqWGylcE3kg+aDNHvcHtEOIlZnpXdqknhl7
NSArD2n+e+PWZx9sN221A2Utdww3FcnyjM7C3DVS7L56W7SrQI6gynOHr4wG6zv0oMltv/qCXVZi
rdmqhOQ4DqSjdRuMvPqHyqTD+gRW3Siqh7jWtD3va98rN4G9EFgp9T5fq6imgGkih620TEd8gttJ
ny6piyyN2OvvU6N23/vaTw1ogr2Q7vYq7HvEfvE48gYGdL+RFnO9F7Rm+ft0+KN9UWUot2disKPj
s1J67MLH8aHhiiTE7rb5QzzxqFa5dS0UqR2wZTZ9mTzVaOHhroEpoqu9PZBft2FR1/aH8DHvIaBw
o0ivcNU5SJNuozBhgkOdAejp04N6imPBtmBmNJTSpBXvCvZK+O3efQ7EIrTKOKZsgqFOw0fyUvnm
uk1ON+T/0wYvKRwGjrs3n3pHWxGmCwyjLsQijCBdVWYjX+nlClkunazG790TqEC16sma8/9qFxim
+ma57XWlt8pYwRn88M511q+mR3wYdAV7yF3pyuBZNfx7TXe1OM1oyk3dge4XusKgD0OGD5BNFf/B
KEMhfvM/mm30MTdKe6dKTvosE5QC1Qwr8bFOFMBSdLVYyye1mMGJAkFPHUxU+LW+WMYit69gt6zs
HgxDk/+hU7zElhlK264LIf8JX05JsQdB20Vs04pPNlNh/B7PIY+a+aHyLPjyl4odVB1pSCQUMFgj
ndt/8ErStZdp7NPcPs4UWUJ6uBd8lTO7YuFMy8cIXth1QO9/t9vZzu5/pGeSfZSZrfFUnvqFIr+a
0hL6Y7+FcEhyk4JY/arN9bpq29k38MtaMQYshrXDGLxyGFfMZS00kQvknq9zlnkc2IZ5fzhh6DDT
ZLyLYtAdq2Z7bwvqIHmxcVnsVMZDqL2qqQG9dZtI9fMc2++lesQ+e3n2/L++lfr4rrhsfLdLX0Fp
Smhiz/QlYQeBG+1qvDzYMXWZNU6+f08RZ2J1q+SvKxtpAsFUxJKmMHfYcyzo2gij7mS9kb95Lino
Ag36EbXWhN4UkBTosd68FXcBMc3un1FZUpQtBEk8bsBubIUt1aCCOwYesmfZGNPMhBswB8fQwKXp
y2vUzrUBwji+X2Ljkt7aioWBQBUydJqy29zi4K/xcKPvH6hUFRXH8/4kkv0LUWASujdTqgqvr7fs
XVZXmCgCreU8sVrcE359s192y/sqk160XsPRGZBHy0JA6CfODeRGKzkJhQwWFGr3Fvqi2/gloQ++
MELLTazQ0ulY2E8xqo9P5V6vXI+PZHiqLD8yPmEw+i6LRmSGVMuIsPAotFhViNrhbz80XD4dU7nJ
wN40c83MrpanfFEOaoetbEo7GJTVCXP3OguKeGYTzfWKql2SGgGhuUJpci0LMKRQzN4/t4gbeXNw
AXSH19fcd8p8/emMul/OJKb90xwNVG0l0hANWRqWjZINlFCRkzCAbsIdVfm2ujZQT0tqkXR30XfG
y9LLrA5nby9d/Jc0GAtKM6LlhplmVwba5JmrEeXx/MoCJGWg9OoXUZo/ZT4B4fvrV9FqUClql8t6
vJhD+s5CDP3a/6vx9Q8PfPm8St5rf1hzFhnETJT8IIxWL/URBfiQqX+1x4aNXGXsBR2CiJiRDXsO
7nQmEQeHkTEZxZ1hcm5Zov8Rp9s0cQI9C21UZpaMoI//0c2YsiKYiAfj2xQyaX55KF26PSK3m3KG
itXD18VFbqWRS7M5rAE5emFNucxw+YiQ7DsvPA+mKZeMGsqey2J0jM/fXTsjL1Qs4oW+akX+rIHD
AXglmlfU+qdEsaDeNUxNMPgtQH7/bqVY4CgVtB5hxTCGPoY2/hVv84kpBvJ1zloc9OsMzmzMXY4J
HXELtMuGF2UFYSipbzLsemL/uvECCYs6jFZ4EsSs3nWho8n5WjybFoGbWWhjjneVHUGK4WJK2sHK
gV3dr7ocuI89VkT38ewzjbGQpxV6G6KXSUN8Y9hbpD8aK4eDjz/N2ZMJbVJkk9aOp267uYcJQgUY
tsO5bfijfqg5x71ZCUKkI6j2M6DNxO139YT8avF/5Z5pytY64vGzjMQirhY6xLtONMjJzubIDX/f
Bh3rdXRfIQMspbGQ4hOY+e/Y7rxvQQiBFwXkfeQaYe4F+aQJbJJxQLXo8FlMRkWAxlco9462QAN2
dp+bGb6mKCYG3bi1hd8YQQHO6NZcS3G4Lm8ps+8rmuaIOc2x1hsdF8M+9jhhqeX5p1RIzs/Z1bcH
q8/Hi6ZWUdZ8lvx7JQxeRNl+CshHIGdSfsmkYms7E2ym7P5zOUCvjW45XDENe34nyO3nxqJng9uQ
lLkTx6IyXP32g9WBy6ZBDzA4DGvw0OK73euy93GAmleZmysSaUbWu/s5aRfQQGZ6EyA0dyqqrO5P
afdSlm4TD19efhb5tU7sPLlE7599ARmTHcUeDyW3Fd7HFWzpH5vbksfoOo3Ljqv6D0l1V6Le85o+
vrX34eprek2FYzuLEl5BeWcogW0ezKtKh/XN4poPbKestow/UAXbFL+oMOErEsZNYZn8laYQcj/q
kKVRTt8oWRL57IK01eLm+r6VMTlCCqFfDjSg7006fDZuzwv5M64ScSGEgL3W1kvcyFOPfIvg1Q+7
EriekSRh8PFAvsSu5usKDQkCjfunKvukJexxRt1UzuKHe5+6uBUb9DmelkXLui7MGTqienbpoEP0
eoeLRzfk1AqY9+keEipr1jGMICHtOYLq+lzhdndb6byOTZN9JPlpk+jxGGu4vqvXmOA9CZek0KIE
rZQcPuFc9MgnZ7VwgEjLTTPz1kELaLY9y6o0ANdkz/y8wtPEpXlbjqvI4uytKt3WzVEIoESE1x8p
OxaKSVvSVuYWVTMjSQ0rkltFUEKT9HioIGLejm/OGAL36/jUk3cNyQaqJ4eLzwLr2Ns2GJhB0W1u
ceuAujoCwE1PgbIPxzJRYMsyGZdjZWcbyaxpbih4H1XUjEHPY/THoTPirsW38WFL7o/lF41Y1H8P
Ui9d/eYrp4Ru2LYHU4gvdkrSN3LhKj6IzqipSZPz3F6dOtDoWfggg/V9ISOicd54lRFbV7PaVnb4
9cu8drt16pdppA7pRdR5BgtqVt63l/j/fDLXppzaFzNDHY9UlWpriMBG0cHtu0RmRAjAMqmFB2Jk
vBO+hSYtxskglLJB5kwapGGiLtP8ZxfErz4kGBqtgxNmQ5KqkULfgZVKLckdP2BEbNDo2GS8pi8C
KIt0E6agA5vX/3ZDCxGmNGYFmxsyqn5Mgb64yO7RSJt9zobTAY/U7R3MC5ZYVF/NfrGGIgY+tilh
NGI6RVCpjUM4RNTeuFgqRaLFbApIKBDYrinENndUUcrU61DLWBiXjrnbQYDBJUEYivV5FKr4B8hh
LbGI+U8iE6WYFK72k6vQPX5HU7ebWfnVBqvEwi/fDXUlXz9hbe9bSAhvi/UgBeV3Z0HybsvooXeF
V+8Jow7fXpL4sGL+ApsADdVJxEnjNCHFMN0lRf5R0cPnGWgzmoRlCePy+ivSYeC2yUqsPMVQa2ky
BysMcjWzpaZHGoyQuae4ZHdaamjwGyfdsJocxY0Kb9OnllvDpgT/y1rG6wYXXS1XOTS1RI8YTiCI
GYjLD+kF7aqrGi/Sde8RR02g0rk91fUBcarzPgnScq9yKDy6mPNBWNIc3uk3BE3BUaDKGq0hMD8p
3STJS6nqxc5inPoZse/xNR7Yn5VgBvKm6sgKEUBz9mQsp2f7uaxPNUsKNOuvb/G/eXyov0pGEl3k
kPyBrty/xVm6f5AnkwrlJPAIzq+SYRgRH2YgyxtGw4wD6h/m62WK5yvFE3nnxkU12Op/I+LbCbf4
g71WhkCjohoESh4bCHu6z0wuEzIPoyYMQfYvzcNC3H5eGMB/xB5I/l6Ckv61c7v/esYDCtG8zTjt
2Ne7F1sSxn1rir7faDyLEwneRUJnypS7Qy1Uq66VM77kEiAI5R+OhcOKQFj3VmN6PxuQ7LuGZcYD
5WT2jrRb4CTjgtw0bmBzdWNchp5CJe+w0SBROUBNwX6Pg9UjlYy+KguwNbPrEYLX+wXdOOsKcwWd
Q3MC9/oVBnr4mWBqpsEy9VolQmuASz3AnNFUdLWTpYxixrzxBBc/c/7n85PnVIOnF/JIJ060hYuh
uFFvyifN71HGrwlQVPDJX5t3DsGrObpn48E3xvXhglXXxhokYcX9dJVF8VWXAb+LvE7NoNqtJhcw
tmTwYGQNTT00qGGdwAktG2I64dsM2vhddXgcMXsq9IR2XtR0QrTMf/wNieiD9Bt+ftT6+HxkdUlb
L3p/fdpBk4hT5nBmy1/gLCm4QKuNrDhDkiFBjqt9l/vlwWFYnK43NMFmXkoUJn6Oxcz1dxe/6OPQ
TSE3VgiK35BQRMfX6+Zqwerxo17gtUFR9bcxWNMVQvHCMsDSTkFSPKasmF2WnzGPC2UKkaPs+7eE
mFrBqqKuK4/G4skoZLAxqG+zBDfiUyuMo4VkhketuDlPyhbSbqBL9yezzQBEiynlR85TlrJIer2z
tNwz8HWpKTxoRH5l5VhdUqXXZbLhLePu4TVK30tLzoSk3BEvXsgQmAqrrz4Dl1dTKB6BKKL2wwM1
mn24S9KVoMPzzOEO2HnwFx7RvX7jMI8gdeIGusgWr/2LWBdSK6BfHgql+mdjrd/DZ1oVVu/Sm9Bt
oR2pZU2lAAGlfGE/t76EzJ3ZsQ4g+BwR0/idxlvdhOYBDAuis8VF60bGvinX2UjY9Do1wbenksEK
Yrjx8nxfRgROQsRIW9nj1kkTMxm4fnL3akXrKW1oqyj8yLrT7btVMz0YWFRGDcW7VNe0yvHckv4f
AYi0H1X4We0oCdNCW8CwKDrl1z1VAJXLWKIf4U6LJN91/lUdRgia/eWYW1RysyVEYSZoNT3C37BZ
iZ0kabJJBXQ+qhQH+p20EPn+mCZg+44yPgMD+GLChD99AQ5gorOYVY312Y48a6DhFfGBVKTVldAE
bRCGRN3cWKEDGYcAzNzXGUCztfEI0o5ZbFhgBohLH5a+SY8SGDkDj+nt1Cfw8Qa4hTO6OUTccvPQ
nae7C1AePCeOI5ESdVkpscM2MgBl/ozju6oYr/BVKMAWCP22dKZBo7X7PFK9jNALb5YBxaSNkxNG
pUneMrTPyxl970bFVPKMdMSX6H3b6G14rM9u3Xn09z8NpU0n0tz+YXJRYzoM2PT+9AEUMfksrplz
cQ9XFElNMN7AqpObQ9tlfjfnZKI72lmPFql4SgeBrTzUb81b50NDUid8kx/I0XXN0YsUxJpYLujL
3yM19sM70qW773/3cdYgG8Nhvm7+zfhsYIdeZfOkFSliLfM2lZrWjeAjMAJ0Mkzw9iOMLsTq5E3S
yn53xJM37o25MO/b06kq5RaLBwOzzzAUpbNsIb8CYhQ4BiEwZ3Uom58+7hl74m4pDxp46vqdYE/v
fmnkaNk27+J0PQgW7m84esvL+3XHmxC8rY6ibZnc2LWG4JK2Fkup1QqUrPDKqSKm+DRVcNOEZeip
rWO2bCwKS5Jhz/S3yRvH/W0PSBXshjotM4FzYmMqOBVybKYOps0pwaUPSCfHbBPUcXQ1YGjy1odA
3lIbQgZ6+WbPATi2zem0gI4xHngw4voj7SAPqYAUKHi/cFTKVZvwScgwWsB/GBHkTcsGmd0req5a
WgTi61EEN7vmQsbFYr5gXuJq4ufP23BcuUrJ+OLW2Ig6jlcpDztil2b6DMgPEgf5+O5VAEnZ3TVb
ARKD7iaH1vZs4ac0uteLv2EGWAZPHqv/S5eEyued+J4bXBWYFN90mXAmgtfpROIxVhMKcHYMMeRH
wiowAgCoDwmistA+UDYbFzF5+agAxGozuIhPZIQyjngUpSj9ueddT5oa4GJf5GCb+nD/grGKsVtM
EvDpq476+5FAhntxV+QJSEquRCNli2dxLUEZBbu5QK5J92w+CSKgHzyqUa5rF5XJtBVPu4zJZLKe
0SMdsOQ6lsykWc96WHIYEuRUWnOcAUx+SirMg9H8mn63hBhlrmcEVPopoWB9VeQVDELKjTDMcaOR
4T6OHmBpYzEIpUbgae20L3OxoV0Cj+IMjC4+6u8pKCDHBhK6X/wYs3bjWc5f4etgmu6Dz1NcW0nn
MpjqT+XA3cEAkmftGJzPvyWxSNM9IZc/iw9ANao9+seTwGOjcV7BxskrCVZG5jyZ5tZimpX5eGY3
eIk5n1vsK4J5czR9HoWB3ZKbf4LozbRK5ZEK6K+9051oq8lYavF/YKAGRqKMpPZCfjvqdLLaXtza
LAxGCk2UN65zqzrZMFZfUMlLJUyF8FZfKkjCERewqj/12HNdf1NfB4trn+UVFL1dBXf8xCFDKHHa
3F0HfqdU5oMjHybBUPbIpPLKPEYLS4+ZuNyc1aiyXOxa14DD9NWdj8HQpgpKqpqgjcNxZPCHEWus
wK02VtGNcY5khneFZmaYtgfPFwSZ8q4ifToCBYQrBzx33CEcUpdEZs4Mm/QegRIQXr2BeuUeIVsc
hx4ot5IFnCfNHRJY4RiFNV3ICpj7vMfJSO2Ut2c93/3a4r0mRqwUKvjAXSlIbU/2Fi3IRn/DHHU8
NphBpkuGjSTYv0Tq55g96dLELjADJpN3nLlt4poH3fZPNxeWdDyBW18sq6ocSMLsoDUNdFYEOSRX
U4X3cWcGpi+uEwJvKtKzovsjX81lbNZV2H88rAa7CyRq2X+7432zAJmnOLgHBVqTtlAcRXm820Yl
8wTY8ZLHYGf4Z4Rbi9pE+KVpsahwjL+1N/QZOeTzKBdTToeGA1W3xA0Sdb0XwRVevOyr5gv6pNIq
KIraY2Eez24rtFLVWUc4SAftlTTwOeoTofyA88kuoPu4ZgiWirdgFn+7rUWX/pjR55T8SD7qyznu
U5Fwxr/ilUAR5AO65TkxXz2s4DOGB99bPF7Q4G9JTdL4WK7mhqcil8C4VQ9JtfvcuwA7XhOoAMzg
uAsQQs9ZhB/uGCo+ipqDtEjhAWY1qeTn8MHlxZumN9ppELgoUvbZagOkvStkk6pu9c0k2S4rm4ss
lDNR+IjH80yOk5BO26e9OdpeTvu+W8TxjbsJXAZAVFLrc183X4jXYCBuo/goIQFo3JXJXJ32KnmF
FBUOrTtZHysqB47bLuA0QVkeSsn8e0C1cgcrqmk+YcPsK2hW8cJNMvUWdZlDu5iCVnBnGZkzfTcm
766J3VcfcFD6tJ8n4m/6M8mv6NCeh2ekfIRkovSqNCWYZON/HjnCR013jFD+AUGZPTrnY7vtkdGi
EVxazCm3vomLCtpXRC4e6zpGyjlQbVdEtE+MVfjS/zE0d/bo7jpdmLMfJgYnluDdLF9wsoq5DxWI
N4USUBi0f3dyNZMaoVmVOlQdDZ6cReNsNPF6L4mFE5zex3Jx2otfxW9o+Hm4o/3pPFDYBW6Po53J
9IKzwWt7fS6ffvc6BP2tN/hRQDpOH/z3F30niPZX0pRl4bO+DtFCrdvtUBoiUwbb4VOOgwTcV0R/
wYjxfsKa2cyxeEv5qqrdcHKwiRCxLsnIA5jmX792Chz2FiVNS4Qkx2il8UJ3L2DaA/tWRGvdONWv
clui/dGIwGKD5Bi+Ii61XOUuRQ+74oUEsk7BcIBp22REHznvw0bNV0HBq76uz1SDb64txU2q1Cku
iET5+VhmhCm+GDc+HfbF0+QHeWi5MyO5YKXcXciYGHRFsFWRmQZN39ahfyu8YqXWCq4oZQsWcK+s
CnvPIqT9spbsAouSWlk9pimAZdm6BEeXHXNptoDLui17NTT0eI5PybMW+3cvvZa0QDurn7I/qBaN
h0utwk2T/559wyMbmy7t+Jlc8CVKzPDb29vinFE+TgZVrPNy4rKSHzMfR6qaX04+Ic/r0kiWP/x7
9xtYWpFtJg4Op9raqegUj38dIuQ9K0KIvVcyCxr4xEAt4eFHwNHhvQG9d4dabAZ9q4TY9rIBwwZg
eWVfbsQZoaS96ZoKMhV7xvRcbu1Q/HfFy02sPt1uLZqsKgFuUNIr8n0cKmlby8udYSkDbWIKMaHO
rJVPPtAMyoYH0qz/yishratIu1wlX8XxweW/6cHxHoNnZjwfqeu/uI3zTtn1nv07ZysiT5aL3YfF
O3y9TppAN+kJ81WCzbmkZ4vxYFMSGOA0MBUdGWZWWB3sfgTLQBZwvLZx2uQA+P2nxGkzr/WNAbCm
3Gv62VJcgpWkI2lRDMO2XugKha5qZNeSIXGHy5sZpH4NfXUSoC+VHbH8ByU2eFHWuj689eabKqug
oNTxe8fsW83JHyGi8ikCRwIrEeMuxi6j3e0sSWCDfLR559QMY5PQyC8ZNdn9qjV8yWzO8kppGOHc
wzPbsnqFdKGAC2KUwyKwVmSdzqJAZMxLQu2vZEomIyUtjjaX5ol9Yt3PnZo3z1of/eZ1HaOhJ9LS
6LzcY2r8yZ+yUikEaj/rRrbn/8Idkiyzpj45RB8MxNUdtxqiGKOivE3TMo83f9Nyf48NOOhTXtww
TV3TfQ6++RxBV8N45s0J3yjQsMiUVEZdMuCG782vbH6DwIMALgF7vmTOhBu5NlCQvIWkwqzLYPmy
WgiG5fk+qqfDBm+t0K0XRztYIB1OTE1Apa3P0RKj/fuPES2ifnr0ZajuW6YWw20q2QU5InacHJr9
YbQLBrJBoby0RB4xcEFUA2LsKK7xIeG7mCPEkcJs6iuYvu9ZUUOyzEWlSnT1HfvZ8qeoeQ0nfBhL
tEkU+ngzavEsagWaziFfKFwBd2Xv7ZVE2JxZ5hj6iZFs88KTp/2BjrSbSU5UpYAAzACcXR4d05Ab
Z9QAcOO8mbTHhnFoDYM76LGZhy+uu9cr8ilkCwXnfDfTziNnVzkDjOXCFQCAHF+sAWzmMfayK/Wx
8rI8Q9Yfxz9I1T47INy20EfXGoB8WAwjPZ2agNsnUPLBfzB/7Kw7TcRYHjoA3Uu7H1ZwJZiQQkMM
MQ01MeGy/fYTneFIATGf2vrRJGlmNu8GZTp3sQ9arIzTKEUqKVTzjWFFOUHTEBau+ZW4wGick/3x
ehoabF/853ZgPJbzX1+qylnZ8us1YKvJpHiiZHwnQh15lb37ICOR920vEOFRMIgWudaeJoq8BazK
rsOfRhafs3tmNZTt/Y5IAobAPCyUOpiLPeE+B0mqD4naOIn0lVCwI/p1yx3hoY9gNq0P5PduhhSo
DXNsOT5mE2yMBCGHiy2N4tSdYbDbww1lPBfjYmcra708rSUQ7k4n2YXWEj+KvfL6DmoLZ6kE8hWM
Ql2T5ALjM8O0JRZahN+GVylg6m/aYMUPq34sdzmTEx1toXvbz+t9XUulvUgaP9yLgHKWswnBKtbE
7ph3SDBPDdxfyrxVdIOAKngNYk5Wune0jbTT1KY9nWMBV9ABIGF7fZC8/Ik/KAZ90E97/Yam1ekK
haxIa/CMMkHY/a29676PQXdiBJrk1+X3QPir6cIpdgnnixanFAhMeGhYP50QSiqRXdOOrBA7q1TL
zdZtUVgblBt4yglelL4MD/CVKaonl0DxReemJ8yH5mmUfvQk5/bAwu9oFVWkJQjRVctFygYhpRyV
52QTlgb7vRY8H5Z2Sy9tETReTDQ2Uexi3Itc3j1Y/Uy+z39Prsc6td87E4ZefgodCpbqsBRcEJes
FCn2bvGJg3BRGlMjYy1HK4Xc1j1/kQAOetKvcIa9qh9e2FXFYNFvO9eYFZ7V8DIue5YzW+dzYibE
RWZAq2Kwv2JR+BOyB/8a7ETIKEzAVYNXUP+/8xjVvFTHTXz23jzq0j9/VD6TjQURYxVbqk1zdtc/
OAKMya1BtHBVdCcjpuZ9/Cfpkq7nEHD2952XQ3ShFIDBhhle0/9dUBMktUnd5phV/apg1dLHcWbE
qdhGGrwFboB14TDmjj0bXiyMfnryrGKbkYZgZd4AyeCTyrh877YSoKopTnGvEQJPd7wfT2Zo5ToO
TMGNcOEL1W4iFb0pQ527WU+KBpBqvjiu1sh3Gc/Zsus5WT1oRR14m0QHkmhArBDVL67Z2JudKfNO
FTj3Kzkz+WpeRCIePSBoaWiaGRXXM6LdEiOswxW3pJ4x2xR1eE1eSXTU6wMoAEeN7wNJqqG3S83A
eBl1iZhpW9g/3091xSOF3lTENfhL/YTl5OrhtZ4bwAIdAHdyTSsXMxDI6xxYeZQkIwPfXSUkDVN/
ySAHLpT8umf+ayEkNIwaFcLAC1RPN8aU/bOOD9n9ykDjy9Rtb50SLHNPfl3jN3ocLVYABW1KU4td
stD6W0sxVYJpu31znggfxUmM82ryFuXvyPEWp+z/MH/ggs7DnzVgukm5o2WsQ7SUyAARMTbA0dAq
FdysGOTQZnWxfQ1LUDypo/HFnZqVptQVJhheHhJhXroyvfxcDbiD88bkFlAhteUTT/0X4FPqrSBi
pOrvabZTNhqWUDw5yTwze0U5YgZ8K/uaFXEH0SI2NNgtAfjeZ8OPjtJ9+HvNSkAuP8BVRsQR6acV
bGx2qVWKABvHYiEL6yMfMj9effpi1Rno8G9WklxipMYkxWmED4g56g5wwb3CVSTKa5EfdO2QqQOh
ZBhkK2kTmEgaf7Gep8K/x65rEt/J9vn5Cz7oEb82OhOlWwKKgOUEI1Xe12QNuCwq7DhnvALJIwbH
npg2UrRqQgpHZvMcoLdVp0UfyM4urWL2yMBkp8RSqDNUmkBewcDNSaWeOe1eo5/HU/MlG/TU/OqN
OXxnP9nHhk2UcDXck4OkQssvyPU4z22w/zd+oGVXWXhgDYofXMuky5/FoeNzVkFNYhwzD68oXGXK
7MaJspxa6jAE0s4T1f401TCyj6I+3oCi1S+0toyKPeHcxg/c6ylGygll/uoxfSq994w5im/aZzav
o5FCHv/YD6nYn9/Z+tYk5nsRXA+R3IVdRLE4gdoHcbiaCv8sXb94Cv2NAhTZK4xLb9CFQFM+tw/p
9KHNhgatS9CGrsrFPvbo9bBmzUCEMYPt2imiHgDwn9ukqV4+nFpEcLIlEeUdgOa33boxxA9UAWgM
NBc3h6GcsZCCCNkYZuS+pIWzhUb7SlP3k8YNCMHzbP+FFTjzQaW/zzVXdoqhx9ely1dM/qo3ysWp
b8afe4XXUtqpOwdQJvungTUuW8L0YZdIxpEEU+H8CUFftsbbJncHn3pM8DhQPIngtu1NXPnv/d3z
YR4J7eKP+OQ1SzR0jHoEtTR78zJ+JXa2b8wPsnnyFMseRwg28sr/xr4gCkd2K+T9vLT/Rh+khMN+
/lplJIaSqG+z6PfsSFh4NYNOFPoKFyl1eDE+02nhiAjJ/7llae14+NxLFK1zclhNE/HH24pHFtaC
/TIUW/m9UJ9oHFFWNLKHv90MyQKLIlq2Xt+cUMXESj909+AbT2ZB//hYx6dsLStbqYKAk83koN23
2XPweo0ace4QUlxYB/LOqbTw0YNfTp0VWPnsjSRV1Q0K+IQkiLOLjP6hi8YbwO8dkJuNQ4qIfPHs
JlG3xSdO7pxYLTsn+XmF1T6MyVa4eng7vjEFlSagmxROQKrXseeVK/ATXQSgOO46QHV+T5JcJQtu
3hBkmGhwNdL/J2dpvhbRTTMlwBg/MmKuGWjgGbl6KD9zTWeZRMvC6OfveWUuR6z2fb9cRnG3RQ1T
ne2pFWklOLdBcBdxKBU/RQjv2qUHjwskBzVZe+Y83dbVleRIHkyJU2nVifAtqdduTDj2crm9E69x
T9/KSetVQ1Kzkc+cAbjTdgdE7xASPXH4tqPqmThlhVIoeUeICb5lnpOnybyr7Xnn3tX1bbVJAaw6
8cGRlcZOuukk/+Kh6MIDz3+DBilTDjAKsj6hNwjDosMEYT8JoBGob9VCI5iLRj8/RXo2+dY7llvK
tpjZJGo0e90MW8hgrgCpjmY2+qzQn3T7pLVL5kIcLqzIfglzwMUJaUiyXONHqRXyKAS7rkjBJLgL
GQ5cZjRDIcvut5O6X1VO7eriZokNanUBnA9QlNz2xeOlCM3+hvON9jUnAOE5lwKAC9jBrhm5nuVG
ouz/uR1Ofi8xyDS2KW4+iQ2wDDJuGldEvxLFARV/dwmRCuTzAGWXM2fo9N1bNoU6ovOyFllfNKed
8JSFJ8klCXYgoqjPwF+d72rXSy4mGBh6kRtVVhMV3zdwjBhXX7CRv9/4vCbPw9CPBzVwRLsxpGrm
SWAkGD20/4P+6MHUqOr8ygZOhkTiY1GXRdrmo85uwgGT4ioOufGha5b6humdJsPuUsrg/Ps1QwF6
nNC4nkNRwh23n38mALBkLsPrOOq/DrDeM4acb/Z4Y0EXpouSOGX3hjhAIABlaZ5dHokVNmHPGRr1
Q2aD6ZAoQOXIsdHPvSHTSuzLS2YohynB941qbcOVCWX9osUeejnKUYe4HXUUsnf89InrLeUg9aFb
4KIff/W/0YzDuy4m8sMWFYcqWvMS4XcJ2sqZooXDYf58I9NDNQDOH5zHqhpyKtTfCQaj9ZqAYlSM
ZyrW25kgZ/0InKrM+WaDf5sDmg11mTcaVxeOmUqCPrJB9xntrVaKdM0OW8owCdProl+CkFtGhMmk
owg7QCcJ10d+oZ/NlnObEGn2dAumY0ZXlE0ZB/YelI/QRqVPauZQy0iS/i6qn5Y3Akg/tLnHV/X/
q8Fn3FLXBJYvPAf6K5v2DefvdmeEGhc2QVZR3BAeWbwSyiQHaoZL255WCyEG058GrTLpQ4oqChNi
EwOHHx+zcMfiYFtDVp6QhjF6yL7eWJKTE1ys5ecvuFwtIGJDWiN6BsxMEhZ/M3X7CQDcbiR20OQf
z79HullR18CPvn3xiG/4MTO7LIGg7KuB5Zqvivxy+hGxXPi6PtToAJFyjR9KRuAWBi9ML5nDd9O2
jbO9AI0eQ8/cU/K3mimb/8ZYsdMipjr8Np4G3y8W0OHCWUk8JFvEVmAEfpA2t5haeyCwmrmGWyaU
s5I3mL8k2QC42XBrDyCv9opZCDpymp5ve7yEvUBeDVatzqmFYkuEJMCZDM2wjNbfVGmikmKbkmyM
QmNkZTm7JfmpJkJk3Arce5Oc0KYdzSQBBXV9hnZ0/uoWTWQ1KZ01IZJjrzMD5sifUukTP5zU8Hrc
DPa6Vpem3n3O7V3fRKpn8j6T9uY3CRfgNTBevewFy2FFCz7KVI6OOyRhSSfTMUXYXoFLXD5G+42I
GtiSZLbCX84it8rrGDfM2xQwWADnrIQxjUOb3JPBv6M9TXGO3kIe2nZsfppN302vqL7O2etk8zAA
igVOve+VQw3geX2hWZltK3DXESYOq1m9wWj4xQ6lF491wYv/FK+AwgpGyun7u2BD+TWTBTtokixt
rHeWGu8ObKWcdDxJm8vh6dyzScfSM9+iB5RIdam1upqXDOhsuNNF+Dm4XTSNoGPW1Qvx7EryZ3fc
3EKiEHcdAOVHhmGS7oiISvbIKzHh4tkaQrVBvKK/GYQp8mq/T0arMFWu2MNa299hys2eYUknl9nl
XeRU0N6pG++LhdDTAE+x204cQ+pSndASpKRRQh9tTcDTNFIO/qtYqiyVE6sHPC+uJS/DvItiUz5J
c5xdyqRLPZaRpLK6qx6D/qxgJRyeRPsYxxrZhytO+0YjN/AZSuDh+gRK0waPsROk4etrxEG0HSjh
kd7g9SdYjY1UlIEcheRCaxashtK68ed37ZxKjvrTv1on/qwmxtA0NVJbEhj2o+/i1nLu0NAe2Y+z
FJXkCbSCBr5Xnr+qHOmZg7z6xVuPjiTesJ2vwubsRSH9BMDsBS037WRqYH2l0P6vmuGHY7/3mLv1
3yq/S7LksREO2qGJa+Kt60CwX1Kfp9/VWWdavlFwPLXbJrhEB4VHGrimPvwzH8LYNoAZC4euUE6r
gpYe0s/I0oemKt942tfvd+T7KogPzo0aQKyvTAkd+oJgTUIdD/JHa5FVN3mPiozKPsyZqUyo7LZD
YFbUVB8h/qeMngrFMwBqPN3yX6Lf7lPaDZyM4JQHaiwKc2OMw196jLQVALg0z25ShljKswdqD7Bc
Ut/3X11a4C2oAtMsqXt6kh9lNap4fKNlAWxQO4jAx2W3nh6nULdFKbbl217PXpItG4R/xQ0DucDT
tGYo8f43wPLTFb19OaiCwSRJjTmfe+2Q9RB9huDoJ2XOnAIJ3Uppw/6vtlM02Ieo3pZ5RB7stPrN
mrPs50GgsedwEvF+UyZ1Od77ixJHgHQfRcSXn0LxFfUMDEXab3/A+XmtZquRyCrHWx82gITzxCty
+WlA2eDz+3vHMpQXDV94TdolEcYzpAcPraLkYRAeHdpSPy9C4dAT6kzjAQRv5wc41AySZP+pQubk
FR2IjgZ7JvbPakVradKnBNHpuMNHySkWIIkViLs8YF+JGcZUg4tt8jREnY8fof8lPCienGQsWSkM
Zv46uwMmIC0hYQAfW9ufAstT+uJLgMPeujBHVvPpO9zPm1zrIddgKtQ0nNjkCrtt7YHZ0FbYx2Sl
UWYUdIlp8Z5jithj5wdWlbepTUp+XCrpmBdfOHsoPgtSilK9l1ef5Q34fhCuTUnM5Ux2wswQpSMx
L3JDou8WJnB+c2Io0dmGSUoxnBLfQl6oOvracEV0/7HB1ZiP/UOxiBcRncHG/esxdoI5IZNSjMTN
13uJx7oOUuAlb/PpPkn32R8dH9UJu9dRkDvINIktThnwNVwrtq8bkq6EILAlvq48C8/UpO56yXtT
zaaHxc5NbcgjQ6mmnAHlXkMl3I/k+xuBdRKWtXYkyNvYS7GosMMNXXnTcM51uFGLmG8q9+xZknTB
p+mMkKlyona3TzCnG9wlfEhman0v2k7KLkuUEbOoHsMihWwm65Pj/QCXJrtn6+sEr9wQy6VF/Qs3
eDL82Wypx8k0glx9+jAdlZfCp848GPieoc7stIV/2jJNTCFp7WVrgYiOGhh5XOgPOrE0n+CfsZjy
nsBQyyMEOgtDkLOeLPLe9x0RnPidqpc84Ivz4I0PPtrZ+C8UCc4FbqjAgpFZksjPOkhnz+l9WcEj
s59q7z9acuNe+M4hBoOPYoZE1pztTu+ETuoQintJBWY/N404EbVpyUBXvk/ul7l588o/9yrV/VGd
PRHBXtnkh2ljOpH4rnnUSUF7891x0dIbygpOq8bTfDLB/H0aBhL6OKcRY54BP3aMCWhZNyKPd1Ws
nmHvZnLYYgOGGachO19q7O5qn8V6Otkh+vsOai9AFOIgWo5Juwo/emvEfMZqBonRYbPVhURFcOQf
EAFz7sdS6ivj0uL5fRUYJJIhwr7DSQ+FDBQ4dqo3VJ64gQ+mF98kP/hXV5hb2xeb3HZd03OZ6Eiq
tHJS+r8bWO4HM+X38Ufm5xlitmPb/4JZXS7fQ/VTMC8edBrFRfqBD4AeTvRogXXhEr/LDajuzgQQ
3qNLRDB3TwYVwNk+9YjMBeGHwBROW1XPI2nJ9/j1tM42ir0+K3b5Cr80MRzfxJwEf1uvgu2ahJLV
iVIut6DRu2r3e/FoNO9iDzRGc/qOqBFnJTTxFhuuzlmIBF0fqkoaBXoc9Um8ix/m0iDjdUZ5vzdp
UZRWivPkCx/ADcoeFxInAy0raf2nZ71dobdG4WG667/FtyMNSCMaZ3lRYRgqBSHwVROy35v5vC5y
+j22HZNct3T9zPeEOIoy0uwdMHy1B+geB/263Q1M8txcmVgBKOaeivtAuXnDN1Vbge/cpLmjGpvT
4HaY/TmnUtTew3Rn8mImgnKv8Lscx/nGtI9aZhxIWEqCR+m5r/3NK8L45mWiKnA7Qivd5U9uPYrs
eWhNI+rZbpt0rPpO0QzJ9jMzLb63ABYm5fAX1sxUdBPQXYdo8HQSIXY4lM3RFBxg13a4maIHkwpU
6VT+v2uOrt/POr0JN8OJ06bN75WBACeXtruOLDK+5MH/fd4sHUVyJ6wIDieYI7UJFIE5hnrXsKTY
MHJf7zPGu7PuzeUQeBb/T2FElEFyM0AIyNzA2zquj6XMA+Hl2fiydYDztXpJVQ2qDy/TtEddV+t5
xcJxPat7BB67fHfQma277zj6xd6xlMGwexewQi4huYiQnk5QKN0gqo55uuOCz4Fgmh57PiTdPPEJ
+LqBhvXUG6/GVMgVnpmyeRMsNT//XW4Kep9dYSiEUwlB/MpwypljdReC7b1HprU0JviI1imfh4G5
srBu141hHXLp8bvjHWf74S8tY0amvOpXDUPBLDkNoQWMJLDsrvXADtM0jSPia7VL5azgAUfgdB/1
YeBlS6NVqb2p1cHE4edm9Vn4nIylGnUFjycyih5hd1uZ5gXC0RVxZ3/mbXnouL72Tgkp8MzpVTAf
RNTtj6V1mycIEp2ckifPBCnhoJPX6sI6DPiaUGUVDhHeGNRkPhuvBT+eB8VhTCByl0S6a2bErO67
6GB6T2mf4c2RXhe0HHG8YSZnmQQzaz4JjRA+d4Dn1r14/8cLkR2aLwZwRjjB0P3vId+lZgPecwEn
WfXS8ns6hXO3oWXTLOz2hgosDisH0iOcBZF0ShpL9mrMtNTf7sFd2O0OYbkaRkX/Iku9VL2lraE9
iPyW1zFEZ5GyJY2IhUfl5a84IaiQvPsKrtOhxBKvs5Js+Gjf2fzW5U0VS7QqinPRpva/Qo/9Qxqu
NGY2TZwuLWIkDdrwxlpefLl7W2x/VL4zzm/WRIUTDGyqV+Z2+TaM8GSBD9B8m3CnFb6XfjdFiITy
/xCHezDJDeqpYJc31hbnhaDUmsE40npkVLoIb//gs79VNYbJRsgzXKJdP3PUWY2bBZq3yNk4HHZF
cddvh90YKgep9bMM+IgUoEidX/mlFKzG0YN6JiMeSRCK8SC2Otq5AtVw1YaMQv5n8isK/mCWjJow
gK3E3fGgHGJ1HI7ESSN3lT/LN3d77b4a9tqXCfzcq0YPlMtS7nLrx/60iYmBX+zCCnT13Bw+1RKZ
SzGqzRkxSHxxJGHrbuYA7f0a5en2e2VaPBPsZzGWnCOhihv+7ojLP7DSUGC6jeOVi2QWAfcGw2BG
qNrIye6RY3mojHpVGQdq04gCvcbiJo6rRnlghgkIFnhMOfiozeFZgA2KGSKttsNoFix99o9topYP
4h+EUvKPtKIJVyBT/SWpdPbl9hZjlM4DQJIRqgxw27KpIRdATvvdwp8yaiKqft1H0WEaFW+Z5O8o
JuQT6u4YZLdL5cnGxw2W1PMbygQqk5ZbVizmNmVOHW5wa+5ZGCS2HIzs8VO9ZNswOZQTryNGG0bv
cNy1Uuc4kJOOlw2Lau8vCYn5yyPbiAf2Kfq2pEQqFmmbwNy9TEzaqgyXaRLnxf/YoGNI2GiR6YyC
yF05ngzURkYGnd2ZVEBTPmzWNkYeCqHad7ISfOKtFYq+EWZb/cItpHMan9yJNCo4iyk8vAlreTo7
Xu5CmG3CcskMjpCfGqnRSObUyhhvdtHWggDj3UFSPbuKqE89Dttns2wREbJ/9V5OI260uqw2qZLT
L3ldFX2JxzA0kjte5w03Z8VJoelXJUhsJs+l2Cjki1o2HO5kJfKX2tLd8Brxg1/N+fIAhWeMT3tT
SbxnqqvjInKYyp4ieKes8GXMnZgrvdaNhqQn2WiBEeW8qvVQ/bBnDtt1RqXd+GOAOM1U0GwFTTTK
CVHgeyxCVfG3MqAbmpMa37sPTIbf//xDuWXWzhVPm40R+5IGyYiexLEH7+UmfGcH5okGJCPjf22V
92yBy3btH8H1RQvGpfSx3gksAw5HKscOCmYFOpJW2FED5cyXYpIpNtL6eOu01CpqTjajpY6YPwuB
MPnZNrEcjbDzzz+oVLzPieFVjPEXb1QfdmqQxjfl1nxb6r20ysusrSe0NOnoM4giV1SNvvZDQMGD
N3yDLRD47Fd2TUR3VBytOv9w560kaldjdZooC0glXMCdx+PdGDEx1DdS7/7odb3dAgya0PcWN2Zm
gxanl8oYE4v8HeIUz+xjYhoqPeXzt7drEkwGbFz8HIqbJHNOv0uj+Eua53I0CjWrS2pyEKA59FG9
IOJgXF2aXvXLRTGkd85wHZXfqzGlAQMC/TBoRiLiyRE3K/6cmjqUzhgPKNWFov52r9JYVeFyvSKT
wuTRG46X5PpiCxuZA513IVnMHTIzQdcwbJfq4q9CEImi9LQJ0vdVgQuQ9lkJAkGsDcvXKsG6bIRH
yxOWuT5OnIW5S4bus1TOFPTC2OJaUfJ1K8FEXRQhWhmKNbtvodr1Qt8cprBBo1rvukBkSAe0xfLY
oInnwf7qY6t01Z01kzxCKddaszD25VK2htXCjC9g3jOCtDSjc4ti4vsHKiF96JA5kXIDSxu/nFjN
GZeEJUSyiYcdmpEJIRHOYg3yW7+qKvd2UYrdTUxQN+9MwL4wOHcaBqVIt4Kyzr8r0FKQrH7bDIzD
zWIlfx9MVCeFGxkD3R2hX9imHAKe+NZIWP5VpkDgupNqXHimKKyEeTJVu1siMcVXPamm6Vzr7nmJ
CDmr6iuMwYl/2bScVUOcCIDPwmSvLW+LSo442002XKR4Q7nnZluk3DKp1lErz8LHb475PZM6RKeF
JEiVIYvHXJqgJ2vCYo/nLjDUV+lf/cNvyhXh+b1QlNn37SnqyQ6hgMxWtbvVu26K5RQVkxXYt7I1
7/z8zgfn7uXxAFPWN5TQyeRE0ltfWNT6dov7vwpr5u/Bit/oJStbI85b55qc991OkOhnHN8HUKHv
sVEJYLz3DW5kiBCGCLNdKnuKTkbHnc6O6THSG/duDTgr/9VpnUS38beaDDiXBn85eojno4x0M3gf
kB4B2WTpSfDfUxTZvaxQJP3mQmkLGicH7X0pQ+IVJegg9zezHpNkNe43Mu8itrh9RzDQjIYUA7Iw
CzXLYc8AhVZ77y4EWAYDis+2LDkW6w1Nv9/xm4M69me01K3W/CJ+02QpCWLlxF2aWO/gbXb8TFkz
LDDAjh/CXnXdN94HqWOvGrDGCJkW9WI9aN0guIehApPltLlwsXUltUyNwocmOomTPk55e4XneqpO
r26+tHeN9T38yPR12qDvr2woDWpOTLiWJKEg6oJryHxx9rvK8LBcfQQJiq5jRcXvF/g4lJcQXeDz
j2VrH08pR2DUYAhOGwnS/Y+fHHreZ/4GnZ4dauuCctKjP9eRz54zXKhm30qwaM3vnkj6LFh6kqca
mBQtIkutZa0ZP+O0pQUFZiCPHAh1bwbQl0/j18I7Xh08mCTPsqQzLGP68fMT6B8xUI25mE+RSE0R
59plesdF1WtyRrJhpr1r1mRYpBCFDNI25Dk2KExU8HzeBqFsyi1b86u9QL2bH2ThCse7ecBpqGIs
eppnxc5OdsecvXBCnbrWmFdSTt4l9FGot5/6usYEwMNsJPm877FiTiB6PP1gC/HJAFKDcrd5QIdU
p29F7dD7CLv18TQVuecdNnlzaynUQuOzL57/l/w360siGJilkdP5DsSghDKXZFIxr8QGT8i3M5kr
53QxDySi1FoA1dhUV8UUfMW5zwXdDiCPEavUedO8zptDgEqRn+elZ6UPQtvzHuG8eZsqiCoTYRg7
HYpX0GyViKayn0l5JvdSZHX6GrkZFu2oIRNNA+f7narq9yv4/FwqgJ+fcfyvfaaYneiwyQnKMAOp
qzp8KLfcLmwB3y91OQxMms+NC+XUnXgSDr/ywiRYBgiMBmdpfggsHMcXjvfJzVXSo/bbfFhdQ/+o
6gIrE9+FhgIMkHxjyXBP62/Y6Mr/K7FUKqg97h/8gLDAaZ5e3Vu2q6v4g6b6ZLuLBUCkGAs0GdG+
6aOqkiJPfSUl/2fu9JFfVbu6borQP1ugZInA7KisHCtv7U2OEtTXMO9kBGwmw/FRLaUw1HTu0vXH
Uq97N3HnvCw3rJgZ7cilbQJpQ1RBeXmhoIekNo5fhc06z1KlSzeBw+bH1wE/m910cHT1Nwov7fUF
K36+bCU7FaXHwc7UV57LC29yKPH24pYwtgIIR9so75+NtImR5gTkx1SuEkZxuaBt3qr9TS76O55J
+WYN8gsmGlfX0ua2ObqfHQUdZJG+S0udf8kLPyCbpCeCX08x8SJFR9L6onmo56WLiTbBrOYAxKSu
U157UaXUa2nWnPhxXzQr24856r3sC06SaxyxKsRe65Yzbz/3hEJxAmz6n0nOqaRYLUR18I1arlHb
xUpKVfulSRJUOVwT/G3J/Jm+w5m+MtSTKUhjoJYWnq5/uoWF809IyqPIbeibxORjigTgEAsyUoBc
0hCEx373d0F1NKK0RwS3l84VsZvP+um0hpQG24mlmNqK4Xa6cB/u8+Pe7ZaYhYeRuGnQQ2IuTbh8
LJpCE8MSVnTXnfGMOYRt5nP/mWHDqGlYqgtbw0qu6mnNPl4aK3S/hoawvMtwUHeZKAA+/LQTc+Wg
y+R1LAaEI3d18ks3uxAHUmXa68wZG9zzEQMT+q6730p/xa6Sw1bNUO8TlM+D3BoYGYlTmlJ9o+ZS
UoHsZeHDp8KHrFLy3+h39YTfY8KTo1nEhsPpdvZS1pbG+trlw7QBm51VfSh61w16kMF940ZPQ8rG
aIS7U1y1WHgDYpwhnq+nsnm+1/IzRpvb+p4h52EeaotSKwud9ZKqaFSkJBGqPxFvz3x8EZGkZNa/
Ohk3BZ7XlXN+1XsjZzpHIaOLtyAyyrQXPjuik9ZrUM4dUJLkBl2j1a0G1RGRB4WYGCdFQGntIlW9
lE030rYaIrcClDZCq81tiP2FZuMbc0bVmrCcc6FhBQY7KqMfviYVA7lcNSiuP5ns2yaUNPaIWtx2
FZ2g1gQyFUCxDq2xlALrKsKYLg8yHa7pZeyMnnR/iIxqIpryZpISrwQRkqXPuci2ZODZp7uMfMe5
cINQhSFZSnZWofzwOvuQHIV0XZTtHx67WQZ4H4kb7xAk34uNx1+VqlwsVdKwTXh0BL8Pa0pm2FBu
fGw2JXPybXSSWs+tLD0iUyATIvttyNdlOnvYwtj8MpnCGfQrZB0zkt+wQnL6hDyyfgG1sjffXDTq
fM5cdIKQj1dlYz2K3NbsGjHsbSFyeDuVnYFY+K5QMpUNH5t55WudNQuR2YAA6TKnwq/VDu+aayHE
HCuWraYaNLqpVUonKhst0zoHArkw5JSQsBDdEr0ha7dd0Ijrp6cJfLeZQFOlZEVwO4y3fEt+A01k
73U0Fnt7EbYMHf/E+mv4dUeoG0F3YG5n4Fn5no3uzd8sJ/h/7xeMHkWOVTaSvz+hTCFIkgf67zvv
3Q+Rc3oYlk5bG3L1CGRtQw051rgJoZw+97HXp37CbkqRpNH2bVbCiQewJVVuIkrPtGzM9QTjURaT
4A+sZ4bJsT9fXWXqRfX+LPhHHcxAdSrCoQvm+BUWA3zJcmYtcrA96GCQJsAokEdetvkkOMwIXi1x
Cie0SovgsI6ttp6y47qJaNoMZdA7bgrqwCCz69hc1V+oHRyoikvI670KfPlHDiUOKnKwG4ny9TzN
Epbv88V3cb4eRwSJSUI/LbGFyjqk1S4DGbp3nKBG+qy6Bkkj0gOKxJ9APQTD051oJNl0LnFgzGwJ
zlsVJTMVquS4X45UiG/ikrz5Qg2D3Bx+lhw7xjRW8zOFMG7dIb//oe/2DbpVtfqmph2rdHH8UU3y
QPDGnUKk6dglqGNtTV0wdIY0SsXajIzJdy+g7w9qrzX5UBB3jsF+dLB8VJ/cRMp1hT9/AqAUN6K7
igHHBfRPzz4VmwVClLbcZfKoHN2WcKoy9KSMZeEc3rPDHzG+1sBZzhX/VXpFwLF1Za/MoYfJ86VB
Djw296Bq28GJMR0/JJ64UdKL7wAE+1p5znFtPYYHiFOt6lS3h4KR7pVCGV+m5+u0EkwMUWsDd2G3
dGT8pYysxCuT4kDnzg+sWZXmpcZC5nF62hACIU4OlJb9jwNe4gKPNvV+Ksp0Mo/+HXjjYyks0IQE
O4G12Nss7IgY+euBjJAMru0kkwISdRls6AjVaT2cj8RyQDXURwN1lTKCJSH465HJcaV8xKyqxQH2
BDfG/ulwFJ+BwCBjrJWlabUzOsF3SqcWt18rVkjK9RhwpSwjTsCrNXcev7ZyL001IBiv7qHAZkQY
wylOPzrL1MFWlwL2835xjeUUMceHSkO0OSODtRqk53nj3Q+6GRdnBIyH2wge5+1Bo+EPrYWrkmWZ
xx4REkvIO6cSA/gWRxhLjjNXUedEMF3zzbxJjlGf2yknOXBzze27JZBKfeEHZaUerAMyO0Jw5dNK
zjYjU4R9IfIg3ncVRbkaCjZKoXUWvGI9s9LCqh668r+3cuDBu8Y3sk1d8fxkx+sEWLHwVry3XDyf
SnbOOQzaHmZ7fejDiVBIHlHql8+mxDQH/0oe4PVjoJTGQEAfiVYuKlKecMPqm81Dhpexpa1zidYg
ftg8e50814Arh7WvXcKQXSrf9jdI4bWmG63QxhsSAau9slmi7aPsCJI8XSzgnCRherqYNtXj6K2P
/99TAzYvz4akWbXLH4hx8elU+D6vFQpHTgP+YIvlTu4x8KvhZzXBCnk1Ch9VjX6/iWBHAqcyUIu/
RfFffmr2ZCELRUFo6qi6Bb+dwSlqQZ5dX+nVlHSp2D0zkbmjB4b7NGjy7Qr5iaRanPqhLPqAjPZz
Ace11USZanjf/AuMKK3agqCgNriLTrSZ8d8N8DXcVY+BVgU2BURy2fZc/ToT17nF+WYgvmGPwnNO
AvNzyxn7rgznPi/SmX2s4N1L6LUdqwYEz1O/Gqe74k4HKPOIVzpKZ8wHHotzU3yOxslnbx20mQFN
KItDcO/WdaJwMlC3Qlh7tUhH7Hyefp0/LJrn01wG2QAFXyzdPB26NYWKhgPw7OXtyRgGg6KntICh
8oXHJGew4XRTY5J+quQC92OEwI2mVTcNYVbyPs4nac57omf+KeIu5nGP1zgbDIgjkA/nIMNHciLz
PPRiNKqroBfbdBbgk4Wp7wXYdOSxraOXxsrZ6AVgXQWEDSdYIaq779aeExlsFh+xsCFEdwTUp1H+
AmAhrzZprFOhwc+yUZy9lYuUBlxhHyavHAsU8i9v8g2ss+WYWLP7xfSK7YgCzWH1ohOc3PICYhLC
KJk8/m/k+v1PS4ZNp46Mh0+QJ5ZORBNcV+cFnYKl3NmH40cq/DaWu8/8TYGl+Umr5wMSE+whvJ1m
Lgrge4mQzvmuYGszOqm39ZfjnLk/Y1TLi5nCu+QTh+iu1XA7r+wBYFiUlSdLf1b91BN3Jw9uDs/n
C7VxjNX8CY0VXJoanC1vNKU0Fojy/UN+qLd8cQ0ATX7tHTRUsmHbjFk5/PcIkxuNMJfdnzdaRCoe
GPK7ixOcykPZYRj4meITs7woYRJz+d5RwT5JOMpTp7SlfOt7n8wZ6imnGiq0aaCuugSgNKYea9T8
EscaLSML0IlGz4CN2dVR15fLtGQiCs6dH4BhV/gd1etMY8YZvHAPrPTzFJRre3lgw93jvEQ+Xvl8
dWwdoEqQ5h4vKFSt7RWuPAVVZIPbbLoHuVj5yCWE/emF4v2GJpFuy+5y3K9MH1WR6/qaXlFye7ns
D+PG4QK3WHM6Iox++asat8zIlFnxNR8cs0u1E/iJGeboIcHud++RUI5Zq+w02sxeX286TyTOzWnI
d+ek0WjtBE/hdeD0N9MOPLbRXctkSsioNyZ1HHkGnbhj/nqXe+1QnzcqHgzSG6FBUo2QkAG/VvJ5
I5q8wFYVwtf2EoH7psrvTYrzb14mRym8rgFVhUD/H96DxOsNxC74b/5oeiV7DoNQXGwimT+apaGb
7RdRyGGAZmKPN3SEzKkpc/FTacUM1JatglgT+r5A4KodCUzo9K4QnVuS0dOgonwigJv+zAXyDnW5
ty6zT11hNw1/DGZS0jTNOWCWVuwwm8CEB/L2KJ/YfcUTa1882kMNuru/Bo+P/aSCVvVag6QCRRcb
FxatTKt9Y5BGUUnDwdDjzAbmmf8JGqGm7wKjSkOJKEA4z7FHVCWR7MZUpaYxWGImOO6twiOAHCpK
yJ9POgp1WzPM5pGqFx0VN8WKWqI/EiyoUORxlj6L8ARKmHbDQ0iVZxwcVK+oCXvX34QI1hx0XsKV
GRyQ//Qa+et7LXVnfx8R5caE5cfCrmsG64teD3pw+fGzAu3N7/CjMQSYaziZKQt91+kRhFBUL5/w
jnGdC3foFq9bxuRjRqEjnivmhK66Z/biiNtB1l2Ggr8xWn5RYRVW4EDWHIazTXb4vFONxKXU4NwE
g2Ld5ecMc/L/9uEILNL6VEaqTRKWYdL8KcoHgr0jNLvA4jZYRbHDZL45bcr0t8KqmKLoPssjjib+
DOSUd0TdNb20MyEuSM0zh2fC4SG05DSxX3AHteAptJa0ECGvW6HM3P3UuqNBfiB+EYVUCcjH3cHt
MF1bYr3eAHyB30hDNtYTMAK8cpJVt0jS+YNfo7NsD5LfKbLbrp+WEDze7Max8tQM9P8fKuK+wH/B
DZ63FOBU3YYxhhIBWVKOthtfmfgWWcC0/A3ip4OsGAK8pP+c9Fre60cM37t37nkLLkMJl1/Bvvas
1GCC2Y852poGVkmgsHi6duVdk5enTphbFBmz7ofp/4B53MiASIlgmjKWujgFjdTlwJdl28Zq5bzz
L8Q2uR7dKVbIypS60gYoKfIPS+tf8cf8gFD7CloKkXnNDuGFaMiNQF+glgRhd1mYAntXn63SJwSt
d69xB5GwSkEv20/NaobXUpAUno5FRiGN4RwQrX/d18EsAkeGRXwmkO6rXlO0LgIcW6Tw0gfxk7T8
r1ea4uCSWu9LpCma4KI6MHD0tJTqpuZBvyW340a6AxO5zlF2eqgwGME1HXMd079LASUZ2veLz9Ht
WoDY1huz/XFlFYMcG3jq6Ihp/xxd6CVxfQGJPTlo++bzksb68R4rkbeG6D2Yv0nk0d6icOUDMl0R
4kxdqcHOzkm9VOX5KYGLYWgKxSkgdPe1QpSr7Io+47SPq0uDsj6oYZ7GCwjWPWpIdS8v1IOa1ech
elFwiB3K8GhdlCq6h+rcmLU8GURZ83ipxNqq1OWRAZ7NsXbWIvRcAxZv4VPFekOahUW9taGGPbds
/x4k3dNRFK8WfvNpSz3zev5zgWuVg5xHIXIkLXB9tCyiBARwWLiSYnZ0viiCZARvWbCTuTmn7GQ0
UNcvNE0Rb4uLUnaJlrIgd+LKv9BvsSLBxcErQgWD/o8el8neRXGkefelM6kJyHGIA8US0LlmV7ri
+0qvmy+uIawPtinUsTWGAScEfwFkx9jnUMaE7JJwyhLR0DMVXvm671OvTNXaJNvaI98Rn86dRirn
NSKv8azD/Bxc6FRcPkEn6gHAe0hXU4KwmnXppmfSdS8mqAfGhu8oe1u9X3gPpZ9O7BTufkblRWA3
tR3+CeaWPmqmdMF+7Zmqpghct6RSD3p7s9mj4o+uTIlgfrCFF+cyuRjF/KwOYJwyUdcCF/yk2UoK
BA9qeQZSMbFN5FyHMVpMFxMQO+xsA2wFzZCchdjtVh6CGHaHk/ENBnQGN1Bj7oWnM7vHJ5Bj4cHR
mDjFlARBFmbi7qaQPV+gEwhwfJJXxCWqILVSSox5Ar/nzOB2Lg8L7D/JHIlKKn7UA0Nict2QTjwp
OlD690xdfDb32k0OAkT0qW/zuILT6sf8Fgy9B2XooJJgC0wpNv/6z3CRcK9I/1flWuq9U3+owhH/
eqUI3tnM8vO8IPqGrjsFiXSx+SxYwuTyUkKKCrPHRATemnvyiqxWa9uPIn75VtdA520LVLy1AEfu
EZFfCgkfYwbhLhNkhgMOpJHpbXshU7QhkwSXvKx2gObHGL6PM9+x1vj1UzAJHbm27i9FzZ5TWfUj
nLfnRI4wno7mfGdjIziOqafOmIHOBoNZ8PxciVd4tnrGmRHpSWKwYCR8wcAfyR+3CgFkLG+iri+X
UnGQ8jpN6U1b7coNBC9EA6tF3CD+yyq0921aIOkq2TZ0zoMRoBi+Ws5e3hdjeeSG+SJ/PfI5Ytqr
rkJ5pHtn5u4dPQ5WHDvkJQghQo/impLDtUnDpzBq6gax/cZVCTqNZyg8sOKIwWsEceESg3ywhkfE
D/dCVrTsk+dgW09bqPR9paUMoc3BstwWUSyw040A7lRVz2Fp8Wjkzv3mbTit9Ym1komKqC/+0c+g
an+A0+01slsPp+lbN3aciebcVHjRM/s2TINlEN6BP+MJWJDWpBqvOgBTIBRA4IsWr6vxCYraPr9d
gGJ+D0nIc21s/yXUiSnnGPNihmuW5MZvES5HvugdNuXb28unz8mYhPpAFVgyMOMcSDpw+dPiGfx2
zWXA4h0gE3ljhdI2dmsPy5vFQYW1foSRZDkJRuxu5FUO27J+G+gQyrDTf7CqjIXJ5d+gjRQKVSQZ
MD7L6UdqmWJM32Yy7vocTKyXVGa/e/nYHaNMI8n4uTdayrs2+negZ0Whx5ARyrR4UarKqMFbi6Zd
YVXIHTejQaJfbvj62LRblZYDpFCmv5gOvIxrDFVwpjxq48QLPL9X0a/rRhFmGvUm37QiCQWQfQuw
HRPyD4jzSS3X+myYNQ43MU3uzK6sYSgqACsfGFOtllAhcxY3xkZfUndqS3JyQju7wHZD4oZcxK6J
lVFVHn9z7KMOuk5c/LI8Dwb12EwUrztU/UTr6zjUitsr4ROcH8XoRnDLyCHXwpWBkKjtEHMzs2VH
SeA7QZM7XJgwhDB247QcLQ2ajm+vFIx7nZvqX/OE4ymbXTub4wYVzen4FyeDksOKaZkI14kTR14q
D3PnmM7C/eJvvUfVvo29o49mNcAZrbNBTUExugnVNsnXXeORGk44mAC1GR01JpZIRCodAdFLeUB8
ZEuKi6C5NDgqNDbphzMUqpNAgObW53uN9lvAwz6bPU21/6e489mygjZ2LIaS1elH963EAPWt3P92
/kpBtL7WREPnEv8FGAexL7Cq2G6+788jJXkPIHT3iF0t8Ojbn9UxE6Wcs4hCXrUOFjsAB1HfEMW3
fANDqdNRQpT1urrX2Jd8SJFEJ+PUKoy2GMCzIvsktznOAmANJ3E2pSZ0EHkqwtpEJZBHxq0vntZQ
480fq7LovXO/OG+gcKDkaQiryzSk8yExI7kulydubPq8Q+Rx+LgGnSWnnVcAvmbwDnH3Kx5D61hu
87NMDfUyiA6kJbV2+scEZcF50B7OxmgQKYDNfOZ/Yck1Y5PBTc0cwPOBvFr5qpyVi9HJs2jBWvfx
J+tm4CyOJeam+DHbMsf0gm9ap1a1VfvJrkmmNbWp4sdTdTudR+X6TmAMwxa+Brtc3GrotXqBSr8M
Q+b3qMygfPa51DTRQJvzCz03U7MYBIgRERc0Iqyrm6MORVOXg2M22fGo8poEAGcozNz/3n6NK+4U
Joxfjx32J0FIJ/JqJ0rirhnk4vkfD2U8ux2g8Nc27NVK6ct7CpVebS9ao9YigCTIzllZ1G16mY1I
0SgF8+s93LVWa3WOWVojocS+YVAOQoPYYI2OJcutae54DV7UNyH0fqoOSo/qqmxs1M9/08oVUjxx
WBJcjL0JXnDPtSbUk3qSNir28gmbe1J/GAE8BVnFedalWCOYziuTN2Dtg/GRFrrSxjonrXxLkSXb
kYmudrn+Srr5MgtgVyFblC97MaFxhS+xp6oqY/4SDwg3lEscfne6YoRwyNypV6mqJVmbDb4adZRU
wlRWQuyY25pmeDCXAcMvOve/k/aMPIwjbFYW+NYszzw4JEbtPM0WpRwGSG+AFIYLBCOiGyBt8Yta
6Bs1bQPzIYOeS91erQihNVu0j+cHu8PJOvhIj3+XSnLWohIs/RIL/gsHcu7BYiJpyCaQ29gJ7SWk
LVnHtE4FDKTLYhT0gQErVrwNVrGc4tb3QHmAq44r1qINLkI+U11rGrVwqa9Xpfz5w93YoWvvrTlW
3abGDtatRVZmM35bW7/OKUBPR3QcD1WMy+98p4pG4qFb1GBsl6Ve0yiT9kVovKkAsUt5UyidruLa
WMWo53m2vXWhNKzOOIErLo/9SVIg8aUvrAaE4QcKBmBvv0GiXmzyxLlT5701iioFh1IGb65EvCWE
4KQtUG/L6U6SOeGwOug9KUfy4j+3c4ySx/jRsmIeW4SI29fw+CEwGwqrvfJPPNFbnBkDBd9gvtfZ
64KN1IcPa8SY9FKysirWj2QKWuYQTBwdKv7IyHOYoXqFUFGSQ9GCHIBIydv3cJPEgykZoqJoQWJe
8GDbJs0lj+QaEHWp9w3z1z2sSAw9YSZTTrDzxy/3cp73ibedw+/0pRc9BDSp91Vt/PEyccefuku6
D92zaFbv3yXH2qL3hN93ogeCki9MAPhWqqTv+fjR7fkoBdHs1kHd/ySQVEwqDpVn7C9Y37+hOKKc
Ub/HU4DdvYuQUNkJFGliCRcrArpkiwntK5+MZcUG9dnSvOUAF9qlSuWjfCNcPCBTAxcsYmCADSvR
nGjJPjoT6o+SJtwSR6SUhO51l0ZyMz+7msaYBT2fibhaV2V1kgAEz46mBQD2TTWlXkyjtYXherhe
4CPo9VVBdjeFuj0z6uxndUQxqklYylKFCaxj1RAweSG6o+xrWyY/EQ/qOulS+rYWev7OIS2anUxh
TpLLjYiiLCCFi9IcaAj6u5obfjp5XtuV996R2TLqi87DvRx12uOEDCxjrO/WJvfTgmDyt3iytgB6
+x1wDGX9UTsvvKWg6OAZCBnDhP2xirgyXCw5dyE+245auDvEIvNNeHTBTo/lpHOnr6R172QGyG+F
Z0B0Qoi1tswGidm+cXheHuLsV2EinMLgsIHa/7Mog1edu7Ts78Do0kYUUk1tpDctgCHW5NbLBS/r
Yd0U+Q6r8ejNuKrCdYC64iGHx4DW95rv7wtswydF0teOJTL4Uqfhn9GkJ+BGAkEOPIAVPDfMELqu
Wi9/Yh+bU31gaUV7UNcnmtSbvcCyacRFWqLPkcHRaBABIdrn29GgAUNYjm/yPjm840a2jB8UqPF8
piogObSeNvDmKb7vYeecugD5AEr9CDAtRfwxpTvIrXjbLzjyT8CTKvrxYzdrzMmdQOU+EK+w5w/Z
O1KTCz7lVrtjqYpalKCE24ZCpnyQiJl6DmuGHgo3nVxnKA4dk6qJTZIw1BtUWox+QAAkpt4xWKKr
ZAdq3TddzojBVl6EG9WrNHqc5RI53Q6yxxcclGDop6FoaHTtuWo00xcpq8QCxIuVrM/4v3ckNIOk
denPHqWkKuSkuIxNEIps8MGS1WA98n8G5kWgA/I/uyxsIbo2DonrrwVveWut8xXltY3IeyCMo6Tv
eGFRj2pvf0OvFsHmBmfpG2rBTRZtwD/US0ksvouCZdn8ZTn3UHqfTqapQEKxU71BL1A2t8DGyqQK
+VwYAWzs5WMu0PCy/MrBWq00F4L5SXLo3DKZl/j7UkpGfICEDYW+lWlcQr9yPxNE9tJC4KpzYZ19
arJx1sO8XMN4fSnDYihZO1q7wJ2wQHgZN+Pqtq2WxzJ0BUa/ebDR7cmCBjzl0SY88V6xkf3e+Ky2
lDnxpFdEw3EtZZMHb5cepLmjczUx2aVwozqGzbfw/95+gUzsAxXAqtzmOQSFJOOZeIbMlqP1JoM5
Q4CpbWn2r9x159S7ss9gFHnO1TF+qNQI3N+xZrQzCpze5kBvOkOudriKSqdQ7Ks2909HyI/DQLyT
I/GfJ5mqMmU10ySfLhYph6AmruCLFa5DWmDeYZvMAxNrEOOpN3dr9pRj5f8bnQTsuQooc4iYlqQo
xn8i6RC+FsVzTvaKgfvr54RudquTlU8bMNIz2WgiZLbG9Lz16j6iPDjpAAh7x1+ldRoKPrRwQf4j
43vY1rlqMUMPgAAyKZSWbs2GKROM+9AUSay6eI5hO08y8r/VpZjlO5O7VAFX7KYRRWYNk5UemQgr
odUHkI8iIExKxZ/epRMIhqfBW11OB7BcUf+JKo9bBcHyFcnYox8wZndKCCQmHbaWb9+ucwKIf8Mw
hkBJ0v0UoioMjJSPdkzhUvP+KayR1iLtPrpvMrobWNq4G6KKUPt3NSPMpYKumnTPDldpT47TAhUW
D3D3PkrGFIIY50K9NhUvaHjZd/6IVgEIETIZ1aRHQfYDSQQ0b3lALIVmjBYsN2rPQ8GCKDIjE67c
tcDZPPtYwfEfmVrGlsTHC20coWBlEhNEPvhjNuYqHk3+/OCrpdGvDrDOQrks3fRPZJIpGnRWevIi
Z5D/QLFo9Ei1caMC6GuNm+3sMl7uLARE8K9U8MczRw7kFXDbdEukXNE4mvIC4EUdUhWbVOg42Zyz
/YhctSsaNxCX2wq3NTcJEc3Nu7OV3VcLhO1znV2aqdIG9wJ69kNrJlf3KFfylhmTnPwAIo0VyRTD
WODhbqemb2Vy/GBxPpIHUPEgbFyAXISOBeTUTcNKzrZYqVzm3bkqovIKhIN16FQSCYbF9eOXerhk
bRz4OtYJMhEzr0fqCJl9r6eOp4iez9EPsNImq2X5w/LIJFeEj+K7YY8wLIgAl3xE7hrnrCs8TDI3
1A4yvLTCvt66sPnW5nAe75a6SPChEWPtUedcCEm6fCz9kBiihU4eUFtA/ZBgVlDhP8KbCHE1zLSb
oMNeeAGQ6vx1qKEVpn7F/uOLvVeRGreBIgUGjiSJW+WDVzZsodUNo9z/L8CUCXcIBh9rlTJSmHtc
LUg1j53e4o44o0F6NVBThrLmnfLVME6V9BeqrEEHa3pJja8PPBnUqpTxyheJ0kDMl7VfsnKfPigQ
at0f1MTV6bwE6s8sS6JDgHgfYU0CnOCkA16PEgx179IKvT3AEohhtY24l9vyNhAWluIWgciL7gL4
lmupZsVKwn/51uXntcNV+jwIe5wIugLrRkWJrAkOvYQvE9UbDvaXCygbbox5alyNQ0G2XOGj9wto
p9v7lRGIXd7rOmclhYPBldaOMXYI6pLRqe7qvoBOS+c5SZBtYdCOd3DgSXnOe8Oyb/nrQgRXzWwX
bnna6lvE0tWudmO1+iKP8Js16MHgGAHN3yoThA9lT96lhiqp9vxpQFZa1gRg9jBr0WAECOl7MCt0
TXbSWQ88lBms/0EIm9ORtkmITmB21/ykJBH1uDWVADWuxUUARdfmNuesAdaIiBAyjbPeVBhE5knA
O24LILfJ5MMr8bTeTiaGt76jms8lWoKn3HGtkeyli20k9m/qqOP7N2gaPnsVT3YmE3pR0/2Hn8Jh
/dFdn2KLKLjIVQr6AEU9QQIr4bmzjsFl9Du8kpfB13JxJ1g0By1dIvwVLmZJR5FrSVpGHdW2zvFU
MYRpy0ZGlhV2aYRklqR0AJS8xrNEjYno+vWwFvRpbVy9EG0bFzhAq7pgw6+kj9OY4lcPMUUmtfcI
ow4H4ir5FDA+TdZ3kZVi2YA/VWptt07PAx0VBCMz2AJK2GuBS78kwrFW7UiiK2yZuRrzxBLBJgm3
eL3YhoCgT9eGswwznpb1FUt+P443HQLikvKgQdUm1xVZYKFg6zh3+f47MDpm2yIMPaEnBsYzFUVj
N/Xn1Ob8hASOIqeQBECRgaSzEFN1i1S5FDen20nI+o6ZU7mbc9lLFlRRF7oaXQhjVk1MOqwNUD01
/P2DfNXjAVH4Ovanpg9XSyfpCQIgc0lfGNftdFzbkNC6Czn8cA1lJnhX0815HDYb3L0R3Iynz8Qc
gbipXcaYfi5hsF+bCOv8hvvVtyIwFdEJfncDHHrqDl18Dd9blUckqoSCjd0pZ0BkjPoxMMvD7D6T
vt9jTJvK8ilAl3Px9yNceu+C8yN/LulGmzdQZjN1OAy81WBsh3cEl/fIANcioPRpqLGkVnKODU+V
fT+XvRbRSp9j8wJIQntLHjapmMt+kBnTEuS+LlEATo6neB5xZ9rM2I51IrepJl1F4VQ1eQdKIPah
f8p2Oq39grShCCu4UHXnzENJ6UMFclKMpnfZAmLZ3YN86R0pGFLRPs0qnRiKDWaVPUI3jl4wY3sm
MVtdWzy00XNCfr5g/vLxc8APYayc1U2QW35ZQy1Mm1sIk0Oux1XUMRdw2YJCL5O7kXq7E9n4CCtQ
wL2RDfxJIpPJ2dhMwnzFxuqAHz5tIWhm7zImoUdxJwj1q+cYapTfwmbHB1yG1yrRkbOcUGfcWs1E
FucXqTSjM8pmYsn/X0tKPUscSU8DslC2unHjzTadZjlD/JjuONaAXWlk+nD/DI6wd7pQhu/xa4nn
0pH1jlV1c7GeSQLK5lxpsjbDWA/6tM9fR6t8ubE5DWK8N98s9DUeBK1Tb/bDPHoHnVM3WWBiGgKv
bAw9bN/zGPPxqj8bvLIop/j543l66O8mOqhQN8zfIht/jti6LhDvrjRy/fUlz40NHZ4R5p0APFSA
Lt+Z1EfGVfWsM8aOtlksD+zJUn40a1t99f9bLjvg9hk+HTt/PrJ1IgAG+jprIFiJEFmFPVQ0DAIz
MY7Ztzko3vR+u4lyiOQEbNzAqCL8MLCWKTsUTA0ID+DgO538l87lWdH2FY65p9AvqJTBwB05DBxf
DsnA1MarHzAaB+X97mCJQEFG6e0Tv/GAUtXOLcsYxsw/92qaEJDJKMH+Ew6Up2lpGnmKm+giEYwt
+6AMqhAjnGsVEF3xtoDJWEYIntCUXi28afIqXw/YI2B0Qhg3nL1Dqv1W3tJ/Rg2lE/q4R7vp/E7a
OgogXOjLD77hCrlh9BtdEwdazuGyN+rtJyDwoUHLBX9EYSU3nMxf1O7K4SRJ51QmGQoIwRCu695L
l6/OcRpKgrey1vQbjWZjiydnwhJU3sQtgh3UPaRc+pNQk4ebfXPeYIump6OtNInh+e4EOBOQTBVx
i5UVLWiGzSt5Juf0UPSKYvxDyRj7GS3fLjyx2CPTIUh/iVrNmaPLq59hJImvEOKlWp2cHtY99dlJ
9+ICv4RTNhA9dob9mZJnFL4UAy3L8+LuR2lMEL0LkYyw0mdNNrv5XY+CcGq/CTwRxJsuZFwMjKo9
VrdXcmdqEJ46vmZjBacb2tav9xQcXWy3Vfsu8xth98/v4CxQaLGfO3eU47BIU33z9hKKxBMo0CgD
G5Qhx+2WUPrd7UbYMpWqyhRMcK+xaSr9xNMVLvCxWx8x+dW8GkuiI1jWN+Hoi6BtDs3gWYvaAb+8
y/sS+0X4IaMakL5vdqzYji9697QrFu4Ei8LCNAKblgQRGMaomt9ebcMztvtaQccuMhN5UeLSBnlG
qIkfc85aevclcj6v58ckC2HntvZFLMFRfK4M23eMIyR70cwIXGRlb3K5qXrphjSWQLg9dBLkbbek
Nk2ome7Nuaq/F7qhCbp00hCwbloSZK1GPlM42QtrsPGgZnaoONcFEEjs0JKQtX9IHyyhu9Zm+Onw
CjP1vx13ga4pTmhf+ikvxQWkInwAKBB0XTXXi3krd9hSkSPTh8NpIowDsIp7vvK7Zf4q2gP99MAX
hTzx0gUZLLmNrz8kYbaGUuD4Ce4pM43TXM0jNnK4dkWhuelhOUSLNfdLz3TOa/GUJEE7bUtS4ni+
+L7popNrG+w5FiPaHX6Yf8aDky0Z/WH+vsJhRJarMJ1dN3nBZt80LpxEANMkAGLAQrrVIHM0VBgV
K3APxgQmlB9QFMEBOS3JVD8ea/3qxlYNWUav4M41eI2T0VJTrn3XsV910sCzYzKi5zwVe929X9dy
XLtJNGfgl+HGKWoLjg2xP/0V13Yb/RWvlTQVrRWmjDPRYbJbNhnQ1DuFOYO/PRfJnBig8J724npJ
f3bzVrHXeDXF5TDnlvlLBpH1+ahOD4UlGBEV7TLUnqFaQuqZRc4kh1Watey25wC+1+JRgpOfv+K6
7xA5foTDtz0mhmj+Aem1xVztWzP5E3siO+cAm3Ia9gdPmolW75y+nHFSlnwM9Ynb0TWYW8eKrXQG
UTODL/UkfToOnZNmjyB3BbPZ5PjKH/5v//Akp9GaPKiQtjopm2jiBip5bC3As47Qa7+sTHnRdeWp
8CZ3xQJcjTHmAGy5HoQ8wQ3a6ijdSV7aISWDhi2YzlXmwP1vv7OA9Q/hPurt5NnTJkqYT9G96uRI
oQubWBN45R+TxqCg0y9jQ8HHP4pmZ5LQKTyCDTSFxsFpmqjOS8esJoGaoCAX1h7aw/T2JdB4Ea9o
4T01T88ptGu3tbRFKYCyGOPssqnSakYKFWHj55JinJ8LizI6p5Wnz28W0rikA3MguU/f/bDJpA+f
3wljWHa3YN3skhmGUzItCHIeRRQH+ELujb2/WYdUckwb2oCsctrvnpmTYhw54vwlsqRiVlCeyheJ
m7NfGRZD4wYGK78MaHKSl3XVlmD4K0g9bCuTXBo4TDsJ7CIFj7WDP0cT3/AET4xgp3QSZkx0UC4h
ShTgTBKsgqUfB7ZDqPQI9gAsC6QXsdKCwycPN8Is1/FNAFU4Wc10k+3nkQE2S3w8lf+Aln5qpjI4
xJEpLIETVYK9Yly/2BcPyAscrnGYCMADM7s2D4RCwn8bm6EK6fLfV3OyMNTHCIUb/pFYodgp+CfU
Uu2O/i0FX166+twi8iyy+2cNmM/FiDCDjQDjAHUQYwl9NiV24/LX+ntQYl1CWo4MSlQTKXRkcCDH
oio7b0vLItnBPMC74cnv4VmvkseQNyjGVBZjExGtMVecVGDsZvv81fYZnzwvmriLNFdxLUl7mu+y
4MoXCzV4OJ8shZ1kdD8C4+REOOZGwSpOEqIqiaSCf4ZSVH9zFJ/cSMDt0s8nKgHsVwYgTBWndT0b
xbLQ3GoEiLm9256BRO7noiOXrzrNeT/CuaAOfHMK6ceLItZTbpBUy2h69zoSL91WUkXigbr6sBHF
MSrvAdlGTEabRgyEjHEu5piGbhVLUcEdFZGz83Ici14XNonRnrepOZNKHIXQLjwlKKiK/TFcgQhE
lFQO128sbyEskUR2ERdwG+Pe0eyHYv9/zMfv/A6CtB0H6Av+fYxPSc/HWSNtR6mJEfVE9vu0Kpf7
QTR5iXtlycIF/yJTN1W44mi2lWzZdLbP0KQ7YwRg6S0PJ7krX5bFvlAQTJce1XscaiuDpXAZjJmV
gCZnA76RKqWLjiucClZQpwE5LwgRQ5GX0dtDoxOGpSILu2GxCpemweT9fK0tRoaO6AS8SbhhIkbU
cEvrdu+Ac0er7DdeIwayFpr4xM9hetz+RLTFfKdA6vd8SA2AQ9v1ZGm6b1VTvcIPeje+5Jn1gNS+
oovVtdt6Y5NVra/+Zt9Gtw3cjwrKJcyKmDQGYst+htVL4tvN8y0402FnPMxWgSIslLmLJGFofnT7
6ls6PEotURs8iQAEk/VIWYG/9QcuGuGapo/Ft1RIqExJNBL6bDRVhlhPx0ah9VpyEbXELsPFTR0z
eBcpH58QvoyKpojtdY3xq5FBzM7bl2FLJH5OI/dMUVkC55BIjgJKtZqbd8Od6n44KW4VvSM56C0t
+sJTToPJHzt1vQyPcdjBAepQCQOoSm2JAvXSxYriDPqqPwekhKmg5C+RKzdSWt2PRebyPwRcWfBz
fPx3z7BZhi3IUv/IXpAzjTSLJbQVSpmm3DKe0gO7gavv4ZK34sTRuUuJ3lFvwakOGCY+gYMfMmIC
E7OkYDVh6VKjYLVwYooUsp+qXaMS1IHiZ/Yr40zAlWdQcjBshJyBNeyNmXZgHBE7WEOLsS3MVTqq
U4fZh88qqovJhSXl1qc4Z2nPuc54B8wIB8qsEgusTfSzVOJrdfRepnJEmVTpFiOme4zg0fw3XrHT
xuTn4n2SunXPLmN6vuefkg8qHKe2BxFBOvZ3btLj0YJMYhhUSrAMaJIjKmNYw3xlW1BVKI7HF6f4
pHcW25lsdZAw8VdPEzuW47yEvnQkeKyZLBvEiv7TmsMwAHyMeXbLPiDXZQPhG7SI6Nnv050ob89r
Eu/sODZCETscxtgr7SUSxxCfm/EOIpVhbIuSEtJ73mtDiM17fZHP6vqfhVyjm8xTxDn/0qCY7Dzc
fO4UVPKmoh/1D7QfM016yquprHj+TqiZp+Nf87vIZ1whEsxeN1S+KxwmPRsiA0rV+It8Yu5tA6HH
FJnIFYGeUrU1icoZAJZTeatDGSF5aogFFPxNTPPwyZ2SqeWQeMl+oo/zeaPrdsW8RvW68nhSHUNf
soah5ru03SNxlWpQffoyhjRQYwQxRzRBMyYMG7vKWJ8ysCIYqzViRXZU3/uoE+U7gKydECkP1klw
oRlkYZ7co0BA5GCEH3WqTb/6u8903wBv7dXrdGg5D4wIgWvZ3mU2zXn8DhTTWqqDqdijKvXqjyQS
ogZ7ufcTIKR2Ihlq5m1bkPqWCzLoJnkLEaZHTldUA4W2eLVULVIR6QktoM1n3UeqXxI1wvL04Oa1
UdJnSdNM2wTffyKtoc/Cigl9zVaE94/RMljh+Uqvfi7LRFF+VonR7gA/JJuinXAO2ntO2i56fVVq
LBvJ3wuOof+3jxDUDKfpzKxY4Q1PcWy3Vw3t3814diVQHFs6xIcNnJB75yL3Sn2QhHLAV153F0la
ml/VlHgpQlNzqnyhUo8LabeUzKsGPwQ4xJj8z+HB9cPYgdFdjVZp8jPZ0ao/URZrhnhtyUN/o48g
KexSc02ly87sDOkuBzM9HF82SXxN8lhiiURWGwMLu2qLdmNdTmFFrGNkmpdUpc2Z9QTmkDkTGwkU
KNafG1rj44REgfOIlyDEXGdaENza+w5Kgr5KCdPuhKle8kfiJB8NlCS3sPRMMIUpiJngtzGa2epV
4pelyGfA9N9XXhfE6i4WDr9zvwsgSmduj/9EDN7/l69PNZbkbU8TsWLnOZUiiseXCGUMlcONsUGp
CpUWbpDu4l7DjlwRk2Vwx/rThoXmm/+Np5l0xrwUgiGjxfpoaSZfS+jpbTienM5QcOCnthHkZzNB
HyjmrFWFB0vnJki/uoDEAkguWfJhyI0JhqUaiP6sGLihcdX2bSJPEeIL/QcCSupx5nQB4ISqs3YM
3ohbhc2PEvrQnCtiYQMh7U57E83gmGBYnriVFJTF4L9ouGdwJm2mo9iYmoedxW8lXNhbux7DZJzF
0ffDUwsIjdBqfk2s1m/tPcZOGfMAMQzNGyA0gHrbVyZe0N2Rk1zTS+dC057mbxGrDbSoHmmtiW+G
6DkD75eJeWlY7ChygzIUyNMwmrShQf96/ekTILTAcNUeR3Kh4gr6WkARTvOb0wTcsKu8QlNnvvwV
4KcGg6Wm91JkQt/oibXNV5YlTNw7smyD59fj5vX6873mVgrrVQxwg6rklXJvPazA9e6XH8ohBTpA
0CpehdkKU6IO36drraZSITeU+Ne2WUOSdbV2B9TWfckxYVaunjRsteAtC/apCfmLEF5iHJfwpEyU
1kUYM4alXa5xHO3Ab6cUTtVQWfUT/8L3Ev2WLVdP9Utb7eKUsJ6f2PijB110vdOT7nlVzmAI/My4
HCqaDw9QaW/UD2HupS3ISzoZQ9bpTDO3bJcSDRa8T717un8araZwh+DQskf0ou4Yn1z1MbNxJyWn
kTVWNbFCeDBXfAbaDcBhCZaIZFgEJo5SeRXi9LYGPj4ZqvvQwlD5tg4sNQLeqrpLpCcfDKt1yprm
62ap0adi6/Z7VhYg+26WOMHgYhS/Hn06HXBmhEb7YgwAlE7IP5ekeYW5wsU8lnG8oEZI1o7P1EXb
p2DQxwNTuwD07qu2Lp3Y4bRN/k3/ABPMx37rsORIAJeVSHGlS8ZFoFgcqAhhJ0jGbnLbfHONAT36
eGnJzhRIIL2ZJpxXDGyWkshVJ2CuWZPPBhhxJTUB2uYSBlj+yIN3wn3pYXQ3dZd+jXInhfQIxPT8
Rl64GaML7dhp5nEk/msQR+M/Bpow7ESq8GW5Gy4UphHK+kzu5V4Cv1h0EMWB4WiYKAJ49N/bkXxE
mkhaWZAlnYG5Uwj9BEepwa2ZueH+0iI/gL18DHSuDMH4syL9zFpxfTB1ToVGOo73Z2UFqs7rMz86
j8+1PFfJrZ4vUuAYaRTt4J8YFXlfCwyLRbfCtMGBtGcF90kiP6sjnkAslnL4LWSxP1+ZVP+4RAXA
pWJ7QYv53r6jAS1o5YOKtvdAvZ7QLlCfT3sQp7ycnPk2gf7Zdqd5g38f0U2gNKZlP4Hc76R4RquU
FZqEvPhElcDo3Zh0rIDK1XeKP/iICPSoW5a8bL456m46bohp2aqXigVqpdWGVumT6tgRmcj9XSwR
vzlIx7/8peT8lujciHAJLCTy9yvQgCJ7X2pSPEp26ccGN05b2CHEBngaT21MxiAJqJvxrEs+8pLc
mimPICPVREPPFQ0+J3OvpFYL7nRAnRvGZSNOeGNmxyy+vbfejjnc34XJ/sL9qojLNEhvJkJpukdi
4ktwEynTCAdqYYiKzwgiMZVpbCywhFzRoT+tvYiiz1Aqf2CA+Fmj3C509xZjEUReh8v961ckxSRB
PhzRiXRWseBqcMQrxQYoWhS+gaCEmUYQzVQ1EzbGBAgBXcyowHsvhA5lVuFzWnW4KAU3FOubKwV8
rJl5VmSEN1YxCcr2UtCD9ywBKIj9zyStUCmMoc8nT/qkSgu7j37g+jn3VvCfRsLx9vTuBrZfzsb1
VfvGjlVl/82xlNEiZHrEXFXEORRqC5UHUY5IDDK6H+nA94XyilKdE1YJALt78ItYXQ68Kmfs3w8X
M96OdAol7OOVF2iCKThe7ZOkWUTx2pyWy2xipyRDmIwWg9SJsHrb7OpkL1km7xBoYARmExle9GzX
+AXsi95ItyoyEH+XmrHcc4akvcFFieFWnloVs7HbYdgrKCwDXLN40GBBU+4icFf183vHfCyeuzSu
MOdN1xxcknZejjtrRpjr5GEg1tHmNKNIR/KnWqKAMEC+kRJYRvTpYcfu1wQcY/XTbAgQADVUbrnC
zVFt8SwErMWWFy7Rde9v4bqx/Z9Dvx/WDJ6rZ4B3Ana3PMfiVP5bEx1nK49h/qZPKc2LuW31SApq
ca8VfkDxNpSKbxKNBFC3QL/SGqngf+QEvZsaxaKaCQ2hy6bruXTNIioxh1Yibv6CTL/Ih8fA2XG6
e8pLH1XOLwHPrBhG+Dnhiu0qx7Yjo5uKJTANwV5eQIvoRucilgiuU7ilKeR1aXvAWuOtiDWfrPVb
mbYwTnwDH9jcY0zJB+CiIkC3geI8tuPuU8djAMDttiihPK/ZlQ6KCwpbTHxxNESAWtahZRtu2E0M
1Py1pxPFoa4z55ZomIbCwNbuCDbjLuhQvDWhjmQ/yqvcVNFR5lz6B2Ft10hYfLw2QkJ8sS0oIA/C
/zlWgL/4yBGMjVOkr1O9JxljPyvX+OfogEd7K1/kVkiEoqykSMOlAmIpRr9dcSuNVcwxsY+0Cj+v
OtK1J0Tw6XP/nPxOXZSWgF27eir8ljCJU2OAJRA2IKoaT+T8C1+yT1r375lhA/Eb9ah5NsN3iEMT
hR4Z82pXiT4xlcoZlTuHqy3nDgP8JiBlpBUQ9PWFJhot8LvsYnsL9CFKDfR0XW+DI8ZqI8d+uUIb
sXGOx30zwwHHXYyOuh9qh4iEPsFsYRudBBL+opjWmZXwAuchIj+eHZRwGfcXVUM8aE3yS1oz8PaN
vI/sRN4+iSah6ZnIvFclyZPacFuIPJsk9Bk+EP1edXtQE7QJcoqks2mN57uEXg+Up6vdl9E2v48j
mkR7XN9u+eQffssl20aJOIPiK4e6NfO1WUO4EGvjP+HMU8f5DJYTg7/siMOxkDpJ/tRAnXuikDJ7
dg8sLHyfrFlpaGjmyq06zSZWk0Vfw/DtHwWYhTG6U5VFX90I4bks8gikGAeGaU9KTsl/96RkQw7k
FTYTQp1iqDr8CNFgKYF1Yy1mv0XBsPnaYmhPCZVPhH3pM5hxeL9lBUeBvsjDXzZjIOemNgn5lEwK
kgytsX/F47ztogO8X9J4KIxh1Ca/jnp3eooK/W1PT3J6yOMJNrdKC4WlokX92+ZV1XiCWILugPQo
YuaTmvqq3dn7KvUFfe+1liduj0lE01kUjSD4FMaguZ8tJP9ERyck9yy7WFj0M7U/1wiCOlKbqIuV
NcR6p3iwnnoeY21jIB6a8uzpcCfdod/A9S1TowipgshuWrqvboblfx9zyU1G9u1u2+4Qb8DAf/ev
meQ92puY8/UqqsKeOGmdtdIEKXJGa9VCH/J1AnBlDI8UcQ+BgHBLcEjCg7GogDuRwPvNF2Nc5UiE
5fZUcGops3Bp09nvY2Hc1Q0czt027Uv+vlbeh+alOrDPSlx3AmsQGmAL2ezjzCm6fT/50U1LHJt6
++eQ12hoLO2DpIcaqCEPqXSEykYdPQtAaHmjLF/SamYo/mP4869DhXRNLe2WatgEmQZA0HLyPIqu
tIjqdWBul/hZfflcS6H0wSGN+9wcb0EMDuxad8zw7RzuEVh7svwGjX+chHjy7/Qki+f76hbFGLIP
ve/q2/2JHdN9tBCJQNKnQEn/JvnmRIxW8qB0h5cmzkslIEXhxgIk/3zPs1acFehKJ3NbumovvkD5
7NHezt9THndV9L7xOnNEJ86X2D0hJiBn2G29bSM/Cqzp3B9xgJXD8+dQUAMjCI1lprZ8HHBB2fu1
34c1BopqOo+oUT7RVz06P0ORQyZz//1LC5HHso77EmU3jOIhJEkbEma4e7W/x7X80rOKBxeBz0oV
nvphEH7ybzGb2PvWv5u9mljQNOubvB9fL8QYxvTWRhH+TiWVfr2mZcq0CmF5sXPh3rCY90tABuYH
o9zEM4GyBK8DKQu36v0ldbXmpk6mZ6Qur3y+ObvaXwvXU1yI6N/QT2mv3Vp5b0h87DMsUgrRGqGy
uttXdBITb3zxk/TIKt55XpXPwMvx0D/2r3s+u9D8J6748+dC9trfMlViK43g3l3+05HyH3EdMWdZ
vx4iTeGBKxXnrwCSec2zjmi2aesjD5JpM69Amy3f7Y9KXUciwZs9CsJN061xJCwanNAhMA2oUrxU
NTIARvpCry8UU4Y4lEAGjgIBNn09bJRjLs3LW1FKoBdmeza2uJAnuBAkACIBQuYDu0+O1ns6mP9L
hyJudOXxB0LL8J8wBLknyIhcVBrvza4FDm6nsGqnCrmfrEO7LZ0AxEbfFskbHtAIz27Lyv/25ARa
WKoKaBZej5zKzPI7ccrbYbvHEG5CqLpv2fbdF1H7DruApwCUhv7xn1HIUTYLn61FoO8EC2gHgB/E
exYxgcJ0CY+bGjXg52inogoJqPXzX5fnNtJfUK5ylYvNRJzKEv7Si8cd6pmVIAHkLrvJKYIreDgS
wJIwmeZI6bu4G0Awt5PoU2mTDdfqG1RrtOmLcn2WEFLihiZVvkQbGaNTK++rQeV64euytRmiSAw5
sYpEdG+p0mlHi9Lv6AbntUApAPSRfTZWjX+chtqQpCbUh216uTev07OngmgiTh10BgsTWAMEIvTJ
RxFPU38mSqqEAwCQykstrVa15G2DRFsuoPu4JBdWCXMwi/d6G9EeBxoTp3PSsGrXi+tuPqCmDYO/
K01jHn3NE2JP/fE6PyERqP8G7zSQ8N8YL+XyQYP1VOtowi0jENUecQuuqVucMYcjPjBMQlmtIujf
7rn0PkajyQ2/A1vLSN8jekOR49j8tSNAMB31lFVL2JwVAsBwAtFT3UvMIc3hzvb2i2Fz7002FmRB
fUSTfRrPjMkCzyJ7OCbPshAVf4mwY5Zdf2KJvhgmuEeBv9AOIHItfZSqgaN+v08L19gWdGfd4zCU
B50ALSzwVPtSsJdNRHb285omw4PNHlyKNOnAi8R0KdSLaXImYiv0TzzbUJeLjFouwl1CtWHN6H/9
60f+04IAWSplX0XJ8YLu75b8WqOK1v8tJ8z3TekS8nzEu3n1tgV3yOhPYavzl/4RQkmJ3YAVWAL8
ghFTFrJrjcLF6tu5tamTOTb7niyVc2YNQO0dpkj2urG68GMDTOly3jnklRNJlksdUlKuTjbgCiWH
r74UH+bEdNL0fGIde+TYK96ErbYuyuuNBmJXhX6PnsK7epAWIYH3R0zwc/gWALyFwh7iQ6sniCO/
mjDi2j+TikEs2lcvDA/blSTP7F3S18hDSK/McJxt2j9quC9dF2u+3JWgAyMUIiVMWzJjZokn10EH
VX2/s4q7kR3P48ooXjrYdH0bUUkb0SmmPrMRgpbOjj5zuMrQI3odsXsT/r+I827/d5FCQjpdYCW7
Gob/07GmhY5I/uEuMZYQ0AHl77GKw3EkF4OUntCOO5bTlzu4icgQtxOeCP/1ALq6G2QrAgVfilzG
KCEzBUN4QAd+p5I1IQQIuRSPjD0kSzz3eVosmbyEkOM9eYvV8Nce8ZkOiURWolk/1T4W8Q5E6R/R
a1abqT74juGf+8bNTJXNa/MA+BecFK8zjmmNXEPdUijgZ0Bb7ZrKd9H9C+jdlUZI4ULgF79hFXfV
MdsOsN0darJWMCmxmmfJYAqSkJ6mTVjwK2KdlCLWQfRyKx/E4B3POwpA0+VF2DOkxSroHBNzRPSp
NM83hHP/+kJUYWrV4ET0qcpNpAVVm2SHiO9I6gIpgc3jZtd/ToihMTC3hMqtAgBRYtLIgBgKTwOu
QBkcjijnWk0mN7YjOZMmevygDwcl7RtsAsJa1Wmh57NTD0RxcQh0flh4C6yOYGBIn3cQC8rrlsli
P3HOFGlmZ64nfSxrfVdpvAkwm+OIgh0zwUJ2Bdq3YsbOZAqWWKJqJIGnDUrjbK0M5/GYICE46ee9
KoQuopOZHStXYmzv8hQO8RwU9GW+SSDHOjf3iuSXkEkOVgWs1VLsUFvRSbpP9MHEaqky13kzqIKb
htgnlebcT9Fbnhjj0SdlJbJ8ZO7OgrRyRZCDaigMNQL2kcGfm7zAMBK4W3/7gQGAfheBijMkggto
AotGd6EKCtnRdl2F6r5WT2x9pe+XNroGsFoLjpwEKWACp7z06IE7MnPfx7jm0rrgIBUtVd9eDmGe
MsWrhyLneVgd7fr6jmFmltOWhn+S8HWnBe8KK2IeG4ALVSw5ekiGJE9i6QYRbeNH0iG3ZUh1Zktt
8QsGdtRQgszkpTqv1qfaSWQiimFJrQnaCP7sK9wSWVHUf6/tESXSx0BGlgPdBCwdIUsRsVG2aHUl
ilBuXG96pxUsXwrvYGqbRhGyvGmsHBvGcOYWnh4wxEGwekpBAOKgFz93wr8L7EIIN+nmsygmcO5p
+hapNDd/W1S6hMIuLmlK6PRRT+F33xI5bz2ZdRs8d4GJBN1WKl2mQqy/0rhqB5XxH3lP7AYQWZcZ
m0eEiFxr/NG2f8UI2CxSAkEhqVzcfjiEtcW0UugLu3eZ2kHybrZ12nrd9cG5v2vfm+dkWIRlJJPk
Q9Y7OC4mldp0744q3FgAxNKticCQdyChr5VCQ6iA2s44lN2ucZD5swKWq4osYNP6svVUcH552w/O
xnYHa9Npbltne94w+6LsltRlbNdY9OOFAhJyxtn9ITwR2ArEt6DhbBBpNw+nVa6C59qUAALfGOfv
XUCDe4v3k2PRPF7k+UM2mSJnFjsqbqGGea9rQPzg1jwke5XOPRc4VUDgACVLliBMzSS5L3oCTkVU
laPFsYH/O4l+HJOJmGvJPID3wK0I1dfynCoYgxa+C/o2SYuy0feHAUZ8hZ9l+p8Yr9p+h9DHxjVF
xeVxdTZqi53dBK3NAty7C2uHnof6avsUOrNXlugRwzRvYRrgyYI1EWAUD2YaXd8ct/voDbIhsTXf
9/JJas/ltWMKn2tr0V/bhHCuF4FtsVRXG7CNtPfpa5x9cccV28SYNhnVJAG70JtTeM/q7kEduyxm
rQo5t1qvyLnx8rf2KveXn4v6tyve/KTD2EGYlJztgzb19wTCfUgBDrQOJQmlcZLsjEEht2O5gJIE
tpc1XpX5SHYKOTARY8ys9Uw485OFH30oQW0ZXzsRzmpRQxgidrhNH7/caelam9zvup031Cn1SGFz
ii1PIht3SkXpa5/DXvOR/y5bpyodMNbbHLK85Sgf1pAj0fEBsrQDkFPiYoQJ0vBgJvQ2OUSbGW1r
xntfmCfpyRbDA2Wqm/bWD6cIYJ8/mpT5q9jasZ7pFaTdueZX4AQh9DK8oKkaxGJpEvXdq3JQjIAs
0DdrNgclSiR0sNo20yJl3AHJfFsX3H7RaQESBvbZ7yBzqYD/sep7W0Fss843v3fbYvWJ6kW0yjTu
+UEXiuQTOcjC2yVwfMyR6oQKZfBiirjw9p7+DOZL8cpWvUuVjsoaqb7S02azfbl4wJh+xojWIVPa
CVr1C85+fOJ51vtxK5Jc6b1MclonnXynN4AWX25SHMAD7FfanbKogXsEtVCYwI3alThbBl0ArVaw
AaxbjQyRuAbddI5/g3X2Rkb/PdlWwjap0IC3OOsp84JBmsOOY8h2FJXJ86k0aebcGkkv9ow1ByAV
gg7D/5S5eJhP02gIK2GYW4k1byNYyJVKt4K1NZ+Ydw+eWgUtL0DBN56KMzsu8/rfa7TcYkFt0/qL
mnfVEjTzvtYvAWBba5EQoPoCozlkQsz68/GnvyD0mXrbnu7DidmtAKdEsdl11fJXagUyeddzZ0da
+6WoP0HlJuGqBpHcfhjnfv306E1xLD06rmcZw6s1s1yART8sea19jxzElj+Zn68M6GA2XM9YJM89
S6f8rfwz3UCv1E3m6SCue/jpZzR1KGCLB4mn2ZqzxP8dgeqBX/VdCXcGPypaiPGf7QMmChQ8Is3W
JVPnSz7o0djzZ8aq56MgAyW6R/KRvt3BlHbvO6yymlDNfa6u4tJC5DQBwrtGQv5No/9pw3aYV7o3
bjBCh8yKc11o6u66jKfZTqPWNHKmAaAwvE/d+HeE837QeWGr/BFSueVVzQjLmQzKngk0qH5yQuCu
eaytAcVnCDDFzIMtNMTpXOdqSsbNPaiueX4VsaFQ4dk/wU36KEijifQNjqZoXN4jj3kAxroWSSCH
8YgPLTeoWnChtPVm2Wmf0x7jFzr/AlowMDTDBrrFB/piT7M3PAVnEFhUsXiEyFAw2wLwgvQlqGqv
mth94iGIlujPszMVjpayavyC1fiMR+lLl05hJL3h/ddrtut6CvUzo1URrPrNRwglB7leKAtvcFXQ
hjofjI9ZL9pM2iyb5RrcJNNh9yFG1GUBt406emDxplkvhazppO/zVS+xNjyjn8WjrpwxMjTN1RMK
EsOvNgizGh2Z+2TM8uhV+xFMr5YURheM+lmP0cv5HI9XgXa7TfaHmzDg15FWZA35jLq/nQRNhykR
wi0PLNRtyTtLh6gRKsfEz8rEZfDBzTx3adi2wrdQQXzfTLFhhHwBU59005sYRr9JAqV+CY5ACEYc
TcFZ2DnzIEOzjWs8L/kxffG940vgytFZlnHb5PehaCTKIfxdK0esqJTprWOFpkh8U24mhMZxAUrE
clN5E+yTPFA+yd4pm3Do2RI5VISx8SGR27y7Z8oDxNu2i2PvYT+jOQhcpOWh6b5qUhgDq+UtpY86
X3htkJUqVwnnTflpis5KGqbpy5iGw2RTHss/fijvNqNtHN69vx/Fg7ajcLlHG5oXTAtmGoaHDl9U
dXY6VKTI1RdDZwGI2JGTsOulZsQUYa6vhZkdqKPLlswDEK9thfAv29ttX0gsz8v7zCwFvpryJviw
RQZtYnbyar1cNMOudS/upawdbR0wPDEq6ySUqeNGnPmwwYh7I/onSo0N+uHosFqFI0M+TMepnQPf
ciJjbv1UZQn4u6j1IsOp8XYGq++bZm7o2Xyc6M5YPfkVKsOV/7Xjbm0J2lXz39FKZLDd2RAbf6a6
tRCnZ+ztWTbh3W8EgBcP1qG0n77qrqTq0yxVr1jjoK8lynA0zxxQAB2mT9KXXt9klHsRvqLIYUPC
QdLAycssbmXvW7KbEGlLfZpHhOin67mKWLcU5tOdgavtMczkG26ZiCgMhpRZ5r7xpyAiwqCj37wR
emdIXPfDIEod9iR/WEwCf0s9v1CiUiCamua/Z4j7B4C0gRv/sylhSRV++maSrFpLRQff1ja2nbXX
ufSeR7lLD9W5Q/E+gb0S7KTbrT1tcU7iXwlJx07wfyY2Bb4dAaXK0RxypGMtnW66PDNCeH6lwNJH
3NYlXrDMkVonOwYA6tzzIIY6vDKzkqf7HKVxsNF0vMzl3Jx+dQdsrUjTXGybFiVEeW2QkyD+0aHq
A+2T+d7+MZYY+CntTa1az7E+EZMZ3W2o+f7OwzsmhaFF3yMx3Iwj3xQWN18DvrkVMZ9UZED4tJRM
rnlJoEldDPZZhe1y+ZOhZZV0u98BQc0wCyxT1ZffmjUqAEwA96xoU+kWs683mam/M3LYc/unVR8m
Deirc8fXpNT8gMad+uOJEFQZ0UgVyTStFBV86IiJLVV9dQcUo6mX6Y6ep9L+eSJ2PEjtg01+z5Oa
gGlK4zkQ0Jg5OnZiIh0a/h514o36ORum8M6/5Ayt1ptKPnm7IdOcvGKn+T1P7kubAr6/UYGn31XW
X+Ls7Jf9LxlcACuaGdQSlA9lYoOZonqjVp/gcqtUTFRNrC/brXVB7qRpObjMs8Hk2vMLUqMzLHlU
hiPQhy0iNhdqEfgS5xS0PY/BM91f9AjtNsa48BG6cUX6/5x8KlEDgKkaCRp8o3/3L3RlooYcid0B
SK3GoceKeI4zbW2iTCjtFJKK3TVzLpAGwdKdwW3XMtD/w1CE9fI9n/TQn4rTU+TCVXHJQCxAcgLW
xkd3Gf2hvAkbNUOim9bKtV3PSBu1dX6UnDNLiRDWWQEB9iJSt1QsGm0asrVjOjZpd+QoVLbfeP5W
hpD/2v53ZT+egMHCOdeB1TRZB0/qTVCwZQgVY8KXBtlnHrnzAmqjCoska4+6F3lH5WfoCeQ8T7+z
RdWXQhMUMqGHdQSj6wYeEogPV7ikN/maTOzvwXhVUBEhHL1ebhTQEoyeZG1bV1vxHVMz6VrqPkwK
hgzCiQmoxkDw3VZQkhxjxbCullAg78yHGtRxK11fjM93RTNjSYT4IFL2fovLlHy7CNkCWOmF9X+D
+66WDHU4aJR+L/awoeL9naGSbp2ZjVQ3sk9992j/xkM6/0ijLsTTYP2SZUc2by1sm/MiYMnkbI9j
GXfIHAfio4xX1B9ut9K/ZABcFat+Kq7A3PK8i19RckhkdzTjrPw5dNv5iEGzg+g9NG8zLZPjcO3h
AZHmxdZt+V+swnUWJqQU1Hlie5kr/5dwHMq7GOY0rV7Q1HOX+PlZU5y02sFm9f8Xk8Vm5mdhKWPp
+oZO1iEFftJbdQbxgfZU3wW2VxtshiRzsXUXkz6LlqxYN6rJIB3Z4O/3MS0o/YTeKIJ0jy5MORsJ
OBBMDYhKOFseOPL/CA4NO0Z/jer3JS/fHCzinmkQZpCHTAmnFn0xsUT7Ir7z11eVREXL9bnr3LZs
Bso5HhFDMJvO8nQKy7Qe4Od0ltAsnoCxJPvjYxDhPDWRHzu4Dpa47l10fyTm3DJ0R6Za1EDntITt
OB6Kt5mjQMwgZDmXqOph6lv5cEmE2iA669UjGKMm0s9awBK7CknF5ZhKHPrikGO5Hy1SB7FNmhcw
JwCezUzBBMIcC1i6Fz3Fx0yJFtaxZ9d7Evr5Rsmv82b5R9xfswU1LETc1fAMzuDuUZJo+JOncDJO
bSqCORJ8fz2w1QuFQHrqONNbg7NsEQP8Blv5o2oI8Jmh69tYpjz1SvX5TqmY1XkIAQOfQJ2XW0NS
sBVLqXEVPeOHBcISRoJaBgfDCiYOmbyEv7jBPJuV+NqWopFWzMXfPJq7g8na1Eao+TMNQIoLmCPc
PqcO8HHHqxeWWRQElSECaUdAu1FgQbPG2SAcC/VLgoupj5aeG/FpqohQo0Az+qF3hqdZJkXb+uex
Z6L4kkFZdt28e6jCyKrg0KWFSTlORjbmhaidvDjMIgXuap9WcxNUAT6kObkrHUm2s4O0s1N+kQSE
Y6sqwN0jpo9MrxU40UdZ9xgVbDnHRfFdEHpgC6YL4HO9AIgIlcbTqbC/S4vokeTyEWgAuEGnzXXd
J9WcSoG2AL5Sj08GmPC2C5SqXNYcE4e2fsozLXWcTQVxwG1Rx7O2nktkjD1Do82cdmGHwMRJ1U0x
pvS0tWfrrJwNsHO/h1llhY5rXvImgVtzWXB0U03olfzXZawZPb/RKyC1B7ap2bru9tww2+RIOVz2
GvgfJKCytcI1r+SnuLKJ7+OBIcMeHNmKIt2ZirznOtqi4o49kXa1805mYaRydmWNKrO1wIaFMFai
rjSchrtOmar9c4Bn+sSXeIQynYddxfMKBLTzx0ZI4NS8Hnjc09AskQBDbZg95zM3TqEZr8oH/12K
3XqMJMjCC04r56MHoKDHUAAq6SLgkLTbFWcAd1UjwF/GU+NSp9MFasF0pOLU/2k70mF9tTk76YLO
wPpsjaMlxy4V60nDHW60IpfZwRAVjbUUF3ZODBhKJ0y8f1l2G98Yreg/dF4/3ryx3tC6qMaMoL54
A1VxuD4pok7fWNjxW7AzsSl/JcGEZqOXKI+JlBrp+bGwpFl1eh9vLOUNY5aTGRM1/fTWND+XCyUs
7mhKajw0iSWNGZXS0l+6AKBCg7EQTjVzBNr0sKt8mulzBbTc5By9tIzwYrEc4KbAnlGKQZUkC0PM
L+4rL1YBqLXWIwRKRGwCMf8gY2zv3gVxsDC/8ozTHeKammlKh/0bcXih89eG+II0n9u2HJnrXRTS
ttk3u08DuwvjJZKBc69XRLNSkVEGuzwo+OFoVkEDC5w4buhOcnOlut2NpnU+oGEfsKQE8Y9xVR2N
IQqFqW322CxMJ6En8UWMsu5lMiCLVQ90Eh3OjDTo7km832foQcXZboi2jvYbNg9f47l+K71kGYr6
YGuKK5MOBgTqMMz3YyBfqFSY5EDyfu6PVqqYqWOKLk8FDJCasLyqrtmHWXoZGk/qZ1NHxjJ1tRvo
sHZSeDLI5jXKCPh1zE4qXn1L6GrZlocfbILEVfARGI0KhHsLkT3nh7WWHpy61JkODk9GzJGZbJse
7nhsUfl7l6mdN8cy/vml5PhA+NVmeRaKRSLVG6/UO6YzS0p6dhyJmybTiCZbKLXPrW7rOeY2vVOa
4HpnD2RpmbVGgluijKv3JsNt7qzNE9lvcC+PYaY4ScwkunaFtjs2qlGuGYbZVkYSGwxa9QXuJkmb
Xeu7k+xpI8zZZYtu53/MWu2Q9IgbhmQUnkHTqa2RXjv8NvDI85MbYY/kKnooGjfc5zh7gDfoU+9E
7Qeb539bBIKsrlDvQmtSM/Oyev6Ll7acTQd/zuo8PTeS6mYNxN4nxrt4iBytJr5zGrTiQgqcI56X
F70DzHVTXcxQRO26EzWbb0hDgwLQxWZppwm4loa4rxJ4k/J83s1UqT1FT4uya9sMyuDkOVqQBPO3
o17GD0BGjaLyyXa4cxZkhfgNA7lURGZ5ARJNPmTiwOE/r6rRN9QqFPYC6xFxCrvYluBnaVOV4kBx
3txHxgJHR/nmpE7qPIC8SUC+ErTsvHBACu6ZiI7Np6j3IIma/jzvuCdcZGG+M7zZkhLEPbpehC8g
Xk41HEdUIFK/3MHQYCjc93iK4yExR7nhHm2vV2Y+tOFO713UCtZk1V0meeFrQB+D8pF4iQL63AoH
PtdaMnp91sMBboLxdMrnS7RhopoOV81xDfsa4LA/uTPSs7S+cwhWWyD4PbguRpyYDyuPiah5l4fM
XcdsrozADxCRRFMT0nh+jePNfDYv3da0bw/jFDN4iRT9wMy0Tr/pm8yV/eIs181A1BV4nj/K4QyH
7+fYkOWBj9G3LGRIioETqIRA05TXMD0qmQdgVL56aihIwmY8eifmHcVw50Fn3deJOA+Iqsmqg0Lw
CPg3BODJA1y+s1mvkssbfxUhx2wfQp7ucEMemJHLHaIdaifn7X9O6rA7Aufvly6DiekN1+Saeat2
I6yfRjdb1p48qxL+zCHzTj3qmpooprxlQXKGMVaPQnQqACHptJEIzifgP2QeBqSCZrWOVF/vIBnS
78VK3+/oaJhyi/NZuViu+QKRAsecu7ffYplozI93zcTxjdqx2MYdahDUFvbbogyNmIClefApPRD6
z1XOmg0Ep+IHCTQoaORHNSJOxdLOisaf+1rXzyoETA4ryoGSK4Cbopi8Mllfby8pXB5Hs9GuGtWz
7cTDXDkd4WE9VkunmeHMNyM6dZhe2h3b3xFeNpDBqAF4AmsrvNqs5DOXZELbnKqxhX6cO9sHl21s
fvFhDA+bR9lKIOmoCaum41sZPISnhoZmv87ADU27jNZHiZKyVMC769tRBPJ7PKE6x+PXSEF+br1O
/sQpNmziyfIEeFZb68U2SscNslUyXP/rI4yElqFVZiHL7cqRWAfzZvBwABnrwdjSgveJ8nOetabr
LmiQ3jGdaYyZqJUNESpN6eMK8GpTb1zfZCLFcdspDkeedimNo72acOpkBed0Ht3GqeojLPyI76+v
Zg+HXpBF3aDLyG+Ycpdtc1psrRXeFoqsIY4mwqEyAsl9o2FoNcZaydxxOBLhKZ4dQJLU6cHKvA7d
ihkZ4v2uzNWjSfXQBjNXPavWEAslo1Cz9DjqMkV8rAYC19dcz2NLMQNn7F438NkrINV28qk6Fi1Y
4hQBfi8sW+yexvpDR6diDPA5dvwFnO8voHLFcyd/dwEIxcH+9b/S7tC2cOsXKxYNYeADNGzOGtqB
aR3U2jyqbsvgvGRt+Kr93YFaO/P8Mx5nl5VVFHzDPQNm3uFi1RNpp4r/81QI7AzHpxeONzzjsJvk
gIj6QYyprmlfW2H0hvwzgLKhl9QNOQNl1MNqZGHTFE7Fk327k27NG80EDeRttdMkCg1lewMwgvk4
+DPG6+mjzQYf/ju/ZNDmyllV6t/08qShwrPpKCAp7Nxk7PTL2kUYcxJWDmKOCqJivjpEhRVNi0R5
BcK/dUi6x3cMmOj64a4hjRwua6IfXydJxO5rb01fXH5j7Exp07l6s/AnYhNduboHpF5/7BM32BKW
D1V/eneuvXHFdRx7pNPa53xkknAmh/b6iDx6JDXIowBiIQWXddpOcXCjn5K3y4omUQ/QU0bpWK7+
c150qlenPhI6db32GpXj5RUVYCA5kylC9EpaPUZtQV2S7L5MeuF4Hnzg27Hfluljzv1sGyZp5OEb
RLLVvSMtyHN6dDkaZaRICA5cVXCS3Jyl2zo4zjDcy/uhdPIUUmEkq1Gkc/1zVm4OJj+dG15FCsnR
+JOh20SXD6AvLZphteDXREN59xJKVy4NkVMGc+qcXjAnUyErsaQx421cNTgY9I0y4K0neeqBGKYy
+9E0hwdau9lPpDcixyWPSuCPb8pkZvqK1bkZRaqkVMQJUMutbtTy3QoRYE6aU81bCZM34JeBfOMA
gIceKslz1oFxvvFj1/B6wb4wcm/kvnDVOyrvnp502YWU/m3UeWnetRbpB/osBF7YwbesZeOXGUdt
t4ZVegdwhJ+nwfq0uKy1QmNHAgBL0w9aVBWEqiwgAmsMxK5U5Jl3gs7m/C+2GL21nJyzalopQiJi
Ad5wAbr198lk7HFxz3ZsF6icVvw5I54VpR7E9yNjgAId1TYslCPe2WnE51DTWG5g3pDueSXKu23d
XjO1NoyMGN6XzN2APT3PeuRC3SUeXElNCly5N3N0xNVb7UqrbUMNErrSQ3nLIXQJRdGnc3UODqQV
gjKFPfsiVkfyn0aKbgn2B0YyorGM/oOzCRArXa561EmHGFCneCrhrMNMLNlzo4RtWgAUHM1QK5/t
j87tK9AjDaSlCHwsawRS3vMAfll+YcXTQwICLyODzEJ1cSqFgAzSmdP03zdSMH3TFwL2KNGeBSkf
O8yhY9yXDVskIh1BekYbGQHhiXjzJ4/QmwJOjoOaYAGl4BRhJbzGJ8H/orOW4c853mBMXM5WfxZ4
VuZ0EC70BdcqKHAGRuN+2nhAPnV7rKdcwAr6XQ6+nW0wgWZpqcsolwdX15sKBjyMrot5YlFB1cVr
Z14Hm16WutUpQkWf64Px3aSum+8VAgRCZJQANTSCh7LmpX9mAumw6+VBawuJOJkox0aESVWNefrV
sBLsUTthpicpJjNpURXk+ly+fqsRPwhR+enGk2IlG6dPlgRWgTzZPECOTeo86qeYwwfIgfi/4Soj
yK9PrHTBvwrYIP0zAKhol3PxwthAI9uhiZ1/+s+e81Ahe1gU2kGGT2FKyJkNTWdqGoVV5N4fmkL5
kxoDag8MiCRCIaGQaxT6X6HlWfA9bpZC+vlE6EJkGDnZpayRRnA/ToUjHF62BfeUSJ+o2NZwbi8c
+IbQQITt+UBwcNC6GCpMQVjnxB3XVcEjKlboxj5lhTPwXJbMb505uJRTf231ho2gbveVOCJXI4eD
pfVRJywshOL1JiNDITOOnygZx85m4CXwHmG6GGJ0SQFNNrxZIpisopI26KK19YB5+x3NjHYQtpGE
XyfVPPUDzmbZRGDuHLZkBiSzc9alC/KCbWp6Q+cYq7/YyYVFcSm9bz6bFK0PrwPnX3R9b7ZlgS4P
MlIecX+1tUMN8e/0mkNDbgDvGOvji7hZtpF4OhwG2Jh1rCd2xTatK7vV9qRg3GviF55f+129P/t6
VbZq1TTMw7AESSQuqBTHwEb5EVkc74IK7EK+BJzFUKQ74AO/uSzpggaLESVJgPg7dqUR/4uBAnMc
9rNTsJyjqu1fKbmc46hTMyOVft3o42fkRDwFN+8Dfjrr0lsr7W8ZFZrb3jd2NxaFvhp2wb44U0iD
z51yTieaRRUx9olYAyhM+9SLKaUoTu8JP2ORI7pLcz6J5pOO6k+kHp7VplkIrx8e5A5KteffQzBJ
y62PBoLPFM52sYt36vGfo3OAh3j4wY0A8nzi5Bg3ogG9/E6Ez16mokxgqu94ytlamPbBAbzYr7YP
dTnKTnQn9u6HqfK2SXUWfx8tQcLNKQ/p+9VVve/QzvUpFdMdJl8KM94wlzstAX6NF0ULceDLjOBb
ipBOWpwMMhV0DSis+Q/dBrDhj1KJhsfmTGY3UZlw2GoVLHHK4FItwqrSOLZr+0mOF3Y0BElipA5x
gq1NOxtySivPycsAwCMESh67oXN+aNhOtpoqGtrwKCJSYpw/4aCdcT8TfnxO7Dm99aGWFSgemBRX
X2mND+ufFZvPd+EfEjxQGvZJdwgaSu9iTbxX7UrA1+sEaBLTQEO3rHOdXOXo1atj4whog/6WXeP5
uYRG+7VRYYRYhzTcnsphBTOCTC7lUDrvy3NkLl/gPwXVoNJ7GuNM7aBEf/MZoWA8K1GvrgiKo1fk
mhUwi5GlAE030kYXYq6/UL0Bxs+L12+rrq3wQLfJu21U1GO/McSzO6FakpzjaV8wLGlWLCmaMwg3
Lnpw/BrvdACDJkTnDVtYAJPb0NsGDRK6/kxXbR1iIqD/BFopOE9I1LYDhoHEQ+5VlqezG0MGEx6v
x/vD5I5tHG1QXYj2PTRqwOmpRqG9lJzioMQF+y7GcKKS+3Z9DQWEErHfh5xNa+zFTvCIEsmF67Xc
ITM1Gi+rW98UHT6jK5qkytDHGiug2fpikBW9BfuboprIcOjWzEq2xclGq65aPbmjI+QTgPBF+pJ9
z7L/PAcFCia/E46/ivOz4y9hA+YxxUVbf8O1XsArG9VEjrGMlpjyOZtGj0dkqyKoxcejJqFoXnNT
pNCO6D9uzbiN7atgfNdOY0+W0NFwt++rRb8S710s2Iw1TzVY3DQefr7EFf4M66pSgYNVG/4111vs
L6wbyfTddcsqOym4eFQoCc+RfRAFXVvcCMJMkgHWQy7zAatfk7OoWwgXZloBVx/djqjmtZYElZ5O
WqNEvS6eGd4BWT5PHFt3aRGI/LAJDm71wKSqzJPYQeiyM1cw7zVof9XeDgJAPJBLRVuXPo6ZBgOT
Ays2J9eCKishIDvl+jOh2KW/7oEjKHFER9WXiZbGv4m41bHomaAfxNtv4N8VXvvrNTkXOcYC2IlX
IQVz+dIx32dglKaeS/5SRqcLrryQ8DmMP3BQhzw1SSOFGPOsZHVVJcvN19ljZJ+kQ2cKqek89f8d
PUWmwQbvJCb5OHJj1y0xi0we3u3bHO+QwI0okEBOzPkIyT8ekj7QEYF7grT+luzn8AOv8OPKUNIf
eNSVIGnhCQFd9T+UCGIuOcFgPW64hnNc0ES8RBBATluDax9xrijuPO6n0eGjfk6Dk0hWPQSdNY07
CGNZ37u2pl7okR1wzQkj2/YpLA+B3/RXrJNChYy1g3V1RqwMyaw2tPZt9lhGGwFHYgoyCz/+kw6J
lhUWoHI/VGtfO6NYxib6XqYGjSbbNdr6VAGu5YWbeYA+tbLdffT9uttqSDzmlB3VhANcJ9H6M5as
oL5HOj+CZ+5arc0TkL76ZbJGnqH2M+bC5hYE6rcW8XMyw+PIAtSgXs1CQ9rHJZ7Olx1TqMtmTBdh
2LLh7/hnFI7HfqloT4jz/yI+sO7oQaP+5EuzMzdQg0ML3MViQ2Yk6TbM8CgcMy/bUbJ+hPJ3q/Ry
p7M/VHVK1+bNMkzs0mJYGtSYa8OW7z3Cvn3MXRVTiFK9DjkJfhK/uNxZzOC3BJN296VBQfnHkpIl
x0x9b3Y/cUMlUghTVFBOkzY9TAPZWibC+eRTmViapPagNsCv8AbZ+X1cR/gES2+uDQX4MHUX22GO
Uzk9i8CD/R4RalKz8ymSopH7Ow7n4ybJgJ8c5APNeDRPpCKQz/MXLQcBnHtBxjWJH/mjM7eD/aeX
zPBDYz/lZL7VMzN4Tb8tX+6xY5f66eiidUfnko2HAWtiixtFiDDgyVY4EqYP/OcfHH2KrzEW9n59
Y8jvZhyrthZvuXgKb8o7FloTfBCkOQNYSNns0sNqKiznbM0r2n7sAjTghM4TRfBVLSyejJD0UN+L
Ce8sZ+arXSWYRQuWh/2KKOsWfPVzJ7QT4lfn4S7BFQ+UfN9t4iMagn3n4/thKfsWbg43r9hvnGbU
gxeB1/6yMKHwJOBMsBJC81W6GHMcRgVQpCZtdUzls9YuKRNf4TACIDPuL8HhUIZNqj8kYI1yCgMA
ob+VLXAXPIkdyzdDOYyoex4lIOWam46LGByjscGuLhkMWnO2gqRmwLr/A5lUB5J8JaWyKbv6dWtE
n3xRxTIFkP7XONXIWquQietE4W0OKj9nCjuSozddtdBbzCE356oKon+pQb8ayYJA48UX+DdFxyRK
0bhWAY+v2oD88oAewhc9O0GaJDc98LgrVb0bMiKUqvJp/yFc37U0xz31AgExAuImRGbyxGCcv5oj
2ESD1rC4770KdBvZrAxsztACJHvS9qwpXey4UpZrZAJdHEvyMa0D0z1hea/SQZ9e4dLmNQNK8xGr
BwbWAE5ccCOvIWnn1VBDPP23KGw22j6jNhrN1kzZLbKoT2Ng6Il1SKZhgnYJch1Y2vYQWd7akkVr
KTMRaGNH4zXKEtdb/g8dYPYFNbExfyw0I7Ndy31eOKGdOyXKzvS38dVSY+L/M/Aq4XNrrkIrATAy
O61mIsc3saOW95PnZcxO93c/Eb+6LcQTmavE3xQB1+WbTUk1jIRjA7t6LVVMxh6s+mTBEAYj+Zlh
9VCtlkF7qlaGEmVr90I3cmsIFx/slbXovKcRGIKb6TxP5gHExXM7A6vfRGv8Dn55TsOPcBXglb8g
sr3Fxn9GSZkuxbCN3JXAkep0BLyLBpNRheeft6LuZZ9rqa0IKjLF1XM/y7RdrrDue8L5BkyKyVOR
yUQ2fgyurytDDoM611E11PKVejUnyS4VFSMFHJgABC+aD7ozPetDkj3HJOjfCFJcItNacbSXAXCD
1ARei6y3GBYh2CiTVW7tBWx9nXMbQ4RWSxHWbQwb0vS1nBfaq6nT+XQLeRB2W252q4ktqjot+Wj0
N5a9XMb08IX/Nl/C0/ltUc/lU86pCPhEmySVl7sHe8Iy0NfX9oY/cwIZPP9Midmuny6aLO292yjM
t3BF7sjDIlQ+MGAu/vB0VVtVFYcbNzjylHj00qbOKvx3V6DEMG2iZRsCjZJdihNMqegbP3p39a6p
S+iyX02xQFdpD+wdy2xVV5zw4n1/bKHEe+ZeYUYOMWDXsOH/JARYH9vlMO66RLrRD0QwGsKxGXCV
95gjsB1TPWzC8duwxidoF6oBxbjAOyGPKR6492aD4P1jcgLBhq0v598Cbb3S/kDDg3NrRJOY7tM9
x1MtwT8Ti7EpNmb72w9qz/wOPjXxVX0soe4b36RA8OtpMHffeq/gP004b4Ups2bfcWvhmi2vzuQp
K03RA2YWTbU2x+IcFt2a89XLb3hWqyTUmgTUSMS/ombY/nbuzL+OrjXQ6KvE9Mo0gOcfqDeYi94G
HKi5oKrYpmkoqxwHlooECsjvSup5uA6rIyhp3twfnl+1LqnwcCLNyyhrehcaXhnAXAYMWcoutHGp
IjwQiO8wW7MJyV4HgUx64XOLKd3VVjDINIBbzO8NaBdMVFSkeL4b3lkIWxBnzk1M6qDW9GNYWyhb
aUJosHDZGgq+H7tZHGpSxrDomsTlZ124R0lET/c/9gMzf6fYbohYXDX/qRYhpgBCaj9hsstp8tvl
ESnk5zJvdO4XzfJ1jhbo3o/2Q17ir/2IdtCnQpAnrPvb5+LjSPrSUhXq9V8IHPZYNVx2gHOPD+Mf
bqpwZES41aISFb7aH47EgpaK9N+aAb5ytA6yf/loAusYfC/yonLzn5frL5ChU6ZWPFNMAOj9fhue
Kqxp2gyCeOD5OUJOfu5jgknBBcbeV3C1c6kICoVcvEcqYA+/jBZZBoi4Dyc89yaS8gSNIzwCgq6P
wtZlxcno4dVqjNqCmDS5blq6C1KleDfhfDaPPHqNSdYTtEXoBmqt2Eze6VODRUUk7T8y2FEgVxb8
mnhhedGg5ZeYVvYq707A1DbSBnhU34ljLzFojtJss3vvYIsWMlw152ZFZJFdFRdNmRDk2p7OSqqt
Kw8MoKy7mhifnDga6kebtM2yPd2A2W1HxoNq7Izg693UgSW8OTfO5DnqltpkGdNptSEeAsqhJJMd
gBKAmS0QOOhUu1JdTBqk8mVliRp+v2wHwtGYHnsA6KMl1zteWPxKQ4/IuxY8lK9zLKw1QL/F+2xP
c92+cSttYQfl/kruS+q2Qo1+sfiHJv85+ryBoYcgGx84xK9cI1XRL+/bQZwOsE2ZcZjf6dmJdGTE
cGdBKOhHIdBtD/qSzKwJU6Eve/PUBYtxg68xuMP7FlPo2H5C5oZubT5xVi6nZ9cAY34JexdWymLF
DKFUq7K1/0OpEtSytfN5eWgsa8zhyFyOlViKqgIc4eL2UtH6aQLftJvKb4HM5axxSTUUfLTaQrbx
Ol71EG4WIpecYo0d08WDwijV4HlsjtCqkBvCAgDh3zCK2VntBs17hzs6WETFtSorSs8QTcnbdK9L
lFTlMUT6hvw0metUm0DwkqsnU6jhLTGMuKQN+//hhjHoVnLbG/sLGyA4ovJF+TeTgdxHmJin1yKv
lNs6/T6xu7oZjkrvzzs+YGYEOQOo5C9dcPNs8fXVp8D+DSBLfNjeiAhWGbHKbe9E9vTepvmfojYs
Xk0NupmPJwAbAMTli/MiKZFNVDAh6fivMbSvHkEF8n2yx98N6BrUfiWB1CBxjbg0Qx9MqhYVGd9O
chHXTFmEvDlzz4mDBXDGLDb/irWf6yGtNqC3FxvEmK8UaCMC7KC3Zn/XzeanXgk5XPOKEjR31g2E
CcO+C04BxjGsu62fzVxyzEOYTn3j5vaBBltLoMo/VqGi+AsEDXJHMWKevN5cxlM6DnDgDT4jYAfo
JffFvHaAJNDgwPqgWXfEOM6taEPfYbrLa1DC1TWFeuHsSModB/qaIY4NvFSMrT7cDvPf0LVUo5mA
UoPHlhQOYRhZsW/YFLbjzyptCSDSjbwysvQ9ooKtgx4fiWwzFM9dXq34tJNHQfU6MekD90LC1P1Y
QkPAKAJWmJVIGObyfbPjYERswjOA5ItM3M/+uhV5NV3A14rPhB+sIaab/Hq3gGBrCMWJKCieD/uX
xvbnwm11kVFVSFVyMIvll0rs1ZxPufKmHESsyRLxl8Yu6DDXCGUiNxe31CysDfLgBm5FYCfg5EJZ
vAx0IVuNADWrEQNID90R4pRfWMfemAqTWRU47d3AeAxmwQDFBQuXepSvxsLyKR4IOampZ2GLUBGs
JMuAg86/AFkq1/qqAh9xrJG6/eycTS6JIrno5HwttvE5MquFcijw4zYxei6KZrTIxmiXpa2ZPfDs
HIpAt3O6A4+oarhTVIk/djWcbGLcNf4gmJSAEsLiQe1c1iI4xUGqk2IHtWVcOGc7Yyksq5dXf9U4
AmEfKyNhjlP4L4F8o7/2H/fZKGZ1x1WEev/u9CNTcUyGWVWz4N/BsnPX8sWebHGiMi5qqJi3THiT
152Ute0qHixrCpLqKaIHXX86YZNopXYotwv4KIOiR0NF20gG/MsXsfc/gpLMgNRUMinB4cKrDwFu
4Fs8wZUeqNDuG6orBIs/TZyoetirqkYuluMb9N0QByFPI1mU9Om5Mti1OZpxZEIvVd2D7Rg2wtLQ
PtFTO1PyHXJFjPaGvdAb6G6i9KgMatjBRmlgOzC5fcUYfP8/xPqIMKk2ZvLXNgslCBKqsFmpCRA4
88FKBSX4J7SOSXFmm49uGWPrJqn8Rpfs3+0QylkZStz3QmOrT/2NgnYGRjXYsKfxU5VcvHr+ASEU
AqKOC5GwwQwcLQJoDKCBQwFM9UZtedeMfudR0pwWZGajW2MoRoGI1vcUaJPq0HptKYHmW3KE/CAK
YI7R06gVArHPN4Wk627IAXliRdbalXePWiEdfQ8sEZz/0TdRTzIU3K4T1L6Ax1dFjWtXfo+ssGv7
rvkhwW+rDG1ikPpSu3K0hurE13CKldC4GjTlhQex0UmCH+uLswqpedEjxLA3Ux2sWL9CiZ/xMk9s
UmYcLUJ7MLCb0VL9o7Otxo6NAEtEWfGZlSAFCBY+3QP19mFZx6U5CP39QHIc5Imh55iPcVLlfxuB
k1g4m77O/SOQ9tmVFyaAInLRgWR2GzDsFT3kZPdmu3x28u6C7w3TIDUCtABIvqcimN5S1Pa3lzCL
jA2iT5XizbdEOGB8aicFmOBp7y/nSL+kOJ2xQP3CztqN+XLLgw==
`protect end_protected
