XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���_���0"T�δ��4!���RW�����݊��9g��a�+���k!����&?��:�\���ת�i�i9�ڭ���uJ�cY�.�,}���D~K� j����A�_B)ڻ^�H����_яq0�3;7UZÛs"�V�(��Ϩ�<v_`C��ٓbI��LuT���!���9 ��ۛl��ڢ�h�Mi�P�ѭ���ʸC�go+x3��'rK��fGgX3�bo�U~�qe,m���o��L�u�v �p��R�!�s�*��orc��M��jΈ����u�#�	��`pI���x��QBKӘrޣ������BnA.ƅ�Ƴ��߿�f���YL�J���3/.0�/��hK����a��J�f>^��!{����(�e�6���y�D�`��8q=�_P�M�@���~��}�S������*"�=�9	�8�eC6��/�hCQ(�|,|>a�Z_�����Px $üp����h$�Xs�?PK�C��|Ŋ�a"��3:�$��'�P��x��M�_�3Z7�4�����',�Y)*���$����2Iaw�����v7@i֨�`x�E�"�Q���D�G]��W}��_# Gߎm�M,Kk.���
F����X߽
��0������"i/EΤjv6Pby�%\��A��jv�m2���X8ZSq�s��^!����:i�n�D~��AN��05�Y��p��G�d�Ъ�w٩�S�,�A@�l+�����+��t����3Nj���XlxVHYEB     400     1f0� �;� W,�ҏ60L��Б�Ec��m<��p�
��ϸ~)]�'
�y��\��Ҥ ~vHF���qv� ���T��F�p:��9�)�Z��+K<�X0��4�V���/��N���:�C��ĩ� B3�lʪ�qG!���KD��)�{� �_�S�)]�����9<�Р9�ohK8G`�����f!2,�h�Ff����S���0}l���:G?O0cEa�֒��3`Os3۫�O�0İE��h�Ds��g
#��8c?�XM��1^�:E��|�p���4t:�_� ��X�����e!��h��y�1:�F⊴�x���T~��N7����aA��-M�-����ԕ)�~����ǐ� g<kQ����ѽ�E�s����S\������q�k0R=YGB;���+�J�q��n~UU��D�a'��i�_^kx�mF��?�����͢��{v�RF�����o0�m����^����qQȗT~�R�XlxVHYEB     400     130�.T�k�Ie_�~�~H>�4R )��.�����~	}�M��2�ːX�36��4n��y�����z��!�5̄�Wa8��H�y���HksϿ�%�z���p��Y-7�N/�|ES�z6l	�8�������M}]V�^�P�B�%�T�,K�̡�Ujet=$��Η�ݴ�4LrWB�=�'�p�V�-���Iϱ�GnX8�X]v/���1yĺ�Y%���#@I��1TwX�l��;;ܓ/$�j�$�ld�(C�rU/���������W�lv��"�'�r�h$΢�Ob/\2�umggUJ��ZXlxVHYEB     400     120x*�I�
tg�X+�,��*�:O�;'4�؋�aM�EJ��M��v�Rލ7[dI�rvC�ʖ@Lm�L�ud`��j�|���]>��d���]�Q��W� �+��f�S�� u���5
G��s��
m덺z>����it�z��UJ]��m��A����~OOF67�$,�W*D�(�	uf��\j���+�%9!��n�|���#6���9��HU�݅�>NU�Q/1aEK2�^���^ľ�����!^k�D*Ĉ[�E_r�'O�?2�M��XlxVHYEB     400     130:���彃�f�����"�%(l���ڎ�'e�䞐����;�C���s
�B��c]wz�D 0B�jMI3f"`ĩd}MZp-0+��]�qZ��m��=F+,�1���%����֌��+�3�S��H�jA#cfz��ݫ�S��<�n�G6�g�R��`4�g+#T���������r�G�8�L� ����#��$
�:WF�a�*��ʄ�9�h��2�}��&�����5�Ӳ�� ��xmh`ݧ=9��@X�y��s�羱-�@�_\����u@g�SRy��=P����%}��bXlxVHYEB     400     140� �<�'p��;u��!/�\&��� �~�G��}%�)m���/o��Eǵ q��~4�"M`��Cdf����ۿ�A�n�ڸ��.N�k�UfK@j�c��<Z	8۠�4�<���/��Q���x^���J����)�ђP��l����2L4�C��O;q�@KE�0��(��#�����S���8��n4#�u�cwQ2me��~b�(s	��8�*�ʚ���_#��*�v����ջ�|Tj��ҽEܣF=5�h�Q��	W<�n!_��AK�&� �c/�Y����z��
���s���+a8K�,�T�Z��z*XlxVHYEB     400     180��A��>�
6�/�GH�T��vg�[�7�a�z�`���>P�?�}v9@����O����r<'��w��t*�����.��sߨ"ڨ�\��<Q;��ۍ8c �[K<�~Q�^��gy�0-_��.�)�
H�8GO?��#���pC��\�¾�➅�m:���qיψti習���y�$�+��_�?@�={��kDT�t�XL�����0��S���|�b������xԈ��`����s`C�����i���1�JPH�1���PE�����I죇�?���_�����[Vl�O�R!.ݭE��$4v-���,���{ab��}�2wj;T��g��Y�����J���{�S0��XlxVHYEB     400      f0��=�N~Ú�&���6� z���D�B�Ss=h�/)}?VD���x�Ö�d^!^�s�����,_P��#�XgBL�B�#Dj�r�~ӹV2��M%ɣt�lzD��N����V��g�(~��n�g`��%�j�oK?���`T(}�S�p�����魌Oi�Mxő�Y-gYW���xy����lf���w�٤�6��zbʭi�"`�
.�������6b�a1��H�u� �7XlxVHYEB     400     150KA�&���B��}*�$B�"����������x�a(�i���bC%�{�W�"��c�9ӮX1ɡ����-o2�6}�.1σ�a��p��(�3�vqMC�	f5�Bx��`��j<e����h�L���>ߛ�7��5I�fᶜ`h��d!�]�<U�6�M�w�hA����{�^�syu��~%��c�Ά�S��D�׺J���Sڭ>���3Z���¼���[/�]Y�\rv�a�/
_p�ě{1v �bKƣry��!��d���"�;�ޏ�����FS��,�)o��s�=�����TK��F|��H )�p�l��"fr��"6b��Z	��).[~9�C�~& �XlxVHYEB      b5      70)sQOZ6�W�D��(b�-��w���g{P<Foc IL�	!&���{����_�i��j�g�~ �u���Ǌ��P�^�Ӑx�FE4[L���lT>����h�� �A&%r