��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���3�VL϶���<�o�h]m^�N\;Gm{��=Yu������[��J4#��&��_�t��̅o^
g>�E��I���1h}�6l����p��m��ba��]�L�TQ{'�7R�oU��D7�_��n~�~@)�7������^h���`{���駰�P��e,	An�7{R��碶u���BI1�+��~ޢ2&�
!�|���ǧ_*i	Are�Lj~ih&<��ٸGT�h�Ɠa|h�Tr�K�L��B�&�
���!�ax�4�DȒ�D�V ;QӫHb�d���,�k����v��?� �O���65�|��Ӄ����3� H�we��~~�l$��Ԓ�_�� '��/�m�����;F�ewb6�	��Ks�>���ޛ$�*$��}���4E@�]�c~��>�����6O���-�S/�̒�Dtx��h����.���Z��Ý�s�3 �`}�fQ��D�e[�`v��ߓ��сocD���5����u�.�hm?�
W�8w��JOhT��O�WN��xzk�{�zA�P5$�[&h��	�9 ֙\�tV�A�>�u�4�[�?W/��^g�v^$�����[��wU�U����ᓻƏ�P��U	�B��eBjQ�_�FKW��i���*�S�������W��
s1	&��"�ȍ����@��֮��\��'<�����!ⁱ-���(��Ixcɖ@訂F+&�]�sqCOm:W'[3"��}�Ў2����3��������7���/p��&��_k̀r#�@&P�2�"�U��3P)��n�.�d�?�1ɵ���/k�� Z���c�ɏM'�����e˧b6�]!h�C���r�+h���?�Y�x}L��Z̫_�%���	���R��*�ƞ��d��.�49�C�Ɍ���߾��y�+r�Q)S��CCA�����"�B�ֺ*�
 �h�1մs/R�t�?�ƧO��vZį�j'�1Ө���t�)_�ǰ�E)V~!��>^"g6w�j�����<NP������B��!�v;�
�3�i��ͧ0?ӄ�ꔑ/n5C�<�8q�"hөݭI1��t0�]E� Sn��M�pa[�;<".;5��}1k$E��o��/��RlQ
0��/��i��<�N��3���ns~��D�r�����X4?Qʆa�t��#:B<6d	Ϗ�.w��I�V��i�a	��J�G�|U(֭e���2�
�`ܼ�L�p���.�K�z��,�]�T�Ј�n�%I%��0еa��$�/;����;x�V�T�!��Q?O/��>4���w��V�d�q�6��! ���$}���!�	s���˅
�袶T���/�6^>�Z\ӯRp] �v�S�i�M\d����� u�PǭXKkBC4���}�6���l���\�!���5���/����Ćc٘���I�|�+;�ϓ�^g*��4��1BE����wĻ����1H�a�]8�Z���v���f���gLU�a��j/�O�
¦R��P|�?���n�r���.4�%bϨY��⁲yy�o��>%2�D9�^�0}�/���qgP3I^
�l`��Z�ݺ��Y-q��K�^�꩑�����	��z,�'����`������/�?	�F�	_-^H��!#S�Ȭ`c_fY�n�*��&}��v�-�L"��Y&N^i�������0V"`Q�RO�G���f�2],h���Q��o�I��34��kM9� V�l�*
jOǗ��C�l�弑7�H8�y�fXʴ�������z�4Cma�V���:�mu`��5#�#�_�0j��=��T��,V��#"k$3��lPo��`]�r;JE��suz��]ԇ��8>^WǼ.=P�4U����譄�~a��(9�w�ػ�oPSKF�WiA�`�7]UpU,j�NHj���=T�@׮��S�K������� �-,��[�θ9c����UjZ��c ���}j	�?�L�K_0@0�8,�WОB�l!U�ى�G~ПQ+.���X�i����E�O�РdT�����jn�&���K4�P�2(�n��g�R��O� �8�#�J,�G�#Ҥ����{7�%Zc$p����Q�GN��3@�����>���*��VJؤ18�8z!;�SRE9��+�z4�V΅{�J�������㧱������ݟh�p����BK������(����l��Y5+�Z�3/��4c_�L�����ǵV��H1�����t���ȭ��#�����!$��a�^�f�J��Y�qӱ��<3�@k���X��90I��˜A�x�"�*),�`����D�� �P1���H-yo�8��~vN��<�#���=��jSl ���WrmmƟ�[�8P~�B��/rB�5�������t���Vd�ӹ�GD��C�ڀ��� J��=�O�0���#U��=���T%���o��@��:�v�����t�H8A?\�Z�ZU|X}�y�R��!(�NR���N\]O�a]$���$���&(��tD�:���~���������}Ö���R�����&�f�]Ul���]�H{g�{����#&e��|	5>�Y��Uջ`�)2iE��!0�lq��	E��=��Z�2��
@�+��b��F��;��=�O	q�j҂ݸ�D����ch
r{�o͚�ap��V��^sפ�)���d���W����m��u�*E��.�(N�$n��^M`��ˠ�N8<+�<����7��W���ࠀ]�/z�W�Q#f�l/x<m���U7�BE��YA�H�����]N�u�z(�PT"���j���V�����T�Mh�[�x�9�j�X�/����h�k6��=�r׺9Jh��������j��x��"�Bҭ��\% ���	�{~���nA'�Ĳ�O�-ή}<�}���e����@�%���.�3r��""f��wv*�͉yVm]k��9���'����UТ]!��x�h��C��B�i��H���;���M���Ђ,}�8�����5TBR1�<ݪB����-֛��1����ۈ~�x�����h�S��[c��w֒x�P?Q�j���c(�8
b��3����