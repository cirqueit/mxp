XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Q�g�����:�;�q2;@7��K\L#I}	�ja��F9����D �5��,���6�F��A��?���߿�����QJ^m�D��l^,����0rDiǧ�b��K~�7OY��U�����=4��S�V����	o�gܾ��?)��ܽy&R�t� ��y�:���|I�CN	6
Z��M������	���KDs
n&��ay����ߠZ@�MӈG=���� ���.KQt����[)<2U�P��9��fD.1 ���\�@�>y��Cʿ�գl���vt�̚7�3�W̭21�i� o��3������p�s
/7���5-!��~_p�٦7ktG@�����M\��d��J��.��z%��̊�pz3���r��1�r�/rJ�Y6�q��;u�]$oi�˫)�\8�т�Lz*[�{�HdS����b&�O�辍�4=�eܠ]�hf���w���Q�gD�3�U%������s%;�jG�~��&�����uj����hsE��o�T ���7����8:}C9�R	��M�Äf"��b�-��cEc�r��Υq�3����[r�)*
�٩L��m��xj
���%@�����qH�:����*�d�P��.~�v�L2��~�(�?���Y�&��?cI�l���M�>��G��:JWQ2�D(hO�_?��#b�=Un5�?�N��{�w�O���^ؼv,A�ꇇ��U�ˮ�Ks��G
�J8XlxVHYEB     400     1c0!��ji�5t�;��h�hD�^�s4\���/_Kl���u�=�W�rS?��bױ���.�'�g���p���]�Oh�{i�7Kx8��	�I!���4�f�Z�g��k5���Z�LP*��k����^ *�q�y�DR1�v�Q��D&(��#�1ܱ�����mN6.�M�м�<S.�н�������O�zQ��RU˶,��J�!U�5I�T�G��x��m�df�!p;��`�$���=����ծ���~_�]��E���fqAy�o.Π@l�V;�V��N-�z��~�A�������U��!6�j� p�EyLr�d	��Az�܈���ø��?�(c(�H2�T=<���m�m��^ο<Y7)�I�&Zc!Ԑv?�c@=��A?���NL�PWC��w˖��w�X�b��'웥�f��Y���.�(N�XlxVHYEB     212      d0��3�P\��jS�3��
���XB@���F��^3f�ql4L�yl�"�d��;��Q>j3�$^CE�ɟ{4�c�l���P&G����E]����ym�r��z-�
W�?ۓ�JJ���y�S�M�x]Po��ezC�X�`���,��v��T9B�a��Ŷ�<X�2���	�'_ �� /�@�e���O({��w)��dW��U�Ծ��nZe