`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4176)
`protect data_block
+w2OqazPXQnR6COO6OQn4Mv5WKEzIs34cxoq5W8NG9IHxstkP//iAsADfZQ1DIUSfLMvjDptzDVu
R3o/ksoS92Xbw1en56N8oAmOxdmdoSQW7VGho14ezoZlIvxXFhhUNXpplKyHGOXLf+viKV/rspdK
n5t7JbJKLXwY3KS/bfXPCDRQAn8ZF90e1rY/YRTksj/3qbk2x48eMwkllo+lybKmXaIx1V9qYo1S
usa2CFI/KQLLHBA2jzY+rBEmBMe1k0k1zUzbLz2HlbKW/qiiLqwO07Nnoj1NjozuGg3ikxS0XqJ7
efBMvat/P5F3PzSp5gWD5sU2GeT/4VH09W/bEcGM+3Jrx0HQExGfzxd303bdxOf2sSm97lNLvl71
vLKG4NLOh0rXCkTmoXiLUHH38TbtXJzEfZVSADvDHe3hbypMdlW2YUURq3rv1qP89JZoJcmY5bU2
BeTI4tvxzmbsudG1tSxnTZIx3Vr7zsXOYPf5CKIcgorwu48EXQkOmeF+5nfgriDZ7jDYMV37ZwgJ
m+jTvayAGzha0KlaAbvBD2NnTzmj+D3IK3ql6d+rJ6t28c+4AcjAmFbxKMpI26T0DXm79EeFW7lS
qf+Or1pRVNbO1SSsykKVDXq4w5FE6urlAXs+niv+EZR+Cc46HhqOwN5J9VohKN88LpVw6Jw/Llwt
20R2Wxlg7HBozxailiO/qUezpDlyDddUd9zFrolxr1zMd2wwaTe0scykUJXzkTQtz8jKNRFbM5jY
NI39TxLhAR2uinrYZmmdoQqNCvp4eRJBlrLiKwxWoIy7fWI9xFvgf+0NZNzFDZrdlTJEeEm9v3Ai
8InSJjldjShhkoMppHUTCJ2UIlkHwH3LRSM7aCuYBlAS+ZnJQ7G120aEOBkEq7c42+JcT4Eoi5xE
DyA05NXWzwtrFSAZV4yu4/SVb1pcxA4xwC0Vc4XjmghCmkDUxpivzrPwJAiFrCS2GdSiA9XOZu+s
ewBOyNkMLQDMbYkfK3sESVuMFSR1nCFBnK+WvmK38r+zlY8zVsbVxO0Tnno4ddfQRTht8ucALbTC
t6NKqg+5eELOVkB6KGaMpazQLByogPER9mKTv2dm6vIbfW9yATVko1+xxePh/iFiJ4Fc69I7Chk+
dxkvRs7sZq0Y6tEWwExWXy6pRAgWRUAzg3CPHZ2ewoFccOwGJwLGhuoHxX13Sa1JVq5SqNcnQn/u
m6MbVGkYKISMqWgQsyJVE7l5xYDpvDylz9deY8gbzpXTLU1aBHlaE0NfWEjCk6SoB/rc5V2GbTdg
BTpPM7ZavhIWLY8YvctDqmZKa/mw/kp7ZcxOkVt7aFHxLWVoweqKaRQMcyUuc3+fNMtUpvKIZkD5
QnIwwHuuYVK7auGCm/X2mv+CyKhbd9ifmu4xi/TLIf77pM4irRudGUCKO32d4dQK0NQZ5C2xDMQs
kHC4jN5Ocpfb4etciQlAxEOY1drmw9pN+eknvcwSRHRS4qyXZVTAn6O+3qG9gexoEO2haXKEwNqD
MRsqF7lnf7zCkc5LL/UX7VPGhxkdR1WKeNa0LYFH+1Bs7uiV9zWSHsdJJwlBOlZmoLtWWj5nOzWc
i90PfYf1w7k01Bzba16NbmMfTYdsHG6IlNXV6FfTEVIlOXN/9Hvw7eoz1hkLJ6HQ2JRb+7hoYWMU
UdmTw+criQZfOHpCsRbVdeQbYI3oA3H6S1jYILM6NFoyr2w+4D9KSNgpByllKE90fmX5c5FAQ4o/
3j9KzTiQCOzWYi6dPLenbK5xrIevz587jhV+PFosr/6lgP7RfHrSOqlEnXE9QB52N3E+s4XcjYq3
BdxKcjbDbhyVa9lVCjMQthr4uxDZRdejkMtlKvP/2XyzFDTGdrGRQzVW/9nIDaGLkIch8bHY6HsJ
u1UxYxreQwq+u+8Jxzk4Etg/Oj9zu7xwvYl4XuGUUxJcCAygixiWN+f0jtaT2rGYKMuAHSTysYbS
p+58g+Lkzsb/wiAML4Q4I7ZjuDAO7iUUY2U+a/2wCo3A68RvkG0gpJi3yV214T1RNNay8cWoxoKO
MZH7ulm+lBI7ZGM4WIZKKA86ArkA/CNzLYRY9Gc9S2J2XfHf+DI08aV45NzR04mpLOxgnShG/ZzD
IEdodXQz/JMjmShg6bDo8s988EddBtjmcBZkZPLCKMRktHZCf90DmQE/mLS/Z64I3M9DkawfHMWD
ZEV06+xOhz0De+IX62Rw1QUp16vn3OCKN1u7CK4zqCHukZgu57aBcGfetbrpHiUJvf0PQwWlNVMc
e118v+gkCqq1p737+sj5Ep3oy/w4kNakMKmW+G4R77Px28Mq5DhFiKpWLzm8PeWblOVPsi1Qd2+d
lTbFTKtMycE9QHwFWZ4WI1BwhYbuFRgQYupOJTbajrf8U4xDQv08i9v5kp9SM9BnIlkHJxKc+Je2
/P2cUWEGfs/yCuhDCn2Skgil9aVyuKQ/HQNr/dNboqPgqrhZalMNyqacuzYOfaHybgSNvsy6IEuT
uC7iy/v/wdjiWkLXFfJYm77XI2OJAzdl/xmRlckeggaHoljEB4ArBOenhi+EkgTZvyFF2OQ6djZE
odHtQU8IxeTG6z72tjbeT87JwMdh4yvVnLmpjQ4BIzW9ebplVVOTAPHku2+yAUrtLXEhEM6GJeKa
lgOmojRRo/jQBziWWs29QtqcrxiQczPOtbFZVl0ZA5ymNgmkq0qjLqdlfZWoL1Vb/m4Wt7iy/s6C
+pXqcnvxUZ4YtZV41FZyYcBCQ+1sgJ8iYEiNidc6hro4bId5/V8/KaUEmJ/fUpOynDIjbQfv7F2E
YOgda0k8eMBEpROG5COaN3GUhA0T3X/WSV0AzgU99r8GE1J3WroREmMva6kSHNiNEd7Gs6Du14h/
4/f9tbz79iUDQfhULzrXK5MBriQHRx8l/GbWvfgmxUMzHwblVd0soYdJNpW+o8zA3tqxnfJ/n1+y
hXv3ILEI4XBxsm/Il1S9VNoC+kQbYsioDzqCa6sCRK0ry60H2bzdpZ7S0VbgRZfu0Hso7/84vzbX
Vz2hb2vGbYnUi7/OY7Rc2iT8NtOmplIXHjjKsWM+s8gGYd8AZihvTUFLwG0nK8ncb0HvuAOuW2Tv
XRUVM1+x3LvkdiwltQsC6PJfeZcxVVvp+pyFg/fMDI6nuz4JZDd2TH/teUyJSO0g+sJ5rm+DS6st
jbFU9MZ1O7/hBAEsnkdtC7M6W01cnK5pqr6XJvwxkp5HPLW3O7KekA/poWrosgx0HrfZVXLm1vm0
aZIDOYalglC1M62slrFLBUeIEQ4bQyfFHZzNlxjrQNuVxPh4GwpmPJzZGAGa/UcisI5RapeaiToG
hYPax6aF9JX9HGq/l2CRU9bnc1sk0w5d8OqoRn6IzKVPQntitokBNAtbBbgVG99arf3X0eQrH1ag
I2O3fMzfTBUNzt0GcNClxAi1Ic9pRIxCg2jCOJ1dm4vWbyGHv2TxNNqmEDDWBWBsphmKCaEPW2nT
LnHNuTJfRhI7dy9t/5Z+/GMNIdJlhaE9MJd51HnDtcxKHRlabbbUi26hn+RNcxMi55BL3ANyign+
O7H1fkIaA4pwziRUPn860ssItpb9fd73vm7NiBCLbVdYBr5BUKUUaFN06WwEbb/egDgrQkDTEJNT
+pOD57pV8X8eP6uwg3hjG9LvQKGiJbAPJwQsStN6L7f+vtjaeqkai1l+vKbGuvcyCkQZRRFTKZfl
DKYSHkLS4hXdXzu0N6+AwLOAcQWF+Kgoy1pPikkMobDY/wtdYlLREPacOmQhrpHWLsE6jZZ1BbJI
1FJPfMUZjmuC9/ZOoyNtYkfu8YXFKaCuMy04i3jnccRVkUvk2LfWkBeDjdj5qkXpzDGffXoYRyEM
2TJ/PaFG4mvo1g4LZtWkU1l/hPEkyfEdNjNDWQjSJzSvA10ZmAdUkNgATdH0ot9z5fjh65NNNVDz
408tdMR0PTY7anHI3A0PGpZBzPsGX5w7trcjq3etVrLX7NFxVxEW/hsfKYdHZn+eOWi7bu3mUWlz
iDJ6pi3TeYO4oU4vXlFRV4U+FPemptwEaTirA3c+1boqDdgBZovWpk3gfdc+cW42HYqf73DI9F9J
++yNgQbTNiQHw/xjVi6iqUODYplbZ3jTXreqEYff2jCPrDEg8yW/EO9bD7vG6aIxVGYXRQMue+9Q
HvifEf600xfRb8zT9b+08q1EyiKpTiCULu/WroR0MlF/e8nx2xLTwSPWQGglTCiOSGVVxV3e61An
q4OodXJ9/3rxAARj8hlO7NScOoi+1m50Ql4Xq5V4GpqiCeQTMbjP5QyJd5fFLJmVV3xkpsKJGeyb
TQ0Htk9OjMZqDm0vHilTJ2ntfGOGKQcRsSCMnFwgS8pGynF8aUHZG8GFzflZ0ohNICjbYuqL/lJe
6lwaJQgh7NoTqE+wSxLjEv8z81MO2EuV2Qfj7P8X61HHEVUvTSpMTCpExCgnRRnSLAzJbLdFYsVs
0ACJp9YWd+rILKBA1c4SUx1t8n9ZUf5EihQd3N5pxCWriOPEEX9mMHwZiymm9pxv5GAHU/vbRalQ
szDczF0Rucf0CAPXY3Qf1LNlpnKn2UXEHXrAFWS/Aq3NOGb3j7kXCYWK9FMRUAjSyEQBqt1zG+XQ
O1uZQd1dgePXKv52GbLiN3CYtIF3xA/LbxV4VqFnAL1OvRnSb7AtdYkbCZluJ0XOu84TwWLl10t6
J3w/s7J4mHmpfnAdtNAug4tS4yXlnNRrFQrMSiElcpVNwBNjKg6bkU992V0lg7VRWOjPo8kTdoDv
ox5NmE4gkmjumXWaA6AbJlG3AsYTXJHrZ4bTs/e2t3rLmUxdp3ut+4VH9/AZkecxV1DteJYquG1D
g3Hfqs2dgwzD/bY2IRpqEikOX2Hw5nkjiEU+WsjMcSYZdj4eV17ck+d4Fphx+kB0gn7Ewow8LcII
mE9D9vS/Q8JB6nb9LwCcf2cJWjkrdSZ2QRLKLpw+X+8cwKm2VxftR6Mcb4OQyglWAaeJ5Idt5hXg
4JAjTLak8ZAXjoFIltrvjciNHTcAGHOn9dDe2q6OI+ZlI/94jbvByFfFkxiOz2vdQTv5tlJzDg6Y
H2kAS6bCr3XC6FHAqkDejI/GgPjOsWFRMSMEdE7lH/VGMxsLPIVkcsHBsto2cNW8yk4zt5IFpxy8
Hn6/b/Ux4tiYFarImPgzioQcGRSniI4vqpuP9d8B+U0iC66LrQq9bNuaClLjH8+p4a1U/f/b2uM3
v7xxMz1pkBM2EXnj2rMqlOgbQW2/yW92UU7j1a9da6Ooryc6mOhfdY9ReVjASObxpM5Z352gGUel
a3HgMlZrZ20vPc2j5rjXPillr7TJVIHaYj87HgRzhpc5KMztuYo176hYnQpSatyn4P88LEQaFVWS
39XOL/sQH7aJklgnAmXPWzO8FBp2dQWKspOgZrzvO64h9OQW0PY36+hVVi5OBtQT0S80COVG3kBZ
QO2dmYzYta683g/q6ucinhDhM9uR9wsj4cyyzN3JkGueFSFAERALt9ABlKPzk3iag8hldPlwgCY1
YVpPOamASjAnqsJg9xqG
`protect end_protected
