XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a�Ѡ܈+�nNX���"��̑�9྿'V���'��G�4���Ԝ�hQ�ƈ�oQ�m
%���
���[ ���xg)=�
y�ďɸvF��K�hvL���N
�|!���Lpx\�r�ª��*�2��8��U\�CwX�%�����&V��83D�@Wo)zd�&Ι����+E���{�VqB5H���^A
S��#���byJ�):�*��r�Ǥɂ�e�2m���U
�S��x�4�L��Zx���@��:��_�o�ARג�xox�'�2�4+���@Ȱj�8�u�i�X��㯆-Y��h/�t~Z>��;�b�����b½�gR�Iunt��c��|�,.�?�t�P40t�Z����9��0���H��g8�"9/W�ŹqJ�?���3�:u�o���ǭI���T��_h(?C�_USj�z?I>/�-z�ћ���,5]Fb}��x	|M�;d������c��E}�nVt��ɝD�3����(J�i���Pj� ɥ�ľ��)�ݲ!0b&Q�7BAI�!>���N���&�@��[D�6��7�xu�a�S�ޕwz�dj�6���GX8��r��|�`�ԫc�Z��Z�c����nK {�60p�F�G.��F*[��f�WJ�@�A^V;��X ��s-+�����n4"F�n-�� �(�AKZۦ�\� ���:x���UZ�?����L����4��[NGdV��Td����	�O ����2(�UQzZ��X|���y��P����0��4x�XlxVHYEB     400     190+|~�vR9��i��ܲ�����R��4���! �0s����yԅgFJ_��R[���U��$�:���7������H~�.���i���3~�J��Q��K�ENvF�m����N�]��6�:�z�.�$:[8,����O����~;#Aޮ�Lbu>��ԣ�
[���#H���7�m:�bJ�s~�0�-H��ƍǀ���G���Mo�xS�4v�_[�� Nim�vzv�Uۻ�.�nE|a8���Z�]:��ed������񫎵��P�e�~U`���$��c	����0�}8�K7l=��@EH�QO{#�kJb�ŸUI����8[�"A)5R9�U+���o���?uRvkա^��z�	�O�"��}
����'}	^��C�j�3	XlxVHYEB     400      b0;롟�m�N@BӢ=�x�,&����'f~_o� {��|p���v}R�)Hs�d ���$��8/�Q~lK��:�B�⃮�(܅��Ors�Ip4��-��#|�I��(Θ>J�c��C��Sz?Ī�_�sL��xa2�����̓�EI
p�λ#�F��&�� �v�|QXlxVHYEB     400      f0�Aym3�q�cȐ�5�>M�PdK:���?��$����?sz�ޛꊱ�\p4A��qǲt
�P�{1��x,�H%��L��v1����:���yx/����i��"K�'[4T"��������׷^�_E�0GLѰw�a�9`QA�n巷�q�7�����'s�&���
lv���(�To�o�>A�U;�K�"�?d�mn��~��t�~�ԩ��٤�{gy��|T�|��`\����YbAXlxVHYEB     400     150� -j^�������v��»;cŻWT�.�J�T�O-��H4���T*v��IX�o��vW`�,ܔ�O��mޮad:�M�Z�����Jc��G=ե��$|\ _���I�'4s�'����	%?M:��֍��q?�sD,�	EQ�;��3�ZP� ă^"�>y����J9�IK���F8}�i��r1'���j�r
|�3g}紎dP��P�'+W���ޞR����5H�������j��1pl4=�}T�c��h�f���CD��Z91������H�s��̌zV�b6�k���5��J���o���KD޽$���u5�X��u��z�%bXp���G)_Jɸ�XlxVHYEB     400     160:�Ĭ��(Q�L��IC��H���ay�c�h �G!�����	0q<�?�D���%�^?T唄)�����'����@b�FlU_��z�g4�:2)a녅
$Ɏ���=mT�%3�*���s����֕>(.~�*u+:����X��1 �6��)3 ��\����W��D�~�Xz���=�[�Ӡ.��cG�q��;8%�q��ߦ:�����B��ڮ���(��n�)+C��&乖�I�S�&�k�E�����Y���BB�)�,/�2�E���V--��r\�C�ʹ��0����k ��N�%o�|C�[ ��	S��E��S:=��]�����η��Լ�!qXlxVHYEB     400     120gmfu+�,/������=g0/K9��_2�D�L�2Gް�zN�����Az��D�!�S�G��r)0����=%� m��r��Н�(ٵ_bY�Ek�$�ٞ�8��;���'݈�%�Wq��Ҟ�Gm4dNI��$�e\��}?�جK���q��Qfi��qɨ�1����7
w}�y���pG}�q��i��U�щT�ƈ=|���C�1�H�ۧ��ؙ�Y{���7�K�!A��!m��c�!���?�����qm���˨
=n�H¶�>`��XlxVHYEB     400     110�N��2�!jp�bp89�k!�w1ll��/+����I������da���!�}���ڠ�iD�i��{VM2�6����2����.cI.Y3�f��V�rHeυa@@xC- B�1����x'v(�U�t�Z1�R��� Jzc#�e�H�����a�
��D�����xo�m� �ʿl4��2��Va��<e��=[��.�T$<��ʮ���,��D��c��Y���h��&m�E3���Z�Y����;)Uo�&�T���cA���^��H��Q��XlxVHYEB     400     1101��3#��+]hk�d��Omk����&bH�a=W�~���o�������}�7�8�+���^�G�Q�w����䘫-62�����eߌ�z�d����[Oy�ƃ�(2�j��~\��hI��~��\G�p�gS�U�r{��� ���(�=lȢ��hꁏo���.I7�
�*1�V�Rn�8H����}rEy���fޑƴ��vJ�K݇F�Y�Zl�#��.���,|�<&%+(}�D��+[�:���]�c4�$�,|��XlxVHYEB     400     130��ޏ;#�(A�/�ߍ?�յ���A�Dά�n���y�Hd:~���z%`�q�w~��|9u�]ܘ�c�d)ՆB4[Hb1l��*,�D�3p��3�lD\nh����8�|,�-Hnu(B�붒]:h_�7��̿P��Ԯ�N���:.H�;F*x��R�'�ˮ�GY ����;��t�K(I;���k<	��!4(2a���9|�_�~�T�}�P���.{&��l�ݬWm�@����t�Ǖ�<���I[�N���T1�2��%t��JX��>�?�䐍ss�ԗ�r�\��]�aeXlxVHYEB     400     140��#G�8�k��g�i?�9�q�fe�;2�6Z�,u'�����f7Cfر}&f2�2Kc��	֥�NA���o����	��%�t����K|�)�sJ���z]�|ǢN�N�8+�t���s4d��y��ɒ���v#wR��1P�b�
������P��j�F1N`�3]lS���ߓ��
)һ�XEܽ9��,����X��%�"�ϵ�:���̶-
졛�}����Ֆ��_]��|gR�0�se\��m�>:� �A����p��`����O]4�*]G��z{> y{̟U�O[S�f"*�I� ��בqU)XlxVHYEB     400     100Wj:���Jgw�'���a����:��`��
@�Y����)q�b���\���.I����D��~�#B��'U�}F��4&0n���ױ\��9�ܛ�(��]���+@$g(��W����n�.��YJ,�Z����23��?5��{�IDE�+�ؾ��e
/�d�/l����(5���M}��e4~�B�O\zm�1)�넹DGhoZ�<����E�xb�,���븉�;�=�}�Ԇ8������4LAat�Yl�XXlxVHYEB     37b     1408��AMω���ě�5N'tM�>����W���ʿ�0ʏ|�q�Jj_A��j>
+�p]��f/8�Nѧ +���\�`�aNL9o�'��%��=�z�Ay��mC3��]�m&���b)`��9Z]a�QN����!J�?��$�ΚYS�w��z�-X�0\2 �y��k����3?Y�"J2U�ݴ�sJ=y*�N��{h3�I�<�r��i���{#,#X��c� *�F���{�L���'�d��5�@'d�+���M̣��R2�:��0�������^q���^�i�Ҫk��I�x�".�AR��N��
]8�![�