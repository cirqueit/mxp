`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
jXCiUucd7tuxdNSToSpLJiolTuZCHIv32FWUduu30EXxyM+hTv5/Kj+625pCd0sXZEIo+OY10Obr
1bvi8MTLeTmudhpRihgS0pWo+IrYBZLK6gNsYwcctZEDqkqsq4fcrPeNlKzguVADIQHnbNqtvH8y
q9HcE7lNG0vl5CJwas+feF4KDmlPOr+UWacSR9R+E2SKrZaE7/4c/9fhDhODkMX4Gv+A3+CeE9r6
SyB1r3ARl5/VWKF1beXn4/8y9g3S4X8KzaBeNcqNzpNHTD8yScaTB3huEewRnfCt/B4/6pAW/BKh
Jo7NJgQxJyM+0LlmEJVJF7BQ4K/NxJjmb/t4+pch+zsQ1lS8fIbMHcGVNxxtwonzURwgppWMX8MB
D9egpNh28yKTBMZOMk/bRS1yHVQ4hnld+uSuQEUi3/30+SXUqKWLrWOOuF7GD5dnjKO0OTHJdlco
ckk3M3Vsw+adVy1wTk7CwOt42bufcq5aUs+oYtjHCAV4TAUAXXGzlxN1OZoJZFLLQ7lE1IL3mfMb
S7uUGHlmZu1/r2UpaqSzZjmBCedc8bdyrANei03QdU9zsQELbrRpXRBHGp0rEPgz3Y97p8U0BYPS
UvMQd2KJyl1+8WQi0z6CCdRM0nA0l9vvVVNjqr9ESVmVkXl0VUTxyg9JVRVnoiOPXTl2IVbYEkGT
kWsWni23Oxa6iG1eEL/Cu0HE736scgYklTqLRe+WJx4dQaHyUJw/fP4hy4tJLjZ5ZAXZljycmtzC
RBRnI5aMscGpuEcalCtaCIwP9UySW1rug5yXRRjbmhZmvWlvM+OjuAHZ5GDV4drHJBlxIz5L3g3p
KDaRoLSYjrql1MQ5Z2bnyGTtUUXP/Yaljy1SW60YqYITfOiXrxj99MwTMHXb8NKrk7RyNwyRuD2k
OLsUgaCZ2iaD4cQJWAhYSqYvIgenK4Z/zv0cQubgBxTbE4xPDEGYrTCwz6c+f3VQvO3Vp/LPZfr/
YojWGsTpFmEMYKU7HTeVlw0RslhdZwKGShOm2cX/qMwYf7UHuvkDZG2sNOJ0v5XOxHkdvgYcsWG9
sLCRXboaMvoAD0/mLFlSfUJrbhKp2EWjqRi3GBTf0fy6Pudem4GFd++R/WZiUPAhRUJj+7i+6AcB
raUOXeBOiSsgpmnX2JfbQNOjAAPfevHljMelPFytg6Nv9c626VpHVACbWU8QXTDYm3W0mfbgCK8T
I/367CyPZfOcobhml37/ph+RedCOOx46u1iRaSog1CWIeCXT1lBx2rhqdDIe47eZ/yJE39xhNUrd
onZUEDs6eOT4L/Kdn88MQNnkoFpRVaqFQjlvUt1nS1AjPT7nZ+6HipBSr5Znwbd9GPTl7OUuSjPk
qxjk59ho15MwAEWLC6BCqu8+1QKa+rv2ed6WqkIKxFAo3u2DLqk7IaxpqD2mj1kbwPh4r+qfM0Hq
dV0ZEqIvoSG+h7A3NQFdmm0ftFX//++PxQ2PmjJ4V/Yy6QCiVjPaxow1AmQ2ol8fOrmp1xhkMrqX
wpF3wUUt6Jy44rmkZ3tLddDHyTUznARuUi5WxMYDo9uZX7bthuINjwaultDxTc9vDK5Yl3nlkIGJ
f28pJOOleAlqV+JBou5DKiivHaiTvzpc4m0pfPMnL2Zw546oMfwoz6egtzNubOu68A8AQbphPbh0
jA4gcmXhWUMKzRhadBVJ6yQ1aqcR0TOlPgz2tnQcy4PjGK5u3zwyBdOgtdIzkT6y3Arz9Lf+M1cE
0kLMtWBK0uX6rPatMaO49hoAM4/YlKXUT6CCWUIO/JwtMngzyuLEWPuknrTzN4N3anmYzVm7gFKs
6vqaABAqVAATN6SFtej4pwePZQxgKMFzCKWEJWXeUaWMnNxmLtqwb4chz8aPaPXH4ZNJzFBHjk22
U7NxPzo0rYmwu9JmISKpXArLwKGtGY+qfo0eTOyzhh/MoJskBg5grin/AquA5bkkqnfAbsEyIBqR
6i1hPwZrEfaacnD7FDqEsjqgF8GYYgfUesunjWrJmKT9pE2dW9vrbI4IrX0rTSLY1eldV0dGyBJm
mwTaDFm5L2q0ufNaYpKT45oAzEcOOU1rc3DA3CCvRFxsBRYsYMv0hZNomjrZeBIEYNr1FLFszK30
nryeuMsHQrvT/ibt0e0DQb3ExMU71KCoI39VQJwk+z9itPdel3cHfXGBRADZGoJn6K5/qmYjIaKO
5X3qj77BtQcGSq9ZnRcZCQWCrxK3iSKacVEk3hM9PlyBXjgv5n/kZ0klfntv7/AI5bR3Apth4h6f
jnHi8ld3V94pl3wv0rgk68GAEK8BZdycO4vHOoiG/JsyJ+KyZk+MwEdhURcZhYdtF8z8wY5GcBIs
FntYpA5fwvVzVZEELEfP8MfQcQvUHoSOHyd7Ar44g2Rca2vaBCH7orYJpZ+ErUQcRlFK+S8pIRyp
Wld9f29p5ZOSapJ/R7bWrCS/9gy/OqZGzOplmm3Ix5dKbV5xfakiuH3Crdb17lMTruM+Uq0/DwKe
f900H0BPi7UvlZ8fFsifVZla6cL1lC0bEgXcUMRcLn/tWWJLV2yDKYcVjSjnVRHJSGmABSPaWzvt
DXRS4mMy7EvkA47nsEWUpw636Mu5WK5OyU3VthJS9+UjeIvFfqYCuVMEyiPt+E4ZPcGJzm2IHOId
h/HErgGGX6UyE+In4Mra5uoFPqe1Ui5k3NP1cyZk55oMN3blPDvr6DkvE9LxGTdJZ6hdFBebEcDr
YXZZpfjJ7Pn+b68dsucvKSO63bBPMS8Bw7ChP+RfziMZO8RWKiyS6mycyFKn5bCvQBOgc6psAh09
myNjVt18Qahh5hmqLVJ89LX2QeCH7fmexS4kjasWv2WdCdym8vmqL/OFoPT36RAIZQchQlxvgqQj
mFGrYMxQZd2Niz7nu61uokHhRC2Kj2m7lXc2Z27aTdG3pbpEgrz61JgZWfrdfO/qbWhJUu7lUpxY
mlHDMqg0usOIt9IyeIyTj9vcSNZBhu6Ldw7h/f+0kXusIX3YegVEkL1h6a/Art1bh9Kf4Z/M3JCW
9pXOjvYVm7SY4l8HBth7lw3vneL+PRGdwiRoGlN7eb4XawUTiXLCiV/KrktgNTJA5gtz++9mMsTe
GqR14+0QLGRnIGW3g040UBU9K6QiWXq81PK5jFRgpG7a+S3aOWqIJPDsd73WAzUXdzKSAcj7Wyw3
2CsE5G+U9KTzMHwfnJnCVii6gqXY5ALlOEZQtn94XBPCjOHTCjyRt7gzJ2P+GCp/LxGvXTMfE0bq
xmq8NvYpkRfIbvxRo3LYH0toVsPFmoRPFnOsynYkRdLng9jwQy8uFEmQXgxcmTd5Fl2Rtae1OsG2
MBqCWPSRsE28IQIKYQDJnaW74qsE8DF9BSpqths19nq6H61r3gLqABXfvqqNqXwFFBNcEmEDuDm+
qt56Nu05hMqm0pC11SVfpDAhzqXxt2XNxi1sftun0PwN8itLgteNUNZ1cb2pf7dp+8vHhNg3BXuv
7yzaOra+L8dKgy8HAx+huZbykD5cX+Ydai1BYUpq89O6ZZ5olsZTBfoOIh9F55dcVRo+kWspNT4G
HReTgEGp8I85C7nEZopahhH3upvUcuJ1ObGT2lkiXwoTil8wvrAQ3tdz16FVPdaAABnLmxD4CTNG
aZPbbEn83KBe/zS7NX+0C19jfBtTOfX3wjGnlm4fjLf1uqZH9XiA1L4N+vBNK4JEL6JFKWdWlV9V
z4mdHIvReYCl3yl3h3X6D2gmWk1HPCuIot/NcQT5meyoQpQtAlIsIPVPHm8+fGwkkglw1YKFwex4
wbzQl0xPUof6MZ8n8LBLv0i0HIMcJ9cy/vWjLbrYNF0I2j6WWTseYU6CkVAeWxuzgSYBZH67jMDg
aPWmddsp5Jt8Y77QszcnogY9/3qqpV8uLImr48kX+MlCTDGnkixgppGWswQ5hkRQFYifwR5FJAnj
6+kCiNu2dH6KS2IPvvGh+QmAOcGXW6R9mtImIHnx5SuzSuvzn7W5BeR1HIusiBEV9UkHlmFGRU6V
VPGhPTYjIQEvmDir5DwBbllTxLbzbxsXBTsN4qTIou4uscu7ChNRP8P1u/VArAkcoWbAWvCFNz+Y
5YEjlhO1Y6WrKwr/Aiwr/1QtdfxQqJ57A3rPFiGZW46x2pshiTMpYQbqM3Ag4KUhw5j7FBbobvHf
zFVZ1NFFL2s98NkZl87stw5SPlsnH0sPWu+h8HvjUbaBWJVU+KHX/YHNU5zlK4suWXR9/1lYZTJ1
mtRBLrCtLH/NPSmpczMG68+2flabA2SmNG/Rveo/LhxmgpsAlfX4vJ5P3ySIW7Ry24w0eFq/csnD
/5wA3xO9tNLPBoasTiYU+BnynSQTUuXKfHn1NM7dekZ2jIpfNjL3k0EFi1LPan94hAp8OhmSgMgP
pqkEw1pMtZBm5XwDrUXdwqWxRfZt7Wv3UpIWUyeNkeNUAaDlX3E49nk8NHUGdWoHLbeuDEGvYEep
ftaoS5iEXFAbqxYW+JOAuC7dhslCVXWbmaALF3cByBA1n1kjTa1MszJmLXtJGMH60vjMMCx2iymd
fboJa/YMRxOwSCUJPR0J3fWkoflPalIyK4PjHzxEOs9sYRPKazBTgHi4H4EUrn1wdB3ivU1MrpUq
y4Sui8xR5EvG7hEFdCtscfAJ+Nu+4g0lv8R5Lt6MiEMaAuoUAgjkqtM1P3IyGFZCYjAAMXHQ7y6f
86ngxtUqvYn1vstfKpJHwpyPFJlw+J+THFgco1wmbY2g5RmnoPImsDjqLiK3SUKxMWxjzQpKCq1M
lqA+zY/FMHBEmkyg2Dr6+ZadS49iQpext1mrKLSWtUV5TL06quBccbaOMdtrrHtGG90fX5uDhtqS
+oxPJbzXRsobcuTrEzE+h6HdKNv6C7K9wB1IOGvT902d+ITiHGpCHmXuCk4lElKU87j//bO1f2WL
8kdhbvhORle0dANFDj3fqMn4Vx+vNK3kImEizGMhMz28Ts9wfzqkWQFN0kKlwQB5nuCucLPhYhOl
8C7cb97iYTRGRNM0swJuIHTXT66bEElun/5hdi+jC8R8FC1/57o1wcaVx5P9gFTwJqXr0lfgE3jf
1MpIVvzpLfnrl30n5OmzXZHYYhc4
`protect end_protected
