XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��f.cV`��*E� P�ՂX`��X%� �i��O,��)��*#UΚ���,�4Ӎ�Y��I�P=��I�tѫ�?(��(KJ�yim!��jȷCLES�+�����w���դ���ַ�g�k4��A��A�$v5��J/�K�Zu��ߚ�S��}i#��'F�~K��K<Ei�L`:��#C��I�
9c����x?}�D&��@8���s�����`��R���e��EfU�\~�sm+���C�#w�N���к�7�Jv�fU�B(<��2����l��v=�*ꑕ%��HڦSӛJ�f�q��l'7�%S[�Q^*Ғ��c`6��l������4�~&>����,�ۯ�"�S3\a!Ƒع(B�]�Vv��q]�K��CX�� �?��G��A������5��zD1��nI& �2�k�LsJ�$�7Ĩ�$�=&�7U��d�ғNJ[��L���x�Ɇ��ؘ�%�8�>�n�.��mS8,ޘF��u.�i���Ga�ca�r~��ubܳ�6�6�G�,RwLw�� &�w���05ۚ�!�8�m�w.�6F��Í,Z~�_��D�Sdm���T H������B�8��P��v�[�t�4x�y����{mA)t�-y	C-���)k�҆
�N�wN"f�Ik��	�Ht�r�EI'�`wtk�)_����zz3>��Kj��C�Rf���.�yՕy���]2��I�p�~�����h�c�"�"J�t�G�I��=�o��jC�£;�+�(zOt:1�XlxVHYEB     400     210'�� ]���ka�aoc�?;+8ꅺ�H�����Ci=��W0��h����9rE"�X�x�"�`s���aco�#�#�, '/�Jf5�}�����g�7R���2WW�73}�}P������GM�4#�����
��r~JsR/�#Y�j��rEv��:a'�P��͑Z��x��C{	��ص֬������rA6����J�lO���Y-�u������$Ȝ��wփ�ˈ�^΀� &�PI9bgʎ�8ޝ �q2P���_(?�.�R:�}�C��0�7M�Ѕ�A�ku!�BK���1���ZeJ�Z�m���}�;���1�L�s���� ��v��Z>�����i ��%���xm
|x{g�<��i��P�kт}��T+ձ8F	�+�^Հ���3��Ѷs�йdF锓M�X2��d@f̒�!p���)p�����#`��XL��*��|��,i���Ѭ^���D���-
yA�Z�5A���?ͨ|~�T�ip��S���G�����XlxVHYEB     400     100&��=�6!"ͤ������*�:?ǩ{j���,[P��)�`�6�{���:-�	�� �Q)c�1�N�f�s��[��� 3'i�I�֥IB�"�<[K+2�*�c}(�4��+�J��hٛ/�q0��?߀^W`V���(S�%��*�[zX���42�G��~�ۏ�Ƕ>��e
��N�š��ڬ��Υ!s��Oz󲲲�rb�,�ӶEb�4A�h�*:d��lyl_�i
�s���U�)�VXlxVHYEB     400     1f0�v�CK�WO����N?e������t��Ytv�
��<U��Q�$��$;C:>�8�T�����G��{�J��
e��
{��/D��6�h6�<�i�!+��e���1DZ���x`4�z��[ܸo�5�}1|�H���+i�[`��G�Ìn����}�:l��̮q:�d00YG_��)J�~�\��>"bF4��tq���g�%��(�����W�x�w��=)VЧ��/�X9���)RW�^����ߗ�l�F��E�6�J0�ٛgsR�ӧ�Z���ϐ{M"ze�ɜ�pw��x�T�=\?gBj5!��x�OfX�mt��k,��b��?�B���<;)�G�t%G�����n���������y��s�8� ]=�x� �z�x�A�^���8Yۏo ����t�VOJ�j-��q���KQ)j,z �j�N庡jb��|C�k5L_ia?��������s<	���B�?i;��l��d��Ε����M� (
Ėc{H26>T2�XlxVHYEB     400     230x=ڬTޜx30J�����P �%'����c,���h��n��~�0x����iO�4�s�%PM�(x��Kq}���z���ߗ����'�<i�H�C$�|�^�T�\'׽� �ڑ����P��Ă����Ɣ .���_��f�c�Hp�Qٲ���?U��l����)4m���es��1��BL��e�$a?����	�8�ǼrQM�������c��?rD+�NL��c��.k�&�kb|
�<���ң��~_�	�΃�W}Q��Jh��-j��������l ����l���'�~�q���]8�VP���О�V�5��v_;��.)T�T��	�� ��8�hc���s��P<�������l �l�����J�Ea��E	(Ik湝�"����&�z�.V%�ؐ���DpP�����^d�w���ߧ�K���rn q]�=�T��F},��!��΀s:��b�%1 �42Q�Ul�ۯ��k��Y�+����re���gg�3�Ea;��p�56X���ot��g�OAP7�;6u�RS� m��.m��|\u�XlxVHYEB     400     1a0�N�\4�,}k�H9M h��?/�X����� 3[��m��n���5U5sW����z���p���t��J�����kL8��!P������7b���x��#�QI*��<FONB7GsWT�IS��
ǉ��(x�c�]�i�U�]���<+GL��'w3����|)/v�UO�v�^N��pW�t03)��<��A�Jv��/�#�B٘�-�U�V*��L�L���[��ߑ�U@��3wS���ܹn �a�zl\���I�Z�8f�e2��_�܈��%��ͿG�'�p�0:�&����}qu���E�A�^�3��ߊ4pS��@
g+���t�zK�ٵW��m�VS1p�1)��m=$�dL3lf��Y$/��T:[Z�$n8�ہ�v�������x��{J�� ����(Jnޙ�XlxVHYEB     400     1a0̬��:�����s���e^�h���:���3���)��`�W^�6B��2���,h��B�0U�s�S�b�1�f�;�8��!�# "2�D�G0R�F�u��)�=���)P�������^�%�a?��D�G^Ii6��4�u�7BhP��a^'FMK�5i�YN��i�C�.d�p2�#5/w��#e6K�^C03y���3��1B?�����g�mǃ��\B��Fv�����s��c1�I苙>�tX���5��l�Y��\�h�&,������a�w%3Vn�(�[|�py�Z��U%�9���b�~q��m�rn�J$|��Q�N\��[��`�q��cC�\��~�XiF��u��Q�l2Z�������H��?,+&�0h�`t��[�&���� ׏�-t�7�/צ8XlxVHYEB     400     1d0�/��K+,��Ě,��K�/�:DY��_׺�"�$���%��}��2����Wdp2].�~���e	!��c�qh�uv7�J��Xi�M�����~�:�e��\~"u�+��v��{�MR�FG��XK�<x&�t�C�|�� ��^bŅ��51�E*���D������;��k�P�|F���=6�J�� -r��e�N�/��z�R�������_,�����2��M�Q'4�U��묹Ck��/p�,�Ebʻb�B�Fx�?]#м���Ydه	�	��
�/﷙)7�/FT�e�����Xd�u܃@��ȝ�� �6�g�Bή ����W	�O�A}��-�0���M��+qŻ
��w[8�Q���9�g<���{�V^S&�  �M��K���W�p�Q8��t�$�U���-��W�� 02���ee�]�2��L�T��n���W��ҢVe:��[6XlxVHYEB     400     170��a�)S��4�翫N.�dWﵳaB�q�,�
�D��G��&qfш� ��v��ճw^)!��7�_��I��ғ�D�,%Ƶ��n���!毅ƖZf�,?�:ô�K�!�Y�%5�o#ی��T�:��Ƹx�	9$Mr��fj�S��M���×,�;�>6�˹��.3�!��� S^������	[lW}���_��]�b@�l�\��-���IZ.@��t�\N�Ō�olgL��VB������?''xT�b�)c��iNd�f�v���p����R.�7��k+�NY�$2�v �ÖJ�B�g<�֞'�fk�sw�7�T�4��Rq�f�}-j�!#9:j8+��pI�y��ޫ��@�2�>��8�eXlxVHYEB     400     1c0��i��,I��o��mb�!tg>b����K�C�������`�icxU��=�p_�����I��~�˾���U����NOF���;���\`��Ww8�QDX�PX��ao`:D�|�#�>��v*�]�Оӛa�:�)�������%�]��6�KCBh��|� H�㠵9�$��=�K���	�}���3��X�2sc��8pBX��~.
�I� v��	6P�X�l�^����cq�[{���wg4�/:g����r�ߺƉ��Z��D���
6k?:�lS2{\@'yI��C�ڿ�����Y�0��z�Z�?��};��ӊ+��ZH��`��%��З;H��к^���ܖ^EP7B��X�UU�A	9���|�r��Ua�gG?# *T��Q�6�+�@� �/�&Jz���Ϯ-��ֆ����M�XQ�˵,I�G���_e��$�]�]n�p�XlxVHYEB     400     1a0�hߒ|#��6�,����S��9���B��2��{��i�iE��I��$:�wVM������'rD;�"���鱎Oc�'s�E0�Cw����ZW�u��� 1@��JO\T=� V��P����m�n�d�nw4;���Uz����a����Μ�a�ی�{�(�D��s�l�g�Rek��g�x�?/^����\�/Rݔ���(�Ĥ��?���v����.B��XJX�ⰻQ��M�Um��K����Ȳ<a�
G��ʂ��/�`��h3��B�C�Lr���5 ������>$Zk����l=��T-T�P�10��F�.�`�%i�g6Y粴�ba���$f}������l<�v�Bq�D�o��عJq����ռz�l�.��Nv�$��+��S�I+{L��*�E׫;�P_XlxVHYEB     400     140 t�^�dȒ��a��`����n-����(�(�^SM�\��sO�������n��5��ii���g�V^��=��I��Ǝ���_�S���W[��h�/K�^ UٳJ`��Y~�^P��`̵��U��|WgN^�Å��	(��-c���x���y/�DJ����)$���c�:
'����y��|��ҩ�R
7�s�
���^�V�\
�W�G	d�J�G����Ѡ9�ր!nP;�D؏߯�������wڗ�����z�������.�?z̐��Bm�%�!	��|\c��.�$�\�s �m�Z�������I�[ȏueXlxVHYEB     38a     180WD�YyX�>���5���Ռ@P �yZ���u6����0�m�)p�w��Z"�è�#"����l&��S8|�8�Vi?х���2"$��9��Y��Us��m7�a�Ć�~�5 ���N�残q\?��=ҹ���'���Ϙf�$W�Al�mn��C���r�D��^E�@���0J�g�ozW���W��K;�(XS�O�׹Ľ}(�����c��V .Ԧd���l�1�P>��p���6֓H)���K���sk���Dz�-1ⳓ�M��C�
]��U�������<a�Pc!�y�뎪>�=�v�{x���D�|Q�CR��4Ɂ�c��ƣ"o��&x^��}��d�.[Xc3���P�	���X,�ӱ��95]�Ӆ