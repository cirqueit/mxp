`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 100176)
`protect data_block
4mScayjGdBIoO5y/yFH5n4rss53PBV92JT9ecmDjBzi2CSY9Prx0rvvvzptV+RdKJKIbqnKYj8o2
x04QyA851+5S/XAtOcptzc1WKggnxmlwyK90+6XRbdYQOQr5EqpRZ6SbUhSsKdJvcEtzmZ5qjav8
l1lFlUA9iHF8BhQ0mpOnGLwxJdG844cLU2rR98RAJI8wegPrTFg8QGa2qWCDm6U1F/KvmLbcCFCL
LE+cAmBKWyP4hPe6auQ6T4eHzZbWoVRjFAWhtSQhrHlfMfV3Ss+blk8LRuDq5gBwCc8gZ3L92UZx
Hxyx1x2JPia9S168fZSVXhVZLKkiGbxDwsmFe5WYaqLSoTEOelpr1aDh5hef+KL+Cv/m+RCKzNLa
EfA3+P2NIwWOhMjJ+pO5v93gp4dQzHTZtM6EOyL00GgBPNV2a1rxoU00IrtW7R8VdhZRNVe5nixl
CfmIM7aamTZ7V7q3lTE7HVGhVmzp5AmTMtOBzAnQbfw6B4YDSurEWsjjEtNdD+9mRLGxhsRaRkhz
g/fnkGXFTigz6tsX0UUPbA7hsH0ebh82zLySoT1KMKbyK281K3YWnlB2vRJKuVaCq/ZU8ms6hm6L
+/Eh0urxcSXb7Vv+kUyaOlsOQa0UY/ThUM9EF8wgJAv/Qnd5luDmdOMTzrcA52C5wi0DS8XfyqwA
gAxLYxwygQLx5pYnLq1u61xbRxql6EFLczmlEjEv2yrB/ZbhE7XANN8YdegXPR8gxn1LGQG374uv
5iruKkqCBz4LCfhZZ6bMnW6w6MViJjIixP63r60AiwFs+FrA5fgdCgtOLvDlNX4MI5WyDTae97c3
ePKTAgoaNLUMO0oh91jMxDVHFXKuL9hw87xnSe/ffxRBl0zPtq1uCkF4gj9ayyqv3yeuCGi8YknS
tvQChJ4qY6V+CwXWxt5R5mQBSA+X68ObPFqe/0qsDtDZV4pmuAq7sURPLx7n/Gxtdnz//8E1awqs
5LwP9OHGnbiP+gkWsG1nGXc2yo0idWEGR0IvTG+vZHrnzmsYn+jhNHkWyw28TKSCNMoJ5u/ydtf9
7hbtoOOqdpTKIeg0ikMJWUPIPU+p+qNRBV5ZFiDCz9O0aLM+HrsGG4FzlHJIhLzlHNFSQVCsU6Wx
OIh+IIaRpOAuVnhdc+8685MdeLGxSjlTN0fK3j8nsAeNB/k8kwEkb4+NkkgTEhMyUhAuWOL+6O1X
dI+A+hg/ZIksXV3WT4wbcC8Gqr9819eL2rmd0hTyrfdXT4sO25BDf/XqbRzB10FN8iNWJnmGYRQU
AAbxFgoEpzl6G423gp09ALqJb/ZNsLYWtApP7cMhFuFgoJOC3VEn7P44YGZOozU2gM5ctF7YmccO
Vpz1PoBvPLNZUu71R9hF5d7FNJuVzqHmvryzurDFp+r1pVqoz7dNyxWaXEcBKzZxmHS6ur6yVTiF
/r4tm918MLqN+QCgTWYHfyrJKCecqwsv7PHUxTX+RlK5RWHlt8tklPIKDKVECkSN1sLqeLyWRfKz
YY1GQFL0za+cDZ2xXDpv6kRoZX7noC+LN0axg2LwjifKbQ6KtSnI9y23qf79uCWN64MGe203Shba
g5+5+gcj50eyGUKm2Y8yoWMphOqq8mpM4wgADJ/12G9zdCw/RKtVN8MmGeau/fSFtIhn7VAQdrg2
KGF3jFxPbm0s2thMibfbViFZrFNoVyL1ar7aanfwJ98WtclvXYHP4+7B2P7oFmXnTSiUB34mQkbm
2RT3KwhIapNdGaoRzzktNmzrQbgkYjHBYoyR/dpIfzu53YKusDZANI31m1SKk3hQNPUluNQwnuBr
JtWRKAUcrvobFNWAzTpicZKI1pAXsMf4HgLUNBaHQpOO+dfVfFhfdlvUxaZXkHPa5yyZh50V9mg6
q9MP1879NGvAAAXZSqlBxyexHkddJQaS6KnbKKxL8oTvOZzgGeqnGwY1adwBVE5pR2v/neNLq395
b41z3tOljxE+aBf0kkHj9muJaHWs3rHlVTQP8tuCex8Wxb7A1w2PAZujEONuVLPlYAfZLZq4/H+q
4MqQN+BIYFO0VWJh58D8oH8MxLDuAzpMwUjnlnHS2hclf4LroKgY3UJO7awt27cgq2U/2nSNNLm7
HwwQ8UJAgnpEsrxX3/cq0RZx/hqvH+AwpVcMReIUbrDMko7RDzriKttGW/Jj4PrY0usYCL4IEqED
RbdVcDxKDdMODfkfi4IstX/AkbZd24CEGKIy9EyOgw/jCXBIlbcVRxHXo4yB5CzTG5615KoaQQEy
YZnz/XkSjCnbSnUCznAVqrx6ejDkrSkhQqZq4ykxx7riP0ZQAlwAtu6Zg4MjtlRUdbdmPzUqgpJg
OLP4rJIyln0qbjcTLVgZr33cfNKx/mYZ0AqfojMa+jea4Dr/b9+6v8JLt5cQZce92hgJ6sU8lO/Q
h/nvljBbcahPGvWLv6cprf3jwRsC1YTnQjYWEUs2DoubMFex++lp42kOOKEnX8TGYzE+qy8PcUPU
kl6EPnBGX4Z/0SlrLPZbOTfHuFTxpu/ndLP7V8RF8QQSzGcKOPi6JJ0Zo23VUzkTAnI9WeXemrFm
F0gGejSlPJ8OyoQy63M/HWtTUuw69UvZkDJ9z9E1zhZutNSe9/EbFzexHkPjswDaebPVVUij3KI8
qZBFXLPzwzClNSatubLSdZ9gjtx/da3oPePU4wxOxCILeX+Cq8wO7/eG1syesBOtw3FNyhlwZSr7
/IDn4NTYm9byfDSp4Ut8SGDWRc86BagcqEcuMTN3LvigA5bnhqqwbtXYr9cqcvnXuC5aEEg6G5dp
Gs7+GoF+FtlORc4XCSL9db0Ggz8OPJpe613dZIybR8osNvWX2xdQwn45S49CWiz02hh1QNh2DMvi
bIEcGlzTb6K1UC36+//O2pr6hGw1UqZYmpBJvOG/PedXyZyAXlu6Cj9ecOX1LBKqLU8rYy8SaiyA
PJH4FjEIoAKclrhPSwiWhazMQM/svjZZSQKcgUd/LrGoI/nru5fLV2+21ZOUcvI3ENmPxJBR84Tl
9YDheD04iih1JQz5yhQXzNQDoXfFEC9I4rfpM6P/EePTILD3oqe+YnGRDkjei3OneckDldmXCTAQ
BqIPRUffhFad1gcH2kQI6UXhmMxKCNMScwiNiYJAwYbbrkafrZ0DFPaKolnGzniPXTANKJgkyLR8
OFv0zgSYJDphcC8qsM21S0hchSc/utZRfXMsvVQRTGhO/Gey73Qqih3zhUBhKjySxX9ee+tiVtZd
N7+Ox/Kt5UK4lb1JExZH4SmhnnbtJf7qosjQNz83aJOLxOtCgVPNYPfFpgLX6H4GbpkBZyZaeWnn
kD9KakRj3rfUWox+jpLrrCsnQfRpHt1Rn5a73bZGFKFQFFxFu/6Hfmvda2opDKnwI/T38WQnIBhR
mAxyJq/3i5mwnyEkSw2fzTVcCkhFPQZgP7nPYQQiBAfmGSRkLbsqHFQdBfTdbUMAtStSGL5JNy0J
94cKzovPVC1j05l5PeRbIPK2sxXDZwGw46WpO2qZM0XCoTz13qfzjotMtwpbU1CPELGWhALJ4znG
FLy9WK8G6sgePS6XiVjeXT62iMRFKaVeRxor2Y7yhpGFVZNtjSHuFSHzgwQreRsqK0hLFxQ23qqG
lFoc6Ag33oERJP6MFQKtWULQF2WpbkywGZFJdIsPTaWUEm5pwXFFQxjiLZFQt94jMkrK36rBZWlq
FLimLV6LHoC2ADPyybmwRQd/m9UJB5nDWopm74DClG8T3wCMC3e/Dnsqmo/i6guX3tpZNxt6wnmG
yRcbqttWBG5yovJkW78Io9FmdIc3hjYjfrvqrdh4ub8C+HWIiKFd6RmCHEa0J0R+IIO+LP0XgI2W
7ZxEo6fx00WkMvS3dEGrBOqonwFq9vzUDL6+FsDsEekNWmvVdBPFeXeDwjG/AYi8Bknxtrjk7isi
gTvGHlG6e+Y03TBgKfg8Aj+7rRHxKdQkPWG0Ljc3tSEoss8QWztyPGKOx1pEqLBa4BaqIvz/6ub0
w+8liyjY20XBVqznnR/dOp1aAzhtB6bGUSEx3BSTnV5xidBhhbpd8BKxCxyIajymweIxNy1lj1jo
6U3DB6A7V5Wz/pkj0aw1Vn54p3Ry7XqrUZWYytSh9/iTeKAbDJgHp0DIJX2S1TruNXIXcMtS+fsS
+MsrEcDzKnofLk9svuiHI3HRaEs/bX0Cw2LyLyXQpnfnq2fM2Y2ofoQQakCXnqsprW8SFMPMU6q9
sUIJgOy5f3P+xKxNZ7nsXvJxVj+qinlx/qvEHcg0N2Wdk/P+La0RDwlpkEssuNfd7M4hlB2tzYcv
e08w8cIxsxWf2+8CbPXRhdFYLx87iyOj8GKgX/5/68g0RmsFDPAlvtu7A3ra0JoIFs43/716B6nV
axV98VVXmb4HTm3lItYvF3RjfIuqx7RJVkiZCB/7ouB9JlF8A92wZarpb/ZFTtmSmxZCZwPXw4Ro
7CdwEqsZx1qEl/z6bG8HI2xF8ex4ErjlYwNQBtqD3MTp3vga9kCg6Q0COrI6dphUa6e54ymvwRaa
WkmR1/IwwwxDWa10AIUnEEKm91AYXHFTgH9IDrHKQUV0RFh4oTwdbRjk4JgPErIeHnPiQ/bPoUcS
d0X7LoPFbo1iGb24NSdzgqHBHd/K6KEsHtTxLWY2hknfn2LwE6CtNpsqm9ncIZTI5/A2E9f20crz
7QHlSLM7PyDsfNn5LVPqGk3ir7Y8xSoo6g5PH61Sex2ZK1cXysjTKcsXaE+a9rAmJWOoo2vOh5MM
IIJLzL5wWtBd4QwJOu4ajytzPNFSuKoEkivZ1DTwj3TI1nzWAiKnHEftWgrXkZV9Qgb6wRQh6QTa
gopNTEhORLv+prtbVCnJzaKgRLwhfRFwfTGpw/ENB6HHu6XFMydjmNM+Zh+DdDdhLJLASL4tHH16
Cj5ZybJQvsDPaYtSa3xyrkWCPvw7hcQCFR5mwQ8/CiEV56Bdh1CSd4iPd67V9qZakWFQkWUOjxtu
quTeQPD9vB4pyk7MTXIkLmwemYc/o3P0BiP9+NgVJwV8rSEHvYHl6WEFHlce6Ty+AAYZA+FaaYuG
THxMYe8HhYN2eCFR15FRRg5URGf4MtmtbYxJI7ORqweTIr30lIpkRiMmjWIpurJI+Er4nd1FLMF5
41ZpwEAW6eKqlwQdp/kHddLaSq0Iy4yM+Oe9OLwIosHMDAQqA2fyY7GEjO1QGNywJskN2yDKuVzl
XJZAApDpxg/2uhcbbel2tUnEE52lZSlPzDoJkPjhp+I7FFoW0y2xh2CheG+8b9nl4Yq3x2FMrLZN
jxpltmy3dL5HQ/Kl7eY1yQIdAKX1QbmiTJVetNDlxie7BTvAv4u+OMFsYYnW5AGd/Zk7ElfKDtyB
XPxhqLoFjlmrTF8sBZGbENxHgZqwKOaOXa99JcKDwweBS0+4M6+qgWK3WqelMDys4dnYr1XP62LE
1UaU3xbBhWgmrqQvbSiRklCOwQjqK1x7swV5W/E+UMg1qDee0OMo2K0Br9eedDEB7b/WKO3Rfoww
c6eejctR+6hobHxmXg6VzDYWnAlO0/UTNNo0JGpQwBIY2o7yDSWmTexqzVsX15d/pdGXWyAwjIGj
hiVhRUiz0RmWC9/EvVG6UPSrHFkdS2weCmyzjeI0CfD2d/pHGpNu9RyxsluvxTnvpxzpajibtNXy
Fvc131yzYgt3kxzdQwAD35FEv/PID8ZRBjSu0iKmu202+LhNHEZfx8/g1OM70/Va8IxBNzsSJv9z
iWHzEIt2cnfHqYnQqBYJ9f5asj5eeGsB2Nrx+z/L0Bo6d4pIV58Ukt19nGiMrggTFTuvZs26IXUc
i1FNEGjnWxF5FrApBQiERG6YSTfYBr3bxLUTNE693DFy57fKtEFO1lw/Zb0hwHqdMtbiO1KWcZBL
9DHzbpMXc+ayyxIDG3leLD5j+pebrGmDqU5I4auLjPPfSmo7qhvfBh8bUo/w+aY21/m2dCVJbcsx
XWYRemCK/uTqyNPVzE7ODmPAMCH1Lcsglg1C73pLf0TAco24HWhA9I76zF9jQSJNzHT1EbFb1g4C
W5toXj3ht5Mxh0a69XevOrVJx8Su0i+pydhTQZz2oWdDcVv/NVXzqoVH6hGclfiIZeVc2RJjiHAA
WnmY1aCgMvmfF9kXW544S6O8lVUnBdvFpN/fjXQ6vIYMDrIaAzqBuXkOnLAU5rbWvw19Q35lJSV8
juU3b+bgXqm4POrZrbskLmnuS8gyXu3qqVvKuExBsnFHoHInJkzsvDEGyM+qw+DbM5k5J+Lsm+Mq
ZRLIk2e/Rx+6UDRKThLG6q3uNm/7rgqyJ8pERnunkbeCLmhMcwuS8Ws17SWpkV7vkj6AAHOr3DDc
z9yvNYHdCCH928WRqHybQgBjED5GdRO0sEFQfnDArGvOiWGkFTZrx/Z8qCMoIeAVNisZG19Jt70I
iWLfL1FbnOTDW4pmfjummiFQLokTT/Egli9bB/rQ1O+N+L415U6N5z1MCHZuQ1EFPV6vxU6NfLTE
n/7kxOCFtzZyOk6yfMnfsumnTJJ7vAo12I9I09HKKFsz6t6NPySyBh0XOwTZSTmCarw2BvbZE4gD
ILxj5MbMUoRK16mPJBc7LIXmDs5aJhxShV4FSNsYyrEguzTcPVkwS5Dfvnwxb7jsbkJBmlr/1XHw
idchiU+SROCGwjH2zYRA0edPTLfuLSbwsHp25vG/7R2ZYTj80Y1ppcgYbYcRTfXsPvUUd6olfw5k
dkah1NpqXgDgcze+wEOqPfLwF/m5jFI+lM/mAYu86wZFiX03pBp0H2cXRY9rkwZ1DjuNgi+JbrLU
s6Zafh2X7yCjZynfizwufGIpoP7+1LWWLTsa7f7Pdy3Hjms+AadMufD9fupA8LfGkvcfkZPrXt3h
RnQVQx0TU4sk9pvV1F3WyJ59IYxtugfWD1ly4YnC6KVOM9pjxtTDVTROS40JAm9TiG8VepDS1ryf
NtFDUB6le00ADHG/gcQeGYbhULfFZhr5J4ZVlYKAmLIlv54aRpDduubEW8zhaOchMQHniVJ6+8Te
StOyp9WcIURdj6uZIUsdXI7jmKJq7UtYT9lefA1bxPZdH43pMDl76mVOvmgpK7zJJSjOgKmzRKkE
IioxfSeyJ6QXI+Lj1YVFdZ6qIEO9IhouSrK44oDJVUe8Ssw2eKO97cvLffnOKH9eZTmEJn053C5+
NRoEwMeeXCuUB4SXMaPpS0eVo/aK3Nt96cIt2tQRrEpWAvS4g0S9y7XDZMayEPlQzAdg4E1u8XEa
db02ngj1TgeIQD14yPpe3yLfbnO19fii/0WOH91VxePfZIt2WgN//HyPbV1CN3hGRVeuQw0NcTM5
/E0f6qzzJQXpCQNHWTGVJmo+J88NTYL6RIRUnKkEmcqsfg61yIHHUXnG1MvuZyK4v/Jo5/OyX8qy
sSCpW2RIVs2yzoL9MEXncv7fCyipcPpZyOHqJuW6B42A7MYUM7F7r2pupRfripmCdY0O6KzX36ac
aCm0QvjCFTpYEhzlayBlQc6zOeLVt30YrKUscYmfnmuJ5sKEEVoT3HC95aWYNnMkYwUnfyBma3U8
ZXj+ru7a853B6FS5l0nagqZW/+yi4rS+yz62t7M9mn2OMlFfiwlcmpqeUKNZzfNkuI8puFuNhzei
pkbltDAxmRr+8aj4f+KzlOQt3VaDT6jU512sgtQXtydBtOdMiRALCBjPhK9UelrFiveWbSkgxDiw
wtww4htllHXdIAqA5cldvcjJ4bef0cKCgzu6/bvrbNdgD94bB1IIC1UXDOyItzr+inqLLwymCOGw
0dUW8jW52ZSBdrsvJzMKWYLd5TjJCxFb4BOcQfqWWq/f+syGgF7YvKIZV9/LNyX7eCOkBrA82FsC
Qkn8z7awBNip+TmjBfHV4wTZtMJLoc4KEnC4dfrX9uKAT40chdyCoSlaKxA/EzYxz/cLioV9wuXq
PF3WZD04MIvxDkUod1Kvrg3/phi2BIz15bB/SFQZNtPQeEfnyFjSenRigKDM2TvWKIbLPz2w83ON
aF6LLfLvX3XvY0p+fmV83v74a3lZ1Q9gYq7zjjOHMnRvAa3HL8p8Ul+p4q13V3RJ4XiB3Iiz7g0J
nSfIXfY0zsmrxg5K4f72u8dVC2kY6l/xoaAPzSt4l8t4K22V02KHNJjU1SMTuKySKJ7PdYQdEO5e
NRBpfor+3GMwjC0gXDXBLmejL17mwM8ISj2wplXfhMeIu3V7Z7tYB1MOOvl9Vy4cpaYEeBjfUL93
SDexGbeRsBlabjTnw0YF8jA+4UkerRa8yKSE2vB+NL/aJKAsqU/A7skVt9NeL0P3iVeZoFDz0CeA
xd70EzntjwjFTZT7iBrMcqzLymsQsnMg0Zgr4Xy5oNwzV9jfoySgX3Nq0eTfBUXh9iSaf7l3Zn32
nQBx0zlG+B8GdEXzesWMhYFiYb8bXS8Q42pt6zTIRa/UQmrEkp6MulA8kni15D96MEuxGFudGtbx
h+OLDnue5zffgpkBtMZcUhZvHUaKxnD5vTBJJ9U1BUSTI+xPw09nQ6KUgH9qbZJ7+VGekOJiqTZ0
6+b8hTa216CgPHfOwYLYsIwNVJSDfHaQMYrI7wPpWqB3UyssDrWdg5KHCgiQgouxjZA/g68YVfCi
Oa87XvztGp79MuEr+Pdawdz5VX4WO+lpuCUfVhykVWuRMwbmsw1j5miLTWe037dZIO2wxPmBtgPd
qs4NSPVhsziF5kq0LC4iPa3rO7gSE7CAbAZNHC0uvdmoevXVEIcx/E/AyZ02e/G0Muod4BPS20Xj
+LlegeWfzUc0blN8dD0N2q9Cy2gAoDjqEXcdM3V/3UQ25lK8xNeRVbIwUFhSuCqS1TEXYRQE+O5D
946Jp6kBG5BoyL3ZcfFYWEifxuvxxk2ZNJpubRSn8Ji8Su9Je/1Lejg4kudBulw72l9ta3Vmwjct
46ozrxdKUC9Fh4Hxg2jG9Dl+tTv9KgFWySwbZdpNapQ1JXhP8RcB7iC//pqc4IratE+YvyapTmc0
NKDLcTCcls4esjzFJIT3qDr94XD63dbgQncbFRNsxM/aQll2gHmDU3rNWNprhpU82DoHHaFcL1ZV
pfNV4v2QAera+Vx0WPK5ttbi+J6iYj42QJp931XNF+jaESKTqJXr8/CAdzcM3numIV1b8mVWZJ9E
Ol4sZuki3f0KHNCui9i0+k1DekohDeC1fpXOzWUunxD9oyF50Ug+SVRPF7pHQgbgPOFb0Vs9L28G
wNlhiPEld6/1opzIz0DN5+NDgnNByZtlQf/10r0Af69AV77Wl7NJ5ggQjOGwj3+ROIiEpFJsbfHY
JShZ3NXQpURqhXP9vHGS870tb/u0fVfy/cSb7C8OfUVOsNKnt/bd3obcM4s6nYpmG5ETOf/eVaK9
MB3CZT5ElSYBVwLj7eq5S/0GrAKpj7KyrczacOAZ/NwbqdGF3zw7b3YNwTbIgoGsBlmo9DektTtw
gBegnpANl7KNXBl3IiKSqhzxWyDSo0uyKan57RWVAB+K50S8MoaWnsZiTly5WLVXkGiohL+Bp7g1
SI1NfzzqreZtm92/1TdOQnr0sY+m+ZBI9X9CmrJBBdnyiN0rgRSmBRy9HtD7R8o9lfqOfx34zKMg
xzpi+FT7ZgwxnGuqm8qAck/bdnTBTpwkRJqEHrhzooew6VNlYDMrV1KONy0+HI1/0gZThyNe2++E
UtmkqVRbOkHQBFJOGsol+GWWW2H3p4a39qfZr/cASuHRwTteuyF1+c/kY+s8DCIf+ceuWYKVbD7X
p0ppDOuhOUHKkh3HRGLDT8IRJdPe1GJA/H1I+IOCppah5J235/JxI2zpYe9O56/gVygfU7LmeK4M
dWFtVZNKQPgwJiWGmL5ZtwI3y5Rj9S45y7HQj7tw4oiygjrxDhHMrArnHwVSOBYRByg6RRczuI1r
YB03361KofHFHLxxxIVM35S8JPByEmNvFYQJmOTZcebXA4ffaLSEcAKVOUAV0A4IHX/wXAbmGS11
88O1Vau5IQvIWB0AESLAxGkdB0tH4V9924BB68MnybKpNzeYYSJJK3y8D+kLcpnRrJ8vpyYukxNg
A/ADd2I02J/Al0Sh6Fm4Un96L6/mltVQD+offp8/To2WtGG6P2SbBUcrWbxf0Eopdm9NGYS5Kx2v
nyphAJPv/hdMUaJWXgFaKJVFdk6ylrk5sYNp4C7bVBsqz8IYFxIsXMLbfUTo9en3UAW0LmdjQly/
sQU5VNrZwDKOtF9vQccxaDuqJESPBSagEmnMLWRWEsY5ngOXmcG9DX6g/z712BvxkFgwYxSnHlZf
dI0raq4LaQPObuiNfTSL849y6Np3yRBLl5Kpxw62AZaYVhdx7W2L1RV5i3a3Xh9LeZHvOiBjsie5
ChoKlmXWDTdoR9kB8udhkiYCBqhY08Sg9gWCWYnSMHaIn0QMii9/yKH7wY5z93HV7wmGVnYuiEzE
f3u8e/4Z/UbmXNdyj+v+3MDCLi3qKMm6XEja/2ZUo7R5NSGGcu+WlEHJXcVu8zWXDnoJBDqqrGJb
lJXPVveOmbhJm4wmvhLleTWfcYqmbXTCfwC+TmL4kHXvtVVBqhGLzfqbBua9cbk1ZLppIH51ef6D
C6QH0HGKW9sefzZM020vUXGqFV+8D8Vw6/Tl48Rw1IXn/mc8XNpJWJnwpl030yEaemSVGifUph+R
gjFKqclzzay+Z5b8ESXP4Zcw9Tk4OvO7T6suof5Ikc4NygNG96E0AquPxpYEwu50eEQLoL1tVyqr
EyPbvsxqMdiyMBw5rFnF+KeZk6ihKEn5fcnCzWT92TKqpetfncEcKSv8lt2m6///D7B/I1atSJd7
TPT1VhVQBeQ8fCDJn/ON12V3Djw6mtWLA72i11K8oG3fwTr25vx6E46pxIARRhhYQCZ4i/8oIJXE
WdBwdfbnXNxEwh26IPgLWpNGB2ZNjpDLpNvbuoAuOC+/Sgq9sLCdEBh8H+5+ZoRw3nMg+1lx4cqv
Biy1yDPI+2QZ3a7pVW8hc4Qa3pevC1unEN0bR4tpwclWCJO1MDLSmbx6sTwOe2imML4VyXtYlUlO
k4z71JVN/5eFiv8Iu5FYL+dsVrSqlnZTKh96pt+9BcvQpmT0Pzv9RkB61CLJs4UleHGAA8/6Vybx
pdy1Bu90MrkJX/VGEL6ujQ6D3j5SUf3JxZbdi9pk0SPgZitLlla4XcuvMLEDHCXUOvTvt6K1tIQs
opFrA6+C8Lu4rsSHYbXVBACOh484d7YkR4fjXm3hFwvHnaYXI5y+vw8ptDdIzXh7kI1RbZf1eOeY
DXHF1gmCqKAHjPZaUaBpKIhbvtETiPcj0jSCLNjCs/YpF/YxyLg3VbqgBTZzl7UmlOwAEq8d19Q4
OP9gaL/adCFH9bzSi2zwTf3dfkg1XH51SGTC1nFwDFIgmMAsdZDu1Hrc4k0Wgma8l+rSxOgqNgWX
3MhJy2/f1Hrtib4IMIeXhSU4x7hjrETgR+61CoioGSaOVPLP5r2mrx5M4X5RLMD1Rx12YkKMlWaB
ySGFIR5kpsr8Rqy52109vKBIeOF597d/pJLT6nQ+Pk13csX+7xLfJxlYMGiM6oYAmdS/F55VBSa5
3ycrkDeexjgNK4/oDt0Ke+FLzlXXvaRKZYv9iOA7/pUiU9n2HpjlnELcxXOoWwU7IO1Yf7Uv2MLJ
LQbPUCB5vxIHmnWQyWO/nb0Zw3SYjQsa/CtVUxjEqdBTOnKYxcVaZUxgifwQFFAn2B/CMiyaZrWw
3enMzWHkoxCvQsqgOiKkbgpVnIrKfwzHR1Ntxj/dQa7ejXNvo2nDe1eDqZVEz4VcWvFDk3Mpafdw
rgUP7yIbhYCKCY4ftTSb0DV6XCogjNWInGF9la3GxavrRaqksmHtjTKAH4eqd4pI0fA3YtZcLHxM
zl9Wr3v2suFoDS3SZWcdLqg4eFQ+A1T4dY5NVwUmbMdIlcUX8LGOfX0HwsPpmMYR5Oj6tBn3bmAl
Wwrwrd7ZyLmS9omMesyWm2k1qQrKT4pmPvMbXzR/cHLIjv4VITC0DuzKowsKUxsWdOkNzenH7XVs
A3x+rkUUD0nlCELDnAaaM2wyiVqde2xelnznPNjMTNx7pbQggQtbzMiZWGflhj28g2g2Lq0qyrAh
gckN/MmugEdG3C54T+gXXPWQoYc/FJDvjk7QIglCEJOPJOdbrLIz+kCAy2+hi4A0F5NYFzKB3L9G
gC9cUppMUye02/aj+2ssudaNAs2/OwLT7OFk2+gkOFfLFyBCjtwanLFq//Bev8KScvreUSWe3pBG
8n2I7JxWn7zd3WDzEVTBqhd279Y9TonCYwFtivvBHSvSQXlheSvMiscs/DegUQ8+eRTKy4YmkzqD
43zabhXUKcU7ROCe2pKTa95xsztAemHYzSei8zMBfY8VMb4jTGuinaHcGuG8FWupVvDEw9UnfxBX
sbWwJJMg2HJPKQP7S+qyK4YNY+cGhgws5SYMwjGWwzj9JFaiD5NZB7bCE7BUzpaLKxTF3c6a8hWZ
KQjKksvrWr+XBS+hq0B/X1lyr4Bd87iOxVxIcHV+J8Es4IA0X+bhXt4qRQiIdj2v5Zcz5/lh0rkH
B8fd1eC3EOGJG5dcV/9Oh41CVT+RyjnytuFDoht5o4aRqBBxpSlItiFd0VACM0R7G4uPcVAjNtwE
JQBTfRNfSCNSj4zYGZGt5L8TdKuv2RUFZKkGSmV7QsTHefqZyEwXrrojUeIOY3t0cAsB5Zrm+STR
F/W01eUHZ14DbA+P7Z5PuOLr+hZFB4zSsNH53jHfcg4c4KXJlz1jm1TBm8VqtW1Bp/rjRthpYC8H
jARMxLfdIHbcEWpRRLY1QQiaf32BFa2dT+av8hRzuTd3iosSc0tm0/KWYDR00gWtMPsoayJzpFXP
iZgU+ykXHfbEGgh6p4bzhH2qijOmxknZYIuheKPQAYz+NOrtputGqWji7/+FbvvYov3bhhXcvhf3
ht4CWakoSTYvhXd3I0p+M3s0NXO3K6hYl+L9BpJVNP8OgxKN7UI8tUNdEhnXH3Cx7HsD+olMQ71u
8c6BNLsLlre3KOOBZQbWdazqV95SZqPQovNdPOCZFOPzanm7Jj1nxsAlady9nDdDDfuqQX9l76mG
V6+KqK1CObAByf8dq7KyQGHIGShUjDI0X5eaSIYrjHSXfk8dRpRWq1bD5DTOhgDnWDqqVVwsgBFq
7c/3C6QVFAoZ+wAV4O2lUI6lBgu4rU9WLISKMrdDYh4/U14PVLudRmBKXvYiLh1ihLcNcJR73P2K
QEfNdGMSfogQYUbQ4h25+s7DWxSMH44Y7YGqCD/P99gfDjAeM3Ts3zApqo5A5DtDrkhoO6dLBUzS
7nCNuXMEzH6HXZo9eXamJJtFIfemeEhoYQi1zw3MGaqE/07tj89eNqgVPQnDtMJzWlg+VFzsy1on
qUfEd7SzXKKONfV3IXD44DOA0xAn0iB7cQezg4wxfvlETF7BKx0gKfp91GW2IztXt/OoNaUC13wS
wro2kzorCmnOfauhLLXKDajS9pW/lxyDshexS+GZbivy2udr8UkxxThvAqRwEZxLPYwWCT953YlC
3CrmgUA3WN7nXAfndUsdiaIfLZrldvJDlFpKM+pVAu/754SCtkG6nzVkShnZLz9FeFQKKXhYYVBp
VDKm74KqZ0vvGTVW/mmX1mbuH9yEBaYzMo5LSBHJvQt/fErVLneokXZ6FMZINuXJaVjBTpLKSUHG
5GW0vSDc6ev45HcF8hwC96N7LcV0FapyPCAn41fTTUhuK/kiS3JdyKxBjkdx/JusrdepfnZ7awIt
FIvyK13OpTRdr8emY/1MzlV0w8bcklSTh/hla3Lu3+1mbJ7sELMiR5RbkYLcqEPBw+iaeBJFotF8
lc/IrlwLpCwx/1zvelQnlXI9NdC2pwypNaqeizpRU514BLyBcPwoKdGLSk5sGnmK3ocYXfAQV9i9
b3xzNRn6i8/OeghKjqJXM7YKTqrh3CK+d+RIULfgYP5JDlXdPW5DMZG5YvLKkrBQLc26egyS+1Kk
eRsD+Fe3ozaSrqfBXbPs5ZdLFmUZQUn6bR29sHLm0XFO8OcAUyQZA0OXOXcY14W1u8BIWdFaGvm2
3ri+23K7AmV5Cl/xKF2whmeLnbPARo5ubNoffut12HlvFeL2TcFAF1r9dkUCUV8XI1q5tqG0tPt/
E4Qi9FTseJQXySjk/SPhzSoIL/qUVhRxKrfIxaQrdbJ7MjwreDzjmdt7osIYI0whi94yfqGZC/dV
/xPF/4XMlOUhgf1wm7/1/hWV3lwJ38YbdBvEU2Yc7+27IwfOsYOroZLAMcBEQoh1DjlOctwSjqfT
D0qlJf14bvJv0yFVeoAfUymzmPIZs8Ko8aTwEgROu3Kg+2Dy+FOLa4zjnVL4LuH1rlEQasJw6WZd
auXCFK0p2rnojkzHS8hZ3SuNKEqu5lA6s5kKGkc8OgZ3v8PH6EWAa63u11CYntCfGL4kjd7P2Beo
m3sbbIsItFU2HU53lNjW7L4XAbVucZttf6nhvlWUpGYOtGNSxV6Zy6xpLXJsyae0jHyruiJeZl/5
efqnvvZCPM2tzl+nYSoQ+3dTN6bVV4PD2tYvAGoCV2e99RpwaKPdEvRH7Ig8veTGBSVJTBL1Ot4a
zr18pg9avYYQ49nmATvdO4XgNRovPUL2giKJJu2/xwQJfmUbfTM9H3Jwzq+LFYblrgLo+RHczpTW
pYMnAKllLr7bYnBlDllToZt5uTwTeZtuqdl/2e95B57Dv6PnO1V10S6/GuWfLQxkHbSjzCOmCKGx
LqwI9UUC4RDFIDqtYkxkuXunT3dU3BiN4hTjtm7T1JIDNBPFM3rOxY2VLdMkUBVa5P6YBqLMFQhQ
gQghFJusGkGsQ1M5MNSoovpjV3SWvA9TG4w/io9/OzdxI/V3UuCtj2l4k8FT8opk3UWFGvMeIuXO
E3xD5NRyLXd/V0e6ZU0elouEN3KRcFL/LUK14jlgfllNGnRQAOdmmdlw+/VlW/YYdiVnD8niBcqV
jjtxnceMENZ1hiRECV/2fMBS3Iv2b/JsQ3JEijXtRvjp33I06B4CiwMkudCp9Ahwzx53MY947Gq3
oDfiBwdnL/XBZdewpPCIxntPH41WXhOrgeMuORGSa7UNKr9m23yH7J0jKD/kBWwN/85JMfNRWjyp
JazrOA9qPAlsxdzA9dYibUUtxvPrywTki5AV6SctKZXne8e2GX5YOxjHUU/aD9kFRKJuuSsnvqJT
INcshJnuERlLP8CKqcdeHWa10fOmRQll1je+RRv94iAsuZsBe+4CBQwPTWVmx+7pEdDIV6KD6DHe
zJVOYPUvDDf7Q81qINFz2jksgCCZGsa7InVVqPKa3cfLaFM6pqmCueBSY0Jd1SO1eLIfnoYveKlO
vbx7FzzgDxTzcGnofB6zFOfTwTYfO59x6wImD6oV6kVX/5lm14N56DGKHgc6wNrhje/BOnaJ0I41
RmpXW2SEG4VYA/xXyG7tsC4AEf0+F5GPYFOMlmEwb1nKTlfuMWexkGuWnyM4IJUkyMufKFDPwrR1
dhT/e9a99kD9Rs2MuL2CNWrw+lWMqqrb5twtHwIXuQCCrzmJvquv71QC14piZUyDXZLsCMpQDtvd
mgR/++REhyw8FsMw3Aest+Ra4JQpIqnLEpwSeKgqigMeJB2GuOwJpq44MzQwKHtPqSn3tTg/VZcM
5ig3NIjZT6rv4PzK9J+j0cu6EEtULz8c2qpRJp96YorbIHVlQAIjz3nY8T+5lIIO4vpITjkSwVcA
B33dM3nPa2g9nkWAiS0JqS+xnmWyCKbfwzzcMXGs7Ucv5QyGQ86p8x9WkuDnzPTDY8ifgHvJXEhP
mCRyrrhHbFx8r7XkRsJyTHlgAWcy49u5FTO/dz8Qo2ZrRifPHuSH5wdnmJi942Q9ZLDhSznynOOb
oBStx3b3EUnhNfOFIxBK/tfv0iwcPcII+rZQ3Wychu0aZNIm2fE2FThtKJoRN47A/w2ELWzITi5Z
20USMBegWFpp5+2LQaxsxU8MlDN7bFiiz1uPpvtLFy5mdmYV51MeaqE8/m3Yxk9kEQa6onyPXZzr
R4pe5JDtosK5YpONsKKih3o+2KRKW7G1RYkY9Cfjz/w/6ccnezb4r6qgvfJFxMhCZfqIfAGasNnl
FlR/0gIaifzMgtHrvlizjrPFHvKzGquP+Ba/p2Qc7nrN1agG8FGRzJNZXtC7OwAbeNAab31qSaKI
0pMYIlCUlwL6bpHCp7VnPJbjP9YJ2t+U1q5GzSy6ekHRxyObSU2MsL5NA1yME/M1/+3bdwAEUbJS
XhtxcxzaLAOltZTaMl/LiB7wG/Nue42snvuNs0M4pwG5vWN90IKf0QTaEq1XQ/vEb7HFo3nFssov
p66H/abgn70ZzIYuFvKQEUayK9sFI/bTgVR1gtQ9HZ7UQaTmDa0mh9R0AYkUKOtDH+l1y8ivxeUU
/fLxgXSdCwSHPalPKHSPv2PA7w+3LCwVJwoGb7sqA9YGT1KYnZ2OAM4dt5PJOyzNj949cgT5pQkn
vDvk/tld1YMmj5tSjCQdrvFWymYM1OqRrNB+eV2sFj0pK5Sw0BOENK/eCeI4dbOV6okI+jAPv3gv
PhEoP5cHrkmz7IRtFkNT7GZM39xdS9Z5zHd1+/m8byJJJx29NnHtCzh1+INKZLx8csEFNzzatEUu
tebTZ7ewQy6s8Np076GhylY2FR9YhEanraB0ClV66uDB6lr47gL3Yj18fbxoAODEcx/3s242INHr
BLUb4ESeo0sjrbwBIGovo4yE9Nko0fxxRVrcV6KAN4CkoVHSv6hElzTqmDEQoXLxCHfRAO8TZBlv
04Gx24MtWK9ICs33anvCbbUm5O1EojokNfA9xTriajWeVi4jT4UHKLFuFfZS5kuE4D3cD5IPyisp
UzHa/2C0Y9IiT69P1qRCnx74lS6vs5nwGN0TkNycXvrhvv93N1UdF3XTLS+xunTELXMWCzxmBQq0
JXjNN6R8cE1X4rDrKhXcMsMWD+yyTbMpR+RwYipYPA3mtsATfBC5AgBsLLJsyWvIEqdXJa8IQdl/
x5KakpH7KBS2xBs3f3Lf41QQEjTQh7vaYA//ChJWQce8m7nWyjWsLMwsvA7N8Ezcd195+gZwoOuD
XWfKcOYE1CiyG0L/om9ySTW1YKVurCU3FKyaYbHH7hAKQ1OA7dcR3Ww1zd3A3l82adVBgdJ8YOOC
Q6ME2Xu+4XFkOTjzu4i3RJqsqyYRLY/KtFUlGn27sZZOJXdaUo1mLjlVVPjxFJYOjU5eBPfxZ6Ze
f60DK/4ze5tXz+X1HpL6FSDMfsjHj4V4UYZhNHnhuU4IdbJjw1a71TAQxRsVu8cpckoDKRIPAE8b
spRKzIEXX+6HcmQDLkPqBzUL2WsbGEOqcF87kYGGUIy5qIEF89D5622eDhzcpwMJSLoFrCNWx6/S
Dhe5Lbq09hFzzNwMdIzHrSJ8hSnPIKXF0Ag9+lybl5AOiDHHh80roP+gEOaK60qUjZyMpPfCH7W2
/pEsaNnLo+SliFAa99kECjrA0ZTFReLj1+tn2q/GRtHmFRKuhO+YcvoMzVagduy9N2yg8kn7lktg
iBfsoh3VSWr+dePDSD49WsA/aVOagOOKjjs51x690RFAdKKsocW0z24Oq9j4WugYJGpDOEU6wGxD
KQzTJUZC/AzYSWCku0JXVCtR7n8KWGDC5GA9d2RjmzPChyzPOHf29jK1BzRGBd4HCotMmE0sDH0a
n+Xcgn8+bCr62O0zbcJUwFyZ2OndxFV7n8V4oCkcIZkvxacvxCMUS7SWuXNYJQ5px/fNfn3tw6Yg
4Bx7/vMeaX5n4P3NypM2N31aSvc2d3nJwgmza8CFcjigCKTp4yEO//oFNQ+JSDmO+qcCSeY/MNh5
qCO7ML96bM8rwzrMrxSx72/zNjFOsI6iCYMqrX0QqoYZYHtvbBfc5ObqvJDKymw2RUITS6yKKI0v
4NdmNVuMx+X5xpyDeGB9vtesF5qz2mKbvCuuh1mLkgQMhtYKcoqfq0RnTFhtT9/f/JKSOot1zg3o
cmjFwQ3Rrj/bYQXEwrpo5D5iBVj7iwkqFHVzP5e+pE2jEBtrQYniEMsGmOnaa070PdtAm8fZ1LvN
KneeVTXD4/XREokCuiOsFlFVCLi/IG+1z1WyiubdP3wHEiwYjiVUT3s+iWOuheg8FDdB5TXDTSXC
AHWjAHxpiOScGg6DupkDaU/ItTXKZlKPv7AgNkBtzwqMPsqiRBoCzGtjmp+FaAOVwOfsXs/ecVZc
BwXxs3JJSd80pTryDruDRureSncjTfnd+00WQNMCCtvEvIti6Q2B47Z945Hl3zglllxf+14cbAJd
ffpy7GVpgeYpu26E4/dLT61wcmn6cxUff4X3ljWpCr5AWDE4nXvy83s6qSwTK2FjjrB1QAnZn11W
OM8M7qdeTc9/4GT0VSZuCOlvEFlsq9uM3HfOHPOimM6PFjT5W/U3V1xJBTI4sJ9geJBFtFR7vTv2
E85pTRrc+Z0MLlLC/7lYYLhrcHPhkIxyneduTfCLqfZc1XmBmaZEm+dexKLBXphxTD1xGajOI6cP
z5AiFe17pzaehB09QHi5bdTc4JKMLIFhHU8Xx90DZMD1qDAnhymI2uuqTpKb4i1V86rb+OVXSmfy
KmucvcnEpDaIz2SmCdte1zQ73oWxUqmn2z/lO71gktIxAFGRtQqqfY5QyLCJC12jzRr2BViJvejB
1mv6f4L0FiAUopTmH4RcUZCaEIkFAl9HwZXEpWaiY761fewYn0yvGOVjry0oWitj2f+p2n83DzNz
WLM9nzUsbPu1bhOia9qsdn460uPhtoqiSz4lsRjBafImMYIusBk3ZfMuolG0TUL6BzELjfAnbgEC
YW6rBfYp8AJ5gTegBUi98UxF/uEw+OPeBhJc4/4EUUO6+RYYmHkN6bzQ0aMAKeKjKYWEIVvyVuAQ
wjHgTFoYlDs7+L5vy9fyohIapqCOK2sGAdE8WvqiJl9JUcqwwTmZkU9KbeBnQcqgUGZDmtCFz6cj
mNXCXEeAYgaFln2FgY9JneJDP5XJDVlCtdSi7j0NdJIvSIhHFXEFTB1O52kluaGKFmz9kSyKXHDM
6HuwqY5VKfZ/zWogpXbicTn8vVZXEJz6w1fFFJL11a7GbY3C8IYDFAY55t+fizrPsKHJ4yrd7bMk
0NWCTe6BrIbmncmmxlQxomYsdEz0JSp7vNqIB/gp8zuYrLA1LXBKebKwRv68+9EVPeczf9lA+j8A
rC5tl8w/bRTLDx4bNNkPpzSn8QpcjjhD/J1aHKWt/tH7DBnv8QLYsTPSGJu5yg6DAUkt1ZBswiIM
xA04Xr/mf0k4H3d72X5k1p6yQ5OkAzY6LcCpdnchqrIpjsEOO/Ky0YBymIozVqm9F9/2aylpf2Nd
PndoPl89v4uq/wRsRT5uT/F1fC2es5+wUejHDmjSCc6MhLn2SGgiAH49xXl9WSKJFipA8+Go3epf
SQC6ikK+FFNiqMVCfonXGvaGvWTw5BPU/lxoCRLj1kj+Nu/Aro3RF3tf26xoTIYFewzGX7i4zOyN
4km9+OpQU7rNSbQUtuHpYWhTm4Nx+qqluxstVU9AaHLAnxniMtUPOOkBHERwrSf5xFUKokXxRYPu
YcWHu8/q/DkSQSV+4ZpPILh9gZlJ3/u7KqUGclk5za8yWkH/CUlS0AYTRa7gV7u24/4UnqX6esbI
GW6E7cgUaQu7JAZtwZcXl8jMUG5h5URS90+B+SfsGi2cfZcsRDsaXO2cCwmRjQl+iE7il+IXNH3+
MfDz9LWuGcOWr33MSBikQiwV21WWLL0kwgPKMvpEoGbzC1eaKgcv2of1q4zlNnsxfX6TobENlFMi
uHBywt9qeKo8S9eo3rKHhamKdmoWdXJL6/ccM6mv7vbCyeVUky0KIGdObJUzbppZ0ppA9d67fvU4
ZqJencawUj3jpPBIh1Ny9Sn7pcMFrTj1YsPYMkky0uYz3m+kDPPGzw6oZo88/xOIOEyXDTQ0JjUV
jqzhDNeT5e6M56Ji7epRTD0CCGunslvuOg2KUgHFpA9EEmkjOlNa0jQYKx7L7cxG0ms/JERw6q5I
pHNEF7gkfJ6TdV+WRWFp8aaP+i2r2OsHEB3r/OMKeHgNNOA7VsXh7mni1jfiBM4KxUxZ5IXa9b1E
UCN0EEwD/p497L8KHzBetW0RQlGqm+X6YO025Ct3vFktFD2/XUvOmB4RiFAs3chq7QOjMCIp5ig2
Qshhdvxoj8lLer71i50zuDsiTVedmbXPkFmWMIOYAu+MAR1ujTXbTe0G4uPNd/VEPICQITK0NNTD
jcQ28KWjzA7rgibuSlflE6PacIi9JYvavgOBGOsyX3cBEkhk/n+LBEVk7/T/OHu0eOjkmPp9l5wE
NqYJAsGVk8IM9KTs1MtvVVumWcQKm9rAS6XaQo9XnOFtdsvMoeWgi2B3xX+tYR+CT6k5KmmlWyrb
y23gmyQgY0bjfpR23SOdckSgpAdOeV1OZyjJCqC7agomN/aeU3iWSlTmQ10We6JLHgtDgBOmFBtP
ywAvv8ATckiSz1+0gK94JUTykcbAHFT+lU5LpdHtibBcEZf/0Zglm1QBJjkBEfUx7BdB1ZPFlbbc
8Mamk50xXpNf9/Q2PiEzLq0YmYLkyq3UciCwH5gIQxp/s2w/lOr2tR7sfBJaMLlr2KkQs+2TkXBL
0k9IDpwsJCdDxEJGs0FJSpFuJVTPiW+4EUlbK7U5xqyGs7O1ovT20i6Sx53PgSY6r9Iuamq2eAOv
MOC1vmnJErZ/JrD84s9zkC+r0GY+iEOb+F7J1iBJ7+v6m0QQDtf1JDvoRfPdM0pPVXGFhfLrTa12
PYTgmcCMfjhSk7mflspGo9qEj70Dh/Uf26rJqdg9HQlN2oblnHZgH7+z5YuZG+X+pKD1QNhjnXtJ
Ud9UK/4eulK0R3a5SKDSjzFWTrCIwWW2ohqahYPaNA3cR5ReDm6YMOwffG8JjnE+f3mSVcGtIW/N
2bS7PknQYYLrO1vgsRsdcz8EQ4IwPDQ6ZbiYJotOe9aN24YElJnyI4oo227aqCNNbJ9On4MfnSio
WfrveDJUf9yIjz8tgW/Oz376tUjTl+giAtbROu3QfwsUNGapp4IXB3X/ZWpPnrsH09OtWCBlxB26
wOdeakwqxRCuU4YNe8FRv5lTPIukuNNL9PPDSSI3fIDVa7p+zJKugDPzeVGn43+xWuTW0oH4MAy9
FCyECBrAtfQkk4kMc5/htt9yEP7fBfA7w6qxmqrsfxWkZSSKXoG5Judy/SRwqXDLDiApseOUvIZD
Pwh/+nMjCgRNxfsITbbgM9KoYbEdoBbBtGJfjyUJGByaXUeBbkhYqkIGWzAFAhpgYOoZgocmSVf1
Plfi1Xgzn7LQClGs0kwN7fPdJpdNnsk4Oojfd8YqN+zxhUBR1NXRtbQkU/euszhuXtZTH5Ogb9dg
8BHrAAQRcOHO9o5C6Zfaw2YvPwcZFvP4SmLunfbZH/VLnMw/yg+drgr37HfkDDyxbDwXVM3mc8Sq
GXm38VYMlrxDsIvLnJlIJUpwTw8TL3J1gI3jMO6DpZKLRyoYMPeeZi0FMNDlENhP89knI4aOV0Un
1uBSEXnyO5du0nzeCPAr9UYXrF6gZO5r7ln1kcE8LXL988pTyUPo7Z8EtWay2iBfZoYdzo3E4PGG
bzPJ8OylmjdmDFwefZ1xT1eL9MruJfTa4hd6ArCBZJhDezEhUgOStAPPmrNNnTWJ0w3U1Aji/HFM
OOtK8Bx22fMgRmVF1+HrBX3R+FoL3fgEPHEA2kGvGmbBY43AVsLof3nE2IXvHnFQfrrju9Dy37dk
9ms1VonF2OiDdSV2TEKZpiqKkK30c2mkwAl7xFGoObtRHXt0noqwLrrBnyhf/lUyXv1/4VXjj/09
aDtknFHK98B+vwgtsEaPAINZyM8y57+d2ds38q2YLrOuPrMtki9BVOWgDot2Nx8NIWqK5WLvGoeh
kRmqWhgAyyKPL7YseabMvqK2WVS0K9UaCnSS7SwrTMo1gtHyANoh6VCoXv8zyedVdmquO6qR5cOI
5qn9wGcCo/6esh2ur3pBzYsImqsxHAxBTjwi2GpWuX4xSXc02/f23fTkIFDNNTyopjxFBotFAiJ4
GDXfwt4zfdD4P+XYXNLfBcHAvcficUp4648T2a9YmShdOV2YdNAGlJjUW7DKsx6mFMADCrD7h7Ie
a8vM1bgyrWW/1GSJZ4UIS55ACEiZ0Pxf97PbhGMTGqK2Oupxedz3Bgnw/t4oYvrTrkuwu7J37EaG
i+y+5n+Y1Tsu5KvQhHplv48nE3uAQJHibpk1fd7xeX8OJiYYiloLCQlC/DyDgMw7DcCN8KE5LWaA
vN+t6gIdDP7d15h6y0LoW2bXg9mtsbFCcrsQ8XLjQTju5b5zE5yUJh9xmQx3aLJoW6qRaj1r7Rhv
+2XYgYuBmZXLW2NVvNmqgmFTTI5Wz8Sd8rchhzKGiIIcxi3mwHiPanljFyhFdj9914KLsdNN5xPA
3IklHZ8fU4Xhkp+sciveoGxRkVuVS+tGp5xOqnAboCxZMoMwRKX8TQzDZzUgeItdwpZuhPlTp4Jt
bszPPsAVR5TpmR99kqbpm65isxc3JbEjzolz9fRp0bb2q7dxAIiqe0LeoHbSZoORPO31i1fdw0NG
FVi3ghpbyt4zpmTQQRRecSpOynHW6IPBwsAfUUFAX9c2UqD0Xxi+qirBDKVmzlz0cuKuF1DCGo4D
1km2tVGaqUXZ9PqlTDN/3/LIkzkOOePJ7CZpS5m+SltetlCxTjNVMawpO4Vf4k0oo+1mgVkbN92w
PsQYGVnDRjQz+lgx0py/BOlv1OOgS8V0RBgQhbCv+8C/6OkFZhNPLPGfEEvEHIpLcv2gGf4bV5+0
3rS5jNFRLx7R234ApplXzq/0r0a5TKaNdj7HlvAmr/CXeciRGCWD8kudCCNj74/Ns1uc9jmwQKQu
3/OvQa49lpdCuvC0+NOL6s99OlrE2r1poK1r2Bc3GHcgfxjH1qKxiWCwroWzhZL8VA92FizQ3uIy
PpOJ1MzRXwFs8KKLWPPh0IeDdirjzoyHYwcpkzCsSJtNfXJwADAA7/zGPv10HIVqyAGJ1OR/Z6RL
TpXuc5YoCfhZpKEqFlLeTuYHHB3QOLWRZrMxRb9Iai2WPPQQhEWKEmKXqwHduKcMlhSm5vsCR5pC
AFZ1Zum3nmBWdq2rDbzugBSsIWrje4J1UWAWLVQJrJisbKCD3Fe1rlykOqDSd08NLM1dL+FRgAQD
ffH7yXI3FvT8vR7bh0x4AfSghUPoPiYYc9QKmpjgGGbP8fv/Uhw3QcqMQZj89tbc4IwsHShPZ7SR
0/ySwygCYXoil9ZoU4bL2zuD83t6azAinuEOx1P93N2xTmLNfhdm1N5SMgP/DW4j0R0Pji+uTjE3
XAFFq4OeoWIHmydwqpz93MvxEKnr1gWBDSYhQ5R9npa0eEAhgoAd5CP+d51EcFbtnawl86A54i0V
ExTy8NgcsBYMUzgtQBSqaNXxP4N14o6S5Xwmxb/92V8E9e37PAssPse/kD+33q/sy9YTgkKzWd0v
c2hBL9YkO8rQyZCzWysE4IOakp68LGBMXKxuNPhHlaUmUOmdcF+DYMB+sj5eFVd8KgLA3ZiKZXxA
z3UF7f/Yulqp/OsD2kRP34r8x0re96wIYXSbCHHacGmQMf3T0bJwzjoDmjr1a4OYulyhtCIpvkLV
BJyFwLjFJR54EQf0fFT9NRDpfdZaENk3ZcnFzMut9kCBw1FJIOq6yKlVZ5IP53/0a3i9ptceS9y8
BIRyS1PISC/oFgH9CkCZc+FH84nPfa7qq05ascwyLSv4EBWXUocypaotFPyCJ5l//vFPbI5xpPF/
n3M0K5KYpbB2zGSaPnro5BrJMjhl8DFKsXQmkRCtOIJPoRUKf4VIXnODP9utLkwg67CdvLHYZgTl
RxR9f6b/uKmAjnSQxWVMo+TMiNWjQlGCNhUoGOp6Db+FxU+b+k8ICzwXtJ+8do0fBnW+nRwgELVP
CaZpW6m3twCN8LtzvmsjZYNZ2EkVfzycsVBaV1qGAmz8gy6bPcglBQQDi3mNHYu0qF/J/RTqE4jW
XB/ORlu9jjk8K+qjFNtxICgfGK5VBRN0pj6/IKKlbqD0WHvthGPu2uwHc5mwqYeT4hv/bfH+MHJ8
Fm+a4W86r20gHeX5yVFPdjuWHPOceu2AIOhka0dQNv2r/+2iWY9wGFAhfWIGCPeJlaYgvcaUWS4G
7GW69JtB4apSZI5lEC3venspdZr4PjGTXUjhiGHi3M2zYG0p56aSB47oDZDARjOIM53EhG4GenNK
U+iblC3Xb3bl9TycUUI84/hK8dQur7ZbfygHyCs1f8UZ14p8LMsx9UzOYRYEkLo1ubki8KProZ5J
iwXLM4IBr5rxcxBZy8RBiJLh+o6A+FI40jw5xFS1mckK2beUc4m2ZW30mGqoe71jNLjFE2WMVBQ4
B7l89csydU7H5dBWiRC9GOIvRmyUpEO0HsPm52j1cdUbU7kmbBHHYESa3mjGSWm8/pGYFPwFAGY5
E5d36zUDEQ6T3h1ePtFvqKFTGZdCFlSWZe+ldO6oM2FqWjo3X6pcdD0KFI0wJhhqRfBagjOHygFj
B3IFk4E+UgmxekWcRRzn4e1N9EbS5nYCgsdgpyoaQeLECOEkWEwXHcNRIEK2EIvrU0KvejxTynqD
6c+E+gXSg7zzax1iGODsyWv7/0xXxNQCtp/ImYOpacPzv5+6fKt9hLycRvA5SUmBA5JgVL3QrLwF
ZX3Wa+Wu/DprdsqB+JyLRWRNkrRvq8p9BD2fYev5s7RLDVELxDpKIy9JlP9dmntWKai3DeBUA0h0
88Pdlqp+iZ1zqdz0OMDwwDPFOPYF2RpgHNfsY3zqm++ENoVmGuTfrK6I05udo8TxiP1PXIpvJNFU
+2T3UXtLsi4kap9IWLYH4M6iaeCq7qGkBLancBlf3C1vGLtat9UtBzmkqy9MjtIZDdUH4AeK36Nx
M94Ca9Qc3mw56q9VnttlF5rU9T5Zv02bIuClsk9EbNR+BIfGL5satHCp+VEjrR9TIQftCvCWU80X
/PH2c8moaKQtqy2Pvpmf7STIUzHXw15kA3bM5gujkoWtMqxADIb2zC0xEjfnIN+txeEQTWNZ7jvM
Z7c6xA9g6EtSQ5v9O8V8iAoDH0X/GMjCfwlj3cxZIse/pZfbhF/P20kEfKdac6QuDtbncWsH9NRz
ozaYPzpJ3IRgJNUn0+kIWXJmOarllGGv0Ec8vxHT/xahuDL0jYgixDxWqjNKFgqxkgKwihXUilL2
wu0rQUwfzs83RVvSIc/B+jGxVTrhIObGEIrjYkVLxf45bWPzPgb05hTvRGefvwkEAe6ruXMtxaJs
plecwQGq6yZ1E6ZZz+AgU1fN4Ol/UKXoUbivZ/OzZ0OycYLxAUS+AFJvLUDXlrWxHrxtJ04Co6SV
xKfOrfD4YmmBv/s/LaCc5jLLXnnGaionq7wM9hfsoFzBdBPa8UyXHOVCgLVX5X5q1T70i1UgeeqS
ml8KMV+S+qNX83F8/GECcAIR5CIp5VWvsua/222i+R6tqlihKyJrM/kZ6YiSHEgsFugRpScmVyDf
3C/Qeai8nL5qCgQyq34GZYe3Iuzu0s0gnmlQBtcy2HfzhJJCeWakNtLmQ68pfLdQ7PbWYgjaDqZb
xdzG9Yk/XKz44ZHsB82mnYyrkNQ/YCopkFvwjSw2LvT+RSpdLjOveFMgs08jYAR+7HRHj3qyEGy5
WJS18l2bvf6I+uYtEd/3e2z0Dg3Gx1PXJKNmmhjRiWSFVZyr76lwTl8ZsgDuH2VtVHxxWhgD+JXT
fD5qKZrVbFZECerXi7MPVaYPoyitCjTKzGODbPjdFxx1su6agt75wsYPwlnwRnvgil4GVUvz5Ptq
xg8qqD/cx/3as6rPhxBKETmgkz4qg6dlANgFTjIAHXPZVCxCRAfz9P/F9QZK9KFixhi8h840s5MV
JKOHPbw60iY7HvbfniwqiAWDZHDb9dophKKpPL3KwMNL9AxQyLkSTxlHDZdbjrN3VUjK4cD73pQg
rIyYEEh9dMdqHcgasBDbGUW/xdw9ZrGPg5d/hZFBFfs0UPR5MevpzhA93MRreGkUK6Nb6EcRSknL
yy3EKAvgpz65ekWn9l3VqQDNSx6xJ9v8q7juzHbPjiVXZrhGTRJP/3TLSszPZAx+9jfGAQcIQ2m/
RZT3CkRIWQ72tddeFinFoTmWQZID166WBe0r/bhA+HMEWOPepUcixPEXgfeVvvi7+SGt/MMgI4fX
HKMHRjGtcav3ojcibjnt1V7iSCUOTZBcrQinUuFzQg8TLuM2x8IJS3Egs3wBtV3Op5H9+VnlBYdj
IVOhm6I7tI6vn2v7tuy55AjSKgGtTxuvbhMRDwDWnF6Wb+YcZve7PLXFoHHX2zpP85fd3g7MxqoF
fUwHFL6pLq+elOozYUwPbpFkSbh9aqh017sRamgHRdbGqoRJ/GpeEVGe+HyHCGkyyWg1dIHZPBEo
CFh130Yq4pFXwtewwDpFqpOBvLi3C3HDxAOWNO5hGYLdS94+N5aQ0HHNO60r6Qw+af2VixThYe83
Ii1AGhFRHuljHY0Xixt8FQERt9pUnOcXNukhU+Hw68WFJLIndnwoNp2NWPoDBA9DgzeLA2Mog2ZX
r9AJKpqn2U7oSsyd/6M12Kx7rLoX6hppefKfek4Gh4k8m4rAyLVW4F/F8907jTw62zYWQI4aezZs
Na+7ZAuKreXwbcJJ99qoWqvt3poP76/DlnWTqvnCzLPFdHh/+wuVUGnXySMK8JlzAc5hWaf65v2g
DsYHANtCoWEGr+JMmndDiAKtOI/1h7uRI8NG14qdchsjvFZWg7TpdqT++0iIIzIZfdtf2xDgKtEO
wi8TVtdcDnygYFSIH/MhAZEkRtcm78Re6F/Ch6sdNK3+h0Cd8963Y/5Dk8RmI6vO4pNrJNoLaww2
KGb/i0H8mULeEXQNudaoJoJKS38Fa83ew4DwVYrMaoPyXNxV+O3a5Q+vtrzeDdmPP54JWOdRwwkk
yHNT5URzuEIrvTdRjC/ny9YN6uzlR6xNOcn1r/F12m0T8INJJeSf3s9Rg74pTC+kcxCtZJ1dveOx
qFCUgfHTGvJOsKqwu3bZREPAOmPrt/UPeFNIOe7u/Q3EqfggU65gx9CrAh4iWk39O5LNPuN4jAv5
aSAUCh8cnOT2DawOwGA2aIMT8zG0WPYXXS4VQbEip91CsnCueyGsCt/ZOtzsDKqKY0Pf7LirAtJn
+VdDSkQur9j14qL8vxHnktRAtm8G9NQTuhoSq6FHb6b1u+8tEw7ehh8XSfK9/FspAbO9wyGAl3gC
XIj1E9YgOFT5O3UEvwylRKrgTxsjG3a7D52Gf1g/+J90fkxTGKIgkKTu5II3ZLpum394jXjMqtP2
pP+8lOJyb0vRvtsLS3Bs/FQnpflRoGBrbSOZCG1YJYv6orrqE64e3k0rcVAGx9CcMUioNYHOqThT
2IBR47E5s9IUTXW6Qixf+RSJ5g+ZUrNghqPN95J4FYy3fZ1VZcJRGrlKPsVpkB+n0tbJj+1jIlLS
A35Kna4R8a3AQEv5XM4fNmN0BuN+DUfCO1myA+LS0dxwuC0SLymVcB/mH2+fqUwC9lJdTklmrh4v
pC3TDPFRdLQshHBBhH829p7aRCKzSYsgrDDWR+kgixAqBK2YuQR0oCmNID6k/NkgTBjU/xmaHwmv
z9ivuB5ojAvPT/yaU4CCEhEJO1nVRYdnDMl5liPBoQZ41qPwscixzMLO0pLWvUv2mlv30Hbavg4V
qZuPMRTSxzV4UiDOB87GTroNCyqoGCZ18rbmzSM8shBJLToA0/Yst+9RMIW45LOv06t8kPARip+w
W61M5zoy8XKfm/8WRa80qk19dIPzjjpsA6vs4kHHlc7lg5S5oykxaPi1ow3Y9ZC0HaNZ6suZnwUG
W/2pjE/Ynrl+f9twJoiZHusG319py3hPeTWd+2Y0xr2TbyYVFXj69vKIGHWVsEklJU+NYy/yrzTZ
2qQJrs3QqrqwMZmQMOaHngU3Uu/BX0OFO7JGnpr1+yWh/6OPbI+agQbauCwDFod5gaQIe2RjhBBB
A9zyyyukXxQAGr6olV/Js7q3ukxzhC1QAgVGbLn3LKCYw9BvMLjkWzgMgIjN+O1bwXKusY4nbBxh
u7D+RwgXF8iEv0insdVijhcicj3mVGLXb269WCl+fbyEm872m2d2gkwq+c/T3IAE771aICMTjpDw
RxFXZTrbPX0skMR6N0nbNyUd8VG7qy6Ra2D2VWiV3jihtus1va3EhQo78CGrHPsXn73jeBQro/Yv
b7dtA144J+5hXE+q0345KBegOlYkljD/v02qBqQKG5UTWUbAdJULLUrcVC+Vr689VArkVLlDoV+5
5qfpUE1yLefOkldSBliuCGRf73F2j8Ol6T7lLQ1lnYAmHB6BJVHu3WKGIsQLAE0hb00NuXRsF5O/
4dElKwQG/c1yW+k0eHIWy4fWH84izM7jZIoMje1h5/xITATd/Xal0LsE6uxXBVhP7MBlaWUS3NAT
neMnNCQZyFNlSCtTV/JpSjZNUiXOBnVzum4tzKHNnulL8GwE9N9LOR6DnqY6XQoB1zZ/ls20j0O8
tfhMzXHMwxTs3j/MmEseVE1JZ9N1FHIDk6FC/s8jqJMyf4UWnqVJ4WMuHCcYVVJBaeEMGIfMT4qG
nMzoBfmxjyV8905+Pt4WAuxz/IDNgCXkezYdtQaDJo4qW3JvVdMp1lqRw/uIw+6KJ0f3G4As6S5p
MMkUQvI964EBScUn2HwmT4BvO42BVWX0Zov9eKP5oSSuEH2aGXRoGSxHIiaL0cZJ6sjQmSBkTY5g
VoY8nDjyQq5kbqH/HUToALJR6pl7AySxPBvSsZ9UMUq87hSvWF/uOzp4WFMe/a7c5nOUYi9jTY4+
aM4KTrQuQ+x690dYK2nFVTqBrQA1DJdoifDANchcTSq+3YQnm5raVrDWWuMUeCLG7+aGkrUwE71O
zsxLKgCeSnMd1qgOzCkEdNA6U+uSKjeVovHHVUECDGqI+8DcGO+u3IAlG0iJQiw0H0rN1pzYI+KF
MCh1lXWWL7r//nfJ/UjUuSNdXS3xKsPCI8DRimHcXiZFXrc3xWfchZPkjp1LpQi9EYMF5N2NkIMn
JgTX0l+uUypXljhf4+4fKNlfesHxgP3BSfsNn0KCXwxg/B3rRW9vhCHA/DUYp5KVs8vIpj7AQC3e
6GPGbb3cwSHSXSRm340kiXEwJTeslB+IC2WbA8MlZ7ZJlZaUKGjSdAtsJKzR5Fw/tVVtU38bF9TZ
hpDI7CAwNc+tJXKvUBV6fKNndmQQAPrprO+uzW4yRUbZ2kyjqo5W2zMlx+vEhLh1bymNcnG+if6R
AhCBEmYISOip48iBpUYGrAHjLhpJRvcPMuIrMnFtRAmLo+9gFRcJZbYbigC3HPReZRWlD/OIbdIR
kDbBRISxajMUsXWMpcP+gYSQJ9/e8RNzIjscyTo8zzhyl7C4tMRkb5cmNGfOPCvIjcp5uZSOyNGK
b98mK3sluB+K+0+eGQOwhfLhuaSsNlnYfEUU2UqzwDEvubBlfyqlkbnsJxtB6LF+j1roxXj/lObF
k1PS0BQ0oLhdSsE+aq5JtW/7jAVrH3Iqh2KKws+2+FcfNkgcvkjvOJxrRt0Hs9M94yeBWE+T+Nne
1RKoWqD8ppLO5EQHE+pQgmYOJdfEDeJGNd3Ks3mH2wQ3T4uKe5ONleyml0sv/MgwdHEcQoyLBowf
JU85RXmvK3cDVO3Y42uSF2Jk26jbaCNMeIORn+Y6MGVpUwtnEZTxAGkM31kuu2A4p2/McOhm3+zS
CBd7cM6YXuXeL54708Fn29PYu6M9qAwrqRXRnkNcVbXyuhcCWSOQZkvmgFvFBYt2lVqZFTzdtMdL
AKWTin12HycgGBZv+5wmgjBsIXREq5da4h2ZWoPtIIwbfaeU/i85TQGtVZEgz8/naaFr2luDQdFt
rNG6jK/wlZDaNe4jOtu7TaQEBSlZqYRiAU/qaA/jEB+HSk/OEwh6j7PKRXDnblUICZGWFgrwSVQ2
RFWIiUXYqNA0FIopPKEGO87Gk7Zecjq5RvuGGbUsd3rVkAv8TcJJeggu2Ly3V+zULV5/7wklW3Y4
rMgfpdhgcH5WJHCiq00qTgLcuNkqRr10HyDIQIc8pwBM4+f+l3TrMXxtPhzH5qYhZ/dDWSUFRLM+
3mErcwA2aV70dxsrBsWOm7yLxWEyLdoaX75XAEGaHzOqwauEUhRMPUDiRbRf1UUC6PH4QchewSO/
HAajTnO/Qc2h2Zs2SZgX5gvwX5lUpRZznB1LUXGto5eNtJ84eOSWsw9vyap/dCDveasXNQWlZtLG
x29FDCcZV9ZdNK/d1lXVfy5i9hT7/SIiC7JE+NBHcrU02AmhT+rzvbqt8tFq+Tm3atXBwcjDrS9q
nX7mE/BPSSvlUzo8QseHjky8GmjFapSH+kdEAKOf/QqS6Kdn8iKbm+JNvxJ6LbbW3NO7v9EgYwlE
qE7I0niJspcvVL/cp3NMKenhEmSEASxmq/GhWGYntlYIjQiyFJ9Fjl418gPTolPhrx76F14RSDAz
XEGHMk4JsgpBhnrSirKg61sWligTBxm3cIHCX4psMwCwXHCeTde3RqNUs5sXkotjlm0GZuGBpGGw
tNF/lU1Jjb6ITkAR9xhqCE6sVwbsBd+RDKzL5+T9eFy6X+M+kQBkaiYSMoPSh9fMLIU+7sUuLv7v
4nQaRO7IGpUEhEwJEIiwkoF2+eURCm0NGzDIkOJMA3RESgTawDCALN/l8iWBLczSugAOReIODyvk
Mc3yTYEJfIV56byvWwApW7TvKvUqj6oknhnveN28Z9YsvqT4/6srmzhW7IBkpSacEr40KaweWw4M
r4HKnFarNiWUxPWnMgXJmDdsFFJQaKJA0zCEav9dKdEy/EXvDXcGmgSEy/jWtvu9k5LIW8nkm1qV
YW/FxtHKK+wZhdW5CbNumoB3um+YFVRC1pKeIkhieVaM3Al9KNKXvnNcPqvu0gjOq2+/3x/Gs9Uo
Rm5Bh6n0tjOTaj0yrs0m17UlTIV6KSmQ2atQ3JQpsQmvZjn45qdeHTZv4OWZSKyDEPjRvH4XR8IM
a6xJaDc0dJ/ET99yVbRZB6xvSQoWRkWP+nfIrgSACiw86wmmXx+pcQEXbpN+BKCll7nRqyfCxNjW
AxuwAvXDuQ83HapGhVkjkuE8tQshuZMs/9z/cF1PQQTBtDgp0X8hehEaGaNOVNwrzaM9XsHKuPrv
bRIom8nSWDSBtlin0/fwuZB7NUg6mGs6mgWwdFAsQVGnBSL5sSv29wFklUPATDMLLBFg6xpOlO5+
b0/BqBylfAsVAIbFPt0+D04A/i7g69Qnuwby0BBTGK8+3Kce02Jl2Xm9zqnu5OPsxye07+QwLq29
dbO3Ai6zTW5ljjimxbLsGtPB1oQkjnC7KytoPyDXmotB+RqeWDiPgMUgUJflsu0LtE5DYfoLWt8m
ALErLUNZph/AJwK9ZAuQnpV2IGBGV5mLDT2LShkJYbctTJoN/A1A0kBMnAQcHSEoFoiWd0yZ0DL/
sFmm37tH82xyu5F8nNp0yG6L3NHcFwPog9w9Z7fK7ZzT8CxJ9aa6RPvGuZHBHLzPbG5ueG0pEChz
fzx5SpLJpxVX8+H3Cpf1ObEe4B+dd0I8dH7B6V4c2644njWqio7dmpuvTYu6VmwI8LGdS/9Uu+jI
YXAo+MxEcOyQCweXMrrl12TQazfyHzd/4QlPHt6yT/gLKJWvA8WW2Bx2/QqtMbV7IdLC4AkdthB7
JGRpOIMA7+TN9SKshspHTnxaBsO+HX+4WXuMKxXoeQ0XDzRLdb5Banh1vUoCUylANRdwUQMAtrou
hjKZ5QpcGE+U8l2kK1u2C8SGuBAduKds0ZUrinEgBEZjt7zXDTRXP+0JWbW9KnURnIelbL8SXy5O
owegOoUy4Bu3tfAu0SEI6bfi/Zcfl9QK4lBLk2kfRMLxUjhMlt2dxcspSMAApE2e4h/5a9c5bbVt
LLK7oh9M4tpPiy/fir/ledV1vMTBq/d0FnnBt7ysRnX2oGDYzfI9RZ+EgaAqHAcyO4e5zCRh9BfB
Mwmu5O//hiWhhdk9/bj2w8DoiMmOmCrNTBWzsnFiWjZyOhxr3U5Sp2k3o03hG0W5xJ32pIAFTk20
orQWIO/XwiegFgnmj9ElvVop/Gkx84belJn+pSa2Qxg/bnY868S/iSijxJzPCHgKcZXE2yqNQv6C
lXkJpWEbJG0VWGBr5/BPBCKBJzYZVefPr/N3gsepL2AUCqOnZgHvtgMKAcYgdG3vC2cs7H2Ym3b0
6sj+nSIY7XSkhEE+i8+Lcl0OeEqyZE3nzCEy4IPgvR0dCTARShtDQYVyPHtUIjcZ+FbgnvU+QLSr
mc+DhhG5VsobHuS3WFxb/mYPLWhqhSDFZ+l3mJ7hgeKmoztvFbYM4/4myV6k1SoKAiYwaGLRhV4c
8OReJDXISg2P2VVRhyrUmyWu/sdd7wgpRx34qknjsXKTH5aTwB7WIxiqQqyTxIIME8Z9ZfUn99du
kACj0pAdZc401QXKVk4Ajh99p3SR8wjuOHTNkezfK3rA2530mdXu+ATd281w8cRfJqQAOSHmXJCB
oHbk6Q3jBZ+hcnJ5K+qfRHghkQbDxT/si89zPxrtdL5lKWfGEsZ7F7dau2t4+eNTtdoWISo7OE/o
useYW9qyN+ocGm3BNcnTEr/XNhmePZ17wIaiq0SQLikVYNvPgxRSrtcuGRGet2byqSvndJ4k4WS4
u8ahGBSRHai8oIKLiD+bDf2zdMIRkcvJiqJx3HjyJVV5HuewzbjvR12ZYQCENxauArYYanUh5OJu
j41T2jksmivxyVXcDxVMrtGcwjO4mhA+h7ZDL69g6AbbC8JmXDX3aEb0ZW6l0VEM8AcMsjR2tuC8
voBFlUZ0YstvZvUwHdMAu1F4bONNKomMNsKVo+wdukxYkldcjbHP0cOYruQALw4/HBtCeKvaiWFF
kfq35LaTUcc8dHpwZYv0fa1hkFtOwgIF109ryNFOpPNaJuIdiTdWz/g+WJbpEqT9pFM8NBUxsKo1
SHD0PDtqshtSTLvXT6+HfbKa3em2htDIk7/hTSLQd40QtAeWVQKsIgu8NR0GfGe3brMHsu4dWpzs
1SJydy7aKd4roubPkPSbofhI06vaNnu2Wl6g9DuwqHum7eTuUkgxR38UsKWzP3EJegXp6zV7C5Tu
H4haA0WP2XCuyQaF5TsyxKoA956gYQrYGgRi52lKnlR50QUI12Ux+mw1QyLVv/DscfPBiMe+qbyr
TfW8GUPlD7RGo/C5mjzhM5QnNBE0e/WUE2VgvqAUbqpg7Ek9dvGdBjDl2lzGdmWe1yjQqcn2T0o5
JlV5b+Fq9eqUJ//xgmQJZAmCxWcIC4w6cjA2GtHvi14frKx/2h6jF2lNeNVCodLt7sLQ8I2S5W3z
7cxiggDZ6K9dF8l52qP/qTk7+BOF3l/qQfv4m4AIH1sv34v4nLLMZ0VOpvZoOXZ9FttqVazgbaKt
isjK2sKS7ByB8k5kILbNYiTE5Hh6qOZETtrdtV2+Th3NaYbvTXgf7xUWJIpFmvw9eAoSUTJrXJRt
z5enFmz7Na7FWsdyyKTb/cdg1Xt/fbXR1IDW7Wt7FWve/3WcU8jBx9/daF9RyelL5mjSfAQaD7q9
QwLY+MJYaLh2LLg5RgfjPk+RxmDGs3TIKkHOoPnHetJqEc/eSTf/XV/0CBtSGlGnErryTc4xfOrz
D82fNaEeIGFNgSV0dL2PYcUozmXSkSUOi1MMr9Jc4XejL8kJ/8IEO/Ki01ssDOwapBWZTPtb7hDv
ogaJ5i+jT2t1BwNZdFpWlPDWfNvk7Lfc1dlvSEMDxkGtBv/jByzEnghG7GtQXMonCmLFW0r5zy0/
W1lqmDR5iGNbH0vFiOgmVBy9mf4A1uslutkO82LqYpqnOJUCqRsR+Jg9muevc9Q1d6xNtZ+PhUhp
PsK+aMTexH20g1Xcm99PxaTk/To3vHoLGUQ76BdPjD5lxU0AjClUXYrt5GPEQgLWGunkUjqb00ew
jKDD40oDETfIaWWekIq1wfAQbrHT5jEXnbGQ7yff5X5etBoM3Owwy/3E0U/JqOeUTKb9eCIU7/8V
a8Wl1beGVW4wCT+h7vV86/aD2tdaZnUfAm7X1uRYb+UOO5wbsGnDr7nzEsHyabeX6S6wTIsiE6L3
v/it3wVD20mUJofnoJGH3Ua9ecTcrVOstJr18smjHK9UAGHvzFwMz5SDLeesJpn5T95A1jlOsmM+
ickE8F+N/7yyONkLESpgYTmbqv2mhcGHVFl9NUm+MT1caij67JROyUNyx8PMF8QhSSS6a2VCsvtL
oLsFMMb4dYN6JsfBhuUaUUtTn8MMO2oK9YPQXMBbROrWbraH7OOTHuzVxSUsFieK+JGhVJVzgYPw
Xo+V3Dne8XOxgg9KD4VsimuOUuvI7XVW0ij8eFE4GWx9oA/fCuzPpVFh+ZMSpxLOq4h0Th56trm9
tfRJyroTRgROYE1NIdfnKti49Odz4joQbnrtIcoooZsV4NDvEOsv+C1R50zD5QXwRTfS887M2kVw
wbA7GsOKvMHeegDL4WTNjM228QIUESfd7wz9pCUcuuq8gf0JJOVOnn6GjTRbdNmuOJnh9lFOgfZd
2TGYkRRmsXYPaAVwfN9c7GXC3AymZIQ9t21Jc00e9bnrX1NfcYj9FprH9QG2niAc/LK051QHoobL
daU18b2w0sObRc2QfDohiJpkGazRycHte4DL0t//jXTLafiV3KMhdZJPP2pLaCxW2eZ8GiQ0V+iS
1QuHZ2qV3udXttRpISXMmMjzfnSReABz/uQvaWS60lJmBINDxv0cyWCrjcgtAUfSX3uCckNQhryO
iVuO13cxfjTRCj7SLHgZr5mjNgWxmr0dwyBHsYNUhC8BJ8gvspW619j8Dkg3VZepC3jPEuARx0uG
JZ7axiLTL521GfVbzINCoLhYEC1+0g9stfVoKxV0l8DANMZHAej9oeUSNlQYAtw6/0LDn5tAk3N9
vMnOL3Vd3501kvBSc0jhooeHIJD4UV+YoZskpDqdFUFt2dVgBFKNtmbBzjcLStXBajfE2VjpOAQQ
FGgxKevCa8jIVZUjOTn9y04o8D5V0MZZybYWx/4CbLW8JeZZksl/nzSrnQEFL9UWZWi7YvVhgmHW
LjJRYKpqhoWY47zXKL4YVtCE++GsiKMnOhj08K/gW8txNPYphpEvstAUETvu8PSOgILFoSdpQoXG
3OKl4UkOgBo2x/l1ddlVdg4dilfdrDmnmjtGOTGUHUvrDdGsR72j5p2ylOWKQ0xh6AfPwdr0//cM
g6wD3/NI65jJYTWWrJlVpcaAWTpS3H8l7uuCtYGrwUYQtUAKA3u9LGnHxu3JxL0YMMdVmQoGSMeF
SRaXiVXofSlMvCLss9Qc7wAEmz3m1yxBEemJyie6dTucPiitszVCjMIrznff2s8EGvtTY+rSwDh+
pwx75uPPvF0EpK96lV5FX0W1ebgk74umE1ntUTUExJmLaTciU+Z/nuqeCoLI0hRh7Kga4XC630H/
1IQVCBeyHZyFpq2PivXzdWfBmslr1Q7QWg8/+D8Fw7g550JGL1pmnzccj1tadm5FdmrI9b4bqyX7
1AZSOruAL85kwP6hABh6KBjdsVgmQTYGEFQfkL6KxMaLjUMd4WCR+gvdxOAuDvXnzdGFq+7CM2bG
qRNh4fKVYgOHtVGd63IVytQqiLZ4i10EGtQQhymRA5/w+0DqwofZWelIEGeNlAKrKPlotZInlP+j
J8z34A4TR7G9iApYV+toVYeFv6aBGYcp2oCkREuJ8xszpi/W1+Z5P4noDFjyZkNFh7Q3/D0om0qf
M7lH5rHGfs3gCXpobrNxMLyTAKUC7OC0lEzZ6iPmVqxMMi2oh6H4lP8TooNmjnMHXTYCeG83KyZk
spNZxGJ2mDBA7moAeY7rWm2bg3Je3f0bHrKGQMSHsI9YVtrz3YUsSJKIdiRKBBg/2KUd8MpACq9X
9KZ51j83/68UR0eQn+nxgsr/AgCMtgxqcflPNb49ugcjOsZzZORNWItJRVFm8kBgoiCRgmuWGrYZ
j6J/PvlcL9XMh4SZhjQhLWq019GUWZ4owF5gdU3Z8zfUkGw/E5+ulMbadxsHgKxKaK3CtjPR52Fe
TAbAf0bGKycp/aQqaW2aydXqx7lj81wABsM75uSpdaJTDy5OPLRlVb9NW4qIzVYv1a3bluTagK5S
2XzN/+n2TgudOTAAZNdOq57Ii+V4HYWpx5l6YNWghNRJv5C/WlbKwub+zPWxOl19zxzahCORkNoT
4ztjCJfmqLZ4pHledYCA9YN3q8TCYVJX6CzKO05J0Y7tmvTHsodVWbcVdTbUr9H/Juh4oLpBwxS3
FqbOGXy4JfxvveDp3wq6NtkdI4oyIgOTwYK43Z3uF+Be+/889p5PxAQ8KKTPdUa3CHZ9XsR3KZws
mVYskqX/Mun06CRy6bu7cDeNV9Ei7guznDFiVhqyrcqmUFQRque/oz/jk3rVV5yD+el6OvxgJK97
6iLWUaXMvffdLHDXbAljORwsfiij7hM2OdS0v3ZqcE5cbH8mO7lvhxIFLH6n/r366Ws7VkHal6Jh
iIuAbgRJ95aV/HHdK277KKYrxS44+ipePcd4YPFOYXBS+eGCgoDxLuh7+0W1PVMbXw2BRYEf+A9u
lycRG+QmBWgGX6Copt10u5EG83mW4NgVAApC7K7sxc7jWcACrn7gD3bEUGI9ubX4VgkQkWq972LJ
IRxxbVAdSG1AJfg0SZMApmgJeYBFIb1rnI1MrD0WphBxR1tL5O9oa+ud34R2fUOmKv9F7GvWi75h
yBEMaf3Ae/H6gynbNfNTHa6EVqTfEu0eOM2vW4YQRAl8E5V5ejnlV7ybqaD2SAmm396nCdfoO5pU
ugpWhS1IM22nUiH7A0xcLWYqyQ6csNa8Vffgulkm0JkP+aQj9GHJpvlC8P1DofAYG+eh11hZWAuK
2acGItTs+q2MTQ79Mn6sex6qn5YBozimBsbAYnvygXDOUuYAHxXm1adG75qzfhnW/FHX2kdwO5rV
caQ10VvTyo3YTdI18veJt/eWICrt0elFhWINCmk1tgezJMBOWnz3EJYr+QI7Vluk4TF6sC0Cq5ur
nCuHYhJKycJSMhkA1W6+Q1GDyU+oxp0Xpx+qhBPTnecsfM/S0z3H2VrJDMXi0F3dX2MTQSRlwZCe
h/TNvQcr+jT0UjZXtoALsKnPG3p5aTxTuKzkAeUX5wr9OzRX7Qn9VNFz68TV60JWOPb+gE0Pm+zl
ecxvAbWn5I4n0kzg87JA3UdmYtdTfebTY7TpS9yILmqc5oaF/D1sPiIV5nidOXBYNkXHkeURPhwE
uyxMBwBDS1mrIEu9MRRVX1rBd/OJ+tQpMhyfAyutUTQbD6Nv2fpUBPO8aWZV4N/F2V7Klf+j2gc0
ESEFzXtMjMPS0F0yNNZ9PMgZhlJhvmW95T3K6LBncMeAGPA8rsFWBEroSDLBTraf8csS1WvidWhA
QRS9lnVMVo5nx8u6S1iaU85rOI1AkvkYXr1pz+nfhL3qMCCXuw+VXOIx7Nq7qjW2am9sNRxaE4SU
DiDi7cGNGma37i76R9rnmM5usBgLEDsRSYDRSBh5SbSEIB1G6ELZVrU6KlQFc1bfyWMcCBWUX0ZU
WSCur82xBdTaIPHyp7q64VFNjkG9t+FBwsauO6jeQp3TfSbNVRMNMpkLxNbfpXYeGb2QoKD/grM6
Ontqr3ucsRso2448T9KYDkYt6H3lMU5gFwxnQL70++T/TUDK+5NQoUkx5d/c60VH+nUc7YvXhSEE
KH4DEHZ3vSrJf5AbG9Eho0fGxK/bI4O/COawGIskwOj9oY+O5wdolbnGHlWyQdWteRuz/Qdp4cCL
oqPIDLDKjIPeoAKtPA3/Tl5eFOpjBWlEnR2Egucbduf2USAcFN0EmXzyjcsGDEVl+K5kZUTjntQu
AnEaQmgG0hkjAdFlk5Xm5MkAyykTZVYPEcp3u1TNr3/MKcJL+dUd22ZqZYHL4lcMjEUKHX+Hxwhx
b5Qy92+4Anjligq4EfmszMQ1msM0yxZQOCjRqdcVlICdk7JRt1x+Nv0kWMhiiyUr6Kx68oRwpSP4
e9DxDQg/94swb8HAjsKovjVeHyNHLmlEnqEa5B65xbZo7OvKHgDyUSnaeLzrAFEAs5jWYR1HBAdL
Ed4MkvvK4uGsC7qHuuBtbtXMPvlsmQmhpkPgHDjkVCjviC7mcPYjCK6eTadtrdseUch3ZoHf4dtK
e01pjIjUTI6Qf9cabqxS4bT2Mi9r45uaXDqH5QVL4CmVSClJC1uQN08/zr/1RcqLsla2ZUs7JapX
4QBgGuoCu9L5SmeqakWI/TKpbA3Lt3OdFGyAEnlRuFBq8IQBfp1gAkpdGcQBe/fLWm730UOfrZRT
ejeg374TZwC8hwAQXMncc05zIZTolnlLBISIIiLKYl5+pyNgEzCTOatVnt0Q4+mMbqchlsKa+E4c
tlBgn73akBHneVh//qfHu/+q5BZ4WxwM5vKK03URspuzpOtB0687ToeLACfhTgx0oSZaiLkqbf6B
6YCYjSxrUIKeSUOP1+rwgmERYvJo7jAD2oTqCZGpQQeHZMh+6xodXK7kX59CgDcfa5gQcHdi/3fO
YrxroxOxVNdf7PU7W2PhumiR16Sj3jLuDQGBTw910oLhfp8cKZdyJMhbGQ9x2Y4Ot1zSZ4qfohVh
7HrYLwddVMpApDfoC2VxGbtJHHtmPO7PjT/G5ro3ZiA/s3FQqpeXfHfTkJKdoNThSNVOUxoeGmqN
O4oOFKIkpaJTWGl0JLC0xVGfNVXowuMrI1AkkVmb6XG88N2SOgIImcHZsOh27ViMwwKqapksoMDR
ZOv7IresasyCmt9U4zYkcbIoAzRN9mIT8m2zY9SvRV0J5CwviboUmNtJcFBcBQ0pEgibHWlm2r1x
uA7BZcVce2zOYV7tXWaYfADnqEoQWYXVienxeLig0UUqQJ6ttdXHhPzEjyMPs6SR173iSzbzpiHk
rnllgqBQ4qDQ2UKeIAOLNZrx4h4DJ/p91+hZSMbRW5t0zK247HZgfMEuuQkdnyOhbSuS4PqfVjA2
ixDeg4H+jpZOL5/e0ed3o/qb1YzpRVr/bMiZSB8v3vhepF/rfAvB2pmHN+Lowx74xi1a7rxS0tVH
0FbxxqA1IuLCqiidbW/uVzQlo0q4X8+UXz2Z2Yz8LFAKgm3mm5aS/hx3QNOIOVyG5lvxCW6UkbUk
np7VA/B75+dCPSDIlIpU/9Yz2hu3igTkXuKOwrzp0CoEDV1yhP9jDcDk0/NQZSJrSn9KhunwEP9v
xKhnIPhCEtL30TcN8Cepgv+87rEtnmqQO5CU4RHaRfvZRB0ZAiUYNYC4qdg+j5xlEkpFC4v9NLOa
UR5u4W79Jbl2DMakGAUKm80FwoZFnuiu/76Rt41p0Er8B9mXHE0pw5H2fnMPzXbEnftyFQzydg8z
Lbj+tMFTX2AuXj53auczTuh0jx8tA8AsLdBjTyCIyy4NnF5f9icfcDMaiV/Fjxixz0HmT509hwQJ
vaZqka90YLkuYLag4isxBsuAH9ws8Xo9QJPv0zcONdzqSQWYY7ma/4H5a3TkKWs9pg5tcqoAm1wl
dCPtnJuLz1efjw+GOeTzP48+7E309hwRqplh81Wm8pqZADDR2lrXtnu0cVyHZzGm+zEFZUtovbj9
yTufJG4A/EuqSMXphgQ3IXzsFqTBJtwjWJzE6p3Ds4OXuOUr4DNqiZA0v42/LLml+oTxRpOOtIMy
0lQNWmWRQb6e1VqdddSg/4vlT4zMqw7fLGOWBQ6oMTKZv7dcdF71fLPPdP0cVEvGFrR5Z5+m7XOC
eCE5VXn3hvDGBeQirI4yUvLcBqZoq0JghHT/FHMdDjPVikeR+Pk/lT4Tg5GFgaTOe4oaMdY/7FBt
QPQdk0DTMvDDbpB66tQms1x6cpRqq+Tm3q2rIxCOR9zGwif+Sk9PAa4+x2K2/fecsjpr/a6tOTBg
ic39L5wHK066lJygkODJGMRzDWYS4fNfMiq8CnvL475KgcQDWAxriwEK/QuLJ+C/RXRIcBkaUwCP
Ujt6fMQDvsStcVEY5PRHEETGI6HsSmLXtgyYgL3ZYoh/O9bj33vZp6bZsaA82hCcy6w7zCxWK3zI
fMZu1yEjwqOn6ct3p+SwoYBEUNX9t7ze3Zeq2NNIirHbcIZsDmYDMzXbl/manVuKek05/RdKq64I
NEcznZOSJc7EEIEiEHz7Dk+FwtINpwU1Cx5YyLpvWGlPsIIY73x8pf1iB54Qjsqdf8NOaKRg92qg
3lTOI3R99gKmwS6G+Y9nQI4SJaPmu3uETXhSrIqISWrJLU8Mm7A9PKr3HztIhxbEfk/yDncHm/VJ
3igt9V2ghROpW/s9aG87m0+n2z5onp9WLXpxt38kJDjydg9II7Kyx1PDFwCRHyI/iAunHRVPf/7A
4O6M2rrFkvjgdc6tQ+/iVnoP8AD260y6kSagAGWaU0zMZG6ZR1LwC/FQo4poiQIrkulHSHo0yhs1
sZlshab1ZQRzidKCkstXm6ZuINVJ91t/zOl4Dk38Udhy9d/Iec8EsU65gBxm7dRadienpT/+SP+m
bvJbXMd8BPkU+qPKsMzouAgMtT2pAV3xJ7MPRh5mLRsarsPB3hFNy8c2esBaS+lLb6VWoMFOzFUo
PxGN5FS12xibFS7a/kpeFhfjGtrUEITIWMI+k0+x/V2sllVvpkFumSXC5oAD/btOgOj2EOciy0iC
3wjvdEFI/eKqLTlfufmjkW83MUeCDgEpsSzP+nEjoQPzfIMzQxQqZuWqwqYRHW9sJwVXCIxWm1wI
21vEgpdpmNmSggPF4ZSWR/miF9a9gVMEhgSxPMFQMyca9hW2EGp+Ptij2zfWNaQHKfMGC52Fv93I
SCKIW64y/6adORc6gnSuZPEEBrR7agkf7vO1/8KpLpSm0f3jpfC6DJBGZqbD3ludWx3xA7v9VWFt
cwfWjfJMrGykbbiL1AXNsalfpht8bLSaPOUFVwWUq6dnD3X28udHtMWsUVv1CF7XdPHwiXcoOxNV
WwJ6Z+e2IQuBMqLDg0VTNRcHdXPTmC1rqOgyIhr5iu4qdWrCIJj3CKoTSHxEh+evjBFXm8e+G4ng
PNycxEt3879rDiBKnoZcmin3Iu+rlEhhEzScEWaZKoMsgmNuDU7AX+uvQ2zilgpdT56RjXf9DTu4
Zp/KxOLpbe4cQSV9JcOF7NUzoSl0pKNk1cF1BtU7MZ2BJPJhwg5zFZ2ITd17WOWWiqlSCgsZGjhN
dQmir2ePC+Uk7B8W7YtD0J93jPbcaO8hLI1gFszWFfL+QqxeXY58rgttxzFFcrg5APcPq3TI455b
2Ej3U7dzR+6qAF2lmWf9jd3zBgMrkjgqy4QZ/mJsVfksQ4j1hwEhDL9IN1SkPRTU9HS6x8Q74PAJ
uP6ExSm44J7a2h0bxdF0TrBuW1d1PxlaaUfylC5IG6BuEYbzr9L7MZ9CXvxfHNEi+hasL9raVuyW
3kmbVZSOM0UBaLQhTEFfAha7V2VJ9dZi3Vzw9i41/hj0t1Sgnr/zF0YorokjCSm3vEH7gWYi3hl1
cs43x+41BWdQ7VwxMzWXj15c/xmFkhkYsncRrDiHj8kI6u4q6haHoLoL3B7DN0fq0bLrprM7V/yJ
RFZyJ8q78qsW2fTqKjV7zA0261ZzmPNgbNntR+4oKjoDp4d/Gihn1BXXbcTVcCeA23Rb//2lHNtQ
tj1gljoxmdfS5QyWRAYG+fYKsbqOBKZcYftvaMd5josY49fn1uTOCN3n0bV8OcKEavVylpL5UdXE
lcPFUjA2+bRiI8CTs1jprqwCvIGmh5Bo3D6/2mgwdRhXafzZLc26FzmykuSxbOGzcRwC/lWosZ+g
tq4HKXJQmAx3BL3pOr8x4jQUU4xvY77xnr77YYtcFiPZ/31evvvydnGWfj9gmTCXo3ld8Uxv0LsW
oud5yOo7nezZMuFhNsDHq7/wDDHilg5As9GymPut02GI7AomEp4bJQaJQTjONCh+v0XwmQkYJkQz
Q19q9IUr1eHqkVGjQViiFeYjKWMyKnxY/+NA0mZqaQwf4B37fydZIgflTwWF8Gh6BPqBSGuJkvVV
7Tx1TmSZ46gwFZ0s45ihADfQY6dJwG44LB752SXdqp9NqgZZ3sGVPh51cu7MLYVoZKc6IrsvkwW7
7wKUrh55e7uRIWzKFImrOniT3+iVp8Vt5menX7oQNT4PPQQjiTHvayneNGWLgkWFYKzOQesLyYKW
Ey89d3g91nVrrSDH97c1FSnkmjxzKcQvec8xlmWU8Kg7uOz8zOtHsDg5kJFcinAM1GlYYv3sqWn1
2RD/0LoHnkPUAevkVDRJjc75V1i3KKOyivDjAvczBBWU9sFfkWZYRwgQiILEHfIYe8DHg/8sBG7n
DRTG/64TSWmKGxQP9vMUWnJK+1YhoCbGDWkxH5VtA67dOXJpvAHwV006sdQfaTezyNF2oO+WWUiW
4BtVonGQ+1zEyk6e8kbLmZNAWGF6j/J/zKWBJD42C37RXfzU48Bb1Z/Vi9P07vWeqLmRAeiZfBtk
fuUzyXanrseb51o6VISMi/pE30vP4b0XWP+monmVy+bMlyMv7wy+NYl8zbkzTIP9/Nj/hpKxr+WK
MlNQuOpcC/pDikypU/huIGlJur0XLjPTTYN/z0766nFO72Qi5q3cfwHAW1E0KQczywWcvZZgH9PE
RSITzVvIL/j+hQqe2uaW88my9aPe/i8sbHToebGWSd/U+pe/FY8seF8FPaM0Qe/wJDr3R0q3Y0xi
MXXhTPwkc+zxbcJuCDx2srfrOGgAfUSgVH0RfalqcJR2CRB9zt7Pk3lAPDqHlIyTj9iKduRyUunF
LM1R4cqeSg4k/AOtjVJxFewY0mAHr0ChO3MN+oNir10CN9Co7Cl/1Wj1UYVdfYUAiRTf/WduOSbE
K6d+u1/7GxBLUzfQpeB7x6NFV2pGN6JpIl+xaJr2Zc2eJzvrYJFMoJ7C//YVl7T0KISqRaAz4a0l
7mYL4n7HRY6nceSi8+3y/VI4kt30pvTsApU4WsGv/Qi6IQMQ/ztgJRZsUPS4YF5L7ouAfcHLpu2B
eyDHmthiRYM56wl0qAu80pGkFhjOljnAwm/ZRxSZ7l73EW79/vU1i3QS4jd5TRkVNUdAPQvHPSHN
UARlG4cK3Wjx3cdfhFEEYDf6xEU8RXoCls5jUcZ76HAejp/7GVJX+J+gHO3hwrdPOkm6nRDITVvO
o/u8leFxYtXKMzyUJScEpPEBKPB9c/tJFB2P75JL36FS1Xs3v1I2Yz3Z1fSbG9HjwGNRwnOilwHH
wfcJ4zQq4MNMZ6l9AwNIfL7C+k4ZhlvqzTC9hiiUk8aoFCuEX/VDdp+5a5Pjtwj3+Y/LnUes3qK/
wjiv7Il1pXWr+UBHQAoeloQK7c2Aml+S3HEn7y7P9Mrf2ERODOlRYr7VqafA3ORnXHNvPUdFdDNt
CfTNqJZ/0A6mPwM7kPobEF7qJHQl0r+LR3E26l5WauSlZC5rw1GWIr46Hod/HJAKSYCt+e9U0Fkj
K4F29ehtv3gFnjDTd4djSUDaHMykSAXWvSlSrcij/UPORysKzdRA425+sP1ucXliY08l7XgnrJfl
W5irvNO4Bnwyz5nZCxIbNVlwulsDgL7Zw7Pi5qhmm5aIh/RHMa/qEQxUyeP8Nyh/iuIXqS8jNS7i
eoKTlswmjKaddEwPYR3lK+/8l1W3/LqwY6USa2r87zyXrUvVgiA3U+1l5SQy0Pu9QseReJ57E5qp
p21J+nFMXvWiISUjIROhPVQcY5VwP3WSq5iSKNxlVOSo1W/du5ttJz2jRbN5FZHpyL52GOHLXgo6
3um/0RiiIXNTVm0jOcMmDKx7PPKYzuIMHb27/nlMzm9k5tsD4Oka98M3jasJdPa1pktESrdll8g4
0htGkazP1c8WHNlPWPL/DdE8HHT2aPOy+mpUVa9NFjJ5vPfP74uK7Yj9G0juy/6DS2/f0T66P4Vi
JCwrtbFQrh31plyxtvGtWf/aXVU4HzBEqMsKMwJaqBur/aCH/QjeFZDJ/FGG84IvEyypf7tzR2aD
VjonAxadCqRf5n2PSXikANdKH127xqT02GiTH9Fh8kftuCMoRAi1bfCKJ1G09bTeBkLpyFnMKnon
FiWGc6Fs6MbYD239xIaK4brebq916OyzZkKGPZVOdYCuAacEuWdKbxGb/BZAzIyxYeJJXhiZa+DU
5AJNN8ZYWf1aoAq1liy+QKzkELJIMkVwbetCnKsS3ooZLVNIYPybzmJxAUMSxPe7ZfV6d4xbfxji
89yyM1ZQI3G25evX0hGR7LW53p4UaJLY0m2aMbhO7o9xdzLaYIsrewYUSTf7leZrrTYIo+MvD7/O
ilkeepytnsss16ggSg1AP+kEd1ys3CnIitSAkK4yYF42j3x+y2OSCtjOqn7Tg02GJQKLC27n1bZs
7OlTuWcOAllT7UZNYPWA3Bk0o6cYM4bI7eXHshQiYmJO4HKVVyB/fDX4AsIaylFX9hU0HuQlyXNN
XL5jDKiUy8vfz/lFqlZXUbiUKxQooY48LF6hYJoSi977GT+3AgkHy0GPFsJUpbQctsT1MH+dRKPN
PXxbTrs/y+6qTYahMEAwy5/z5/bqNE2ybnpYYUpExHe/tmZ+geO3BTscI4JR6f4dS/bmyvEfhnpb
86hUyZ5PiaQDINTUyGdjm5/EAgOqBd1EnfYpvR3fJME+xm8F940vLntETvbrXxZnRKHkYCP7/TJS
myJutP+U9Mew2r99+HfpsHdGTylchslSLJQuqHtbi0q0d0yc2gP8EJRpwaMZai5Ry9lnLh2QUfnB
r3K66cq6UJlv9Qes1z/VO7TJuhlaT0WcAv6mmx9VLA+9QteU+VmYv9pkQwwHHbnk8Dq4Rr8B/WYt
1ysacVziuxvTpKaaJO+6VCihPMb1dZ73RGkafn22j78L/FCTAmp8mtnKKzhA82nkWbQJyctvyr7u
BbMSa3TKEReYRJd4xdgEpruzB3n3LtZ3iTaLLS+2iGdmFOyOqsfRPMOqgoB9w5vF6w9fuJL1ltyY
37GjBSXl8AStxRFpraNx837fRghpKFxfOvU0+Yco51fW1UU85SrDarqoXrjMD0gzgBtZS7y2/6pa
QNAiYJ2WcGSM4uj2jtlxHkAxkYrSZ3k4lvyZEku6HzUcRAuQz0id4GPbJErIN5b3Mt1RKdIkAYhZ
hoefco5xx1zvJJ71KFfa7O3ry+/gNa1LHeJSHO2Z1F2hNh/nIHzshhiW/U1Cjbpw7Ycf35JbVZBJ
ralItXjS1mMtN4rH9eiZTU7dcUflcOakYxhfgVIZWnlhphuxF1OEOR6FbnWa4dEabMahJH2yIox6
xYmsH4P1MBJw0IXYbbiwPdAqoyBlXpMYzZGE0cWkoyFDONTYXQeu6TY1DgUmqWRbljVFR7JoURHh
c2yTTiVKOh0WrI+S9keVYCNAWtuv54aAJmGSrXlmdG2rLEJ7jfx/HwInO1PxBvSM0+tM2wayer2S
tQIQIpbmkE6Y2NcZ/3vYigPgybVL5jr2MaestQ2maFjy+IsW2+cmgJsVO6uIS35oZAqXk3UhnMf+
RJjLzL+iPc/1Mk1m7G7UbXznpMU8qvHco+6bgMvUoAHFWmuJgMF9TNzdPdFEFjL77ICa6foCTc6k
T+ostw4u77Ol60YrN4S+UqX8IHySSrDzq97qgb/+c9jMkby6KCdlieEdROfyet/dP0OyJOv4UfnH
Zjki860T4OxK4LSAjBwJM+aYsYI4V0nqxoLPCeUth05k7t6+dNBWK228fU0W7OUm109dqQUvGDVQ
PlIkq2hE7Jq9hSK4k6r3poo0f0NTtKp7BVAsm32XaPuddo6Ej1bMUKRWI0sHLEGMNoFI1T93aEUe
3xR+gC4+fgLe2FiNwPLpN7M9foLITXIReqQmmkQfrfOtRgQLSxqmUr6TBL3AFNHkXnPH7IXCNNdc
VL7bNuks3XJdwXTpRPLTXDarnCf/ZpdUFdzya4wncwoCU42XrMn2h9AMgU4UzQSz/gsUhiAOATHV
eK84f5fIYbgYI06QA3vof9xktu28S+znoe7TaBTikn7DYp44LrbSC/yXtxGbAQKyCZH2LRyuRw9Y
+LWVeaUTIeSs80doDKyiKTkf+GXhAxt+u+hj4qaCsU5Imeods0Si9BRZ59+JY4cPkNewRq+LOwiS
6BdbKzfLipHDTU/9/XoucBUF5jIugpoG6F2mnPmvRTpC/7CO6inaD+Ih3poaUPfm6y1NrKowm1eA
Q1kbjVPxx3aZuK09a4mCBF9BRT6SyA4tirbpq1gsU6pCHzvDckqE09YehgXE4QUJ5jXansgZY8gP
yakBPfafpr4G3Vw9/MpdecoJ4z0s1kisFbyHXJAfZh6K++KtL1df4Qq0ef2P2pmgDO50uFbBfSad
+gxd2lkcCU9B0PIDO9/LYb2B96B4FyPz7lafCJOANcZnARo7HMnXkXU1CUtsI5U5kcEFle2mtVXP
2HYRfQCrrgcu9dxmS3BADwQh+hPW57isN1WHZt3TKeIOwBB/RLYJPhBMXxYE72RQHZzAnMRjojJZ
5NCDwDK+40drYc5ABLaWQF0YtzN91RNl+FINNrOxAo5i8PNubBlnJe1UTrh8HRyx0/OqaG3cXRHs
digrryni34G6TU+T1yIeblpF8UH+0/84D8bD0rCEW7fo5zescdaaxyXgoUs8/kGCKTy8hotwPsBO
Qtc1ue4pL3Q7KA57XXVb6kKJeTT7M9NSt/PF7oNcjAZinBSKjJGoak+Fd095feDsT277XqHncHpX
zSKgomz6YNme94wwt1zg4HVU9NJE5BVSOY/fzU5UCaopHxomX+rPHIWRRK4ah+frVHvzS15ueJv4
4BcMnYFg3po/ypp0SmauxTXB5Tho4i+2xil7oPtBRTVZaM8SYPbvxEVyWiOuPZ+pi8zuHpsH0yr9
h6Qlpm2ruheMTmQQ8ZpGmlvVsfvCJSi9Hnpi/YPBGWXz4QRKeQ4yGkvVNR58HzZJBqjf0hxNWPmn
3zhqnHpvIC3xSL7WdTvba5wP4+lMIFMBjG48+hHelfDZOE1yZiNkYGJuB4uqGUCFYTk7jFvt7rw7
C9ynPQ48W/bOxeLAYzDd7lZJFA1RItHKN9UrEqlYG2qyhz0K3+PDOWxHUzUb3Qx10sZ/5NeGxMTN
MY/R2oH8qnUZpCbIHCJpDcmH/lktNrHMJE/NqVFaqkBi3ckON8DQriuxrRrZyLZ9vijSyvtShkVr
JOOKdD1rmwnzMQAblYr8+EjC7nc1fEMHjH1Z9JOa1CabANsxeFt4XuazXTup8OenbUst5ys6oJoY
y0tXGVJpNFOFTi0sHsvTp5bEd+eKUUlvGuaEYZj2E0WIKTqjv0jBZKI/rjozzRoQTqWtNjQQ0nGN
cYljYRXmsMStumJQ9NHz8vW5jrkXOWy2Ygt2l5j8tQS8p35z60IC37eDX1mLyrOHU3MEEd3p3f+R
CCRJz4pvSRrbunrLevuukUQnfLa2BEAX+6B+p1BjI6AMkKfzy+EeDru0l/q6hFYFFu8hP7s6j4uS
UnkkZzxUhoj0gxfZE239Gacr47uC27SA9lQXEs/o6YLbCfgDqpiAIHpHQnRz3yLGkZX/gOnIzx9l
eJDGqeIZQuybiIRWnYjhQSRwyPRzy4mgua8AW6B+oegxlIe2h0enCtpNl9gsPdmmfqNO/uElLQLQ
1I7ZaRhFHojS378/YJ7n2msKSYn1GjKfuIaRvcoL7+vySSzD10yy8o2RmSEco4ZSsEYZkb6vg8fa
Rv5azuMl41SbdGldgviPR76qxAXaT1XD2N/RUSTS1nDYZf3Bt1FjJZ8sBO58i7sMmqhe6m/h8nkF
1Xs0XN9SsHF/MZRb2Qfcokvr/0Eq2uC+LMF+8B6F/bg8XGDuKLzxzadP6K7IbKNFiWHHKo98bY+5
Cm/w6cD1hnyMxak91jenfz/cspfCl0a/y4taU1p6b9F/DD+wqRi4L09wXck1yTnaPxROy80CWgzb
lO6F90BC2nkYNe3DUBqY8zdeaRqV5xCLgFyb0AVuylJgF0Kso91n1EXfNg2+0Ud96seAhPST+ofV
G1qJjF31EqYIfynabEJWx5TC2LcohAJjb0XjhjB5hlZJ7BNEDvJ/0wn0voaQdVdO5FSC7L2mbVUo
shQWgBCyzgKyLGqYI61vBPQ+eYbHsocU0Py52/izA1g3mQm6JqCPbGSsR9t5JuJogUY1dhQ8QHcs
lk+KJJFtDY6X0vCEO9aiAig03yqCQH+5+43VL2LVoNAdR5xVYdFb2Fve4BJRBVDecJOIegwUnfNl
WgWG3RxUWeq2uc1e16iUqyC/lKfa8AN5KsIpeweA2RvcPVe2IvJOEVOebpqzdrQThGz4PL4a+R4j
OrFU123eatp4ly8Jr/FBB1FZDzrCrOFlUk36pyD0LllecxyHSqEdcyjoXGOJl5CBhbX3g8SlJ3Cm
wV4mJTdT0cAPW1j7dbL73iFCjcctF5T54It9SNQO8TgzFXA6eq1NWMIy20/CaDyHsdtJ9xPvHpI5
ZQB2EqP5Xssdj1ZimYG93eYqVxwYTRuHwiXnqDPEc5qg6x2v9wAf2t4SqYGj/YR8UhxpZZ6PFlPX
AMNYRRs6Kjtex8AdKW8Pd87NLcvW6jq9L0bzAu5sNAhQqOoIhIYjVrLF1zSYWRGhqlnupBlF+QHO
HMBemtdjQQusUOv23/KKbc1e664KEK/TvLa4f57rU1FvGqFzfJJRKmskLB7GNZMY2X/7bwtIh20W
X8N1JdRVIIdPV5PEC/DlRNp/mWrYuZQ+cd8a4UYXUsfNV8JZmy+oG8Tegl67P65qrhmxL5CdJ0hQ
0IXG3XP+LejHnfe0GhJo/scFP/IEv2gMCd2DD12VRbcIqOE7F+Q41Nd/XUrUW6VY6A79P+Da2qmG
pt3Ug6dyyw3ePmt/a0B/CiUKvE8rCPEig1HE9TQdHu1ue0szL0xuUQTOJe5FSHOBMG51q19QOcYC
jgvEul6xt0BWKb602IBNOldtuOfFK8mSXyBgwj36gXyi/JzsXVtQABjR59X1LjQjj09WjXn7N3fq
1gbcJVUR5/kzVPI/FCNxIOoFwBik06F4fkRiHFo5gVWYHhgTyTy6JUUrfQFgBDaSOSXvTEgGRsRJ
ml4Up6C/Uu/tia7AyvOJeX6FTaXqDiLqu1o+hzl3enj8DhiPu9DPhJ78nMJlcTI5CBlgh/AAjFJL
omsLdE+HHgnaWwt6i6+d+x9yrL/3TXkD6vYSfQUsKM7E7d7n97RnM2mBKsCQNWn6GFh5pWLCy9tl
4rLniS7GDtOaPuWL1x36a5CcSjf2b2XXgWDVf/f659xbBuny2LwJaPmh1KKY6s3Q6mPJ2x+ng26z
ACSwUDZ4ueafan0ctkQlS4jF1T3iYIx1iYIW8ahMsLA481cOYL6KV4/5xuynifP/oArvYSGNeSzv
6zw2OVUq2hPH5CiSHmkeEJYeX8FbIca25vNnYhK3lEUckk8uuVUjGhwG01yGMly06oNWn5TTv1lU
pIWVQw9bp8YkilOlIyQQbJMv3K94367etP5ot3WXpfh3EtFqiyCReeuDBf8Rqd8wmbGyrzO/BPdE
I9eouUb+pur3zTFAPM34WMSAYcsgLXOc2njJ+CMQNDofhx3SjLwuC/ldyHrIZa4YekVIPH704QFV
QEPRi7SkR5X1fLKJeCHuACma+zZ2lXcrtPxzjgTFaIutC+riLmy/sdSC6uTX5B6u4gIZKYO/QcAx
p6/sAaUhp0HWbkm/Q/Z0lWz5arRXoMAux1e1twcO7XT6duKHtxw+77beDKJI0D07LZp9byODdtfe
5ir2sqxkPNA3yqxzgSz63KkkrGbHRXGy907XtgQ1p0VHpwuR770nto53iPOoE0uq+sBJgAskCRqM
008r0VsLGGIWm70r3DlMyopulbn+4JTrAXkTP7x1fi85iVBeEnq3mDcMIZH7z4gJLNppN5xPGqz4
TgC2AYKNAMzMdonRfx8yPOguCnwK+nk4Ln+gxCloIELXJgdaz+EbBc9awR5jIWO9Ff7drGik/XlA
8SQfwxVnNZquIIbbiA+C27/qYIdGFiOoCx3hk9UMh0Z53Nd4a4dbuYNKa8NrYqQ9wCSA5Rjd3UbG
vEPZzfEfn52oUX6u+M0ctNsE5FFe2JkjfzCN+lrBiEkvBFcJhEXXqiAWNpDXKrl4GbH1hs5GNzKT
nRqStPnJyifR/yJw1XHBtytDXr1FChq3lAFWL1RYuB6CrvC8i0Lnzp2h6q/ho47PE9ev9QrsxqiC
M9zGEvtlWnUMqFYr8iZySMC3VVTxNefOGaQOfjvcEKr3wyS/AtJJiIZZ+REctJ7KlSCQl3Zwa2iI
483LfnsZ7mroI20VH/gSPlrLAOXGyrTamQSe0nFtuA07nICcBwYj7DQ+gtSJa/owHY3XAd0bd02V
i8uMS6tTFuxdu4dVONxnOzdXKpdIgz586qjI4Ezj7UvmNV6uqx8xPa/KMUOkkZFJmn3wquhopqpq
fy+eky8dc73BmSbj/et2Hi2NZlPGWXx9G8Yt41GRbgWKe330qNmb7gDRDB+hHNmDoOT0XP8UON6N
nsozs4YcNCgDqp1oOoctnqCcc5ucXf3S8W/FqBmpEoC3iFXSen7x4MHhn+PIgAGXnbx0CFONWzfi
lBBPMU4+nkw6Y1BF+iiM7OBeTPabssJsS6TXd7oeOhIZvhL8dnWilIdMVa4+fB4Tr5o1xr2WwW3x
dBbWAe2Ec01cf71MvrScoulIAsZ8j0T6x66jrw4oJIORiMwOztGAFg2IBdLqGPNrCWrKHRhFHdZE
UwrTfQJZNgBPDe3cs9E76Jqg8/MeBGrNTVFCPwBua3i60Xd0k64gDM7MQKiWDeQpFaUMEQSLtTNk
EootsQSmfWUeCgqfqyTmG7r/ZaPUDRk6P+9z+9+hkqO3/e0M/68lU9tmXWzk2YEs0Z71S0CDbs42
p931nVrDvRin1frYaUvtT9eta6zzHGlUL+rE0dH9lhe5w7gH95zBmt48WFQVOTBB3nSUSWXn3QG4
ceGotht7qYp0oC9hq0BGnnrIWggKWFZUUEIolR0nkekfNoKlQvfONlY50nErd9rgYbR89GspCRhV
4hfaYJ4QG0MyHE5G2WxMKQrbJSO82Hmngqff9SDxOdqeHon9sxI6o26enMzYT0SeUn16ug2iYf/q
6Gm4rkMJbVzvu8ETGIyinR7AKWesjVjajZc2/eP9io3j4ifIO9MrMTclO49r6eTymfe2M606Lb1s
vH/VtoEeIdalGbTEj3wtlDHBjhDU8egZ7o2ZnbumxkGj+AVnleRCmCJwUwu+P6guVdSy0RuaBgGi
hyjhDQ6OfKvyLHr7AXjLPg08JB/PHxl5xzlpven8+WBaTZUgAHcNyXC0SemDL7i4VPLqic8ir+i0
F3DjE6Cn3UqiNvxQeWy/hbBVt4YuMQdmdH7H/rjYRvbpqWF5KiQe4SPODjOu3UsjmeCLMATnBvnQ
cNpxkOYd/u7WwlpL9BXJtryWkIil6Top3eD8SW+Mf1URN5nMszldZ7UtDs/vqC3eq8YOrE0IyEVw
z9+eASl+Zd7uU68dbmzvyGWXi4aW/EzprHOlAzDmAD87QxVzERqETKpmgNk1D8Np0Z0XWxlIfX6y
/lmJFTNFaSXdu2CmTy4km5/siafTmhJi27MK53JCPbdnivkjGFbjWlNKnEtykSMy87g36vDVUdxK
TxtBKfTVkbiBg3t9XhanpTNFIdF3i8vl3TTT7nrsYXUw/wxSXEP8xBuxNPSHxEvS8z2nKk6SyOTf
VfI+ygAFyWgZsUDir38y/BIk/Qo2n1PsfNjojqJznjtkAQE21qJ6Jb+fSOdxVmy0j0P4Y9PXv+g0
JSTCWfjn669CsZ7S/zKon9rE099SBWCCadluTCxhSzFxED8d29WECdZ+kcQeklKuxWwj/v8/sIMo
KIjkD1z4BE1ZfkBJbkiu+OGpyX/d66lFc/IpNnpAU0ErZiwWcg3rojtR5cUyUnITTUhiyb9IbAZl
HpKsEISqA4vPQTFeaThmlR5LkcjmZLOcrQGuNO2QpAJaw4KI2pyEyaF8cyXrns0sfJdZJB09DMNl
NOlx2AgWQ9u24QY2fPPmUeSSH516JNBQgjDgbd+gsVeEzrOlLjjX1+Mg6YEsU8DyPfYIRyHinUeF
LVEYqsjsVQpZ2CnrvxpQgvKQfDz/jS7jx8IuqC/33yYR3+ZiJAo5GFZc+S0bpF0hzBEEcau5xmuO
15cjgPnM6nJey5sUXuCScJp3qCnWzG93aKh+Xbfy/uA8D6LuLGgGup9G4o7+EVe6JMo0Gd8CRd7M
sQeFN7rSFBvWtDJJqJkVZGoWXngIEGyHWEiko8TSSZghBoRRVUCRrEHDV8H8o4xRR7R0JFxv/f4W
RbpAoQnhmDbknx+lVSoUxUJRbuSMzKlWYo7LpW5SXncrNVpuk+LPvd7rSo+XpvK2gaXoj692AF60
5CQ18KVPMqQHORwrj0KMKv3NMy0SxiRcJ0zVLtNHVV11e5xK/+2YDkl0LrAKoNlNP30VU/Josv/s
XfDuxn/jA9AkN1cl/Y5cHimX59G7hHHq/g0YvTg9Fe95We3+/qw+OUcEQY/XFRUYcOR9taoi3rIh
vHp7o5WBZWzRCXDpC5oq2kg2EXVs2Zyeqbg+jE/YFCpWiapa4bzPKRm107+anlvGCGVrlM576GR5
6yBDFTbL3nx0ZroAaVXF+BV1yuoLZ07YczY9tdiL2Mlvux0wAC2Ii77AhAqhT94y5UULhpenPaw9
a9Ku6LWBjS08Hl+w1OOIWJL/DS+DHGk4jFqnL5EEwZSboF/4yXmDEYo9z0EIND3oSRrxfAnvF7Sk
kNwMOS1HDtmfZJ7nCTSpf7FwyYRfPPAlcrj7JfjjMLhK9ssU/+OJJtBdVyTRj3vHmwVJIal9fjOX
lLhNNGakPX9YUUq10ljyIuuyu+MIzxcz0aXw4o7bNyujmdNJMIGS3Dn5WyF896IpJmAxCaGj4UCb
S4Baa9qcL0IVbRDNPOMVWPPMfG7rBVrDTMnULNu3nRj5l8AXiaHp7QYso4hZV3pIyckUxmE7sYVw
HDvhoC1bczL3goCj7sr1lJmCInGkeGXz3JlnzWmVrcuPmFoZrvgzry1WTJTwB3SJ5OTXsqN/Vobb
YvUlXuA86EG03AGxdQqAJg3kC1rTt0Jaou7+Z5SteqgJs4TV5zfHB9jTrhbN8xybsrVkIfMHSZv6
pZM/dbVNtJlel7kBGw+gfG8QQjxjVb81pKYQFgTicFFcHzNmOa0lT3LhJaPfeBxFvkpaVrgaHwPN
NEGtewb0CM3M2mQ/4jMvW34T+oRH1IO570Vx+MRhX5mqFSgCObHbR/EF7lL5HhdDJeg/vnOL0H8+
AF+Y5JVagF+feIsH+rVJ5H5KVrLngwivW/18L9XMFoAxH0/RpSoobV3wydZ8g7LCJfX9zwTv4C++
v34QV4Mr7GZtBw1mxCn9nvZo/fWn31Q5s6UvmH2xgqnqstvZYjvLpacsISrAsarJvDchx3FbVNtf
QXh0XgFSwuppxrBNg2Tdh74N7rJqAdNDO2+JJ2cUSYRElTaRyvnUL4aqvRj5UMUiQf+9QG23/hlG
tZUC4YZcwO9++znkRqM8EFQbB6DtWqneUYvN/NN+qXB+nUnLhFkukcL5iBc0sm2HvNmXthMkWmx6
uFyUrITWP4xgh3e4jbMJTTat2v1fQZfUgyf6evsAUT9asUmLQTUoOwyEPDGRA/J8EAOgdq/q8EQ6
e21rOD4kgmC0Z4BSdk2gOULq6l8+61MFr9/DRJwTsNhy6S7ptZeq2rLqMtplgLZX5YgeK0QZtIqi
1YA2YQcQP+TdOqtEgcUZbPABiOKN3lPB0TiguQf0bxGG+d2gzgAZbTy3ODbmmEkz+BxHjRt02xug
TdgMVUZ60J/jlkI71CiDwYvafzAN48AqyC8WBlFM7/WCAWFA88gB+ZxzUJmKn1MH6I46qkqkq9D7
64LZ+HKzLgLrX8y/K3jtyJdOkBXKmvPpK8+M6zSKByy80dE3HCrHaeSYUS3+m2kbbyrGyJkX5vm4
GuiDB3bQnzrqCHDhjRxxniY0z0AH8JLIGl7lYhHOpmbhhqe8J/komsqPG4wgUqVpKwnUB6bVbi6D
RO/Oh3BS4Avx4zZMjX5o2k1+1anGryv3CAVMzjZvHqNeU73VoH4Mq6cCYeAUMKZBa8Vu0wzrwwqQ
2PeiglrzNSuKG8pzfok0PxGpU5MKd3HTjbMdQMqAv1Y2JLF0QUebSqwkg9VTfPuZac/fT0yBcGUX
0utT4uxgUEY6cIJAIvfVHyPzJSHvAWbzo23RESog0TePfi0uhmHS9Z197H+V03PZGJDQJigxl9Zp
2l6xgaOunDMpP9livUijQEipJKf9o/0uKkocGlerWgUj8W81hYP7oVbHpiAhk79zSEBi8gxNf8BY
OEzaxpQw5NAjjx5HVshwlhO5MOPmG4P3I4QpsEeU6NRhssND0DqEvoXipvfHPCBRzluqB78pZd3D
ZJs8iGlcypsx59tSxsqqCXJtw4g0FRq/U6wCnK+BnThKeKq8RyCFQS+hsudrW9sRhZDFfaHbUyGJ
JfEGPkFGlYxWIMswA2aCkhfaDbjckKS1Gnkjikm15KaiZ3wgCL+Zx8XFYZmUv8veqneyBFvTYDDM
UdbkbVABaKyHVEo+kBYNMOotk4ArAIfUeA+osyQUDQUPfwzgHVoxVZWP5Y3gHY6AaLVS+7k+OXVq
coPjwuFYCkDl5sHuVslm1TZ1RNEQuJlS4P/WbkgqFlhQz+ztEE6vmVLZbXLhVPo0aZAaHuzst634
yYiiDWR5O0kM+LHMvE6RGXna/zBRcrHCTZj8LZRWmc8kJRevO22AX4AfhxiYZgzOMZBlwqqR9voW
gecAVfKu3iEovDirD1K3uxqYdqZLyL9L/KC0MA93IEz/tXzFDDryjLXo1vBRZzTmPGuuJGBOAbmv
qZURsTgTRxkT/w9qZruicpq8KkhU4hUN0G2c0Mj5dUIS3wsQuiED4am1eViV44BNbKI2PAKxBv53
XAvIWYvQ2IK5JpaB9imZCeLjLBk123YP79iSnXBClUVOkWmE7j8Qu2EBuELmv2i5Uxzhf12WklIt
9JDuEY7Z2xc5hnX1D8Chf292g6txI8ecmWuaDGc2sXYbH8eFRsuW+dY7TSGEnCnvEFkyLadss6H7
ztHpNKG1JRUCHOo80y96t3YKb7jzJ11pRaRVNP2eqxlm6tyxchif8iaQ1YXOZHW91UlUCT8J51fH
fd60gxWZ4r+P75MCEwm8xf6BuULZZqXiiBAjZkp03J8ikTwkJrgaoaPPzI4VoQ0GdlORsPj+dBTq
ccIvp6ugDyxj2V+TqZOG/hdENYcP1T2TE43z5sSPZhjNsQhV2NxyTWWSnoFmdIfXCxNPmly1vlu3
nvtKso91A/aRihbj4ftt0b9TO6wJIOkqvaY91VGzuF+GwDd1xnqaSc7rWAPcJ3aol5+71pNANSVb
/GlpzXZULi7aFdcdC8cE6aW2kDZWKraJD/Fop9RogcI4Y1VTvu1ZbVSxGLpZBwxaQ83YYjjbxdge
elZTw63ACHo7zHt1mdmaV1DwB0FJuax9OUg+JeHRoGCb3FWV7POu74NzVXvjHT0gGEvocTDHE4re
vef17GFRNIDuRLuguEfXfMP5OxVEGRtKTwwq64MXpzwbbCJDb6gVvjhmu1THviDXlQMbbAUy7OqH
tH0L3HcNRjGkHu5/oZSPmqcmUEoUoUugtKbMsZrdXyY8IfL6tRXdOapuMXQgFpzbmbJx3rkaW2Bd
oLHVgHz7iWqSHz6JW6XnZbvIAbiWh9p1PJcal6RZ3A/5aIDWtLReSzqlVg88VC4I+atTlmT3eB+i
qxiCJf+++/jYqQxKqk34roTe2F9qGVbPX2vyieDj28HB5HIYX5uBhZ67ocY1Fp2W/QUr9TJRtmGb
7sksCIUl4sdBVfUSmgMy+KA/VlmFaNh3ezbNwNKzhEV7dh1MGhqIGMHjaZI6jzXT1nAibli3+0yi
8v416+6dUJrQZIs1z0CpJQdTdq3E5iqeYJvtGGODmMS9MpiA+sKAC6Ic5f8g7zqRHKT7ZasYOk6e
69O/2YRr6jnUieMKD6YuqIcWWUxAMN8SC/L8ytUoARyiblzvAYailmGywstkfNNHySyfwuEjmFJJ
7wDgEoHnQHAXSeYIcpCus5o5kMaHPMdfNZghIQ6XlFcYLw49V3HjUpHPaY/GrYje/4wKA8qx7qKJ
pBg4fJ3DTYlIRKxNPwR7amVDGUInor4UrQOqkZefFw3z31a99UguT58ev6lYtVfLc/lu4P61ogmD
BerZfgr2ySDb71BsiD0WPD7yvsaqrvBsOoZafjrt2ywTrt860pnzVl0loccPuWfjDICUZ5ju3RT8
R2VOgMIt1TcApX8APpVKREJHomzEqcUcCiqE1OBm1sBpgM1E8vCfHwVEVyOZ4psbggCTK4+yqkwZ
u++4XTuM0Ilhh08pgPhsA6WsUcLGPwFjGOOjpmnTGM4A2PFMYO9OI73y2v/azKTygSHOPB0u1FN5
VwUdDqBUMzJP+JfirqaHztH68fhJGanY7AST7nfljdf+pUFLLlBgEdS4sWP8JIYuDLw4Qmpy/SDz
yx8B14btIstO9LHJfnUyoUUkn1OuzkJHZwbqyWny5VBFePNky3Cow5wiHwo9fcypPi8HiH+DGVOv
W+9FsEDgcSr6iAOFgcVS0K7ic5cO9uQuhPp4V0c4eRfSdTphX6QdDrwLNT/i60sYm9Wq3H3W/KgK
zZS7YKn2/m8H36yFmyRBkTCOK1TwItkfFXFVaz4sOok38ZJbP17W4VZzaBJblFhpKJKELlQbiSjR
VC61+Dd/f0Q9tjiH34WoHgMF/QwQ0mdigr6cZFV2qY/9s5IgqwHpqeGs/D9FNhVozeF5vF1OEJ4u
KwIpuiex7wPgpGnI22JDN42WaZyPYQpppKTmHFgfviLhbIbqXpHjDHN4ddH5GxbODIt3fUrt3P6f
x+Crnhop430GA5M2G1UT7SdHH2mqKD+RLHLjrDbwWNKLwbsedcBZmhPaGeIngP7vzgP/uFiT94bd
mQU2a9pfgSE2MXGkllprectWq9+bUyCBuB/217mPh/NAWvM8eHk+3C7ApWWiPZMGUY0FLXSDOFIc
+fJhdhJk6Erim7oPKQwzhNGqOWGSDMFRQqwjGwzhdAQJO+gE2fW+JnvDTD1vU9DVVl70cS0GUekJ
f1VgJyBiUf8M9zvu+e45bGlA7GciHLmx4XZZUsW0YJKY3XG9WPu3tN99obKcTPMKLGmF6V/2cBo4
QnRsTpxycVBeMXxeIZ/f5oqE9cKdq1xDKtHpSf8huc9h56rzlcRf9qJw6EHtgoUo6aL0Kb4UibEM
ckc3EYDYj77W1SDsTANptYvA1OYyRQBqA9eXlEcQbR+ktwFfuI5oGD701A7/t8zBOVoPzSOGQyOo
/U3wbR0WzGw3ltJOawJXX8b/C7IQOnECYkqUl1JYVhvbTqgd1jPPpHtm+n5c6z2NHktOueQFMEUk
AXJ00J1lm8BQljeHJhHhVWILArEsP9dnOQ8iANbZuB/7xcDWFZh6Tx2E4KNX2w450QXUPysgq+I3
eiGQPGnJ+EcVBeSC5m3PPNhM0/LT7U5I07I7EwmnentW8PjjUmN0gQbGLSU+zxEJdlVsf7OVNLAC
3WQoem3WSNzx4XgYe0MZjbPDb+jzk9SkaRS1YQGY8lxnW+EtLuTuQ5fZBRQ703hD4isorEyUGahc
Ru1kF16HLCTDPU72DMOv84cYTxJyP1VylBCllSny2r0wf/Lz5swo8mSrebjpBZHc/q554SNNTz0K
ABqJzFdwa7i3glkO4do0CQT6WydGJJYHRAohOcuKlngTN8R1ho+T27ASciWaecpI3vtp9Hr9gLTz
1VlIGvkn6h1xfM8Fv13is4SDeMLFyeUSTAkhe2ZA5lci9YVJ4g5Y6ggFukiXLIp37V6wzI7CEyp9
MXcd00eGsx6OuClRvlKKi41wWuSzCiGey0q0KqcpXBQREmsfjJq4i7SIVKYTX/DIK0gekW2UigaX
mnmb8MoIbPQBflYuWGAPU2C1ab3cdsvnHLO18I82lAaHBHHnAe8Lu+9+7mAPDSZWs/74mEia1w41
RA1Zl8gywJpXZicuwfp4yeHBREox6G5D2+0ZzDs1ujqS1DfefERe9U0BMLHmoYls84w44gRaRmd3
bOZNoL+FVHoVIF0xmxJZXVoEQrIrSC8bH4mZsEWZrZnA65xt678T1NkeXTuiaBeuViqIg3Nxkz5o
Kz5waLsPUNQh4eXNx3iu3/NKTcMzYAHTDT4zO3kJJKFzwoHClKl2ZYqq2ylPxCgVkvyrnc07dR3+
wM+ZXZZFfgYJ+l7OV3+vMcit2kykONhWlYjursiu2GMlg4z7li1B4Qp+Aq+PpzDS4nXKOXuwrwwy
KzL2N9W6JOBFVAgW9JrupjmOgR2tjQpaLBI7esZKLtW/H8adfN6uEhzLPy9gReg8KCJr4rFZnNx7
3yYb6Nah174GNa6FJMD4F8ursn6MTUXbLwj2ZYQxViqR8pdqdMbnzvZexBNweNr4L994ZUGdkLc6
zSVAfeoErFiKVuWudZkMm1iWz3xwgPk3rexszbuvhRDrY2TVHxCohOlTys0vR6f572QaiCLmu6oD
p7g/2zl53tWgJxlgqczUmFZVgYa3HY7O6ErNhoHWYGVwetnb2r02ih9l5kIIOeZCTYI1xXsFgGUS
eTsKZnc3xZPUVo/eFbhey/UEc5Ya8iXExL19JhcX7gYVVQw5pZzGd1F6ZcC6N9gycuK+14pU7Gt3
6XQ2OaaxR7VdEkUUQX92VGNMvU09/3Cn2qOp6m3CZGEWKI+vUiYX+xwnMNHhL2ygBPNU4ZCIAKUP
td4wsnWAS9NyMZaBLJ4ggjO+rg6Wd7TLL9ALzukfZY+2WbMvEawflg8LUlR6hs3+Onbze8W0t3dm
woIAb/K37Sy1keWoUo373/19y5sybSszAAo3ZeUEsNTrTi1sBq4g3BEet9/2vqYJfCSUbwBqd/Pv
7YbTNXaK1viQNNjVojcb98tM/LKEgJsFOxZ9JXHdMeQZEA+q/vn5IG7bPkmG/QUXTmHAmrov1ntY
M4HIPubZT+st597Ky1+xW5fNe92twBIJgBb7Fr4hcO1uV04d0nynsIeN3PMebk2UQyHWLAnaRcpy
qt37ah6N0mKGMDgIpeJ+ALdr3By1pBfMGG7FOucJvpGaTcOOG2abAR9Sw1nxxHf59mSS1h8ZzXLJ
HcqB/Z7V2ynfvUBoCQQmCI2vOGZeYPVVQEQYrJjq19mxeVsqo4CgurIHYMJnhOhLedAZ3lNZ5PaO
4vmgOl5CiZATYfxB3n97qumAyh8LJax5SA7Yp9iMmhRG3xAYAN3ODOpP3DhfdKH8XuzNk1BkRm5v
h6lpx/ZlLiUAtvmC/yGc/CXtJoX2uktFDMS7MmUNR3h+ppguLFb0w0ArMqewZ7UZOwJUvqvLDpSG
ACQVBbf1Bus824V01M0wg0TEKDuY/1fZCiJ0gb1YdLvD7KVYRxZLBZL+ID2x1YjdwCXbqajY38xs
MkxXNJmDWkplSyrnKNFnIY8xT15Cy3zwJU7Qk/qnokKjtM1IVk5Wdk571sXkf6Oqg6Imeg5vEDNT
GB2kjWYZOHEdftN4yUf9hwAVfYKGx9/F1AIeywAKVNki0UFtI6JEQ56imHLKMaExNINJiuLOwp8c
SPzDg9I+MqYa28WIMzA2KaE59aql+LZy4QqaPVvJSVpko1enP6iZP0n+JyTnxLckgh+SD+bI1C+L
2WQmpkYuBX6lHoR9PpfSbLbTmVvuvgwmvFgQogV5NpnV3JyVcSOMEVA7w/zp9wC6IuaGwA6KLUP0
UNxA1/yf3eZKHzFh3yvpCLEL8AWU/ToxwIi7gsO4+ms3THzlijcNXbx+ZHb4Y1G8y3FmstlwB3CC
p4QL13cabJbz/9K4B7UiaBOs0SCNpbIxL+32kVi5pSko5TFH/Gj7ggreT6OoOP8aXngJJ85XdyvY
/m8bsqBSOuGETYES0Rgc6Aflpgtgf+vNxJ6gS5+nBMIfXUVBJIXAF5o5x61hL9d2TP0CbQxj5jp5
dNXZFBTOmU6q9/XMRj6m0u+N37EP0++Z/3taz+iVNebDIuafPnvucRqtBd1FebkWwLE/P3BcEiTq
v20tZVXydEwWx80xcuwlUQIKUrT9zRHbRM8/5bXtDpXRvmwjOelP+AWNGkgqSatO9B48qKFVewex
1Tt1nlCPTVy5RtrSLHxzMAhJdqEAI+vMYnrKPouTLa/MywZ6YuCb+mGr1/N68wrglrFccGBWUNVJ
Y2mHikSmnGZjTI16+fNwuL03Dfv3ohrLSytRzZT5Ky+mw0l/mUEiUICmjorj+G090VF6VVYwn5vx
fcZmewJjKF9pD1KzEDk7b5DAm8eNWpFgNRL00t6PE53Pn44hmmDRSHdi/igdqQtdXchfR/vK7Z7Z
rBWpHAg+CbeSoWqd9LXTWaMvJAnXo/K7C84FxqFRXuMMiN9xr11q82gS3acHnl9elooIrMkgJWQa
fTzaNfqPquVFKUW54sNO578Dk9BbWhT+N8mkI02aCJ5RYVJSeW3xcc4fwkevPIdHVsaB5Hzb2LbK
4LitzbfmEBwsNncFl6q6oO/w5IcdgRfVQBci6jOlTLGyF/fauTD0SA+Oe4BVafDIl7ZNM6A4O4ti
yRL41RFxtJtL1JpZQ8xGYSRJLvzuNH64HseQmtONKkrOgRpPUW2icqzNhUVu2DN+0ivgzXWEbWAr
PHvol8Ws759M+9hbUV+SOrjgpJZ3F6pHI+ucDO3LWN6M5U3rmnRP3rRvPI1Z0Mznd5tvh5+CPY/7
Pwuja9M9DzagVV+7SOa6YtPb803RYh52K+PWJr19uxOJqCIMSAfSnlcGrSGBLbmKd37jw5lsRwWV
0sKw1HudbdjByEmQVcYSPPEvo7i6SssPnOfx1+v7IcB2YWmmqefD9SWGgqQhytJ8GNYLo9IrlGVR
4/c7EBHOW4wltI89UFIlUp68swFSVfAZv1fFv22ODnFIPPUfC9+4hvz9VNom16dFFyjHWR3DaHYu
W4eJtqkdvORsSRwuvu0i80OBzD89zJ/8dfsb4/Iiq+gWXv2OVqE1PBbj2lpeFk8DaWfifqejqn5G
UWG/ozSwdfMNity+YdBmcHwKZY7W6+kchWu7SliroB7mEBH/l03Ys7E4J/O2cpli4HLgTIMoyX/y
W+v22tNOlC9rDvFE/hR5D6THL8LNDXmq5s3/mgebNfw2rDb6SydoAM3YsCwMwMklrZLegYAt8dO3
t1ZSFxeNaFXLnKfP04NGWYrRuSPTpHMDSAcVdpVI0gKnwblX0dtxJK2Ae2dz1nmRNDcIG7nGBybz
kKxIVnC35XIFi2rEB3uGYhyWHIbX5pfTicRpIcRlXYH57FOwYEro3vN/ydlJlgE0RgN2WAoHsMT6
KTRLLz9dTsSJXXeBh5SbKjxdNb6k6Kj5vrD1THLu7LErRO+2Q6/3DxmTt3eAA5CKATRNzrWvvKXq
UgJ3350ZxlAoPXlzQyTKUydYGRb0exmcY1Sxsz7/1nOvHLe4RmYubh7L6GBae9qkshmJPYSuFo4N
MlxGaSec9w5Qx6v8RpqpRAbexUGfvqgsdczCby0eZTzr2ew1SVNOXMiHT30FB/tJv5pCXnI6dUtC
d9flgmc6/SwkIPLpqKM3QhuRr7t5O734nDvk4OdsHNTY8hWDEZxu2PrQPQz8YnxYwKxdFVVuI6zD
g5YfWrpWxdEZMJDdbwtCizsSSTAqfzC0NZBsZ15fsi8mR/YqXJz9e2GS7ScCzwgy2C88muYBh0fa
l1Qe5oYHGbX1oVhkZ24YCOLbAIi6GFP8fDkCttV+tdpJ8b7suYbUS+pUV45nA7YHHM1z8EYaAEgN
PF3pvB7BC+mA3UX8fulZ5ifss6lyQMLD/dsCg8twzgLZhEAkcMIlZgSZlzKANGmeRTf7sZ2xiwmx
i30ksGJGjbiABNMnaH+Fp3o6wO2s2aPHMSwbv/D5L2yfH8trP1cCw3gtPVtsRjOIlGZotB7/ngPE
l2KnCUbI/qqoCndBO7SEO296xC9Rxk+pdAdHcr2axakQS3KDwz4413CHqAxZLKIj4gKzYz3XBkwo
IlxHYTRMIyjilT4rfcv+njVfg4MyTYYNMgsDu2DVex9I71xV6eAWxu4Br/U9UyQ7LAXDxF6nkt+y
fwkcTTrV7Yu7/J0PUqAmAFSq2N46AhPuHEpGK1lwcyaYi6RqNn6+EHHW/M+hu2heC6dS3I+FbF0D
kKdaGHqkdSGoEEwqXSAvSODJ6L/HDuFPgFlu4UeLzi3C3MCj9UyGsBjUrNLxIlFSOIjL9o8s//TK
xq2i8AS94xZQoxIPiex2hoQ/MVAlTALDTMKA8h9OW6y6uxYzH8cu/65bC12d77gnVxMVzKLLDmGG
T+qbsem96qCkntWqu8HxgQsvFXKi8r/q/+2pMAEzSLJyOhvM9yrhW5kipCf/ul1MWp8vE5CVc4SL
5SO1tNLzbeVl+eZ1kuIMkUF2BUFchkVWruOrOdPP3b4mjj+2YfExaVBuG2PQFkuJRZp9/47m3O8G
c87YIRNhjtc//7zMd3FZored9AF9rx0G36ItvTF2R7Lr1Stx7TmPw25Uqkq1X3ES6MIWVUfMZJGx
6YRFjrRkpm3hDVkbez2TbmIQn6vJuOu5P+dWVhr+QjbnnN9orYwDR9C96Bi3Pr8HFGDZNd1Zb7M2
QzNEW4WQX5g2cKVzNeWXEdXh/jAR1NJ3xPZcFJwZYc2K7uz0/lPlJjlygiCl5G6oZIGJU3mXpG5H
cXY2SxfJvyI6JTiwPbsN4F78Ou/iz3Y/CiE0NSt9IQwgvNeinZzGJYUfxJUu/zSR3YjZ1lLPNbCB
WeT37MuBAhXlu3trlJ3DsU6NQFnOtSL/6/qb8WgPq9gHRb7qrXhaw1X+FpTf+69vlbBlET+18eLg
RrcnybELupaRjkMAAE7mCYMVImsNNhLg3Rdb1YZ/4b7+mWOAKFvvAH2+6ME+70JgyVBwpZp5UODs
GemuI8gk11w07+leA/j3e40HZgTaJJtSiSWjIq+arOV11uw931YUqlHEPWRjzX6ybnfMh4RQe45n
0IvoRcGlUqCI/9GpSD+fMq+3aYKL8Kw44ht7nhrZ88ZbRvfHImveSlLHqsPL3nl3qgRJnDNBT+Vk
BoTjtl9SvphfuBGZMBZ/b6hSU6DxWJmGLuXGJIhrEVM25NCsE5A0mC9XktSJ7i0fZHpeLubkf9VH
lVHqY8HaYmCtMFWHmUM+a4IU0C1bu2SbS793xjP7sw5xMujgPc4hw981TZUXPgJ1k0rpqrqSfvLh
pTmuDQOsiw5+1xItqJ5vt344AfYC4R78UfZzzliSZ3029GvwAj6982vGPYJBqjbkLqDKCdSF2rM7
T0++0kr9n+9Zw5SCUN2p+ba5GIl2G6Mi3k89i5dYRTZWywXPY+WGoYvYud55um/SJQ9anH8rONlc
2XwpwH5mQfYzvJYwF5d0UEjNYei1SNGFy4o2jSbSlF6CCzQl4JY0FkEFEraG9WveT+srDNWRCEIl
uoXgoF39SHG616pUa+yNnFYVvJ7pOhRFRPG/o/dr0iuf4yAEbytBl7LacuXPdM2tL9w64bPhO+2c
UgQmlWbnZ1izQOIdnknMmRufdF/GL7khZK3ezgPg/GfSwP1jIw6CFI8zyml98pkDXAVsq+cpJ085
PWWBmmJF335uCGfYWvamR6SC/Gry6HfrUKrrySP5strBnO0bTZdoHGPOTe8TZTNK8mDHrQXV8Dq8
s0PNMXSWW9pe1e8h0sHETtfa4dIq0d/5ZUltJ8gSIO64mJniHY5N6Sv/HUJMwQG4FEiVppN6x5fv
p9STWfgdyK/MLNFGrQd9Wsaq/hcnN2s5JByTn41e0DXVTpwDhfJQM5tQFq3imHkxXMTXhY8ufdku
1RFeIQpDX5RaOQrS8UabPL7M8AhIOQS+3MYOK5zJyjt3zb6F1JhO5WtKSFb/w+TG/1AE+us8p31w
vu11NJ63H2rBzi6dCiNnEs5BHvcvklIZGmXZUeSwy9MWAf9vRZ7frN8e/qYUhu9L09DF8XodsF5Z
8qnoNSTxRGfIk8mGJOycdCyVokaYjC6mHFQZ9nEagRd8fIFsnvT6HdtjEEvhgJ5KUeTRZAnmHqba
chRDwxvzOKbDwt1wgSeARRQSq4+GUDaaSkQwvrVmkQOv+CU3uMjX1/pP27ANIlAO0N/A4jyVY8gG
gqcGWKojoFlJr4lZaM4co0jRYuYGMge4Cs1xI1Q3VkbAP+dOruoeoYCBNgW6QnFxL7iZcw9gv9el
/aBnwvaZ7LKDHS8hRydmrvqzhXVNSmZulcmZkpJLcv0WwHMdYNEJtCxZ5CTNKpkDWVUySZoMXFTR
hPxWaCvTO42qwwXb/AZ3DSW6ebPW0jALO+OAIP/meFeMuWryQh7HxI3uuOhzW2MeEzILcDLVW5aw
IxmqswgKEYF0y403zSuJ0vPgn93mbWS8vlpxVr3/1Riw7ct0WJjUnIsjwVRApq3DAC8j3p51qrXf
YKPSLXRn1pVZNWi5CH2RftPV+qhpk8CYh/JHDarF38orMVQW6hRQEKJtY9GbKT6xIjqIYniKo7Qx
ggeYBXEbdJugJIwvnqthNChWKzsW83YYl5ZaxgVpVJUKRX1HGSvGpPjERE3Q3hy0NrfD9HSPf0KJ
RbXe2figOHhm4/t957KvPW63ktHJg/ZXNsMe/caaAVfSxjgMKQFrQ8qlgXvseBs0Tll5r2kBonrM
Hi3csZgzXoTwASVGZSYWIVieDhNXQzvDscmX8yUpXsFkTZzwEw16oBuAPNIy6kngiwwzxMXU4cUk
HLIW5nk1ATatD+FBd6H2Tcq6th1z0T4jgPVhy45aI6RLFMMd+430mmle3jnPjVeBL64JrUQMzizR
sx7I4F0HfoJQc8qGrkyOH/cWqbKWUJuLvOiDk14QO8KU8B5x5DI5q8hlhBz0PsS6fYeZs5pVP9Yk
4pxcC9Cl/uqVTYtd4SMwNIxLWwRDne/2HRByvnvZehNbERwl3ZdIyt4tBx+Afjanucx48BvpXnxK
o+GeTrcTID9Ar6AJTnfnaveDuPSwKUixqrr6x8+gKEsqlZkZTZA/4C2tRiArgvrzpItVTcJd1gfz
hf/y4ZJRaXyjfin6RPUXl4Vuuu2Z48SuMU1ncT7M8Tcm9ARWKIEf7a2oCUqmVrtfasfDGf9nwdb0
kmgnqI0iInDV5bMNTtZ33YPIOGUkygZyxB3N1UJxSJUBgqZYw9P3CUz2QZqYKjwDSwF0oL4yCRX2
+IHL9vFjsOgTz3gEOMCP6YCYAGY3unc4Q/3eC6rwgn9GVdDtwfKaBtpvcPAM3PgZCJRSVdUO/vHT
2Ms2FekmHvV6xSQZmuTtQPgdP1IyknFhoL3Z8zJzk/biTNBQYAvCb5LXVf1j1hQzMY3GezCvOK8d
VjJir+warDSW4yanuXX+olkqvM3W1QUWGUuy2PKugufTZYDqEZh9yIOdXLkmaaLDXmwXl2MMdYUG
LgFNH9GxvS8k6afsAZv62dLxJAIrmEeV9SnVID9g4yLvVUJivd7pGuOdcCiWwJ9PFtxTzD3cajNs
eDK8bUJNJgfODDBQ5EO4nvczd2RCH6whIQk8O6VT2yO5x7RpMhEOQENeA0KAfudmMs7rjLq99Qc1
oYUIpztXu6SzOE3Ot1PfR2hy8Azq/jStD6VXG6Ag3YbkUwEoyvEL214jcXRRorjZp32Vz4fXkGr7
Rj9jLWUaKyfVx7edQWTgf65K4h6gmXdeD32TRtLjaokj5pk7VfgJOcxOeQlaU6D+QvsJxy2P1iOr
ulRlM22K9NwKsKUxpUR2bzLYuEPuq/9pRymtdULeuO0BZKLSGdoOY3SQ4H76IUH8KF6oUAASbsCk
RpBApgqrWZz4/FMzi6Qb0AZeiUqWWDPf5xXhr7gnLZzA3TbW6mHwYFUNM7K54V3Wak9IwGDTCHrO
vJU2qqePQqh7qULFuEIW0evK/tgV8uuCRAH2inkz7hLQBMafUuPYiqUOQaBpGO+3IAQGSx/lAc0R
Ww/nw4uA59fFHTK/zMv3kJNSoMNW+uBryPGg6mZAsPQy9wxiDQUWLGwMxB9LDk/xn+OkTXbv6Lc6
1/U9gdUz/AaaUu8ocFsWLIhBn7Jso4sVgMQk1tWZqRrvhZ3O140f46CgxVIFsoHgXmwlQoVYEURV
fcF/dSpHiexr9gj+7KgHX99fB8Y4fK9Y6lA7z+26WZnJUcA7Nbg/8Y5QJ8NcvnEIMUmZpGODgNxj
j1M8UC+Va3q69WgBfaEE+oUBLwABiIZaTL5WSp6L29ntWLhC5HhELJH48o4GlAB32E2ou1AweaXZ
6sBnWi+KY5jwGOnfh3pJ8mNC8wCvIbI3FxZ8ptIuCbo4ZFJarIZgTRbWzHs8zJtXCoBDRi/RNwg5
l1LpjC0CHZy4UxPbzlxjmLvYJwi65+3WFDo9qHammjf4w4ZHZ/Y9O1U0Sqss5Ied5STdwRB0a+Y0
bUABfqBYvwd5Q6P8XQOtfWCbmwckqGgzlrGkT6CFN8WXh2X/RzA9QLbBuI/TaRmpOAwBJYkZunPD
DyOUG/rddbgrnjWSpLLNBsdbXI8ZNqlDldV+Smq7j7qW4GcBhyIlbNZCjDtpF2XDAXCQ79/dIQRE
/IhE9prNv78aI0BsSRYDRo5XPc5TCUKsxbXgFCiNnleyXreQZSnZ+9DMYqEKLmMDzOHtoWFY4a0f
pM4YLrxSDstjQhuGfgtKVwjqdb6gtQ/AoZXmI495z/z/+4nHzf4nVpSvu0WRlLzFDmzh0aoUfXsd
30jKhxrpBeXFrHF+I2/akbGw5l+p1yM/DeK/FsAIwLBrOXOvC0XNF/OKfwvZMzFxOLEdpOLNPyFE
Nm0XH3Wnnwh+i/NJRA0DS6OaEjvx0lSdTR35jF99gw328nZwCxbE1d/gQqNSUNINcKzrzL81KoGk
7/FCAm/8IDfzfGuePySJIsIC+6AS3YBYLsGp1/yADfuE7NZENc00v30/ITolnP3hFP7h0N6lXH6Z
f/3lhEgJP+QG64Ria56MWneHgUXap6spbAHANS3SlMQqj3xxLdQ/Ac3/ka++BvvGquGhiiuTihY7
TPi6iwtI90X0V8H1rcRoOEvoJw53fAgf2sztMbqdgWLwJ4EqK6aVrAr9pkhAEtHC4a1Z10+34E8V
frUA6yDiswx7Iz3HHV+7Lv56Wmc29srNXwqnfy8ZMJv66eKHnu5yoEiJcrwfUeFmdTGCceYtzwGC
o4+Fx8431mQfFFr9sA9osDQvKqK8Y9x7rF/zDLCri12wyR2lrl9LrDcGbp7q5h1zMkMSteFhJYDN
LK0lrR7jQYlzqcm0H2qDMZwGXttc7/i6PVA9dThmZEIG8Smqs74R1OVDilvByljOUXgMsHSgn5CY
eRZlbTB8WbwNVuMwNZXq0nKFntB4SQKtCLs2I9hZJpTIvyKemQXEkYlICvqxzuJdFs21yqrdezBD
4cdyKvO2IaE42yyTTKJHOrMiaCO35RRDseSZSV40JIuCRgWvcdejv3EKiMBU4yYeXqttbmI97FyX
NzlMnw0h1Y6XvRCSl7kZFloympzpWVLVWXhMqYHmeORxh0E87NHXOlOuqTuRDXtllOPvMWASNP4s
THtPNdmWJvSaP4GOdYA9ignUgMIikZGR/sxRM3lj6BHCaoTPTKszSMTPRYjFCQokzoO1LJuwSIud
XFJ7Um0PNpOs/lQaEzNuNay6AvziKgZ0fP0kt1CyNCZbcXaHUHuwAlZtADImHenqP2iissy6pf3L
4U2bU4PIjscoiTS2mu/Sz9tTJ+IAjnJqaH/BBXKgACOR351IT9/MSFDL9t1EKSQr6Rmn0nulcXKp
MI7+UZT/VPezilAp+y6zbdp0QQI7LXPWxuKrdAdgfQvCQ6fBCwla8BM4Kge9fncfOW2Op3WVPjnP
hnkBKxfNvOSX1SXt8pV+JaKUj7CjQeRy1/37Egzcm5yHechDAjjhZSxjMkDy9Tmua1sQ+jYUlAPJ
boHjr8Y/eKVT8WBmSMF/G6m7j8VQxTRm7u55rGLe8nCaO732L5FJlo6OLvAj7AaS7KEMnoMEtxLC
Rim4+SmytLzH8QefbuRsIeS+DVg0ur0Tg/qUYDsQLRrX3+y6ngH3DIDKpixhgffQVHs5ZrpyVSdf
Dd1ymCd8Zx+TwqyNGOFEhEeQBXCFraoJ9RJFUGM7nweOziiaydt/yHY5Hg07H55BtrWv2RK5B5K3
7PgYg931Q/r6Qqi4OoJPjOvFL/+JXtnjo2wgiEBINtMmAE1KejeMGdiecdQIOSQp0Q2JRiTWDJ3q
PFGy25LDGzmCnGP22SO5uHCRe41rnku07dxOkg02siCaMdMM+RmOSLD95jijYMQUeEcQ+JbRRkDh
uJ7vZ0ye7qOkndEFOJYnqnUNnMZ+xbFW9ERQ7/wS6p9FBbAQV+oe0GcE3a+L3g2DxHLgGNV7xUJ0
ElOZI8eH2rzEXRP42TXvyto4s0L+MRk66d9oAoaUas9XaSq+51Y1YPE0H9uja8YbnmmzYKhuTt3A
z+F9oiW7H9oTrmLMxyWJl/q+2091mB84jmLhHK0Kpd+LFJ8QX7hKJv/WSU6kuUZ+qOm9q886ISwB
D3t19MZY2uNsGRsyXhnAQKBB8Q8vCn61IfPFtqw9jGFy+lPGOYn5TFMcabnaioaMWqH6yyDTq9lT
SFOBNiqJeA2j0F26gvw86BLio7gYWgQ+LpMsjMLiETMvsyMV3xeRmhZ+lvHS/CB54nsCTClG7cZc
5Z5RJviUj51gnnes1pPjp/7p9nk2B/Me9O6D2J1czVOc+r6RE+FxVu7vo3E1ZZbuVP3bEt2AgjvZ
+vzpc71w8aDhSWjraWqgbcLCWK2k8w+56D0a02G6G2HTJuFePB5PloFzfrc4uCiJEo+GWPbMOW0x
2ZiySCdhIl7EyCcHxfAhKhi6YRVGjtAZhsAx4Ucc9IakrwgM9Cbf2zr6lfV/D+9bylULw8C+K6nU
za64bSIoTE1r0QQW9sLMM3JB5ass9ybtYAxOqkulQMJYkpT/G1Wq5+xAsvoQhy2lV9Ur3HT3rAUF
CBDTi3k2ZahmE7YY7Vf/ZHUL3sVs368xmvqBJl/Y4tt7RWTmg3nUXEAJbpwhZqv6pxpnfNUjIPmB
eHn33+mlSE8G62hs7jFhN7E7BD8ASbONU9bCIZh4TDow2lsRR/M+yqfFHPepr33kUvwIqqqDHtoI
xeBidpKwXIoATZqWWdOLrlja0jobr5VmoCWylpC7Gx8V9LLSOsVa+yE49t/Ox6sDqvUVW6A8IC5n
IKYXh2wq2hFR02gNnlywtR3KT7bNzcCVla5j2dYgEd1kiDIBN22xsgbUzy7mLfOU+pHpSE27u7S9
Kgg3jf9vzK826bPqnUzr3OZ5QwXcuJoaFiBQMDDivIi3T7j344a+knhWaeaDa6sVkkLfImJJMHYD
1miSGYUqu7J/Zes8vTWCx7jSkqKljUWW2Q1SedpHx7KDu/cwXZCz8i1Wn3deSsjejrn549vtJWzA
paCbGMY6vQ7FLBc6wreYyq3VYjlu/ZVbtW6BYiMr6xvRquowYBLtEjuRTydeHO0eQp7NuNB7CEEY
WgDFL21bEENjh/KAiCpQMFeEmdFDwTFrYIoQ+UbV72blJhri/ixF03/f8KKsGrxfyorURxAPbHJ0
i0lTD8e4dba05isZT4AzgdCgpeWvy5SmOFkd4EJaloJKYsu9fNVtMww17KJLdyq0VWqTXZq6fuCT
oMzKaugbebUuX9/myHdyC8po1fxDrfXDnFJpJ2gZhaUrgJvrRwzRvazGuxaN4wcGJ0zz9t4cq3z8
dCc9hmzuzdWRQZgWWL93gSRfWQuxJzu/Hmzsfkgs4HT7U+jUUpY8SHrWI99g4OxDbZ2QR3lOQodP
XLa3UT9J4GvO9WWshkaYpzf/7ohNFBO6+zr8o+a56JCd6ggERp5G9psPLMQw5NmHpTB7OJYGMy0q
UWWPLB3x4ltQ/2VqjCWZwyKCio/ozbJ5zS/34f5KU/w8pFabukW7ndgrXIcDpeQOqp21FKDLGK7M
4G1rqJ+bnxVhbvPEg74DbbAChwME/+htluOi9c6d895zqDncTD9dKnfMi7lwYXtFJjELw0vsXewZ
5qRgyYdfNTmr1xGvgLyPgArLOe7fP1WcdMKfWudV6LFMX+A2OrzJV6WxZBQUDZ4CZFgeOrugvrzW
ob6EbgTYdfraZNbhEGpbtu7OysdkbwbqG9f+C1oSDhqECsvp2z/xxCovuuKSC4KE5BCkMGC9xktE
Yr7FkjrXj/bvhZZz3oSeJ+Pw3wgC7gJso78Jqea7kZr8pS3WG9GJpqhskewdolmbjcCDiTEjAN7Y
+yfUTDQ/wN97uS7nCxMIb/QPp92p4Cgui++lso0TxJ+jrsLucW8UZo8H3jeYWHRBouWB1NHPpFpP
hk1qIBepXC1dTKiUs8WFgRvrJg6vt88qW5wLLsoGxNbNUu1Pn/nVhFNNpvoLi6WPl+6uDYUxt3g9
3jeizWLGtnl45+LB16SP2PwGXtvhYi0v3sXblxbiOQMqO4tYkxLNP5p4M9wubgE8mm2mZAAQ7rKR
ybTScmLXUx5yUKSG2lv4J6k2GepblOS5HjQi7Oy3s1MtZLsqIdaMB9/PrMTw9/te9n0yFaqWM6h9
/B3afewpttmX6Q1e9p11iojuzwO5F3CZhsCzNVohaSylNHr+4bbD6t3HTLgVH2UnJLWF8tmz/vLq
LS6HpsdrV3hq69g2GOffG9MC5NtmAG0RnunMWRaa1VwACQg/74z2vFwxVJCNcx4iMfOTrigHOJjC
sHcKjy3k+O6BH0fn+GMGjTHdo15L268KjabTlFA6uELcwfUZNzfvZhFznxbZjfEt102gxszl4DHa
04km3hRHKkNPVeYbhNpUYBqV7XmiiVzK2nTRuuVE4HJOnOmkd45zZ81nP4nent5rDB9U2qY7Gf4F
N1ZDqMLdeCQgqMC3F/c3vOEWkHUE543EFoCBVxmtvuHF0UtcXqq70E0HAI+zzEnZcomS1m+HgTTo
7UNtZmNK0DK9+soGRuBNDbmdeP+G++m5x4i/ChCzAFdawpESl36ZfVcy/vIMOriMNFwPkoTYfZvZ
qlNG1csoT+8j7NZzrgpv1Y6r357J583NTcxCAT3/hHNxZo5qaNJm8OkBkUH/jdKhBZ5/D82P+lPM
dMsySHM1UO4+ozwTH2YMo01tU6QVANK7k6X754a9LQB25o1hpM4GwZskvxxBvAYKVGb0gO6uo+KI
5lJIUzcG001Bqep7UzlwH+j0WmnjYV+MppXDwTfWHi/QKnLKbGyvbGDYZLtxMA7QWPAootOYOMoa
eg1nbh+8Td3bsS/pZdjTfkXNfkQZm7glnIK5RCHy3hqbAOf5SLgSOaqQDJ/P8sUVo8FL3vY9QtCM
PWMLx6FvcQ/JvXAPjMRx5fsDRa5yaH9eljOmCBnlyNxj7f8s69SmQ0ORokSJW3pNf/JJs+vERuOa
FYEmJypmTcGkhyznEQlG/V0hpi8g3Fthq3nMUB3z57ptKbGzduzp3uw0yVpK56WknMELcF+q1DRj
uko+YCB7gZXsqDqruLbpoHwVveJ+KG1HfF+2rps1KUAI39upRUt4NhFfWO0o9QgPzWsCcl81Z6Ob
YrKb+g7n9Knl0x7XL4QxiHdb/soe9KLtf6RiHLR6wxlDC3mJYLrye6drOSYcjuZIg8+b5beRKkQn
okXEEtEZP9cqoquWIsT/rSs27zzD4RBRVG1C2ZOV2HA8DF8XKrxI1mXST1ktCKO9r1sWsV5Ki/Jr
NbmQe2J4Y/C/sQGE50SbqrlAuxN4RAeXIPykFiHRNrfDEzeLxoYUvob846vVZYRic81m7+sb1FKV
kVfSLSayXB8nAWtCuYDeHJr/ViuLi91qygw5iEgHz7R3mlLdEWqlyBECf84nEm3XU8d3NTs6E0tt
ldsPAefPr5qc2ABHHtNhydWCABTJNBNmvoo2ldjBslxCux7pVQQS6F37ljP0VHmZiUra3lNtnR3U
NglsFLj/Dz1Myi2mFnY7C9ZeXL78Nqr33ih4T/9/Y6p2S5aY+IyF7yIPKxv5YGvGCJ8eW/b/tEM/
lAC21hKUe3CZXUCGvJARy/ppaDnVQAwCyawD1gWc4gKOWYk9Fr6VyxMqukTgRT0pVUQyM7gzhcV/
ANXio/hdSdsjW6ZDU6+Hpwcq0x7zZwFl6DuERiqRkS4yaONZKF9pwOysGXNzY4qShsR7qI5kI5+7
zeHxgT+VVgBvslbVFdmMaJWcjsIU3wIoV6tpvIskC+ADEB6X3hTxsNwN6jPQtrDp+bw1fxiKcQQ9
G1id4LKp22v9VaUvOGCjX86sv0XRGPDsyh/jKhHQ7XxTuwtt2TCV69hjyXAunqHuIPa8FWIFHd0u
Gik47wyQlJ/B6+wDqW7Ci25aTbydm1gsNKf4ad6cW5eeF6tBtosUwHbUWZGm+8ICiFwEonxsS7q7
W8o9qyhTDGoE8Fd8mlj4ZeyWaEiofqNd2ern8cYAL/Nu1LbV1mCzC1upBscI2+oJt9gWSp/cdb/E
KMeqOdgZKsvcxSLfnWdah7MR5pcV+EZXqTurWrxvOZdPrhTLOnI2ndPRbWcEl8ZJU+J612yMc+zq
GiEEfVRv4XRohfFWoa0FY6vh7yN7aqm/mjULmCj5sJmrvXFapThZKGAPqpdMgopUkfE8GmQNV0ZM
ym0RQD0wUG0Iu2irjgj7Dykz4GiIMPzzRJdCrIUt3wqt8AgIm85GyMNDemF5u4QzRl2cs3q1UuMk
G2QrWle73zwxLHwIO9os5XyShFh8Hinj8FGths7AkrDDHmqYNlteOkuYn5UP3ngI26e4kcqwR+HF
DtmpVKwMDThOndPT4PJG7ez6xnv7OgOOy08yn/vUQAaFw2Vs239/OYRpqlxoBV8W66BpzWZVkIXi
/qWUxzymWwMFGTo1LbqtiJxphUWftc22CkSh7ldVC9B5/+NygmMwKkyGCYlf6A6Lf63gIx1q6mzY
kgFHd/ZAA6SRTD69bzSMhO9pAItbssYHAAgUUILf+IjA1hn593W7gsudJc+iVV8YBx0pRTFRhxQO
TkP23lG8kPTPti9SgcoLhg8JJFY9T4ve/WqvYfvbOj0VRHyYSj6RSnK0RfES9AFGmywModkXJOTA
WKZMQuM5NLVtINnlUQpdYTwt47C41AcDFqpy3nCFpjAAKxzmPj3jkqz+ubpnNzZF2FdsnhUNb4sM
FYYneQ3eU0ZDCJVpgNFq0zPlvWCMqV89pbuaqNP2WmrSvuB0NtEiALieC5haTSqOJhCuTdQ35zlC
L6EshxGtXPuOPRuzTh1PZlUDkm4RfyDRz0pRlyC2FCIahcxXBJujA5bP8QoUwMrkouNrlz3SGATN
Tpk4XS/Jg/4pvoHDOm4aQfg5xKFcHcYSZoQypQc/kZG0LnBBEt/22SEVxpJ1+og2YuykydYx/bjC
FiWGbm6e3fXU89bESMNZr8oZfush/TxdgTwi9Pk2LOGiOVlVqsTrqXlK9hgwER5T9H0tS+YLYbTp
tbp3oPAD9x4EJs57Tbm8CixjZBfngmaZBw/OZBolhIkIP1l/HcONWAj+yENpfkSuKezS3w31FDTq
y/ZcMWeU6qqDYq8n/sMBrZ0D5T8khLSX3bAlbgrzb4JhqTmgeFSzfnf/ZPMNiqtujB2dBBRKrYYp
KODXNgkosUKFrG8otisMs+Bk+gsSbbiuleEyNWYi7MoX4Q+CeM+MlgqkW6e1plpyEH9KYbXue/K3
UT0wYHg6DV4Lt9tVsBwl+t7OiKqvCxCkr3sq5rjE1/wQiiBEH773OuyeWXjCw9SvN5zdPRxjJNT6
BDveTiq+CSNWI0WV4kKnILqIMB2zPXpFHDJ83wfMzc3fS7WW8kmkc591T0zH341WhG1Embg2tbq0
GTHtF2Q9zRxfqME+atkDL7TF2phSe2++X2P/WMI7v/ZXsdgJcBtYTMjP8MolgnNJH8ktRZyjFoo7
rYhX6rQAqtXMMyyIJ9UNAWgmHs4ZfnV1e63RM30dQd+19B7n1g7+VAnndq/Gqg9KGX0SeOmD7wj3
Wy5fQr5uFJ2VVHkpBxbq2iR+XCHiCqofzu4o66SfghrT2M7w24+wA6WO9qVC9S6Lk5PvS9fbjo2u
Q9JPjsycgABXFRTduPFngZyNdf7LEQts/JFbhiMGNRLOx72qBIFaOtnq2XBDn1KnC83f2LUsbwYH
nDQh9UkH1SIvOqzfEmK9kJXvbjaYUZnUgfGJsChL6cB/W/gcanrVv7U8HP/zJ1P5J5JyKFgvpr45
MumQGByWnSLy5J4AitUYd0LE6138NLdz5KPTZHM+XOu/JcWa4OjG+XCDhbpqUG4iPrPlSinB9AkP
97mBjILW3MmOSxRFVt7OZbOtF+HV+slgVEfitAA27dPPW25SkM25f2plNskHOc4N6jmIV4TECeYf
z55/97FDTjO3FoA7IIH4GWtQOW8CXKA0xYVJxNdYthZsnnkm/0MfSp33UtQ88U/mJVIwNeMb06+E
mnms6TVBsCyvjcUIduLIy1gEa9KuXx5ZGMhbqbbNrfWTJddxkS0sjXJnUe1yhRjCgVFzj9rO12vM
mJlJGiEoRcQe7P2VMHDHRrca4pJbSAHz+seGm/PaTF152CPHA2cq+QfT5X3naFnaeCmMeDacbqH4
Bh4t/YlSxnSN+/xJxM2ARvHvxb5GNVHGcO4ib40MOyewtozC8gIie0wNdfkWgvBrzOWwdUriJXhd
rIaRsGsvHv37H1+D8GpBi5EE0bD290jPkiQygCAAPLD++rU5QMq/v7Rw1OamEzAZJsbVPliP6iDB
bhTONCRT1XBj+oiqUcTM0riJYZDauzZR6WKFPAL554bf7xuz+8f+1UA/Hg+//BA3KHlObK/KqAj+
w1X6mRD44rhfQgEh919XJKcjNDyviccJwAgdAbTnxiI9O/ooEbafxvqzcn6Pa4o9+vb8EsuA5Wkd
o10gf3YQDz/7LXZLRu0DYJ9AJFdvlifzJVVjips9tBg+WhFPlUlNMOy5bfwy6Qpf6w6I+JsodwwO
O8rAuP9t8f5xbjuQQKJ6KVq1k+HPSusOLe9wsI4CuIxYCk8XHKUCbr4tJ2g5BuoKsQkAGIbVDjc7
9p+zzruFS5tD5RphDtTcRQkEHeH5nSbK6kWRce2leQJTIih+Wj6M0pg4vTFKn2TrgIj0hzKSC/sP
iU5kko+4l65XmJvHntQLcKZ3k/VHFBdFNYJkyeN7iZRNVcCp+te/BQWet0EMwRXnQYfec7KYdkrB
NEgm1Zx1s5bGMmyLpIOMclZ+/gBpxVpT38726RZ0LGm3oibC045C0i2lh1ecWYtrHy85bRtzt7JC
+NJv+Qf6iKTKGMraOhW0wbge+BUm9sP7HrAcWB8lITysVSCBHoQLZVbnkUTeTWDzvG7zykXNsGop
1sbbk6HBq94+sovP9/zJMINV9sDWDY3cdWrmgjWhTxJcCq5lAqC0EWB0F6paUAlV6LseDLuNexqs
kYD1XuCw7Qxji4tdMPOzscLTjpnmPRfTbvH8aSjDCEPreMLTu7hGsZ+rb1mJqegQECsRhYINoVUy
QpjK0yAfSSGvlqW4rim1HUU8vuQhYAtu1gfnCtVmm1fPInunwM4QnPL0ac5WVVG3hKQ5Pj4gfEjY
l0+oZ0SmMM3GyJ30FyvSMUK6JlTkCh+XBc8HsX5U0+ZVNQ2TU/vmOLOk8c7Yszo7LmBSpDta9o+X
bZ/YY2lXA+I6aAtsH1kEY7xcrQIEXFBosuFewrSJ2M/BHBOK/00sZFTicPWVIm5KCVYVL+qKPxBs
dC5u8Z8Ix85NMHhEpq2U0ox+X63SIcz1WJaxRoH39StitW18xtMPStaBiQ7OioKIfAO8TS750u43
+E7CYyUJhAds3NWv34qQYFjJWk6dBdCVuoUDgSzX9XuZUVau3Ms9+rMjOwWzFzgOhv1s5m6LsdVy
L/retDEIQ7bAYdSQhNVxvBl6X3mfqrlR/aGQ5JD5RXBpcaHYlZVEd5WniQ4/H7hUeeBCnwEiO/sO
iA5202f2V2JNvsiIiUd6aG5rIqpIZs41o/G6X6SVa021ZjtpT+jbe53DEdwDXFj9bNDd6MZLJnGS
QEj0VrNiDmJLoYo5KYjGIEo99njmRw4Mex+5YdKSNCISU1DG2mb+Dy7KsoQPapSYyop18RE2ze8P
K4i0tVc9LlO1BNwaXU4TPuKbDUZSsR1G1USUMTgGuFg6+P1DCnSK/8qnZrhMiiqMrTdxV87PZLwq
Jlv10leLPoX87HFWZEZC1QQGV6aZGyuItN9wc3I+HS8TkvJxGjXOr3NQfY7j3gEvPwA7KiHysOiF
mMy7djHQlR4IzVk2QK4ulT0FFHL3ksgdzff9uhTMfwuwB0w/Mv6QiEBsSzTvAV5VIQ0gbz9LKmcY
Y/2zMoWsVv1mzMzW3/ZsKeDhPm8TE5ssq3PcekdOMsSWB6pNOG0ATj6KKiH+PYDGAXp13yb0bKLP
9v4WWfCleq0zTuRPWMeBrxLih+kDlVVljXUxiKq8jkjmZnP4gcS1LzH5Jkl8AxwY12F0U+7f5VHI
vQCxWEr83d6bEBRF7TJ2A8XKoBJCAH+8qm70IzUtj5H+cxFJA8TsxKgHgM2v8KPoqgRcIBwh94dw
12XKzzTtWo93+qrJiZ67sw7Sj46BWmyv5QotOMQKslMxV++mG1I4k7Y/ySna7I1OD348HQ/m85OJ
JwjCrVDEWm042kt45DvuCChc1sC4dn5tfE9f9GMv486f6VuWRARF5u7DWNOudAqp500I+OMZeI6J
kGKj0+sGtkPdt3huExUpUETaPbkRYe4H6NXOerLbEuQclSeqcwyFU5oWptvimaiXCzLSavofDo3U
hLJjLYRlXRjyBbdxOvig5/q0sfMiliycAtu7Q58niqr3Dcs/piWR9ByJfuuyMHZtT+Q+/Rh4uTNt
GniRNucjlBx1eygkBIi0ze9l727THCbUwp6gTHbezGxv7wQePYXcDATWT3mwuPeKbDIUpQcwIcvk
PAJJPCKZOBy06BpINFsZWAWlbM3i4tXV/wEtbshhjy9FKUPQ1AYbU+xT1KrcqZt4lMslM8ASHCNH
8SjNU3vM9ptgYRimsMqGlJCSHlh8rEA3hI6Xl9obAOMtuRqjelOdKrTvUOBVhElAXDzCojyWA/kt
ijRRypbXaY4pb22jL08AUHatJeyXEs/jt3OABGQADRMjtuGOvXnVFCTpGqWNvpje4z8xbaigH2M4
U+xyuKv9I/zvnUZ6/SYTGKBFRqc788Urc2srbIi2zGfVdRortlQss8IsGCy8MjYqBxKZSx2X3+Y7
1Rp79U0Evk06KLA07vfHmbL9XRGWVbNRl2QJ1dRh3vjmZp0cSmP4aLQvIyDDjqrGTWQUGqnoWqnh
ru6SM1u5fjDBMP3vsajP2Egp1LDEKlFMMeienJZm5FvIPkANFaNU3BW03L36iIp/1bu3x7Q6w7e3
LFom0n/yZNu04hWmFyd9xEQzXuxIwR+5AOKUPy4iLbq+094UZ2j+3FAf4mwvbFaOYcnQ92rvABOZ
lTkiSD8h4ecX0+VDLUGtOjW7OgLGf3hcGgKBliIkTD2oL/+4JKcmDfWdqwfd1NfqcnRNU8ccxf2s
BX7KXvrzjA9hXz9vpEPMXUZwPUY0gyjrt1HyGInxOGT5roH7D8ei2NZh7jqvJDJu+PCliSWVMCW6
UHKL7EZ/9ybnK5GJFq5Rwqi0OrLLU3Ui1qeAZc3JnaX6FhIUBBpk1+ptvJ8R2M7QuDKfV8do0YTx
j79qpvvMH4L2UXXC1OyPzyN0i2toq6RZFewolM6Zn6BPQi7MjL5WYSaCpf6i8MPIzpRd9Pez2lTH
xgCW4aYsAbbDyBxiZ0lLwVCRiITXAXTiRbDvrMQfsyQl1boYFsfwNlQDs2uYNVs73ovtGUIv9pXT
byiTWkOcddYsB3aam8TWrYOBUrsiy3LQ2fAT+1vMec8od/Cu6zOBED6KbV6c3bvxErPnNwI0yIYJ
vPdtDZVlIx+KMuGMkJ5IZ4lln2uci5jtvGsTeDe91iUJtns7Da46Xym1p52iPckho4zXFC4mBFZ9
MBtfGP94QgMJbKzxKSHOGw9gcxeVnZu0djeL+razhP65IHbDFC9LgmjOYiuSjjLDkC4FyOomzy+7
m+pvA9zh2xClr5WvPk2O/zy81tnbbXJiKfocKGde2YHgocghlc3MndgtF62seVEsW88SdGVDTyRH
nHg98m2ciXWwAUfhoDXH1Zx+9oAhvG9yMMUJMjp3E5rZN2G1ww8hZwKU3kq9B/W25DEqq17ECrEv
SZ7AwZzaUROQIgo1Ng9w1U7tRVHqKLwe/0ENSu1Hk9RoPdThcWlvXURwg1R16IE+BTFN1eOL6QB3
VSiUE8cCv/97VjUlakP5M/Oyrnq7tiXaUegM2EdyE5YVX5tO07skIWKy23cF73uejm7ZscNmPa4z
lDkI9GyYOUQN7HW5nBOWYZpGNsYJCvmYXsmLiuCIYiz7RwNk1sekZxU9MMPfRHCGLxyHrIaL4h+L
/ZgEIX5pNK8pODzgWBCPk5wQmgAVEAMf0jIgKjFUkvjOFYgNxiQVaF7Px3mOBWVD2M6U5RqBHzy3
Fqg9fA/BoolsIm4WYw4Y3eJuRKCwYrkz75UkdMa64ajag1rXaIsOaQoWuCucMX/FgzSv1DDq6OJv
gpDzLUb3xln7Eb9jKRjACneKSrgxKna0DR5mI6dl9lTLMMrwhdQ5jkDknxHRlRozgCH1w7B30OAV
uC+2KngOxCjdwLkfugfTjYF0Zsa51euXRzDO5Csn8cjafZS2pJ1+QH0xdNZ239m8dmkVimq1sdmm
KbdbLeJ+Nbzn2xFc7N2UTMKUibrc35KVY8JrVXiSM31u7we7j7ABF+Hx8PuhkNzKtGivXagzgPlF
bTj7HMPX9/xh3rcGKe7vPMWVFuwGsoSVgFvmasfL2aRyoyzCDRcSMSUuM6N6RmKYBfD0Ae2f2p73
14ZXPtepm6Zw0rbnHgNOIzNdFSaYPcDY3QKvGVx5tk6f+JB3vMH/MX0Cv6VQOqovBXaLTb8RelGt
cmwqoGrlE1JtF9mqs+KHUtIwJKOvZcE/vURDefc5fxqe8k+rVKxG8J0tNjMgkEV3eZyf4dAEI02n
J5nxBPHOkAMdr1A5itAYe2gleMmjoYbT4W4wf0i4EH8q/cPx/PGAv8OW42HBfSBBgzHAFs6XZrGx
XFiMPQvPa+A5o786PORigVbrK313sovspR4fMtO9yVAbPRd2OnjyJAE4hKw84FlOAF+Xm4E4EcX2
YQRoMEZdlZ/1kWKH+KL/duHFk3eYk0qtNl652AzEiK2kMy5FsCl+eDURMmkI6UCgolvgq8Keg1mp
bW154iDnYVv8CZUIwJTnG9a4Kmjz5TX5Y22/YWYfKBq3J1HWyWk82Y068K2CVeUxNmonxcLM3ItJ
4TvgRwR87RLTwJTm0K7nQS+xQ+1AqrYeqtQecfiHuHifGDp8llSD2wOXlRoY2Mb9OrdYYcvo3FTX
xICGfOh1Ikyfh+ofSM/zljIWksMvVQ1uOq2xQ81sTYNxxqA5r9soqrZ4dUmPx8nF6YmSCGdrKCQ+
1WRMY9O6as+gEpY7LVs+thOTi1GHD/z5Kzfi1SmA8QWbcuR6tAlHeVxPgKaOdtgsJXuErWfUL5rK
fSxCKqP9BHUva/dgqRIzOnj0VmfAAK8ne0c4qRlpJ245xqk59blerHhGzETQCkavLplqYrHqYCa7
nVNNdh1vr7w6ZcEBIhrGqqQ1c8LU+JdrItiTxCcLcevzH6NQ1/5vYkhLvpYgQvqTltOvh2pY259i
7W00xN4zGoOEffNaewxxi6jajWq/T3GECVetfUsb1pXSBIFTTNZNaeXCc3XywXNaPMA353mDRB+X
CaQ1NKBcPZuR624YCeHlly/jOEx0phOfu2Fi7Qxxw7n/Vv3/4bBBwcex9QoCxLzFrZg6983fCrG1
g3yXxN6uZj71wPH4SueRZBFh5uepBIRIlIidncfQg4wN6vc7h5G8xsuymHls5s6zLBINMKS4eFUf
bUlGz3V3iDc6b6fkvSPwM+7IbMw9/96tDmN5GCwsGvzojySyBk7Ex6b/SNMOZG4+7ZEFywwHPEZ9
oMZNYXCcCKsodLYzEswGA3dudmk3fK++wF0itc8bK88GcqriQPG/NV94hKH/yPANv1e+pzyU9N2h
SDvQfn4Jpt6gXRBFCbX2iA62tJ6jme00HtYUjS0Zu2fxi9guV+OB1o9592rvskI+2AVMrtJ17W9M
Ca2bdyig4w7NZ0+yCVjBIvmrF+40NeN1ycg/0XcwPEz72twwNbJD5JJZPb4QiL37tFuRdKzJUPMh
iOi1bbm8+HiDmUK4pLoiYBvSorBDmLb7r1hrWMW0BA4p6hdPIV046EA8l4gFVkxG31GpcnftxhdW
0D9ytRTugRSy8Ke+TdmOKiSHlhjTdX9JqXVW7BLlHbbvWRTDIMG0ldK4Tfwrq5JuP0pid60uaFWf
NgCGNS5OkjHfZluPEJ8jm7179P9zv0FS/B4dwuZ9cr0hOg3pAIdDTwPwzYaFo+Kso5mtslpAgzJE
sNXbKnZHqKvLj5JOtoOpOEZl7+8GP4xZ3IDbArd2kWYvBaN3KDOBBPRgXxxAmoSn8AYdU5A6fL+Q
QSviLUDXT7Ig++K64oPINIYdubv3W+fBrSMTaFdvy5wJovnpemE/zHu3g6QjEssVz8+Doc9hnHE5
5KEwrF0Fc3gzAeITP+F8LD55CBbFt8ceNxoaF6GWYFmL9QyFgCHYu0PmsyVrMmH50EYqAmpJKwko
7F0qNCJabX8Z9+sKQK8sB+joG1q91xYMT22wV/iV5Qxn0UrJxSnEXWQ3HxAkZqOEB3b1leOVRXI1
eyj6T6vEeKQtFgzHfHCBui+tQjIaRiXdu6ZMa+KzxAW2Fqk0RJoQ0VdO79Rx18Z0Ax/vutfJO6Yy
nmR6Kye7WblNPxpRZ89jd7bdT3TiBTUYADFzXAiK6IzHc9Mmd2xf3JB5zLm/TQ0xrGfTytW3QoTB
hlihKTQGnWauLvyQh7IS0MmUTMGdHZhHzo6UEnCG2alJhGUEc/kU6L0ppYkwBbjbRJd7/EjEiZuK
XqkRFNir8TjxjkEsoZG0vt4sTHGuBoh1gMCWR2BKW15TkmKwiaQkKWPwp1/8FQWyLfcp3dyo1uL5
Q1oqc8dREAk14fjAgt483vXLatJVMDG7dV0mudAjE0c7jEcSjmqZRrXjkvYht8SMLp4asu1zyDGV
E7n+DmdiJbdh7kxAGRTvEog9oJPRRZjXy8itO/9JnUXUrnj5PONDIslVE6qojt1l5hb6p7jN+hy2
2r0VMA5DECYYrmEeV8SGeBH8F1n0qXBGxFTThih9HRlZ1sexFH0X3RuARmX5PTT9IMsp7sND2c+S
7ytfdtJI32bMWM6oSBdshIqU6Z4rN4XfWrKIPSxrW9F5Hq6ScleMe0DHHFr7YTOjmHL3iQkaS9D1
7ymPKPQl+9peYr+mnV905VPu/vzryGB9W0prQHM5cfHBV2UkkmZ+7F8ZXKwcW2obJM7yj6fPUnSw
tnKoyVk+HuAHEnkJIyaXzIMuapyBdi3eZ2Q5MWzHlm/7l7DEXYXD7sgkM/3AoIvDH/v/alKQedIk
HqxzjOwuf/eYDrnvZkqcnlVVkgthBxMENtVj4Y/EM8oaBWQxHRsPKZfYmAUPM4l3PEY1IkrgbsJm
41yjQ2Z7NM4DW+4EBCXn3dNddDuZv3QFp9Dbsei3TD6ONnwsebmanXBIcvvrt+5vyE1CS1DWq6Gr
m/1RtdDZg5+6ROyRNID4GORkvztVhjTiAXqoXLs4RnkZR3O0G/0NwPwJN99AIhx/ZjHRICSUqTgf
V5ESrRfVx9meBOgnhZTtcSpEncgdiv1iVPQevjevmGUK7f6FKxNBQMyNB+ufMZarnP4DGYTCIl7V
cfTGRpTpxHmJsesm8NBTQBrVhg/q7L/8ioTuKlvVKNx5Gjq2w7BLAPIuHeOUbNmOjiTQYGquUjj0
Z23tf3GVPdZNA36GY/CV84Qj0O4M2gd6Zq1j5gmaJSNy5ydeKxCbCZqYbYA+yJEXTXIwdr6LHBQK
+b9qBJlyzdUfpNVJrFNfwr0e1CXS+HZ+rVk9exTCo+NL3CFhLvv99gyomZ6LeAw/7ekC7Nv6XF7Z
uHSGlG/t3c84YYuDAs/lWSvVQysF63LKiB8X6URqcmAJEdbesZ2aX7jGaxO60jIQ/GA5lsDbLy+i
VXiTPIcJB1H3SIMinHsVHSiWreegCgdKS8klWlRumAVFv2qqD15II4Q5ia2sScGHk0Et+QHAo/XE
T8f+rHvUIoXE30FHlsUfCnMuALWWZoAsCXe5UuQIeDikxFAOky8NIl2JnSkmFNtdFf9tZV+tsx0B
SGjjXYzPaeLKagZzvoM6HBMVGPy1X9yLBZyVl2KYWe8yAG5uow//kovROkChJeueJ5nB2kqnVa+E
/hRHo04QmMskifBkd1ztZQwpjrEVfLbShzp8RXBUK5TxF5XUv42h7vW5W5x7VxEsj0Gqsy1jgDbo
n0aTs4J2qOsgsd7m+b/xRjbMV4tQMOtoSMNCSBsVHqxzZVvlscgdRwHnS1VvEMQQRY1XTqDuTZaz
WBxbGwM+e34FyCjMVB5REXECaBCuJ+I87Bb/EjX0J//2hZNNCODLuIwwqiZ+EkdHkd+weI6eSWkO
+xlQyBQzy6xcj9Ta233fUK2LuFUwCNeh9uort77TlLbWBKgeZrNo5InCKyWbj8LAMwvB/7xX8lB5
RGg6R0gbv7MesjWAPq27Slkc4IzzOD+/PafBSaAeOTWXK2BZgAFidmY1Cw/5s7AGejaielOADHk3
vEkmes/yAZNcR/4FdlohnTZBvDoJvneGX0NeFm505qGOr8LNZCoXZ3B4+zFDmo7xL62wlJ334bTu
fAs4OTJ4MoDPV3BNF00UNIwhWPzoSBBoxDCHzLkde6zuTce7OHFqmtOQ05w1GQg04LXVDK8PsQWO
VIAE1X/r1dgJozgUOdGdziuSircwknNnAjvLm3lJnqbS1lrGOFjK9PPLexfk0nJwl4/N/O2WcrVH
Vbwdck72ZTpf8S+oV5Y9feiqRm3BHelyWqAkpKN6yS4RJRPZ54YBr/Wrpt7LyL6WaQXvvR6Ozudg
4gmvV4kt1ywbTp0M5/9xPUsGjDC8FFeW+Y8Lo58TWNf6GWCvB1DFXMbOYpwrhjZyCPXOgFC6wsif
85mtGtbTdeNI/YBkJnloPXVjAiw6PJTaiEowduugZ2bBIaLFPdrS4e1JCJjcrTJDSsAA5F11w0C1
Pc4qGjm8bfUuZGARvQHTxFQNFdKAe4LNvsW678w7FBBEJPqc/XCN47AI1lgyz8IWQasWln+fr9Vs
JJk1wUeJutR1o4e4IwsLhqj9XsRtPMWCMyp5apXxWfiG5dUt8Izm8KZEhsruLUsbKRrRsWdRQFwP
IIfZ5FMZJGUffx61bIXTivdI6sfCwExuNDU6+yVJ0NpP3nGba5Hwc8N8tJsxrXSC02LHrj2O5zw2
gHIlGWZEPXMde6GSjgKAR3e7hUZ6DJYuVfaarcOLTey2B9OSZwPOS8/rkE9aje0YpPxsHJzrjvle
Qklu2fQh0H9QI2Z4gHwu76YaZxUZ693M2V7htaOWAyKpjkXibygnYoEsxg8hHi+iL/IFVl3Flgqf
J5esR9NOIna9inS0pheCwcxrGb0Rn84ahulcxytm3xOjt/gew99vfbzOpn+aAOW9E/IM796bwE2/
yExBI9jbdaNtq0UzBwBf1SCFP4VV06QLq0g/gqGdmQoVuHbvT6fScfflR/PQI5Ej7uunPphu9pzS
YCvTxTC04eWDvErHQ3I+qR63RXiCz/UWIIqEqv0DyuvYOd8tLonbkiBn6idP7JP4jLqa3LvY+qnl
48zW1iEnqqF6IN/oip0o7oW0IQFQefAkGAMH5V9VDZtT/NPqyU2HuvAbx8hiUcSp9WfgVGNyieAq
yRqXqgUMB4yqJ15ulZJz5Pt6nur4//7MEXj/ud3gOIWOjA9ypw9K0U1qiGSzw699O9Ynm3BL6Ety
0gVozaP2sgUoL7VWe68BQBfCuxVPpyb33n247QoFuDkS3T5W39pHZdcLty6UEhdKFa+5l6lHQ6dz
6/MJH27+PIiMCfMJosV7a2Sw8c0She9wmVhWMV65RJm4BSppwjgF9oqPu0qcdVtrOcOkfTRQxV+3
chdpP8nYjXkh97R9Jy4XbNJ+3WrKOxOolm0T+Wo2vANnwGoy4URmCXQCHyxmh+P3ifh5KP+9SS17
1l2jm8Z+oXOlxSp6FGPGLtkMIlpRXW05ziAkIFEN/EPpM/ZI7a/mI5p2iVtWxdmXhjCm7M+6gItu
h+suFbDBafXQic47V9B5slHRiYx/FJwi8RRNqgcqcD5RBDvUwZPBBm4Y19d1AGbiX5ORjPpneiJc
rdzzdRYIbUWcvI0Ynr5ZW2h4icQk7zOJsjlK0yf6DzfW0iEJtujHehiV9w98a7lEKJ7RjjD4hvBn
CCj9NryAosg8f2migQ6Bn+6kVQMbfEfjm7NPFHFLjE4wj9CzKRVOEQBjawzNESACjEFFGP/axvYj
gDhlSbRTy+ReAocCoyb+ixactHdGuGp7QjdXW+iCbcUjH0fK25z9YkU+kivNimSFgG1IrgEM7+wm
sZxTBIvwMfR5IJOaAfL+99NQLPAzcEOfiOomLSlbUw8VPI2jmiyvV5foyC7+Q3dQovKKrqeFwnrv
+J/Hh6Ttt+aXnZFlghC8sJBq2agVMCOT05HVIfIc2J8XhpuGwA5/MqulKf4bhW09M1jvYWb+wZjh
2KDik7i0AFbjN/bzFLFixg++7nwA3/WAq2NPSmlCgNLZDHBpYOU5KSbEZIQU51ooq6yQMXrCFhUa
k4BxPcysw5zJB3ojxsqLzOmwRhH7d722MN1n/rJqiSPgeBSuk2Nk9ZkxXjbZQmJoXS6Re1tWGNMZ
nSu2zdCWdXRmW0hUxaPdYYBv6tCdMqMzWfioqrt0K4tKyoa+O9QaeeZ+ZBLTkGxEcjomEgd9i+0u
2E7RhOTrWsidd70mH9xL9e/SU9ozt62Y5ClDeXqeWA+jzQ06WKrdAb9hYRNg3Tm53u5CIAzKMcCl
RzYC55ulgEURDSaoc+yqtuHN8fNWrWL3ju9Z/4XTylE4y6JSGG/Pdx7oT9bKn/xp3Ztbuxe9NX19
/qygaaglmU3HFIqgUvywDZQeuoAnmI8PuyyfpvQqqYal4MRatZBeUN94xmfS6R7R7AxYbJXchAhW
5lGRbk+0721H7jieHEuekRTq7IhSKr4uQWsMKmV1MY88zQ31m0RR4s0OxagA8Ey+3yXNREwJoCa6
8841GPBxzctcXxt6wVFLwMWsajCTsOMOQO4reZ461/R+TqUE1ZBy3Ba+++4EkFw75VINxmrIAK9e
fuHTia3JJWoXjiGJD5MkKKHB17HopgLiN543e+WWRWRmRdTUxR0H3V+jc36vaK4ahq606li7ySJf
X+XP3xS5Z93IhGl336ArGCLrfIX/4yp9hPlEWV9TFRvC3yh719eBxGlhyM0v15foqC8fBhlcYYf5
GNuh5AGhuMNKUVTv7QSe88B1f5a62HN+gngT71rAByoiQSQXD8HhvjposF78AiBa3cIgLT1qq4p7
GD0GCqMz2KAskKp72seAhFoufRBC/ZQm9jxRAYEWM2EhuvrBw1hFRwC/df8YfL8ZKeSDK0ioJSSb
uR0iKCoKE+DcVyz0nwGOy0QqH+kuS5AZpmVRNI/IEBn2oc1axn9uiHBj4oOgLxaOqiLBGHjYXt1V
uP2D89QqXRJQYjI50cQaW3TBS5tFLVd61zcqKpTeLAN19zNQDP11aFPI40LZxQFR8yzbomCCSMnV
OpcCV+zQ88bq819XojRm4aaG9Rvc3cpk0Sci1EA8dx3iCHFHgnD7M9ZhuAuzEoVJ0oeeI9rPvdBg
9oGLsowZcWJst1AUvjxdAe3gqIGcmCzrVuQTItt25wwGwRvuXD1ZLoW7n+v547hOHUCFf+XyobjX
32f7N19YODMsdH5Vjnp7oI2K60LWbVNRxbQ3AdWZZsxCMavfCKI20WXcWjZ//cRO6vn1icy2P+in
Uor0rq9lqjt4goHXwKGmjoFB/QA0xMmpb7vrXMrFC2lPfI967rW4hrubjCl1suVWUaWPq+QZmLI9
7InKRsg29IZg2equEIsD2JxSG5m+nezlA/rKtWPI+frA076pCO9tiL1Lv+s9xqZ+4XPSW+SL0LBI
yBMUEu9J78/OydIxTC56uM6fwrnTyNmeIdd0FSBXWVjSf//63WbsQ7ndx59aLWqLDvR+j2X0mLF2
DWPAa0mrafaJafaWJ4M9nIc1MpkbKefPhKG8S6wNW+5tpiYnnKHiXHbXeqFW70LU4SPY6nQn/xAO
SPtp12f3vc13jrJDLxfrxYWTgvn4QK7X4nGUqPfhgHEsc5g5uWgubLl6dQPGoD2XQ4LuainX6OAJ
MM4XUTBJMo7CkJwhJO+hWq/ddxWbS0sybRC9wjUqY2sXRFK4SiWxsqRPbCIf/EmuYuqpS2UCYaKg
NSui+/QWL5DZs3H40CucyYQHNCHYZyRwFCjPujPZWSZCBvz4a1IBKN/3gWfdahOuaEy0RMDukrlu
nTbLjeu872/cJcZwGJx94+NmNQnCw2kLYy8DNhcLS1JPIbWXEM2OeODIJmY/xiSXvFi3o/JOM70e
/BewZW1XaEAN8qXhFq2i81eYHvNs8klyN8bddERoleriDsQuwWTGAVow0qBrWd7JKgwigjYEhw5h
Xk5dc+DfBKJlYttoyCX3k51LLCIzv1ACHxwUL1fR+QWHeVTlc22/jejvWd4vrAarjzCLttAAQxjo
pdb95U0Ql2Kp+3xuuCV4PGw9pl2l/oxbZKY9K6KYPztUASnYUYAKAepY7U+qRE7S6uLiIxJ4ko0A
rfEq61zHFtZZV96QntJuXd7bXp/BqPw20B3vakFowoxd9MUQa0MUrZc4MqEK+7mwYxvK0gdxyM0Q
zcTfS5hqaU2JHE+A7HLp0SYTPo5XHkbn4WrpIsGhzIXi6iQKRgWdWB6o08i5Q7MVGWZJIa6ZrfiS
0Wuk0110ce68JneXDhBnBexX/etVtmxHcsiyqNZp7DCtW9e4ftEAQ+ui/KsKwQtYN7egoN4IgZwH
B+ZiGxoMBbbl4wMg3Eb+K1Dl9jGgPA2oGsBgn0t6MyI6l2HTx2GI0EdMhOhp/+w14EGw7Mkjgbg6
BXYBbnfxkdTP21SdtTeKhjJED+5YeN3dEs3dgkefN5JmfFyG6SQjllOBDWSP13r9DWksa1xqvBGy
6ZfLdFpAI8wXaSu1r/nLu1oRMn20wVebKbg0qUvtPlFms/ok3o1vpuCd+3ano7v+VQTSMbhqXfp4
aQc4A3alt04jrUBe1N6mmv3Vdbbb3Rdg6JhYiFuFq3N5JGeoY7sw4Bynxybo3NSnPhyyCR2bBLQ4
PQPzo86imdTg5y+bLsPzCJIqggjQrObKV2UTb1wSQhsCYaKOfDzV6rhN+onvs2tNRW+HdPmYeS0E
BsWczAJlvIBPKYqpUEGHdZcC5ybg3frEN0Cbq9OljCuh7gWS/778HuGjNfhGN+4DUtv3hUNJq+C9
e+5uj+6hwIHHkfiGDq6Oo8RRqvTkDC6GRQWQ7tbXq4WIEa8tWLQd2++Qh6Icr7Z93sA2zV8A6MIZ
9MDtPaLLbx/mKwP1250KLkUT++CDdbLZ3WrHsiNVNaS0Mxt1yvA2CZYySd4DsyIMGRjgw0Rb7caR
K0jx2t2Gycnkv0mdsO94zKOm95YRe4ZGqX8GYuwKE8r4cBGgGmE3M+GGOyyLDzNRpZOOFWslFRrj
I0bZGjhapvD0TWNWM1izLdICkSxK5BXeQ3FChIAWe2eqWnUPGLF2+8oITZs/65bx2w9ujyZmBS0J
lisYMfvWnVZq/u1x1tRcNmlx/P8J4D3N8Y/hpzpv/cRvG717E+NSsXi6T0xQu+QH4Gm54zQc/LKG
3xAYh8VxGE17VkQbzExn4H5sd7kFSiE6TlhoWFvR6N8+xTFH4K1X3+ngKs0EvQt9qOl3uvVBXbRy
NzQYZYqd9TeXFam4YILX3tG9VWCgOQ77YakB0EgLl/NcXbRyRT46H1V6u322d8cHmU0JM3EcaWOt
ZnnVi9dO0+rplpqtbIVRIh5JRnck2TG1fYnd/RBnfvoWjJ84lQ1/ni28HWdkizsCRJxWey8QYvy2
5Lfmiu+WWyVf2O3r0MDRHFM0VwCAjkC3xxgh7WdLlRzOSFnE/8IQcgTObtuK9k74aTCzK/UMQOKp
7RNV0wkxTclcAZTBZfmMV1dHSaR3QUO+1xvCjFDDLMC70DJ0FAWUdrCr2LltYAS4sZKXUzS5T2iZ
9SC0gABGLnWEYxBtLyxvWoAmuiiMUeNjgfXfUU4LBfw0CD8IKCc2/dB6+6JFRT/5SkQc07EgS8uP
8YX3Mqo2IiuoVXjYxGu9rEVK1CPmJNZSYnM/aZ8g89q0WBCCWVoEZA2GuTy8QNeZ3Kxoew7iEjen
E38H8XYpNPLjWKItL2q7zotuPf3DyuX71SH0c/MpC7TeaUDhN3TrivV07+W8XucF4gKY3WuT1Gg0
a/KW9CxqmCmX9JHHM2pvKFLWIHz+9kRJXqUWwauBevm7VnILB2GfQ7GuxZ2D5o+af0YpbG/cfo5y
jcAbRreLYCZTLkuUb4djZ2ahMlKr0i031yGBDRrfDacTOhU8NYZONPXlKul9PomTLmN7FlOpkn3c
XpUhH62cWh4MkZL3gKvsSew6hXpJiE+8CBmCMYQ4Ele/p81FJtXlSKJH4zNo43OSoF8qL2Bt4A59
HGMva33HGhVwIt4KnFqfwAVeBxTIBU2O9Hn+Dhk2AdFTepjCq1xXw7b2fomaA2xUDWM32jsEm5fn
QUCtGoALRgkZMGB26CQkOS0PZeYyxJ3M0zXlCsM9TFpGrxtMBzftlFK3QfcqDgzTrle4u/SuwLTT
4255eastzjgU/lsVT+N8B2CR9hQ/gsSG/uZkQSB191RviXoyA1o5PXrfALZjxDTlbifxt89KKnUf
adH8hwunjTXO375g5SrFz3B2Yz3LoK58cQko56URYKIEyVOW/tQdiy6iIKshXGsNOgb8fIWmzvAW
nF+omY6AQVH3LjXq1rpfH4T5IhL5B94+MqrqwJNhLJ4V3PkRhE4BJswlyIbnyHexwFqisJaRDBlQ
dL/2VtznYo3ka+GLUfwpz53d5RUvmdrVY04x5FSwL2/3qPNoC7wI3jhBl6PCZi5BvLBjyL5wzV4R
65/9kIGs/WEomipeNzuai9Sg9d7rGoOCUJGfmBF/rQrpB04s+m/BgV2ZdOvkG2w0VBH7B66oWCqm
9SVgnfg9XQJpCg5KBb5QyPIhZEVoJLAgTAtu47DwUAAnO7PbjbdFBJpFSC7/3BkaZ38MDGBzKFeP
ie+PE74DH323GXQiSxz9C5xFfo2hQvgCUTNM7ikNGIIPKLE2PQXF5wRgX0I96ypz2hvcS3Oi6MGp
+31KiazY6128O32HrQB3QATubWWbTViqzoD/dxPJsqshHOU0ljVO32cTiD7yAa4aeMRkX/oe4AwM
bCMJ4lHpc1T0OA0dwmkymPSS6FIQwiiYXxWvEBn2wvTiyVRcrScPqD76W/m5/oRXYzkG4/xyVjCr
Xvf/N/3M69RnZfJjlh1YbL0mPJJbfYfssjbwynmBM8yyfRKbYxQ7ruBJzJFPkkhFF2YOa9LiWLK8
eIHLAvAAbNZ60hGPJkZjwgm2U8Agk0jrFhEWTsK9J13czoXjrXzdxNhTHO9POAg3+hmYeSxJUBRm
EmYpHZe/cOHeQiGZy2rhSzosWiGRc98OLjSUnwt6hTWraP8b6FzW2xe2gp7bPJyd5ZWWHwNwr96a
D9jHuly4EtuxEn4V4q7RU2IojVs47kGvrzNdAL+byW7MBL8tFqckWlq8cw2Fi04VI3jhpqKueHX0
m7dJuaIox4bA95Gi1aGLXhW5rbKNHkkpNSRJvIcXOaNqpn7EdLj6amETbeh3AwEIF2QoK6wcmwmG
biWIJ6qppDjsT23Hc/uAEhFJqpYEQUzZoz9b66JeEp7xKk4BjWURzCQCN1pEWTKSIORdmWTyuRHe
7n7VfUcNYVW5KzxSRAt7cVTa9KCP76rdwPZwS+lWCcLgP5V5i/uttUj53Y5NO1dIkbNIFmEvVzwG
BgNmiyDlptF0400Up06psfF1u0pNu65suHAIPcRARGNEojiK+l6GxsaIUMdPiy/yHh2/f7DiOU2r
J/wOx25vYx7Mu6RRl9Yx6lBLhI/4ALpnnq2HF7+Y0mDBiSOwyq8R2j/u0yNbM4ntr0RA44KxJAHq
OIV4eX7Fmht1joEtvYukx4WyUFH4k9/FfkUHEJ5quemYQD1j0qHVsxx+ohXc8ooHS1ryvcB1jluG
8tiRC70TNQsIOfWWiAgUKgYplxDOEwCsO55tE9j1dSHEY5V6OP0WY9LiatabGTf0KOqoniYsLrUn
GDHrPBC7iw5TvL13jeMuFhNFrMxwS7qqfjIAz/7ixJTtwcclA47OjSix24SqUECkIQ2YEIn7Sis2
xsoeSlSnhdb/5guN8LWBR6vGRxwio/U4gSRzz1n7WS9cb9Q4qmwreKtU1YXEewGvuoj7MFNvkCSU
rJppdC6xrFJJjGzLPWr6U1+YCLkHhwp0SbO1kBAzjmMPOKQpf6Yqe+ODGKUhdx3kGgxGyMI3Fu9Y
P3W0ThvFDcxfKfhYACHhYQK/9kjvbtYj579Vzy8ZgLFL4NnnfpJ67qKEbL0UkQW+RZKVyncU+0RP
JikKWVPVH6yTLT6FcY5Jv0KbtrV7eyvW3ww6NPkuT+olKRZ59Tmln3QXYZf697bzg7ARvzS8GnYH
Wd95K130jZge5NhucFKBLGGn6t3RJ0M36GZNw+vTxJ3OycFJqHaKiABgr344TvB1JTNlDMvR+8bq
etHTk4uLaNQzG67TH4UkstTfTGLcx5DmFpD+vWhXnykSzdUgZoBPxTjAqlesAZR4h50pP9ccwWMr
xyhfQXwjRkbfpXzi38vlBoiv1qUJfMN9xBzmctPXSfT2xRO2yLl+e3bAuke6ZRXCwy3iy5qFIzH6
znD2h24+uuz3pHr2vEUA/U2bFOyh+vplqqwIG5LtPa6GR36Cm9FeOYPIwbyzqdwrJrqWqrv4PDI+
hGSTtc/taoa3/bK7XEIypsJBJMRdKTFOdaU/q7mj/rvG2Dw5uxeFwgo2rfrF16XweDxZ8eNZNeUJ
3kLDRAo1GUjfyz+qakuWFU6l/tY4WhkwEvRcjS2NKyR6SBAUbPNLQy+SNiAG9QWYlBnbh11A3pUg
YD539DYgWbvo66Hxl9tul+kuZ7+XIf5bW+HcJ1DFEGHxHPv8wlf/Kxmydypp7sWegIHGG86H3WS+
JCTGeb2d5d50OqRMFLdNorb0VjxgoYdtGOEnqUb4aTwascq0mFe9S1SVnWczw5ufrGiGzPMOUYyd
zCBuG+N2Rr7CVU6NpsgUiPeBuXPu/9kJV/LaidD4zSOZuvVhtk/bL0pwOTHImtsWyGzw2gweHBAA
E0mqoubKZvCEVfmoYF69awbUMafAW1cp5O4umnsdE3lMLp9JyxJZeZ3M7P4Nq1YXsaxFqtQ3LofL
5lTzY1EsitKewuJlqkOzrnKhsQS7/yK/+FGXyhfg4bJA2Z9GmHnTc/qNCoMRwBJlL1wqxR5A5h5h
M/DPqi8dLt1WvYkUMowW5va28eajm503CaWMuBnnZeDJT+vxrFSuq9cs59rxJOmZRc2wj6ylOkZQ
vrQF1s5R1eBUXyjF3SEBuqpSo4RDtQlq8odNL2DlprA6JgOYuVDSM+cN58mOxvWVNSjIxf0yjWyP
+5BHx9vycVD5EATELiFnqg6KRa5l3E/RDbrNKsIQMjBUWDqOUqk/ZY48+5qOijWv9+8uWRDgzPHo
Y4PldnTZdJHyjvRdYqKo4GwHhjj2lD24Pv194jMK27Pz40s8ugU6Rtcs6l/BjP6yCcKdD3wx0JB0
sqLgvYp7KktS3vDaI6okgQ/o0/z2OcG6f66CPsmQ3yZjxd6OzFtECSNoRoozaUVANrRsENSYhRXp
6fAdfJvR/eJyRfU7YlFzyjvNKE2Rarsu9gYzIMnW37Y8VuRZfYNWQXoMlMIlWrKKnylfxCJPL2Uv
5HXWR0PRcC99RJeJtdGaZhYVLQeRyjZ23keLaQsS8xMNljMOaBB9hnQMBGPwSV4Jo5SbA8Kx8ut9
fnT/eSLNbXKN3qxfnTpMXm6IU5iZ/s2D6JYmlFeZFvh3isoyEWllJIjIA/Lq2GUj8Fh9bQg4NMjk
c04jf7FxYjfG7/eWB759l91uLnoQ6bk87SkVLYlUg6Z6METLJn7uSEhKEryPihutPwH0fd0TL+Kr
/TpIsaejb8tT4xxHW/gQh5vEDlf0QEK5B+IPvg9wDUKKsELXybwNTwq+Q5Y+mY5ymc0FiTBXt/r1
6JBq+g+B4a9sLRMxG1kAdr5h0cu2jnDLh5bLHX6j9JeiZEBRf5zoJAdh19UZW4px4x4EHx6qMfaJ
NBPfFB4qRG/qu+SXzdDGIT+EVyRKLiWV3u48CM0Svfr/pq6pZPsp2CCEYj9YtwhZ5JknI2K6RV9Z
NKCcPDycabkrERSm5PeipzsjdnCyvGSqNEhM3O2h/R2NQU+zflpBp/mKgfPIEUm9/KVXTqCgzWr+
C4JGyrMMxT2F2byIChOeUWj7CG11NfR0n2xxqItKgfsiccEd+56ycPLDHhWjVDEWuFCbMHr2wuXp
xnXU7mNVvI8MNonY5LTd0oQgk2VJ2ykLNDibXWvuHupI2Cc4LU3q1fzhlb2CsGM5Yf+6owjvMtrO
fpsxsIOGNDzwemjitZbK7uo9Iw7FN004lao1r6NQAN3tvjC2AZmDymwTVR2gBR/iLK5uyVtXLr7T
3V1YB4VU6+vOVaScE3Df8KARrbnguA9yWCph3X4EKjVPcDE+3pvZAgAIEKL6w+UktTI5GezLtmjo
TAJTXwfGeVo7oeE3dnisZg+3xMHYgB4OTzkQESQ2hQUeZdP6c1zz6u863dNUEYFD9Mgc62RCoRZC
ZC1HkmPstk8noRSGCNQvvHbDrBGuU5QDL3FhjtDIN2Qskp0eY/MZi629L71ZMkPyT+Lt3yQUAo6K
/Ka4GZSwOkYtu6TDiadWtC8fqaTGVUD13oT2Bl8uhnaF44q4cRTZjc89dkPo/2yR8XLTxgb361zb
YUNIctAyo4qg70DjZNcPt0ISlr7pkRfUQhphQB0pkWF+XCuooEAtIvAcPC6KM1fb7/BdTpux97Kt
Nh6XofMGjyI9RUfe+bk+1Twh/HPZpvsN9e9SSuAifotJ3OZuvIwkt7Q1pXBJRIgDYDc39tgtoc3T
JaZZ431QvlwZ2z6IW5QTwRAQNyHdPU0kL9EdMzE8hVGuS8T8pzLO/6RBBmFhad0YnE0LX+1q/bzf
x5SOWRSPL/89HuzKXDg25SD3UycNOpaU37czmzJnN4FAnckB1zHJhP2SMgFTtRXvASjxlXTiBuM1
KqDlx++7KOuVP3Z4Vg4NqGjbfOou2+r5W0shJgIcj5cwnMJ/NN7EGnz8PY0RW3hErb3snh/pOOa3
0TN/qX+fUf/Y87pVD1ldLHYH2blmnuQuwd/MreihvAkxcrfGQ2rHwwNeIpZBI2FH5xPTYe3/LtEX
JTOM8HopxnLd+WtBJgQHGWiucOFfkrPV3/eDBedF2l6DOlhK9ZViqePRz1tWlS8AZW08GPXxxllf
I5uf8Xf2+JEme0vaeaVGodLJPvc6sSEr8hfFl2hPDDAH3JhnfhpCE0uYjpw9yXho1CX10tD/6k65
oF0h9euW4QJJ67Ek1K3Ru8hWPmg2qmepCN2VJ/YgaYUWEkJG+Ox0A3YtkASQf6gOAKcKRUmvxOu8
R9z3oIn0nJQB3DB252G58HzdXTOasrxRGaWSe+2hmp4Ks9F7V03TrWcwuWenlxeqxupk2kGOVeFp
LNXqLjeRIpbdJhXn/BvhgSjDH2sPvhUCgbYsH1uSz1FoVpS9WdDl9Gwrck5c8qd9XBqSYNxvWoWD
OY8WYGSfDmLzXtD8b5ILNhNcRjbZkuqoSM8kNRtiDorLCcWdJp6uJZ9Uxp8On1XT9vx5SWh3NaBr
1TjVVqbmZKoYRqqyb6sxSdYeJZNBAfTI2PjJcrVkOyQxwMyOZi5SJvVFOoMAHm31JYvRChnx9AVB
yiAEQ7ZgtjduAs1joSFv5KKt64RKKzBc+vygj+UZkOCyc9co24yHwq7pjF7CgU/JbmmXzpXWt7t/
SdrlayISxI7woy3/70dpJITRM3OATWs2ySxYliHzkfn7CfrXcgwJsG5FCLXU4BdGNyo8gAYTeb+5
diDJEyDWo9cjIx+nbpVJFnip05q17QwcielxZyyqHcshFRumC6n+OWTQI0kbQQGU3Fyj1V/JxpvX
YDWXZVUr2VGx7z18Dh1/lsULKUOZQvwIhCKPa/HgCkHYsKcE+wMG/vNk/MLhWKpIxKax+VWzPYs5
gy0SShU524rGRE8oBLw56vpjLcp2/gLnmqmXM+sRwh2mnb4kbheraWstN+nl6EZuvRBAQdSVrWnk
tS8n9hvyzl2iMM4JhAxwGMc1I/1mjQfWm+/aBU5YZ6ZrFIwlO8zr1ayvFxsriCTIMkj2RLmDeR4Z
ICpTOens0Cv8HEzItCGaNzKl4nw+OxEzKE+X/pcQfuDuea3YJHGp5O/1dnVEi3sMDPPzPzQrnYHx
kj0inOkJEwBaGvoJmLdL7358z2WWcXFmmkJSV+R0bCzxaNLpnA7VP4zqOhKdAs0+5uSzC9Dkx/gy
ZV5cGby/1IL6j/ckEc1wra5zu/mZAO7Z5UpTRc9cEDkPz1XoT/Ilno2QkOwCb7wOoxeGa7of+8iz
n1m57l/KvZICUpU+QX9ufuVi72i2j3nGM87qY7tzkrWV0HhZz1jzRYKy2dR6yeiJVb12kYCjus3g
7C+Ns3PUB3dp3zluzubfoADFnjHRpSJfPAwMZrfGz20CLtaD2mAJNM9QhCAwFagM6bxC/apBSq5e
ye8nEW0JrVWu/69cWHrpiqWa+/uxxiVg5wazz/yaClriLnuiXDg37RSR5EsIIQH2JnBl3PK3X5qn
KJIMD4VPj9LDuhbttHMnrJMITOSZdCIWiHftgb/6Vr3EM2j63v2eGsyzgud3X+jYcVGk5Ra3hVxj
H6WFRRHoRVufJ3YdQFeWGR7IyxrsBUBVYN5pIlEawCqDJ1YzouUIQ734gd+FwPmTXRe4YTrRtcqO
9J5SwrfcD4H7k0A6Md2CNCGrlgJlykSeMO6ENKyFHLMN1uXzTvqCpIZ9yzui9ezKHHHVpF/jbm53
G0M7plx6KFzG4zFTyO82BSflCSUthbS239VPd4SaCx3n3sOx1/zBQBXnb4pIxe6BVYOQL4/HtLLX
q7jQ1k7ebab0luv5ih9rGgQHx+fX3x7eKSxPJ4ujm0EF9IRW0DmFyyZEA9/2Gvkb8FB4KGmaYRNl
dy8uzAs8G0/f82TijtkNBmPg3GBi+sMrKdsF7jT8QztdAnwkTMg6T+eu/Q6Q71WvldKnvO0qUKur
C3+AgIXI14T7lkIPk6lIwVAp8ENgF+Df+oPIhX6VJ8C/RDnboh1Z1lXH9D+vV67M1Tlm++B+RkxT
K4Cphn6mVtkDRVKQ0/VHttf7H/bu6fZdm2Qsu8VKrgy2+912zTQCcbYgCdt7q/dUQcnwBkVxxaaN
w3bjYPIrdkZfN7OY3xy4RGszbaH4oB8S+AjyPsf1P/et85hEXxQYt0Be93v6PSgZB7VAhI9GUA0n
uvoq5St2F1bWEVKzDLrpX73D13hPRnnXAjEQMHPo18VjXGArlleZDgoVKYAvnbN921Y6Lpc5KPD8
B9QB9ymhHWBdBW07h90bIFubAeihw+ebjLN4NkRbvq2lJsV/bYvccSyRlo4IWpSnTaw/r6Lv5iwt
TyKt6xuE6FYzASgQKYPReEe2XoM5WezxzZK0+Gwob0LJTk1gNNXKNLL+yDM2Ca+zwukyAIymaYqU
1i5n3ZT1FvvxwBZx0WG3HjPpGGiX4YyGbuUQDGgzjOEeI+5MeUyzWku3nYOMLi7RIPrx29FA4/Du
T2tnwUG9cFQHv2eUvX6TEkAotdBpLIRoctAo8oSrX4iCOhu7dSPoy8FjARDNM+XotXntuPS4O7dh
bzZejeV4n4pWlE8LB8r0Pdfb1IkL1lw63xoRi3hV/XoJMq3Sz404HuEzlZELj6Hx565tuMiy65Dm
ZXV5HcdNv7lH/EzZlWYvKydYiPbXRglnay+iJz54ucaW/5wOX/VDa9vr7BjHwW+HOoAvUqMkZEOV
QKCAz1TJnsoZYiInVQWoHj89fEG+wTSaLk2/dhkAQHYMJ8q9OfhLWM/Y294+XhNDfQDUFvVIBN9O
KCVjheXKGkPysS4qnF8r/jAxkvlyIM+mZnY13EilmqnD5GSArWsX7YvJ5i3T+RaaD8FTOEHMerQ6
9Pz6sohmDL7pCY/dV4EAYkxeGWp4DDmGIbrLGwgKRu4bPZyVJJ3g/9NEk1tL86iNIPOia8jtAHzK
LTA095yqBsLvBUSqqGt3S141c3CgnzMSjxt4k511giO0Zlz329PrnFhbm1ap2aYS12V+NK3zkEM1
yYIYvaET0U+hGYDI30PoBIf7tNkYJI8g1zs4e8RW9ETnW5pNZxhYptoVnTU9GUP5Ed7jj/nbr7Ub
lOYMRFErH/jLFKu/lSBF0OYxZmqqlr8cgvgeoN5Ul4Dy3pBmwIGZ+jKPIIwCD+czdQTfg/1DrJ66
zkSyfwQ4xBvqWphjfeg3c6tquhdt+jOjDV7w1JVAiHuDojIb11PL9pW9023gtiDrZhVR4OIVYtLK
uFgpki90Ttwv5F9lZaA2kd2ogyru/PpzR2TovG/MYolxnCqK+fAV1v+WldB6nhuO7CwezvNwBOx0
7H+h7qfc2sQZRHNvx6xQO/Mu7GbPXGev9g/RR1QC1H6xah5Tq/tegdQI9SVJN7Cb4vB8/7HKE/ju
99RCnObZHcIs5xaxVTsTcLh9cjO5FUyhWACW9R5unkVdfB6i7GOkmAal11oNo3VGtTrmvUFLH658
IvhmDkxV6jYC08E03GSCNqkf2HBv5Aq4OBFS2YoYuVsScst56TDJ9O2GwZwJAEfdIR5nMe2UE/Cw
W48CAHo/k95IRFTSdN4UjR8zcfuaZxf26JH008UsF9M6jLKr5XxKi6+Sn1co/vLJ0ajKJA+UnloX
774mjrFmr3dBVUVBvMYNWsuanMQnkbwIDhx8FJLKYZr+l5ZnxExlmxZ/Q6yBYpDp05M3YrQsz/za
DwYe5wIcWfYUUHWBBl1gQbotfTQKG49gG1Ye8QvKMBx16qqi3RiwT0ZBW9F26T96iQqXJfTZ1vJs
gVnODzMlbFmLFa8QXObGAjoLIXOFh8J/tOekb5IKHKLWDe2Xs39BeqAtCarCaEXBUFgYhDcSZo0J
c6Px+v0EIHdp4cEnITQNRjwtKpt3Ral4bs444F+4YXVQSPNSjCWJr9KDHpW5xYrSOasUEeAQbLM3
gePiEYnS/2PvS+35OS9zNYGlUrmn18zRsvs70+EzZPyn7xANokls3t8iL71HFXjYWjy2TajvRxA2
N5mkSasZt0FCK86QGgWkgK1YCHyWUnTJMS9kqoTvzZiFh9OoA7EnnUTNzbSeiRUWEd+FvPSFg0TH
Xd9ENRId6z7pAbWMoQRVkcCLvvHR+d0bxtS//W7jD2ifsLgPzd8z4kHBptIgsB7rnzRKCD9R0lal
CbTcKkWJNwZD2qcip8iJkCzpPrVxwUsio8aYpqJuz6soME5+BCE96te5j3Z1EgY7yq/oETGM3jwf
g5gId324uC714jvr1GczQblu/ewf+gUhYYsi1Fae+AiecMFMSfdzzJ6zCt70Zm7fs1EzlFR4w9cf
xdJ1C/IDrCI/ipekgKUHD8iwmGvdUNrcMwnsb+lKXN/aLCoxxBGoN7Ms3eNdyfrzJLR3aGbxpUAq
rudS2PQPMzrOl3/n8G4hqExpbbEYDkK5nxwh08wyW1lKXYXcuTAoyXKPeRT4hmWtU5peyHZhOlRt
dNv3YdyJ4UY2ZhrFnkJxJiZVh3k3wHeOs+n1ozuk0csHErn+I6UghLdYykzYa/Xv4XjAtwprwBI2
BdUEyG08EivFclBtSsuDxjB0rUh+nMBCbUTHpgfzuJ4LUbZM0/eqUXUqjaOR9F32oKR3SnvLAizF
0MeAmpOZvru1qDJSdhKGB760O6507BHsxi2vwyeVXcbz7x2nhhE7MMKCxJTYd/K6EowMbC+RvtM9
A1SCRTgMjHWHSqEPG3DELsQNTklSIYqxRoLO0w4eWGPdhCWPKnY1EDZsj2xrzVPBwEXdDeA0xDYH
svsFoUssRz9QZrUVGUJKx2fHfVIJNgFZ+0kCoRiuI7eLVu42vrolG3TYsOxkkCOCFGcKX9WEDUGm
kN3pUzWhcJrOkWFV2FP9gIe10kqY5pAFkCIp5EfFsSg66cBofAX/uYhIiWBYjGsYlAMKg0IAQZk3
4DrAXTVsu/JMeYLhFaVc6wRubsRIETRTCt+O2oaZPe5NNByuMC0rah3z4+DEB9PWbRb1fnpeGaBX
DWAURdT21uqVS0FzoKUx9HVF2D35bMFeSK+fQHpk4bKbT7q8q2l1hdL53lVeVQGsYJbK8g4GGAt2
WFQW9009vDfGk2yzHYBDmq82vOMi7q4qrZLyxWxySd505hogfKux2c40h/4ROXGa/9FCH256JnJ8
VIgq17+iX1zorw2KK77TEbotsZ+8fYNx3PI7+jsbZ9AgRPFqnFVTQ22t8eDm20H/UT7He7p2P0cd
YREA3tEfgVejaWpJh5lMbRpcPuiiJPnrwxmFpcXDf4BX6nI+WCJ5jIe3o/rS+boXtPvpU8kkyLZf
A0YRxuXSz/8Hkzi/cxzYQH2qEudvSbaMKqpCEfUCkQmqeXSNwrZyk+K01pVt0vqnkA/Vl+XY0cGe
1o5v61BLsmlVLgr6b5FdZds7aFfbr3U4TzI8NhPo6foUaJZ494sLiyHnnXOfsHFMkxNFhqywS9ek
1z5azLbftZH6o/hOZY/Jkq/TQhdoJ7xa0+VHPI/xZIGHmofqUb9ApbTrgSANSL3Z971/yrNn0ajL
LkHYvO8+1FB0lXHbwsLAZxGcOr0qQhXkAezwe8r0QuKQASNbhvEWJIyzFPxJCGXbeUwdMW82aGMg
Th4PIC/AgovvDN6M+hQii58Rh4p/XI3hlqYdT0ErXQ78Imc5MEwtbJ/VlSUppFeWF270SAiRmM2X
mkvgXywt9z/VA8Y1J14jGzSBgK1cg1hKdL9vvAnZiJbIdxtk1FFbSN+b7dkMCE9oZDOLEWb8+8cL
/CYNcAyA9wP34seWnWa06HcumDlVPdAQ00NKuxBe4//YGF96n1wymeZKxtOLMcoKY0oUUzm9U9j7
ljWQi2oHXfQNhAqVeOJEDZEHobObxcdFHh0iVKNzG1vUM7yhOtl3F6vDAhzLgO1n8PduXhdofXTA
TWZZ9nEPrWBgkB5SMIysm50qRuO02lkSo7RqdpEdOZklCXrhGgceuueG4VdR3KwzsjnJDTwo1XHr
cMxa9E0dY1KaVDDaJLOdwZBV7qn8Tvs2ijHRMFOBuxw7o3QNZbeZIXpooZBOUluDjmktJS1/dgOv
Wrnt5/fEnknE+dKXQ2MqHPCZ1QlC+FrncZTkAShKeV2g8hs9CBpkwAVWkv2oAYtsXnMCuMGMJJNF
tPghoAuF36PvXY2WgMUCuh+ilXehLFOFSbHlby18bTZhzzTP5X+84KFwspcYL+iHshpPvpvOC/jt
/0qCbn91vPEjT+769iRlrNjMnmDxZ+VkufYWYwa6FgnsinpADCbI/cGtYoVH2xE2e+vbd/2iVbZj
bmuIPRqKwRPF+lR04HRRIsS9KVR62Pl5wMEsFbEdj4VXPTZf6wo4CoMK71bojgNepbLxmN4kuNyU
eRq0SKhJhSDfwtNQk9SE0fNyvedeyCz7fqChVPLnQS3HfKXSDS0m47ls++pr+xxSfho7G/SgIKdc
MFpshwWnpB8rfsPK7MxUUYIG7TbULzECPLTA2Fl4QHpAG37xFrBxJyIfsH7GnEOgylvJmwgaMFs8
CyOhnkoi91n+cUSqZR7/ZnDiFerd4jxvyXqixdWVGXW5FFrGo1OKxVbj1unBCqca9FStwO6pxAEN
iE4OVV+dwx4YvEuwNvG8QDHnB9Vs1nY52V1ZkwTA9Ahc6yMtWJmnDGQiZKBsm7kw6AEWSM13kap4
jpddmFOhJ6/20hVC6nQmmxoVwUlmFEWTA7sYYi8wJWCWYYLcYBYlQNlO5JD85MW4iSAiA+uVmqCG
HrMhf635xj9es1gKNM9G8IxLyqfj9pd4TrdbmlmuDLgV7CjFDzMywigfkekkYGEsgyizmu6WrO+v
TYjxPEiD+6D+/bbtQS6eB/Ll1ZJBQMDt+cPfwc6W+ferEr66KU4A+lIeAeqxD7yqy+CbbWL9Ld+B
BvaHbSdPl5z7zZLIQgXZhZ0RQW+1sFfm42IHyL99IXhpUV09q6/CpgDF4np5oJLtSpguq5d76Uyo
EfH/q3RJV2jj1u2cJn1i0ky75T4vHDUfLal6eptSkWm3qvRrT9xDjRCokQjJd/DFwoOafGTwhrba
5QzCdwkz4SfLypj3Sma1OFx2SOJ5oyHqX/zCzfDcZe/mE8vn7SVgP77wmSR7uX1lRiZ/kkUiHo3U
R8OPREVvJTYdGpeIfOeWfQ93grHEplSf4VKUlOaZKuf0/WHloOATWE5d34+e0wwODh0wxMWBrqLP
OC0D1FyVhghBS9KSaHzBILFKhz1G3DjcnDDCxcvBGOKXMbsFr+FpU/kL6+AFTdWKunAThwh1TSEf
+Z4Ms+Bkq7D0JMPAowMAfaSb9JYySuSM1mdd4FfgWlzSJo7YxDtE9ej5+DzXaNmpzc558TKEHS5c
is/eXWtnuCpUI7Bn2SK/3iHfp8wc3NoTFhr7cuFWeL8sbr9vuWRHs9Zg0ssM+iEV0LCbZondgXLr
1QEUDDymC5Z+ZCjss541+28hEBO8BqMNCOBqh8Zm+JUeLEw+uEfEwrvRo3LCzWNurDMDbOy0OZ2g
YKI4yyv2uvu0IUlOPdCWXk3eg5u0wNcftVlKgSi9Z4xzYfwCt0ZePo4oNbGLA692qqbrPZgD6Mrn
hDgjfmTbCezzcSoCOGjf4buw88Xu6AfrS0rSQERZTBgQNVB1VKpHAFEn8I8Z8Kl0pbmXgGwZ6TVU
JqS+zWvvhTVP0kOew3zJctTHMPu2yQGuUZVKbGkVSPTeGHlbz21ufWooWc/l37bOfNbTZbOwz5BD
tEE6HphIjZMEfKUHN8VyKgp/DOPDwlbuvdfT6EVxjzfnD3oLUHFoOEw89+4um+pWrTWl1L+GdJPY
rylJ2NKTDYJ0+LuQ7LR/kHTjwylo5xKF0AzyQdywHYaVlu+vg1aYiOnElHWenEkbty13xAJZPlZe
QLZJ4WZuZpzJv+vC0+xjf6oy9eq3op/Ac/oZCAT6cmx3PR+XlFccJNWk56oeB1LKSjZeXHU7M1PJ
pXnHpgWEm9l1q0vUMUaffqA8ltehJD0ip6iHywlebviKosd0Olxnqg/MyrWZCVrrM79c1KQlR8Vq
9n973GdjBWLvAMR+KEzhSBQNrtWd1A5YITKiEiibDsDr3F0ljiMpWSoPQd8qpIJ/0/QVsMrrlHm7
pv4cEtwtSHH7dlAUhFQc1mzRCyUIgzmQ9fiXrR/aXkOlRFHhtb7bwLIHR6poWjCnPnDWQLYsdMSt
Lw/7khNtELbaHsrj/lfjzgTDYUNvkqvNzDRV8rq6SiQ27NBbv/+j/GwLoJScdIV4BfpM6aH6As2t
bvh4vsXyrxR4nhpBl67QQojvQdN182j1k9ldMAbJpnqzs2YeAoR8jG43wPbRDiyBorOqgKX2Q67g
IZjVpH2zf7xGyK+cUe93Bo4K45BLbjhVeafC24boauLQCjanlFip8aXheDLjovlCQaYUDlnzeYsb
eEpA2huOfVwjI8/ekKRWSHhOF6bIcw7rM5b+iJcI586Pq7vldme3GZRDYvWNn4kulOyxRuP00VAz
Eij5/7FW6gyNGCWKbm2LSZ/zYexFjXUYEnit3Qocyx4pJ1tbqE6KEojhtL/2CVRRj6UgvCECVyYD
hmiK/OuO96C68X/qGjq2FtOU3Fe8jiQ4uhp0oR1HXDKDY4B2shGvnKjgFKhkY+qhNZMuo8GHGvhA
iFlzDYwhSJ3rvPA0MpEEzvKegJ/AtjxjECprbPAbYTOuazoSl6RnlWBtBcOmSIOtRN4e0NWDQJM8
QleNyCLZffzN265uKCR3XJ5jS+8lWxsDqsf5sBq03YQChC93G21X6Mq9j0obfq86Oa4jfonEy23l
cgN/UK2p/WecIZBQzd01OUGdXkr69DuI8ACU3qtZsbfSR0GMSV3vKbg/NyueS26gdRwWHda4TJJO
VOckQ/3q6jPvsFPFG8zlxGL6SF9xWmOQQ3jYbx22fRFh4CkxNMao9hKjfnaEbnqY/HdrAbAeZxQM
3/4gvRX0xzXlK/GSd9B+vZhGLASwliaiXuKb8nIFzX1w33g8Dslv+he3lmu/a+4EY8m3qqJBC7Ft
ecFrPwQaVS2kJYTzox1LtQq8W2l+F0ynR1Fb4WqeY0ckqR4htchKWZXU0CJIxIWPXpu9L0+RDMKB
lYiwsI48RNf3rKyhQ8Fn9xKbTbNQ//Bb3i1Wiva2vDEA2QzZkTR7JF5HYL+Hu4n5cqvx7QuDivI4
D5pifJ2BF/3YWx20joOOGtrkpY8iaBqeJdl9OYoGL19fcmEHNfjsTJMn3qrE7tCixl0IPU7e92oB
RbLC+CSuaVzPGnojdfSiUXlJcPaUqoKZHcUhZ4xpKjcVSgBJh88qtiywtXD9qP4MQWeWKAd2FeZw
jv+mEJQcZHJpXnFqs75NY7tkDLbL0EMmcQmdGuE4pYd8/WchBAw/BHxa/qcy5YDuV+gQ0FWHTQsZ
gqdpV2rZYu/ZFetA7iowWKe6DWeBFD8z6V/52QI7SlPDyU2g7oxiqv9pc66ZO26DTs4fkr6YISVJ
pShXJIkVmNjshtKqsgkNWzlBt5isiw//FjuIawqa0Q3L6Td+At6C6htJzLTEdmRwiPhfb3jjc6Eg
Y7QBWHfIRkrIvhcJhGgfUYLxdL3C8mieqg8lUyDID1hdtFxl5FGr2B44jsUzhFyZgFr14XBOngpP
cmr7tzuewkzciXkeQjHCa4odGPPH7eoLwJ01T1o+E13OBHCSd+6Li7YzBY4qlYZKO73mE2806Ybi
OGAkv2S9TbzaV5LwR+rWNqhqZUKoU0PB+IBIh0SiE+dUDGBXtWKrARms3RE/AMYHGB6uQlWqDxtM
4Ox4L4BQAXx9rD2HVibXrkr2RwifX39aX+R5BYm9to1fG7plcRnsul7lNV8HI2BsjmEf7Vz1J09d
nC4lne1oOM1Bo94gelxt/GScSGmS1bp9/yCTh1p/V/9XjlZJ/JkNYPVzEvhLscWJ0cBMNeIiXyqd
OwRo2AgCrt3BSmWPnFK9msQNJYH9Pa5mXsFHf5RMvYvi+QrS+qReg9njKJtm5R77uOEunBbH5o97
Bb4Kqdo76BHOGlFca5E4cbuJaXW6I8OVdXCeENg4hGvqpvYd3NSesEcsln83Gk+JETsGVyvxQzjO
+gZzAow6Dncn45nyAFw3MIW1BQWgEGyX5ubQsqFWXxyujC/inJRyIuJGgTeUVQG9JlLXUkTTAfS/
fkiCi9JlgscTLLctFDaFcwpAR+EJHjev2lSLE6kkXaE4ayRqutB+jXPZKniavWtII8Gs75NmAuT/
gJyqqsg4jzLHe/4gRtTu3E5jkpDgfQxYuhdrG7OhaKEZZCJ7dzpc1LbQcSzwEVSD2GBxiraD+jb2
d6UTXp5sAuPNhvXgUHC7TsveN6JEMKZid6KD5Vid6h6SGlNqhs2q5UpkH6378PqstrmfkLeWYVU+
CpleFKKUZBlm6J+N9UmtvjQsICib35SL5SuKXsh/4Nad69XmyGSloGVnYtjHpqxf+w/G5bRzOnfr
E1BH3jz5yG/W3jwoOUdK9OITtVVu4FA63ywA6FNpV9GKIIUxvcm9AMbMFlXlj7knpviOWYhcsSXC
Y65Q6dxse+TTdu6hrJczd/OGsKbhfQkUfoMDssbsYLUIL8vWjaNKaik+IFg8sy0tOpNCK/h76eDj
yw8TALBhyP9fbpTUzco6ZqPIo+oREEH10jhyV6zQ1t9o/PeQ05ZnN4BsCPjQvXOdNt9d3UlMsPYd
sTXSl7XsTzs45aXIDLvjZ8MNwgeFv6guvIVN6TwyEUwIau6dcOR4ORAmLvltCm+ukaurRbDduWW/
sHQFsboHDhTJBzQl+MzEU597xPrcec3USAdlkQy4lhvVRDP4ptFWY4Gvp4s3RZPs0w2/ZNyqhQQl
orIb3fZ653KGzts60WuF0FapgyGKJfoYMHdBL5okfj9vjzS1KEDq/7rP4C0t1whKWyPgtMnm1Zhd
sp4GTfNhkzCvxhDtIlf07kpQbWAoXPhcifywQ1Pn96eGOsgUVyTvxZpIxx/EW2xhNre2ldMnQxMc
tQI5CFExzzh5jJJHyYfrIviR2XflVRI4tmWgqQxeDIVSeIS2wr666mQB4e/T1FMmg7P7Ym6SEm4u
NQkVdR0+2hCSNGVUVstEk10BxQmLcDJpMfBTtxn2D9VDMZSMYpYy6ZPhUZoNXS1R0b/pK9Ci41kd
GzwvOHSFohFCtVjr2STwnJwUrxKa8Twe6r90+aPUz1jAng5Y5GzKQ5LW6//MYrC8DNG2/8eSBYt+
Qp4/HE1p2ZcD2Olt1s7VYCgE51A4i9wtw5f9XVV/9Rn/Jxkt8TmrIckR6ILZC0NFxpZploM4fRY7
M6fmghdE5/NK8hatDplusOZn9FilHxH64fh6utQf91mfVUzOQHwm8WhAXnILLhDqvCHcx1TpImAN
v79pawif2A4nyyLatR1j10TfVQOV5dzD5Q/HsRUVCX5ooqpLWnFTpYSygj+2vhHzyfhFEGfPnM+c
Hy/ctYCSYoMu6P4EEvqHU8eVO92YotJt1MF5Lwy5buYpcVywHxniRty/JrnEPxcou7yHC+xbx3uI
n2xMdLjINchmb/k1jqbswXozTJwWQNWSrpgS9ThXTrwzqD5xNT8HhBmf9sKussbB4do/uYziUqfG
2PIt2rSuWmMhEij08bYQMG0uTmWu19QAK31adZEWRiyX/F4OJKikbssOR1SoFtreIUK3jlNcZagV
bleT9n+4JceLdy2mVpOBA9LNEAipndmJK+KwUuCFA4BKZg4Jeg5NNzoQcYV5sNy2VuCOA4uQRgVc
9NLbcOxM9VimlgSBE42u92lTaVa0Pi148LR5oyNQvcVnxTcOavBqsX/UC4jB8uF6Ld4v6h3CVa3b
l+b9FMZmODb+n33y4mfdUGcg8/teZXgB25TxtNiC4Ooy4P0Mqxy+Q0DXS/0luj8Rg+j44C9PI8kx
VAdGGRR6POQFTCas6zFyI2wCtYzRuRzUd/ogeNjxz9OqafhlRkqYLFbdKA/BgbqyQCW5USpPWup+
9TVj6SQa9jI/XYk+6Z8BnJLNzByFQjWbae13jIC/trzOX20uGucBHrsvStkaxHil97xysDTgdCFa
wolsD8IvBp9tr1wkv0fTH69CjVktNWfRtKtw39XLscnP+/UmzSLljZdDnl5lR4NWieMdlBNjSCrn
r9sysLaejn2RJIiAu6IHjcmEDjmWT/Akp7Q2WZ/RcUiEe1tQgHGU255XHSJjUfA16OWfmw9Xw7Ia
Zg6nKhw5HKCmInwuS+Ys1svBE+UoCgRM/WXMsiyYUic6GbM6OUskUCWQ/QjLhN8o0PDDqrHF6pW6
2B2HJJxoH/I16Y0zqAFWVYTVITc3uVJ1KLr0Ril0pi3YHWFP2343PsdCK9+mvptZEmHj7pALzBN8
kx/ma0ifSVIGJY4OAvrgDN4Tl4G6PJhWp2Yy4g2wL7+0NJM5zu2Du5FRitdqQ1xqP8tMtPjyvplY
S/3MOXlWinV7b4D962QE6OTi2FYzEMoUVkdXV869r9ZhCTWNdoeOUP5AI9iolap6pGQmIeJhvGYo
NoGmaJz3BGYhey5B2KxB4GrpX67xkfXrkIIJ2AfuQEiW2STPq/oSzAZ7viberYLrcb/OLTCn7GyX
k1zyss5a5LtVLTwbI9/+0e7yI0T/nB9+HhXiozJ0bCbZsF/gm35c+jo0IKrVwdfq5ZQm6ThCjgcw
CBXJytS3dNqSSPaq6SQMGh95WOH4zzpUDYbgatYPuOewDm62T7Mnf+ohVNmRO2bufQIyKBFnfwyJ
wd9S5s7C03banXQpRALQmML7aOILqQouK0CFp/wap3eOcds2ewHL7MAg6ZGnzi4ZFmp30bf2AYdX
B5DfCZxHUEQITQ5OvNbp1rz8xRfQ8jkG+2LTcCxo0qnxdK9nYRghjuwIxDljmYgH6zhEZqgJLP/J
GNJM1ESDtGdbZ7pOJlHb1M5XX75Zbz3GcdpOJi8EpccIEnxh+HaPRor1uICK88i23OFPj3e7ZOtB
qSvPNEv4n7ZQs/vxksQm9ZIi2b/OY6l0cFaRNe9SLPgp9YonZgQsaohyCBOyDBJ50Y9yhx7fR1yh
rxqtU0dBvhNjFlgu9RDb3TYHx0KM1+8vSmqTlv4+6JpnFkhwXK5ODNHf9D4DZcjWCWZU4PM7HIbd
WtZOiFfwCMh6SZwnCN1qtlWZCMM8D2td67N3YxbYTdgY6NEU85mjTqQEmgYR6HJuUD3J3ZGOfJC6
D8aoPioMzDiWDWwgDHykzf6AFLknpQueAn3CMFyfp66ZOQWwSOlYwSaKQEJhU1/55YNdJc2Ccgn7
3JnjYU/jnBzS7niAm9wrBGe+b3OTfcBnria+ITdmwG4dApqsyvXtKNZA9wPhVs9BllDT1CwW1wEU
J+2FxNZNZ8DW2Hf75PR7MXDLDArm41vqrNaGGFu3siBsRv+rZ1xE5m3Kr8XFlsgutplO+/6Dhsol
0fUPiwS1jwj5RBM9XqFgbweuUuFQNLNbb+JT2VkMuJYTV+siQdZjtNuxM0W+MgA0u64gsruOoCgm
lwV7lqEQKM5qxq2A1r8dv3lDh6+kTA5kCq5+O5HltlrSJ+KK+OEbjabOnO29+R9+nNVfzK49rEP6
bwd/b3C3OxnzfmGsclDPh4c86BcR3oOf96Q8EsU9g6Ffi8fpQTRzt+5zN9bI9JWRw4T7P2nGMxVI
J+/4odRH0dcgM1F2c/7jkBJDFT9OJ3Sumf/2JCLvWVe32ihx0RPg1wa4wKqI9G0rYMnBbLT2neSH
domOwOyLQkXB7SU0/Z77hX8+MdY11sCc0Mt6P20fpBjR+4QpV1sttv6gm1FKQpH+JzYcuxu/Btow
LAi8cdmOU4R2IMV3fp+BdQ7vsr67cIovWuLaHEDqop31VAH1CEeZzcoikAO+zgeP89Y10CcmsPIt
++cYssn7hpp99xVfWL4iGni2AQQ7ZlmbMxMw2xXp+Qcn9yEtdCqQa5Sh/WwICnxyzv59fHQ2EEc/
ECgr7LZM4qy2WOrwMpZtGTGO7y5lCT7fUqpkJadOJNuskLkC8yW7zpIL1ue9wK6WRAdokobu3sk1
0JhrmncFjU8kj+bDxeVBoF0vFKkrQeHzBiT+rqZjbnX3+MG8SKO8toyE0pq8o9UmO/OWFTaM/+w0
lgJTOBAZ4OlG+aM+zlgVCOpA7yRo01+nJTtZ82tsn3GXQ34AfL8TlBBUgzFY/fXI8UqOzuE/EXrW
nKPkhXaXKoYq05Hey1KDk4fcu/o3B0tAeVvQjRkXEhmwOjA/eGRzluSt91pb0KfnoN9Mhmpl1Rci
9UbgWAE4UTXHHyJqjhHLUoSn+89lQOmXFa9FPGckQbdtxYuG7FAFRDrfaZGkMj6D4k4/9VP9SDk2
3T8uD5NxMoHEPh8Vq9YrcQdgMgG1KLZUwT51iVjrP5t//j/sxoRecVaTFLRKD5I21xRd3id4NSeW
sU7qhZcmXvRyJ1mPrRnudnS6Glgbj4bY9FjOWyU0o7TxIvlEf2bgoQt+x9g4lK52Y8lOHE4khDJm
lywyyKbsCwo2FTjwXUxoYA3Ja/zEXiRpw7inGxUUfMl7UumzCseVHbhrb4Vs9r5gGpLove9+cG7M
/PwHl+BKnL5DBX60aXq22BAJvU2E3J+60vFv+QclqQp9qfpWydw67fbYqNcLD5WEkbcyw/ZVus23
pE6tWMQpvWcgpzWI/L5oUbsg9G5madGWV+xziYDR/ogMTHwohS5TOnEw44bfdg6zXdbKPUbFLLbg
wq1rGdyxb4C9xZSl7QNDcnlxKac682cjiZEuzZq1sS7FofwASmuNtKm6OMKWNkMRvCC2NdDlOD7n
Z9ckjBFy3jVe9ml7h+eqxh2Knyx2TjHDAL6KzqKRe1Fooeippz0w+B9ZAgbF7d6LrRl3AM08KfAu
D1/Cog1kit1ahi5REYnOVaCm2mQbStKqjQM2YyYaXVhvO/PAKo/s+a3UBeUcn7i2P/v5hhYEd7ob
pHgE9+TdB+QxqrlBFk6Tz6Q24J14SDV1OMrWBkG4MLH05y0z6Ru4PSMcCmobenns+HuK0BpfiKoW
Zm+wJ4O6YrJgsnY1tBdWWCWEsMpiMnlVo0lTEeZDgUC9le8ZWv6sUXVkOxGObcLDmV8fPnxy5i8K
537NndvqKD2CY98dlN53EH+MVogNqdA6JSChqhgRRJoRa+MqN0Es/AI8do/I7aXqMeKiHC654/M/
4T7jivmtgsQdABUYHHFDP6yD9FpLiOo5eDTw6EDkMy6kCzuTJPDW5B7H9pvVktAD6Lmp2UiFWosX
PTj+wszrrkQyhOcmyfTvB9Y7zNBYzWvu1QIUsa3qo+GKlvecfkbTunVf9E1OxNVGcKFm68ZujZcU
H/ZJ4fnqDcxpcs6CLLE59RK2SWh9vdL6lJFziqLV8Sh4by7gaRmIdWspBXrrFwAZ0MeY9g5GJDAa
+uUr0dStf/AzwxcSJEeG4e6CahyivgOohxj/kSTl8/eW9eb9ijgUh0TltsavIPIlKYfhaBJap+eh
5iyP0xdgqC9vb6cyHHTJci4HqHAtbe5Kw8RClj2E2ZwE+/xgfes9lJRPSZtR5Pe2OUbhPsqWzzYS
ozR0XHz81UveZjOli6R9tu3HsIvzrtggmh1cC5+GO06XkjzDqSsUOXP7pg5ghcuLQUsCb067+Z3E
0I7k6EZ4NbcA7Hfbv39pdH9O5RKxyd6caUJnfc03m3VO4+3bY8oz7gNhh/wECsZZwN/gpYBwLjlH
LFpTwhHz9cke3GPc2Bwy6A5SX7KgOyMLBmJS4I26K9KZG9/Js0Ze6I2I3wsT0ztQ3j16e06ehoKP
mCtwqAL+aUf1sUqet7ljjO7RD1uMEczaqy8V/9pfdQTL+9b/9xSmUQYa23bTk40HRsbYKjfLy1Z9
wwnYN8U61ZZ7V5NRZRw1Th4KFdZBDJdOytRkhja77DJxys5r5xrKtn1GgWt3qKlPrMfb7nXtElvL
VABnuGlrnd1cm5GrwRDJFDzWI8nVPccgBlXyf7GI4odoTphVGIH7GpLobyCb0CD96qvNSo0CaqNd
fgY0P86pQXymp328wJYpMy1mmd/lV+SgnmPBaa8QP8vX573lto1ouFhnDcZ+2ZTVQX8BpAbWOeft
epzh6uIGFgX3Jgd5MJPjJWAY3PbpEbOFxyOPNIqoDbDwAk0II8MYgYuFI7oBWhHxKkAyZ0xXJEy7
v/cJEKxn9HCeEd8aJ7gFLWj/njpkepv4a56JDNrH606wOWAIyFo2UdcNsG6zEo+5+zDPHZ3QNqN9
L1UnvMZ3/UNOBPJAbeJmcIgC99SrArIioYoA6x9AvGc/txfrldV4nLEXGtQFjv2zO5bpcDWLqRXj
0H2YGFF8XEOJ9tI3wmdCJgORThvIoxpqV74yqhmdzV8IYkWx03IS70Dnj7tqs0kZEnnHUYfrq9HU
0+MKvZAgsPZuLyvQZci7hx1VE3m1CdQr6KJiap4RTyimwIxnChviI0FXqnKAkhSGhVTjuE1AZm1p
YXt9vm/+kpQH7Qj5M1Gi8mQngLARCBtFUMpBJGpQHMxS2LfZCQJjs0b3ZWjzbKewTzKkRCn59NBU
Hzp+93OSvSzZ0r2mRnKtJhjz2aB7pi32icT73+C2/X4cbxPN+Nabcten6taxVYz5DsmqgbXFnBaM
y2AeRHEAA0oYD5kbKfMs6MpI2cEqfWEk+gbC+4Wl5ssNLWz+2ZgoFR6hUH3zItBaOGC3E3/ZgjYI
dsykoa0cABXygn+IH4q90skRGtx52IuFEYsyZyZ4jj+/4opOnC9r0md4bBYGVAYZmKZu5lSpFjSM
lPGRe28rX39hsu+1zLTi0T2G8QktQTaVmLvb+lw0XfEYrcGmuj9aWFFyvlZE0FpbV5unNt/jWB24
YBodFPX1wf6hAYRDljkIdnalEoTCJWpid6UTEIrTqIaf7X386DH0vCfByJzWduVukG34s5qEXO2r
/didl0SswYLcsI9GnU+UinVd74yOfuPN6KyQO00NHBG8aaUahe8VjCoi73rZRyAxFCNO4BmgCPBq
kaqE60E/zktGpbwRynNh5Lf5M74/FOrCaiZd0b/+eCg2j9s1Bt2BZp513sVf3hBnZdSxg3nd7wQI
4scMzDeZnv4FM9TMQP/NmpeAwPOCoByR5wJl1gBiU64JFt/V5CbetTZeXflJHZz1qrcpis8WaAou
ROS2TGLaQ3qSL04BiUU0OAPSGJ3IkCxFbe22BNpQtjkj6Ylh4RcoO8ZFqFFFScNEMI9bIhRd0yx8
RPE4lwkSbZ9KJsr9XoCGgAXh3X2IjLj2mHg75wKnx7hDxYDi1bi6Uda4ksaUgHvbNDg9N7sj8cK9
PWIcI7nn8X5BR6mLnjySnnqk03NWsfL8d7B5VoED5FPZLH4LTLbsiWEHksB1DNP8FZw4cyknev1m
idCrNY2L7RNHX86lNrTB1wIfz2DKfYzzvMkiNnfLzKqC9JqdIaBDPjGx7Mz1lDAckkCLEzdJo8G3
e6JLUomZ6VPji3YdMC5875CbdSSfX2T03BdY2DsbBraDDIK4sxaTULcXFpJVFqXjRDBXxHW+Vm5i
CyOo01pVq4JAnnjhz20rSTzP2Iuoxgu3rXlcIbtT897hSxz01wvJXBM77UPAWC6K6EK2MsK+dnGr
erhJ5G5fR0Hw5YbprC4DviRD+xfRIAkk6EDnkBmeuLEACvVUs8EIHtj2DRSfu8YjplmrTYLBcrc7
jlvt8bKgp0EBaG5NAuwlus7lMeuhdk673rwnGcndotxcyrGll9SvN8jK86wH3AqeR9RQ6YGhVsYV
SqqLQEwSpeGMBuH7Y6rwxfETLumB3WQzvXXS8sEDVDYoaAXwxFHUS9/15wsuclEBmydX8JtOOQid
ZHmhZfHbe5KE+FL5NJA1Tmf2udQfOJt6ZlEiPGky/3i0126+3gVoCEHoXfRbKgEpOsZKrJPvmVHL
/AUD9IO82Apm2kgeZsPpmJqeb/yQ0Zh6ieaXxKrpMJCxOqyEC67geAGzh9ab+0x5XFPx84onqIQ2
V8zB0G4aTu8SeTgGheLW/uKdDynrRMF1h/U/5nEhHKpahmB19mbdAurGmEhoYicfO5h5qUR3XqKr
beVxgR0z9fFU4huVa1VUUv6v2prbxb+53L63+g2qSqe0k0eobHVf7S0/5eD4eRldJfAkGW+jtkFn
tvD3TZesCk2kSqHl6XArOkvK3uUE0PFuYxTrCOXzAPa7tE4G9uysXNMLfm0b1EBc3gqseACnyp8Y
iQTIwUFWLp9y+k+ohGv3Jaohyc8wGQm433Zq3nFpimjjcfGx3VIi+o7FkhBzR7UZrsBRpbDqF+Zb
uFxBjNSYo4oxAP4OV+GmeHstMT6w3MU4HVsFiGKWC0QJrwa7ziQ/6icqLimkTC2ohW2ufIlzj3jM
ydfoPxkLUio99WGUuRWiSfF/bDynvYua0ainprx+64SjJ2OnAYkTSz69LvdpuStLCErwIbir+6rA
fvxK0HgAS1bpaZpsTnsavwY0ZPyjA9UHECqZX4OhjYBqbweYJhFpbdRPMOJr7j5fuSPlgvY7E0hb
h6erWa4yhrEtoAfA60LiCkbJIHs519p5q5gWwcT5GCvnu9SDqcCw+6RX0A7CT7t1tZ0rpyYJVIJE
DlBFcMOHelY+WrGl8/LvdN3SmPZatOTFudbqQ9w4RUhlmdtLsXDV6QRi0sAlIBgBdR3s6xMIuBaZ
GIX+Hi/hT5G1w6AiVaJ+YD41k+zA79K/VTBwP55o0Qahcb5HX767HxM3z0/+eVB72nNaJTkd/toQ
ZDDQ7AAiJ5Qa44XQcNaGY7+NTVFUc3W1WrR/HCI1uncB0GApgk8TTlKx4s2SnuSNCxvcMDmL6qtZ
ncGz2bjx5bd6SmbR/o/h3+t+IZnbbUct9YXmroHv9aVfznX9WTSqDEuLb5kQcaP0xk/iWrpKl/vo
FGwsuphKaANfetfG01R4N2lEExtm199mjiyo2whaVdaajtCIm2jITGcl+qlwon/83cn8d0PAa0Pk
hoKTGlOd3FvWtlESOnnC1Y2/G59UbTJw0WaZcXg9gRwYQVqvRkkVOC9uu+JD6lUzWddbQB0Vkl7v
1w3GSKZw1MeR77qfYcYYZXOMxRJpovllFOXejtFhx++3ghQDsaLdxLOLoO23jFE+GaQo3u4Ubtc5
qrZgB/UK4oX9Nsr7aAHKw2dorgyT6AHHpKHZFfXWA2QV+e3ryzHaUoxjvYtEL8T7dW2KxkPxe1J3
e+PfVbZB35w+uCLK/fUGhNGhKfF6+DlZagD5v/ug+iswKEbF0QQ62McfaZpuM1DGW31VKNludhDp
5kOw7bs22Dt5JuWQrjooJ1uprFgtu6JySRulx3JIBufxe8os9zNazhBt1Wk7U5emttq05+GqFOYd
paPCriEuo6G4ff5kKtgRKFGjLevn4Sv23uOY37dnk86sSCAdrWM0IUMVVLf+XKtCB0ljMF1QG5Zm
DB9Sc3gUXTLioped3dXd8zd48vTsAbDSTINogrFLGIga3/qnfb0rAw98w7hjyEAoEcD4rKPxZzyH
kOXq0cYLb9LyEPyZ2owqyXOzMq/YH5mKmEuCbc+3mNmeWci91Y57Ox2B18D+y2JtZPYuVfd8Nlvd
IZp86LOeWVskyMnZIMhn8g5PPllOfZl9/T4ED3rLhiJRx5LCm5K6vVzMj1GxrS3NcrSzX4MCHi4Z
68ImXCBmajHaWdaqo0GpNY868M3tyorkrgW1St185SKVgiozCT5FWz2PNrvYklToYcG2zXRZzz6D
uo+2MH30QnUMPwAR0FFUlGtpd1nKTBpWEJSaNh8BKB2I/+sfGAWgPKkLsDmQvonNl2NLoq4/MTnx
YJt9WCqIIe6kPHGYg6xDasPUl5Jnuun0vx83AaTnhWf8166Kg3Lvx/LX5MzJpv0E9P4G+9vpscoz
D+Tp2r/PdbDfrVfGn//4nbB1QmwHA8C7fEgb4pE+QrhhNuDvamSg+s+wzlVZuDmEwdCa05ZiOc4D
4rJsVhDjFJDHFdXx9bvV1pzRuDuwjZk5SMBizYlujLzP4j8TBOBfpM1uqW8YDoshNX0U8DUzFf2y
JQtqzL+W0mXOuy7aI6M+uTyHgOV51Z8bx7JI/9Hdpg0ISua3wmxstV2eGIUF28XxJXFUtMXRFpNR
r2gn3xNbdtE398dFuziBWSixAl+JcdGtUVPInVfQNn7/JrawkPAsCXmcdTheia0DOw/pXiZZaw4u
RrcMxib8Wc6tIBp4qBK8W0QFx3cpvIZYzoVjFUNmg+iVqWr3HIpsWVT3aVN7KZUW/p8/rLU7rOp5
ix9lj3kYa7zA7tDqw3EHfbr+2r54yvoNZNYgLOu8yMQWADSoAe9CE1pzXyDsmMH69jHG34KTrgrl
fxfpKkI4IzkxytP88WtY/N8ZKhxBDFGOvUiTc6Jvz+VkSOyqfBPx8tEpCXbQ9XhjBlvw6FzG6aFH
DCVZPzWdENZWtGGVCZEOl1iopSeKnDIyZeK9oagR04iTRMUbK3jOmmeY6TUoy3MY4lJS6tSCzHf4
exICJ3LCy1T+roDdhTQkV8L0Xq9GSmokVne6n4rCHU2cxDLoIUOax+zDl3+joqGvxd3ZhK0+bBq4
YUT/JerOgKkiPy3VxiygfJ+aEKXv3joZ0tW28U9xZ0/o7vDxSCmvHOxCxcjUyfKqEm+jjnGgdcHm
vc43zi9NSi/maKLPztNe0yfFJzCn9KfO9Og/yjyW5sm6Lgr9OV7r79a0UhOmPrbA/OWLwvHdsREe
BkOJs9XX6QkHT5seHx+OO9HjfMii5BikmthqpDascI6iQtucKjUw9/vr2toaib4zK7ZvU4oxSRnP
2By2TJPB2TqstpxzwjwZ4y5jvVitVZrqAfyQmm/O3XyeYC7Fp3pkq4d/vGhD4Gh9rAOWOcks4SFN
UKYgjGYNiN8ZHh/5mZi43YRPuyk8oQhSCqhhCmwPoVUQDjE3j8ESmVYYWYsS1xB8r/fxwiYdIU7P
J8Wl2XQmHdHk8EQcaP8T1FQLp0xkM7A+VMImcC+GnzX/2QRGjR54/ILnfiVy3n2kcExWIQBY9FWO
MFDHSk4emglibMDRHbWxEO4yNlvHCH1/95rBWerfw6R7Afy/SqAPNhaQXu449SXYln0IRyfOZrAy
aoUlbrgTS21Kky8J19c/mGzfDbHb8lnzvzVQZtSMZWGh1LSEeodEzwOica3D/TPVDyqASXgX7kK+
pcdcOT1rB5EZ0UmQHGnTOfdYuvJoQnWk0B+2qLfbj77BYptwkx6/Gv7+AK0ArTWnm4Kbs4Ix/oCX
c6K7gwbpvIYE9whpVPtu9Z66aGfypdH3SFDHfPiGVtqlEj0Oq6VpF9uvzCXu7AaTYEnadjtAzaoR
TcO2HEG4/tcw4V2t9LBkQa5vBLZUg0hgIkLvzduN/tVj4G1YO/upsEOYQxnZfeGO1UGLAK1oGfeS
cnPWpstotBma5s4/Jzhv7zXVUyerSAqBO/Kh5QlEvfxdubT0SfTLyte12INtPA/kN/eFrWEdW3wp
stAeseGrPhe8w8sOLoi9GQyJgzQOqFRzzG2fkypAhZtYN0UTMoxevovBT7y11vd10ARIXKRS1I/x
AzVni/h8ZpCrokqEqCQkrVkc4spHkd6Vm8si77lA/qehV55P8kCPn7cz4bie2q5glsRmyy6nrRco
aV20j41Yd+fA2DwocinVud8zVrkYHE+l0qD91ywK3H80/SygpBt1ozaDYIBMz+586p0jFv9FIxLy
4QoBvnT0OvcqS135rmtrSvfUnMRpUdPoFt2NKwRG0eNNzDWakK40pmDylBANflRPP6rKEvF2KDoL
AcM8kIwaU/FYDA5oylJbG5RpoHzRiRME2gn8CXhriPkcnNfCmEWdbtax7UZySjpQ9T/LyzCqGcfF
tT3ZxZzgZkMl/F4htC+X2bRU+Ppwk98bUOgoDq/OEL7PuAuYcs16yWukRgXq04MPDhmioMzgNtNc
oWPKSVgPSxyV/xPgwG2uwqzpg7aUOAMiBkzWQBHO2xbexf/SDW8qdMioqrJGF/UPcrymKM+g4RIG
pGQHP3Jqq/2Vuxad5GnIEA+dgOKbcEFJlgyF5/iHZQULv2IWXMkF6WsrQcYwY+XuMj3GGzazdwXG
li1ZEyuZjGqIBXAgqf2jidVgYj4lDJB6wZFe6aBL3gN7i42oQKEMvV0Em9O1hfqMEQVSiRzFF4HQ
jzcoAEp8Eh3/3blKrX6NeKh3HXYWZ91NERdxrZTpiobhB/1gVHbRz0d28BHKNhSkKuq735oQCv/1
+iGDrzmgiwFtDHDaIPJuxy69KEdFsEM0dYyw6TmnGcCitTXsIUL+B/QZC3jqbeUDNGbCy9DypbLH
q8trfA3hnt4P/yMKibDJzJmNYctsTogm48fX2WBq82Q/i7izZgRp0GO+xt8k3JllT9z5ZhuASLaw
/PX23i1E0Nd0CLyxCE/xwPEtgRSkyyn0zoU1QL1ANuoV3H5zHLeJjyZpcZbNMU6GkG3xdhnuVSnS
mfRX8BERslj1uqrGdH/tuKykkyj0tb1DtzDs4R3rXw70SZBZk5M5YgEcZoc/X8dkVuI/suLmRkDO
SSOJBe6TvZ4qHOM6Sh6InGuLW4lFqLsDfHy2LC7aLujWhVtzc4HkkB9/1j2kmowFzG/8HcJOB13W
0R/3jodeJ/RVKOPm8pzK7U/iWdY4PwDvR+w4zHmKkh9AxkC3TSW0sfC7PHkq1u3qb7EAyLn5MvRf
Jb40M0gDr5DP+dbPjHlsaTFWsnsLenjA6F5CD5QqKUz956fFr21xAeXCTsqK59UtGlKaXCmiPPhx
9F6fM2v7wA36q5ROww924i6xaSlW/w0FIM7ft67Sk/mtLK5Y4Yexm1yzS9kxxISQvP/jI8wMl6y1
FisJGH8o9LveHUAOyLWZhGsJ6rnUXnJoGQ6DYVnSbAClVB4Zlyhsy/hKkEkZl/a7LYkOeIriwgDl
/CWV7OMI45pZI+HEwetUWcRURV95DbQjFK8SvTZeRNoHRZN2guNLMrr64Ue8uKLeEcdRxWUQCCtc
KXlq7Z2Y/OX50sSrrOpohIAapQptbbhpLE4WvaFL3P3AtHmBpm8p7V0NKFo3yEK6eIzr0a0t+lgy
fZNUU/vQvVSI96XAiV31j8oHi4UJF6xBDhTxRhzvdYozqK/ySqyhMYrx9/HRP8XcTfUFZVjbtS+G
mGKAA+00nLRuldaQU0Vd3zniZ3sdld86o5Q7HbBbuG/IM87bUmlh688WSMvFRjSGIREcWwOwXo8s
Y9C1tA9ieE+XPdm0V0Oo8tBSCrQsphO6yFQ7DVcYcuGz5SUsRBfIYk4c8vt1eF6g7Xr3C5APSgBe
tqQL1gmXJ/cZt0kFyS1c+tTWWq6yLtGQyqS0ekyEYenJsldY3sdjKEK90ny/ARLp2AZ7YVWhM4He
0FWzs2PHqgSxryuxcZl/Tyvddbaw61WGEn4rG+1uv3iG0H8IvoBNcq76yHd09UqpymdbLMmZbDuV
ebNdH7276uAGXrJVhA1jr5dDJHu7BOGoci1MkzwnMetVIdW/xwMJ7oJ03Qh7CFW45QhAB1ap2HIM
tR9rWvpEhfjWK93l5yrsbW3TXJhqNnpO+GQbdqG5uJ2jMxpd/DAWfpN/DgP7D/BXULZsCQCDC4iL
qD5CS3J0gzrIR1iuuHEyLBIlfI9+051ckX51FzIbkidOhzhWvb3uWfB+OF/Ga/Gm+zucm+Rc4RAM
gX5dY2GsGKFMOAeoS2xDgKb6uuYX+0U8jLgcn8htDiw8TdZ72WqJ1Hn1NhlmHq4SN7nM4nCcL5uE
Nz7h8Tx4+WdeaovnCK/mOqW9GMbAC5PiueBD5Xk9fQeCH+P4H8cPEvtPgeYWWH8kctetEmeMe8Ev
FoBz4Pnam6bIkQqXBQEIPTidKlpRf2Pdit+0Y3M5B0nw01qa7No00qbMBJQUtdsiPv2oDt//uKoe
O34CFgCp/EfhAAeRxP8Ard9hza5nBsDYWSosJeqbMUobnkFxFz/NDXq295epUkahCpbzOdv5eEI/
eeM3FbN6hvzbmvy1H5bva8RaA8rMr9tCd4KYHDT5+oM8NXD+GGTfPm/psWED8t3JdKHgW0r0CNg1
eT3iPST+QswdhY4sM71Sn0fBqOLGrOABXRIw34Gjib3uf3n9muuw1HhJy6R03t4Jklh0isT7Y9HB
amMO+aSwRk6DAjmrRhI+5Dck/4u7qv6zx88MvMs0s74m+v7GBILn/Xdc2SOVnHVpzbQXQ7ZfrKr+
p/doxmmqIbxD9wqNtKuylxosIzHC8tSJTZUK6/ncwMXorHiSeqe6EZ0XELijCEF8+E84JeDQcxOH
P2eaGIyUcNR35QTH3qbvj2SQJwyv7veAZFyU+amDXWHgmkzpc7ARVoKRgOZXeL3CueQb3Dmfe9vc
HXoa+uOB4mhioXBja4/n8PkVHeCHpnWBwbbWpMWOtBKYW2WD5XYmq8O3zcjj3THjxolh7t+kH2nu
oPnloQOaDnbxZtQqG0mGJA+2FcYY7dMHRUNIcGM3W+x7eIdQEHC4Pb5VGtl6mSUVn30FAwQm0rUj
2ctfaLdKMNnUtAETCDP8M44RJqN/mRcBY/b9fIFJ1P011gZChVj1SXnzXMxVB7yOL8OVJd5hXsEE
EaoJz17MSgTMnAsUlT/SeKOW0BFPjdCAptNYfxhKNm/WALOGZye7yLL5K5pu62bqCXekshDNdp9/
7CkHDxTgqgRJVMy50413w93bqe8SZLrJbsJ0pghUkdgjoZXAmGQTCWLc5E+6/SWbjrEVyXt2Ax40
QtxpTb3/P5wmG4SzMGLkmfP8icdLbcQsH2GO1baAXGMSQvlREcnbdKR/a2uns+LfWk47jAfcQB+W
+c0kAF/f3cYiiOh7WSlmVPz4B15TQY2x7rkhqBQVtGuqIeO5KSKa20NJHavapanJZytvsyfjhYgD
rJV7FhTtTnN0uSTJtpZona1PGPy4M2Vy4rpErUEjOmoxRx39E7IuIuetoP8H1BTTEJ4BYTFpqCzz
dzttVNHNUTBrAW2MiJuwf8WUpUGQbLAimA9pHs79/beDq8DJtKmHmi4V+DEAyqcCEKL+S5kO8IeV
3N1SMVnxahon/muWZasLsBhXLdLhZZKiJiP7TCkNzF/aEARFdzA68ZCXgm4tpIVN/KhYnT/YWWaa
bxLwfIxU62P9Zn2HEPPiPFtUmCyTqFlxTBEkVIHJfK535IYW+Qmy6Xxq/1g0ovG0mGr/8N8PcM49
exRy+vr0DNBRRNU3mXc0CPyd5AUnjxjkskL06CcoH+odwjIwJI36tg6Tx2XQ+LJ8mL/51OYL3dm3
x4vPLrP/zp04ppBZyN6bJ/VQGe+im7sE3qBHg5Rtt2w/rCdmm769mzTH7qSkFSDGc0xZo/CWX8XQ
ciIpYYqF953jxEhCfPARqiYX3EGF7BU4JAuyrzMJbiNxr5pIf8O/HTU3YxnclhEYGdM1UMJ+IIis
RvnmvGa+H1WJer12P+aa7ISXDKQwzM8xeYwbV4yH+kz8qEdrj96EkNoOWy+F1pf7MNG76W3v8tcR
dc1bd2hFovY7PuIBwvR4LzKWTOhstsd8SW4S6fZQT8l65d6wE0ctsjZ50AOugPYdo+tlUbTtQEpB
OhBaCPwONoyQh5ArKyRFSfM2T0Kylwi6piEOaRNJbohDSjlCMSPk8cFeVjK0z79DG3jqVIwZdBRB
6cU2fFhkdBWoknQtCqj10fTyeAEs1qep6okO027h+q7YUIyTYll14nEIEFM9yTwqfhuE/6dZTPaY
6uedA8Ydeus1bbisZH2m7jSMxAA6DgAUScOTsn6jGB/GTy38n1L3/oh/xIUESIPrOh1z6q/Xu6GA
OOWPfryfSUeeMEkXF44rBRrlDEl/3dlPuvzEBMaDG8azpZpkw6Tb39evb0ywF0XLJMegiYon9OAV
4owx2+x+KoWD2+WfgwcNWvubfEX5bjcG0gCSRnprSGO3SqPiY7p56E5kMyoFA1Rh/tTEDqAQlK0q
GSe8n53jXau4al1GK278aO2okBUrkwrCm57DybflQLNHljmmj0l9VBaSEaFbEqdUCUksBdvs7uBY
HflCXr94hHQgUGrRVyK2NtxLo2BkTZUa/p6xuLU4FvzBpdZok2vainVD5toqlMtcXeRuHINFlUHY
NU1POntekFq89gCs78fUw9786KRRtXz3JUQZHe6y4EOfnU3Knov3ePmrJYT1GvXTNxPBKTbsjHJ6
KNsGnjTa0x/OzFjarYx/4pmmgUliWKPxCf3LmZMQZ1rEVbCG1iylEEARakmqvp30FeVgg/cDTA7E
3y3MDy+y64JQbvrH+EzVh8e2Qa7tv1etldk0bD3n3hQAHqXDJyNbm4EKBJyH63Xv48FP838M6RPr
5yL9ITTLxzu9uXxG7+Y+A1HMES3DUOei7UZ9eVc0HcRDv6ku3Rfn+bP9tRCiguK48LDMy+jEHba8
iK8d4LdfWvNi8zHlbaFmGiQWGY56208WxHkiHR50oaKKxeJV0vWYwzoP8RfRfYy636DFK/rfJ5lT
Loyn+aL3XYB6i6EFZxU2wRxcemfnvxxX8Vs8afs/5wYgJ6IrjiQDbqelzEyF8SqyTc9JgQXMsze0
HrzGyybPMntCBO8FEV/3od57/0g9ubkYhPC6qXyLttVJkDVzb+3YwhwIOpcPAwislkQZ3BK1BSGK
islndB6runzaUkHq4SgAqbNJDUoJ+m991D/xbbSCIaFRG2nk64N50b6psImOFsVxy/ofgXAk9WvK
p4+gV90hL2FUBT9YcU7lHaOBIltcxp0zL3CJgsRdqv32q8IFso7ow+eRWwaVzy1vfQiWA4tccGLT
rB8Fc4ojHqtstMr3WypKD222ndFyx0HVRwAGlD1gsbk9SQlcADhStrjSVoPa46D/BkPPu956Od4i
2lFZ7imE98NWn/fvkJH/w0ZOiEr9quZ4SPaAq9NJYK+cUrZiJHqCK6I8a2aQYVnBxsoxRs5K5cV8
97iB7uwcG5UlSuBPiIX1d1JG3vQgmeGGeSigl3cTME+9LDSYnihCXaeMw4QZgQUb3cht2sfTeGMj
9UJ8TFYDY1Dlg2OutSRFSCL1ouetLprrf5hieRCuG7Vd5oVw/MImFY1ELIXFYOLhAhB5La+vgnTp
h959Iv+o6aYuokJkmzL/K1JIX63wHwB2eeruaBac3Iyt/+RTiwPTW9c/TLoJzvJ43s6sV3P6Abbj
zrPUBufkuDcsDKmATCM8mF0/Mr+efwVzgHAmZNthoL1Jp3SGRN49CU4EcztqBUWoAjLg0julXP8+
2+zm5dj5O3clriFzuuLREgmMh9XGxWZmGlLUIinCkGXMi1Wb1RuYd70GeQTz8uz1UJBuvsBpX6XC
gJRzRKKBizsXZ/XamgP/xDuWoRA2rKAlDEER6amm72jSiTMR6WS9PMc6M4T1b6sqDtbnyYkcBZHG
1/e7wpt6Zbuft+vRZ4ulyrE5ctqNEUknjuf9y83MBEusyeAYw8z72SkPbPzyhP3rCR3G8C6RKeH+
/ppBnOBINO7I3ox/3w3Gi354R+1h4qvGzeqZyO4J+/zTW+v5TeGDm7G5ejXl3zcnXwBSOs7yuOzs
dmGlg5kqTm+RPHW3G9FnNv/bgp+NmRJeaKo0ajYF3Ji9mNwXmQCzsJr8KvEmBkXrKk5KB21EK/xe
onYMBpfv2qXzfr30r8adouqD1fid7hWN870F7b8NcFIXoqTw6KN824o6Z+lqezNLDua8qdkBl2QO
R5RLyHr/TK7BngH7R+GbvCTOIW+52w4PLnp1ymm2CmyVaHwaQHOVDKZdwGbGkchieT4D9aFwHZwo
YVC7RbywXOpToUC5rgOkRdtPZh2u9XuQ4Yrf4p9BOhEtx0lohCMvNIk9e0MDeOVlchbZXWv8zijB
/MkwCgN07nU3ibqFdGg8Fgd3MlBkxlkmmR66j0PDUhp84ltgbqEmSoS5na0kP4U1g5bN+PhxL9+Q
nGcrAhoiWOmhFpWON/5Kir/dIgUTNtP0CvRRoIxW23wFJ0LA0J4ZO6P7/WmYxw+JloXJWKEXu1Aw
y7oM7GBctgtpXu/zUC7hw6N1bZD7jSIsub8nFlCimyvygAozyMr/243Vv+p9t+X1WtCl+QFFEXUY
c9jqSrfwbE4r5AMgb4zaDSin5zZwwMPQ31EM4krYfusTs6Sk4yl47BfBgI25MqQMTitsClXjoHEC
ZiZ7fAIe0hRYi00STexwcz0ObNjy1dAy00IpaCVW+dc8LnugQH65CVApMuptGj1zXKhZOzW16pPz
9jTaYr72ig2+YcLRxeofAn+7w9W9xDJedzhQssqM59jkGAxMmLm/cNkVkMMDbCR8BD44Qlg5EoMa
Vk+448ToF4OR+qQsgNe6H76k/eCzyc19PldJdAJ13gy7BwX+zRn1GUSnkle1tFiDTjbbW4457SDM
UKgE7D5Tax3CXcQxMJgaCa9VnS0rZg88QZb9bySpGy1LwO3M6SwieyCB6YD4wk0+DFvpNmYZgseo
GEraRKcUbS61K4VYGPG+rruJcq6X13/Ag2yv5yB5As0C0NmYJfhxTT+0KmMsxPij7GN3NF5lSxlI
lRYumzVxEw1+IwMF+ym63DGxQ52/ObX0OfV9KwGEwO7Qjtc9SxkOSdU03eyI3h12DwlluaJmsw7s
lGcQL8xNVW1jj7grFmW/zoQ4T3o9CjSIfuojQEeriaSJyM/VdzjTz4QLlP/dNcUWPdqN0xcYoP7v
YBt055eYMP5N/CcTx4yY9nBYSOLKtSoWUuhtkpj42K43nKMzgByBG1UKGgdl8MmCuxal1JneIxit
OD6WB367wRCsHoJwUj4jmAF6PNnL1MjsIFsISvpA3GVX0E2MwkRMSfiyolMI4ArHzkWHLSxPiwfY
Aee2NyzIOrX7mSlVI4ZycTtNR8MfvXH7CW6oOoxCalpsgsdN2ZqRfvmKBvBpCGoTAi7ZwGV8oL5r
ZEc7rhJGKcicAzAiF1Xb7Wtb4VJJKYwU+5vDcnFOxTKgmIVmP+9F8cZHyv4Af0QEibZ1bhUP1mGf
Mr/CVdjq/bHwspEKcR4V4Dtfz/gde/pIqOULXCwaZOOSfMSrIdLPsGNnK6i+dhhHJpIDKeA/ujLF
BT7l8UOW+3e/8/pgD0bSGhI/BxvgCyeDlTDE3PwsxjFxAqkh2bAS6gS9oYoc4fQD5dvQ9BYub/MT
OXfvAILBQFYb8avSgkVv1kW6W4b5VCtTbthnK71w6ahhggwHGSpbKXhJG6GMPNhwfQak12eopaV7
8dysPE0cOLfoAANwCuzaLfjJ5Gj3qThaqL7jUcjui2PDn5KTeeIcevBUCjBzkAkDKmx0yl6KHbCp
NG3nWo0VYsJlduzzAwjLYPOGtkraQ8jWPhFnwJ26NIEZdhDR5EN4nanH6dXaYmmW9/eL5qZmk56G
k8oPgrMv3hHN7cpS1vwcOSKPiDIm1txVPfQWvBSVsfUHcKYJedHpa+Ik1kLvQfdHFt/TN1/sHun0
KU0mQJrb2wdlwaSRtR+35XJPyyUIY09elergD4gOZoX29U0adCCWZIzkOTlhpobBD5AqvudbmLpI
8XpbqafwF17Z5/9o6CxPOj8Q/kStARGAIcA3v8PhYyaVU2Ra8wu3Qp7DBQoPrWtFv7JrxoLGxLQ5
iJ6a0NQZIPPOgzEjv6GTF5501mn8wr8Yxipb5sQhCLFKczbzzn5sTq3RUJTD2tgtLFiqTicbiXZX
QjVmQT51WNnooKbHcHBL9y7c8owT0PxgimYe2XD+kW3eh4dl0VxH+H1YTCj7AfaExJeYKHOw+boh
xbtPqRenJwkOMdoLdQKgtGWY2VPni878S8RiWAxDseHot+pZ3vdwmdfUcdgxnet09foR1820NW2u
4jlkpl1AhrpQzS9QKg+/zNsbhDg9d1DnqD1hNXoBPiINaFi8IteFBOCPpQq9N2yTra6HlU4qQskS
YbGB4UPsKV8xq3l8VUA3XdqktQKvwfoJnfUlHX7rASzfLbXRWqypTjs+sEjtTrlFXtaWYXbneOm9
3f1t9s+cIoogDdQAF8DJ9D++szIsHTgZE0it0U1sZOe7v8P004W/+CEjSXe2WgA0/S0G/XSEZ3VY
Gc++2e3s8oMCFDDse+S4T5ddMwxkxRrU81IJcpI+qi4yMG4GHcogDtTxC/vpgMljLRADRtMbr3rE
nXU3kJOOO7g0kuTxCCaX+ZNkwx6T0j+Qqtsh41mQuc5FmSzEevwQf364rhRRJaduhpr5dWIGnKCd
dt+S7Qv2Z4O+9cNZuDy4VwY2XtBtrOLBNBs2MD0spTRHEXpMOtjmYz5BLw9e666UnMDM+grNrugY
zl+pXX57pJPxYgsmeEYhdHnbcX4Gdhq/DvJ+iAlipNb3UQ+A0+TnWxd6jLXtkOnrV6ZhX8Ym8RRQ
If312GLttkMTZjANzSlq+Dgabe7XrinHFZf/g3J7heRUDNZKaU+d7qltgaihkH7KJ49+Qy2aVMsi
VoMeSUb/wuZ/cPmHL+DEB+uWkFRuZKC/H1Da3j3fG2dfIzohVUm3u6z5mbHHWyo+90uJl4JM8PZs
TWSHS2Oqgh1dns8TE0UWEjcFM+PAA66def/lBwWt0l4gRFNrvKbTcuz68UdHP4oO2W3ihSjlOfk5
Rir3kusvpFGqqhipzlmAFsh1N6N9YjT53FHT2a7GtiuoRSJrb+PzynGXc+BQVdGtbadsorxb0aMT
WQN3XZbEvKWhSGI58VMD2GEVki0aoS6mbvggplfoXbZG9DXqAEmSxkXr4U3luC22rf87yGH4nudP
B/XgixPodwpRZ/ST9czdxFrRsXNyThlesIHa77Sxgnily9zLwUC80lwTl6b4lqjtl86BxJRTYJir
4ztoMiD13R/6bpabmuSOamcgie9hpmTGbZf4Mk4qODO7Ay8TN7x9PHts0BwJ3peszn0AXidbPN9J
8cagv3kZSO458JOV8Jng9PfjzXNvrpLWv2s0DX7IFu02/t0Yb3+dVIWkFt7115/+Sf7n9MnwVzbV
gIn5xsPHzw8Pt3eUv2P08zZA1YKO/JV4mQado3XC3qwwzkmdoRuYGfkxPAfwfswCZSclJvvdXpZr
iMUATdVNROLyJgmcsCdpr8wzTuKaflwyEFjNaqXwbGNSxvdwoFb6nsOfmPwoWrlJky0aisRbcL/P
VnGknIKVRmsuEGhBHOhl53iivIDFVbwwprZxt0FifCuvPNfu22uwyDwvUruOLiScaZQ4WsLW9i95
E7W14ULpKLTovTPk4PY4J2E2XoQdZBf1VOyUEQLHZ8xVZgiKXKC6LCqmRNARBoyhwc8JUPTypgJR
ycEgS4s56CECH6jXZHOWbVtvP9WY97HgmLQOfuqe7ZAe5vCL/SrJBCuOYFgReIl33JBGLjjeoqsP
05vUztTmUX8pR5MKJycabLRPjWVkgx414dR1emL8FvvizODS4zBONc0guQGKAzUi64cH8lCriwRl
6GqD5+22Ui1xpUd2QFYARYPF/P8D04Xqwuq/uhulsYi0Eztkmw4HER2q5FhMZcbXcAJUfkMaUdfA
m8B5SxXjn1Wr4R+yi/EpnvMpYB1v43ZzavFssFse4d+oT7qCnaNplkHPtvJIh+bGKaFf0fZNtVIK
UxEiyPqIH5oSY9CnjXdtloKuVaMExZPpG8fam2CX/9FA5qS7ZOUvN7lhNQc2QBVHTZ1ZwVliO83a
XDPMLTnc5Ndwicxemm2uomeMuGEjlvGmsT2Js1INyYniqO4OFNWclrAqYgRGICRLzS9rTNKNqMXM
tOPkeirrIdu33TEiIBvymnebB2YZOB/yInibFh2gzz/+zB7o5nrDYvCNCow/zG1bb/GJsHv5DXsh
pMjfwGaeCyXg6SJUL22Uw3fGbTWar27c+kACITVbwDuEv9DzI0ffDf7/SlwpHJCxHa2gETR5zhpe
LOEN2VgnJ18oUva6yn3TJT0aycJ4/HIHE7Rn4puMfV/3fgibAu4aUegElkBm0TvYrfL+fA0RkY7F
9CWqn+wCvzjahpiWa6zfdYsTbLZesxSKjshDctVdGjNaVKZTILFQ3EJsehYMR+1Sxs8yWHCkx3Ef
yuTffbTgRtWwL1U8fsi9Yk7raHn8FgjouPlkXlxUCRnYcgnLp7lF4RUHQNaAGvt353xCNYkhZhvG
+S8E5F5K0cCkBOORSHzvgOdjFQZhgIJjp5KIZyYw/ldgR8PljieelM6M3uMHXtHw0du/wm2QFGmn
PYhLsJyn2Xy0zS01JIY54PsN0ZhynF/ldPtHbF0+yPHos95EAKWSC6rDM06GPOOa1qivWzVyUPIf
EVuT1p7s5BzI+DxNZ6thJe+q0/Y4UUeztV01yWe4ofAFamxC0grWL8RD79+qh5vDd7VP6ciJjZPb
ghVq7oRHBuoZd2HBkD4qNa5wK/2evDsjFcC0nnQBtryQpgl01en07ur5sToWrL+Q4pO3AhI883sv
1wn24oOmVkycfYukgvOjHJBH2HXpsTRz+vgdamPoMmbnURmxx/01+O4VmGdam5zkWZjMvz4UHxVZ
lxQ8Ad1H7UJvTBoTFdILT/0OKhhR/3MuClhNxm2Y2n7WPA6UU+9eW3sDHDjC3lRdrlxnP+tDDUbd
vcAm5YYUw//D9aOexnWuR+3726OBVtVKY8Q56XtLU4E1mIgpY8bTFIHG60a9wh95qZOEav6tCEeU
sfC8UUk2LhxYjofyf9ZO/9EAZs1FrqTmWub68AL4ftHy2fva5T+VYVJzMfTr2Ro9hUOg+vMgw7xW
vf1vHlOStvp8dFkSORMIZ5ZysMJ5p8BG9XZTpUvr2YdajtNuwSu/kMK4Kl0HHCTItJ4DXPMJc2iK
18Hts0Pcg+NHkxpm9FDiFIu9KV/yjaJFc1n28qAd/PXP1NMtNYVyoWJq31MOeHY9LwF4IgDnF9VX
N1ny59Fg0t/uONRFh8+qXK0BN0pSRVMuYA/pf0vxyb7dqq7lbPJ5lp82UJ7x1bE0h5TWT4CMk2y/
VonP5JhyQEHa6sckqWWUeo66GaWoM2WHXKrvTpKa/T75yxf57cZqyElQ7khXWJch8cOo+BFtUOiR
8htglaQOlGuIQo6VLrpQzZ8ppOzf3nTKkqv4ODTT334m6dMLkyO5qRJz67Cpm0J3fTvdJdCLL0Dc
by8wbLJVNTkW5ye8ypYRIrG7pQd8b/ifuEKSRfXPKUVKujkytc6Se36UGaP2oW+g6D5K9dcz0cCa
85zxhUW861qW2oIFxZ7NkJVKY9pLegkL0T82Qv6OXDFFWPxS/5pVLfCg5IiXgqaoLBKV7EtjFZYU
YJGKygtOtZtY8VzngWXG8TSFQbcuTjAzC/Mlsn+Oo1khZhfGbfJqofVAg2Dy0NUbHt1n3DIH84Pw
1Mvvkk9wbqsPf4RDva6CbTGa8t2R15Wg/AYSs7i0o6BiZ5rBJ5h5YEKeR5IdeA3E5maUQXWEp2Ri
SEqDRne6WBF4ustzDkq9ZAavhdL0kYTYyXfglVL47d83VdsuDytOoQj/cUY2CPl/lNO0amGMz2A0
dVBxh7rg6Yw6aayn+mB6efiovjKQQrjvGoQAOaPUP/DAJlp7V7n7hpbjonlca+YMLBTwwGuWsSB6
TdD0dngW9DjWPnwDM7wEIsqjoXoF7PPZhByQ/nXMSFQ4t9qBxrqpnu6Xh964TM0UIrN014TdMyAa
55dNFNPpkqXlI3lIEa2OsOWVuQ0q+iH29GCQq+nhqbd3KiKyoVKXTEzN8td9CT7BaItet/ThJTj6
KRHYCix9kbX58q7oq0dZUjpvUCX/8SiBJlq+XU8c0c22b6hSJ91ZqVgtf3h60xWKuniY6ACx/rLz
rKa3fKIij9dolZTnxsHzq0qRCwsGMeihMw5IHR8AG4QDp7pV8/t3c3sk+ylf95ye3cFaxRwLOkCZ
78VuYzcWxOl0NxfWaA3SDU/QRNoJj38EApp7C26XohjX2uckLmB1PJAS5keQjYiJL+WF4pY2op/x
eaathV23YQZEFHxORu5dA0o2XviMEHA3djR32pBTugmAez+3PPW5KqXanPS4o2XrimdfU+cCOCdF
6H65xrsfToFcV2xn2lK2AJon6scGQutZ0+d5FHplSx7GRqVC0ZVuLBXWcvGKxM4SkkIc7H7j095w
JYFKSn3EQ17pMrUY3pE0VEiplSRt9wC8R3eH10cdHbD2sAkxLJJLRgM1SyTFT+fLWdp6sLW/BYkT
YbdiawDXy29Gzu9OogQFg/Ug/R0DmFzsGU3o58E+al2lK/3iOVNg+72QH3Um+HVI4MphtTKaauB1
dpuJoTYa/aLR2YfLXxFvWifVzj4sU8wA7ixwNArvyfwr7XPg1TJzPai6y3JK4WwBf9HTodXr0hb7
D+Z4U2UxHALEm9iQ0uD6id+TvBO82eISMMNM5p+09fleG5uUrq7Qx7LsRK45l98igcZbRqMoJOz+
ZB2pw/ggWKI/Wv/YXVLzMhmgIUbPYeU3g1TlzLxiTuSQkAGKb3+UtZis001I8QMfLuP5HEUsIQEa
rSExcreMtSiAE8/1336HXDXy1D8iZ+/eL/uTir3zokqG4fSu5IzI/Qjo19Yk5miuZoe5l2Mf5A7M
bUJSAVQSx6zchjWYgnitrplCCrQVtpyx1jcpNWqL2QIDwBV3dCwQEmtM9HnOUBajkLtt7ggseHqe
sprkchVN39vJonbFQ4ryBcJH4f4JRH99iMF/gYwqTX2b5Yj0I29N5CUGhoi5RzTNvw0kZwXVJ0Ju
dq28yhelmGYqhcH2CfhOIvytysjWN/qz/kveWhumm4jZVwlVhX5Xd+kDkezG0XrkzNSopdMqiY70
jqsIXPbJk1uk7UMjjc1LAr8kGUrO03Ls1lVsEak/divCn6LuhcPMm14AXXugolZGD1PrkKYdCAUZ
/ax2W4zYFWHq2WbLOq3WO0O96nEYBEJkgAf14G9I7t4TWkN2tEeZQxALY8+J+vNTaaGFJlfUFYAZ
ih7FsTDVlmRunAsAGSgJ73J3b/NZDuPwTXkyN0rb7WYaNLRVFbJwej5U/RianzglZliDSs8Xh/yH
Ag+kSrMRp/uBgB2w/spJc8EwIQBiSh4DHyEmX2GP0Lnqjg7rf2e44imz8vyy5uZxjwCnSHeWWx4U
Ts7ju1t0VhiUlDwzl1+CMY/PoVl7re7/QGU7gvFRZEgotvzbluHD5q55/my33w9dqk06KW5uIw+/
e10Z90HyZu/JQttNjB0xyXUrEVqOaMUqxld9lvGQB27Lcut/UKKMOYQYWRKTuLPKdEW88KJpK7+Z
bE5kEiDqtFNG1JRSeW73qBK8ioDpaj9UPhJfjiNXG/UIYktv9hZkrs/MVAtiHOGmI0htqpub0S/m
coHAY/tx++3Y3ddZ6amTnoLTmiyBQ3WHGYKAnDx3bbOU3Fd+y0vqZQA8Ucmya26II5IcDB9t1l9y
Jhchp5tDFMGayy1CIRtNH71MOmDovXGIoof0h5IXsNuZW+cc6DVR1JUdmt8EKB6d7OH9JYsRBTZH
XKp9EPKlSt8buvXhtTgiYdaouZOrKZmaz1k+QrT9cP76UcUlfSCR5FNYNFh+I4HI752tDdPOsnCR
FV3aRZW3r5YiZqSSSeA+ZkGMmSYZr0omE/kf/EIHcPsUQ9+RjR1iV82/UIc7poFwKIH4sioIi+De
g99a91zV5TWKtaGdsjTQhDoSOnOi555R2PT3jfS/B5aQJlBChTWKBbPVFSy92sgXeYvEg6muLx2z
dYlOuVdWa2eyPLBu9MjdFNi4Vu43Zw+oSRd+VVtHAVan+NgE0vIyUUQzwiG/LM9AkoFVl+JR8vbz
f+zMRevoCTrhxdbmBuwIJtRMCnk9ztTX5i1KoTCVPuFvOaTLEBmFngfZoIloBW90izbHVTFHdyln
22BsGkAkEJxgT4ttw3eha4wuYNn330mgacIUGTNSl8AuHvH7hNep9bcFwOjbCo95QXQmfTRDXov7
/K/gH57OQdI1t4Yu27opOModqKRAhZwpSMcPmP2aCoAIds3DcL39uBLR5b8KaOpxJSgJq8r1eLcl
/n7cE10HVcqLiVfBnO7DMkwJ07GJSCO3L/bRMrW9suZOfHlxaRTWIkqXH6MkE1QOW1aQBQfgR829
/DxGT5ExLwtjXHYvGrydic1cW9usfZ5I3PVxzE2e2LDawJKv9HMtosVLCO6KjqkRxJVDyY1KuYgr
CTvjuazcFP2ZD/VrLNAPBG101WUAsf2jQXSHB8Imex7bxSivAfpVVKegwxwlBvPRA09+WUexy5vS
arbwDvMr1+QyT4ZTaIN+6B7qztjS2y+WhidJTaQvtdRQKWGPW1grSZ2VhZZ3hDx4adcjFZZEpgUB
CKZRrZEdNTkw9VSEddJQ+tvlFiJZaij6Xm//yNYzX6vU7YtNAg/r51cF+BwwqV/ahjo/xl/LFGYy
b0vV5qCSYnNuZg1Uqh/pCFCKsgRrdoDu31UOT8+Ml/7x65JDfiiiKwSz/Bzj8vzixq9AyczvQaKr
r02oVpwn0uc/q7Z935RHBzB3Fisxh2fYZbE6p4XBIUc8tPp6N6QjKtyjKV93DrwBfRG7Zp2fYiUf
oTQbR59eIusXG+L6TQvK/Xzp2Vt6YM51nbUtkEI+8g92q8xB2pZpNgwAPpQHOBqlWWWcuh96Sl8e
FIG2GYwGYx3rayZHloQh/i8nVjHncvafPs2uIHdBB9t1VU0w57ZeJFCp7/S5Lft3MuNX88YtVt5M
PzzRUcYG0N6ZWtpQYCBYMnqJJRtJdibUNK7hjqLYlc5o0hrOeUziAss7wAmTZUM0Cn36Xt23PLUx
hEaC0X2LftfxFQvMhvqYrVvTA5T7wBFUI1eh1AerVNxq88cT1x1Sf6gbbvosOG+KbLmXFC9H3f9P
fwZCnaW3iBy0dd0I8RdY0mBTU5wk3lN9E0F1Kln6d8HpBTduBKIf8meEw637wRSn155VaaCuTgOB
DY9AjrJYUal+2mE4921TWfPHQU9U2hISFxF+63lqVM+s92Y/D1PhNVM7IhH4XkR7NLKaElHzHjoL
DwYIQScGK7rXKUGEFDpRkbcFpAj5Xtl2vuGjspVHT2afmPQJBYolcM135qTFrcMsruMYEQn9669x
UMvil0w+GfWHNEBFOQRX0r6dID9pDBg+k5TgvlnplzaGRwUZ1JyEG+xbR8XtpgNX/WKQaaGhm7xT
M2UWbpowGWmcXlCi7MtyU4Um6SXPhZjFO+PuLof0I83poSwXwg/PTyE7nPgrqtNbUCOgz2s2hah0
OTI7HFx9TH/oSdL9IogmtAHtkm+ulj+89zWDdbJVJw33rlumxfwsW2hWTGkP9Cj4yDjFcLjRdRux
I2u97I0Rh3Yw+8XOyPUuTvazWDc432mGR7DVLhwhO+xnDbGZw+2K5d3eD0mBrLPDdLnforEMJ0R3
C/UMCMdpYbGwiZbl0VZJ8iKTcmqLWpQ+j1sPe4cCs06FUwkTGbrO0A2rWHxBMABOJoCJOVyvdIUN
sDRinTeZpAST6ZbBbofudA7MP5afJzg7B+0c72BWFwc1YEjW5E0U5u8yJ1magfPnum4JkTHpFMTL
0R6W2/U0nRyEfVjG3RPnuwWkuf40mtrFcD9JUEQd/VoSAXqI/zmgA7ThTERN2DU9xFYNvtYaDOOu
UUesCkJg6kyKW9ly7d5LZpQ2O/gMj2BNch5glxvYWSXpioal2TNpVZqlQbjn4UJb6xFJw7NHnAjb
teAHnhoAoak4fiE7XnqVPGdrQwpvGtVvpxwmCvJTsYHltt1eqkdHjaiGc0C9J4zxLptbTb+H7ncO
/en2C2Zrx05oU2HDdfHfNH3JFO1VAPh0kM3t2CYQpcmrjFAedVB/O0BWHwu5dZ/gwRD28Krattzs
EoaeTF1EjWz3FcmDZ3jRisI6bIsskf+xJhRTLyrXluC1NPO+9cXrJMgt/ZxQER3HSQj/HPsoQUeo
BqfyNtsvh1V5TKNXWOW4GXXFrC+BubbBxW3BlD5uDEjh2VXzuVOCV0v2+vEmIZpbT5B0vVetm1kR
vbcJGs0YuSJw0J38+rUwL3RmWrAf+TvRvZxdQj0ZFBqWc1WLDrxli5rAcBikxlLzgppNKWBroEds
bjfUEFU7wwZ53JtV38L1qiv9zQCQbyU2FiLxm5MISn3JhSAtk7s80QnNZxKuqaA9L9wH45D7ikN4
sXVBxU3MRgDavQVfFyFf0tXbUkxdd71kEVDZEOPja3jZWoIVnGYNntt92To1+XhiDKA4yMSfegcQ
vmWVofgTxL9ap8a4icIUX6pXEjCl3M7z2fmx/+3bM92sxNdMMhS9wCg9ZJKXdjwGY8sL3y3BUGVL
RYJjmacDpMNv6URnGGLHOP+9D28WqYgSN+Q/rUHsnc+4SyjM9VqBZnrMFJaktbti1VLPYAwKvc9h
hXP5pEiOSQb5mzjCFe4nJvxTc0GRup3AqJCPfV9iJy4ZOF6gPzGbCImxUMYA9pc/G30TWxKsobpo
A+sW/ThJgDgXmNleM+w0019Q2DObciwEW2RWaRKJ1aDFsSsy39CFv80vTHBi3GO7TculsmthSRCU
+IY5l9Et+KgzbayUyKzh9qim32kfu3IzXcb1JzniX+8nNJLeW9a94XeIEaAqcOOKnaS6Z3NTF855
yn8Whz69cpmVpVd7lKEsSV9KkA871//jtrgK8JcWzDJ44ELGFXhvKKwpoF75XAZ6lM916EIQ5rIj
UI7GkLHEBP0XoYTpYEl0KV0Lkv9aTcIclK8FtQqHWj+L/tVvv1E8WZwlPKEEWVevMFzrBGIONZ4p
MHQ+CQ7H8q59sUhCpYoRmLLw9ayLor6ek16W+CPycq16+h4p2z8/h/+hn46WEQ3DUCM/foxqkGng
gcpF2NutPUpdgoel7fiZEPzaFBRLFaY63k6ZsFMAggx0H75fdxy/p1Gx8Gw7S9yUIwrFCKCsrUGm
J4eJhMyFE4idfGJgd2oTKFAoPepxrRLyVznYC5jETvaj0Y/+TbRRliNvGJyYm+nv3k6RzrvEwXeR
VnFBfn+2plhcLyNH1zgjiDXICRyuHnIjX71i4h05VYYSXeEcu6hwU8dVjYCYA2x56eKS9Lrkajz5
8+WE1IL4FZWS3QaCmJdUmSJZT3NYoM6i4YiQiiqm4ujtQu48XVUAWRAsfHrxw6Uu95UL+rf40WhH
iK5NaFrq84zzdMZ8zU5sef5p5MoGs8jBftLrOU0A9LrSm/Op6ny/BlfopeNzewC6k2hEnjlV9b0E
fuYu5NxHEcIMcZcjNDWRVMPBDlrQyJ3LwfBewR0YVBf/mEZ9nZdFpExrwGUEHnKzwCSTyLO0+WOg
ZtQS8nLFELzVfLsdLmryoI9btwRwbDMRA4R2vFSdh7xWs8JsRVNrQmVzOXMg2fSBJPKo+8WRRbqf
WxK8+1lyO3Lo6iS4acfkqrIPSIMmzrEWeaNAKflM8ZprgPvt/BM+q8F+y1RlN6swLMH4FGy2QVAA
nSLv8TDnE23WAcqUpv7/3aJOB5dpo9RQ5Qfk
`protect end_protected
