`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
QayNzbaZc/1O2OKrya+0aKyauykpFD/Tont3uuwxTDTfkpHGnihinRXB4yFbHVKO4vru/ND/lpXv
JL1cDkcBvdbqJieyTu+HrZetUvwPTOI4kywJkQczbMj9f5pVmGy3i3reVvf9/KWI2K8nFNKCq99b
RGL43JQOx/dVV1gKqMBM7NtetkKnfoqbPKYOAD7sLFc5d39Nq/jBXIzzl4QwThBO5tIDTGobBYn+
Brc1UkJagdetR2uKIi6NbsQpmWpp0Zo+Ik5yvh4GhoefIKqgEsyk8NAIR6OeUG6oPCwU3WgwWspv
GnmjsMPDwKNYtGlR0x3eHK3Nqmw/sJ9xROn/gIPJVikr0InczwPA7UPcM/kjYcPgh/KkL57y2dP9
WS5AtSsK4rQqx4kUY8G+ZJThRmThW+xNEb9TeAOLfarMb1JAcsuLApf3rL6UK+6uCUnIqt8Hm1hy
PYjzsqdV5nWEkLZ+0aazVsNS+i68giNyoN7ucXMbzb8Sa1YLLDNxwhsOx+0wSh5Ka3JkVeB0pKx+
5KP2KpfQ0Js9gejDOFsyT5YDNfF30jYFBuBP4TE9yFsZrixGAgdrOxjahTSkJH681VCoJAHyq9yj
CwRHknFWFQxTqri0aFk+2GHv0IRvZFuFfGDeB6Sdv3feAqgIu330txHmaanWS/oW8ynm3YBs/bH8
ZLbJWoPPaNihhmVdBC3OGvdfXFTY8Y5GRhmCwqjVg87kqxx1qtEmNaCp81Mh1Gqxybi5dRe8P9Zs
++AMyjQmmKzNc5Dyq2VEcEe4xtb9Nabe5xB/uQqMOK8B5qZ/q8K2IbqvF01/ZQj6kQrQBn/XSiAG
5KlYpFJ78GcTt+iEijiEwUJt4GNeH/cRxnGdvsATjEpwJA12djfjxidyFrt1RomwyxyLAy4jvpIO
iIMjjRSuHzNQR+yMEzfrdyQLEBU/XDF37AornM5X6N6T2PfIElTPn2oRSuiz2SBTyQbwhORheC5D
RTr1cQFp8X7J5jiOtE2Lagx2lVazXXquDpDfs9yykbQj0aC1nqsZvy3XEGWds+QiclpdhIuyYzWb
epMRIgjSxL9bjkQPNFjoSoRl9NJToVYZp29ZUFHjwAkLd0yXygPki3M47VDcLcmQp/CGQ6J8+bV0
aajuxn5ahVFFc23s/+mVqZSqSVN7tLeWq+XoBF2nccpksG7L+2FQYTg14GA3zvFLzgEDTBFy6Fk0
nvmyBmiDIOOsHVz+vmRCvu1F/hyAfPA7YASOz+5RPMQe3LLYxh05AZKHuMnBPDr5Xh9F8qyNNzRy
T2UN9Qz2utC/8qmUMO2qR1FVsJAKkSrl054uv0Ea5vOvjCUhwGGvxZgrXzW/E/gn5p9E0yRWUfcr
51OuZv+nUO84FOQ+XlBEVKoE6ug7In9duxBTzcGB+P4v0+koa3KM9XLlRq+QkDQ6zAZBx6yHZgY+
hzupm8TylBr8ZUcr+Njd5uRl8m/jZ6jRRsiVJXt7h7++RjgsgFKoraYeOvBlX1tVYNxpkibtK9os
I7CIk6NoZsk9mrC39jujHD6wSudrqOo0PUuQZ4/7PAQD9e0kOJYI2RHeO/GPJn0bxpUeDd0sVV7+
k3eljTXhdZCSSEO9f2O6+FTiuT9mfLtxnkIIRKGsr/H0EVnDS+RqFHnl3Y6CGNnEJzBfyPbBxaSa
IaLuqTm9nj7CE0YVB1mNiWmo0cu94odnAsi/JucJw7Ga2xn5zcqEP2Lb3RZREHa4KM3n8op71kkh
9Tvl1cnGcDRbzlbNfo2lO++JFgTUn3Gox12spAHr81FHffi9/Q7Xk3kffvXQrUlik9tgRFFaSDmP
ol4A2UDydZSxF3b98a3Mpt+0kAZ8kJveTVkFv+uapRH+HGFyDZTkuqGszxmqj8RSlpo2KbpFeCgS
VWgnDPzKN7u/OrgK2yY2D8iThcohHdXoAaqKtP2rS/XoFEiBJTROWwmsoAErfj4IxhEB3K/zjc4w
gOiGJItV06FXopQCmOCu+4n2iu2qxhAV3N+X1tGHboY3s2/e18K1SBPKd6QJNm1wN7TrGPSWcpTp
TGJeZgddkJdL47LtN4D/aW4jeErokTNPy8jZHXI1RfPd2g3pYN1/BnCRyVHJLYFQ8BM6OpRQBaye
eapihHB/P+z50yaTayrNJbGjtEkDQc3jhSxA8eI0D5s3dA3wXLIs24DgTOcqs+paJuSWIEy6GFEr
EUZZtfS6TUeGgqxksMt6g/ZM/67oVsuqo3auMKCyfYhVk7Wb8p38jfLCvnLn2W23BbnDojzCTNIs
bn1H7vd3Q8erF43k4XrhA/AE7GPWqcplSxCYoHWAk4UUwHpz1z0wT59TdOILpQRysN4INkf1Cota
pdhAYBoieXk1CMk8fDLKsaJAu9aFJ6FxRNmeB2rqnL9Yxbq59uA9a5OhJB9Y8h0MU/2LDhYsL5D/
rLveK8L0/Ekud/gxaKvPJgRnd78H4cAimRd2buGET5R5mgJE1An2nDa2R1xs6L9/a7eXhegb13Wd
5ePK6+BzE8inOxbCSGnt+Y1+jO5i6AY+q6Iqbi0YO6ol8ggHCcN+AkLk9moi7mKw77dPGYbwgI27
tGxQCHusopIIpr97XAxsPR2DtLRF2yQUHBRIw7eWvPrzF7+X3oLyS6m+U5zI5CKEJ8Jh/ouCOzom
+Uj4sPuNQumncqOnu7A5GkHd5qoT2T0jtH+uZvFBISEzdZRwzhTC1y+o9v5vEmTReU0EdjUFmz+r
imzRI/KG6Bd0CVN7Tkp1td9XSEy2rhWtSGxDAGyfDu6LYaFTiCEDP/GTevIfvuFUlM4sr2yylUyI
Y8vhgPwNvGQG/VjBAjLpP8LGqxgtNBjM0XJjzgnUE4CAmMJE+nmfkWg4DWRJVrHi50UOjZVPXqWU
UdGoct2ND1+9xw1GXr4tCD9+wBnp+FxbYGBrs44WTBrSyVFx3aYYv2KPhnv9nqc9iyKTGmHUbkiT
P8pdhWEsPrJCq1IA5jLupRZxcg5XM/ZjQjSIjaZXgFZSKldIE94pc/5T05AfDDkcFnD6nlpM/W2k
FA7kCI989Q3PhWJDdJfujzqvWaUTWhG6tp5bOAr/DHllDxwTMl+aj/JcDJv/kO4ZYmM4F6Qp0Yaa
Db+iEpcqKSS1tAimpUDlaj+5posrSzXBZ5Bn2imIvVcU6WTOihz0Jlw7viOtoFy3NimC0Tb/FTTd
Ur41fQ0lCo3strTGW/OxrIjVHBkbJm4m84AbNcXCwXBAYUoiOXUh+gsAGJAbR58L1g+pJrHmjz75
bmngYLxqABKKukrC1q/eli3lA8fWg5YoPFX+DZP8D3GAdk5tfL/YwJCVnMiFbfJX+Dj5u6W/z9nV
9jFchg1UYW4GDT7HURvPIsxX+QaWq6uyE+wIz+u/Xf8Rt+AWm50/miO0Zj1N9tPpiihY4kH+VnAF
tYZj2ebSAQlGhVEkT+IQcGAeb3lExv8BdWRZQqmQebuuDkx+xKE3JNOIIrtGWcPNa+swlJn0qzfP
1krLZnwaC9jL9GUq80qVj+KwojjWhyUvSpvvBEvVX1V4uYYslWfOvhUMUcnaQUeAHT5B5nOW8M1p
8KVjcuVYPyV4MZcO+DqcJDTbVANkA+1iMxxnY5Hwf0wZhYJiurMMKyU5BtMZl5N4nMJpF3Si6k/7
fi3wkPeuDcD/wuZjwOVdCLC6Fjr5BsFCmk1/i/2r/t5mzqZld3osbvKftTJ/K/SAXSHaFmYzpj3X
mSrpxlCcbLzsoYP2RRpLvtHmJOO7kYoBDQ5m3e/iYjS0U6KpsCf3B8StwvvJHOHjPUiZrca7AuY9
beiH8sbSo9xxE8Axm3vMA6vnNQSqAG+PQ34TJVnkkc7gBTtKzz8ejqvXrAoj2jmY16zSaC+0mico
zSL3xHieUfuAXRjPt/FZevJYQF2roTLJHhVa+8C+kVsoWBhrDk2Lmae+4/dib2ZlpoounxQOvO+J
YkqVczTZWBJNaYLXM944FPepq/AdPvPUE6aOsxXJrwoZNQBaPrLxXZqoczzBIpKmaiE0UR9Kj6DN
C6CHvtTIC6U7sDsGNrrtI/6oQHXa9IjDElxJK3yiWtNZpJJXOwWPJsL6mq7jaTfG8wxtzNz8/J7P
Cn13R76FdzW1YJAR72vltSRE/3FXD/92eqE+fpbR7D6lkjpGtc9LWkTP8lTwM5d683Wkk78c3NW2
OXeWn62xdZLWtiMjLlzEKGZd7BjtZUrh9ZPn4kJMvbDeeLSVv0qnh5sPTJJJt/jWnULlicCJMm1c
gcjv7WzIJM4Vjb3lAVOEyzh2leFBf1P+oWV9VWiLFzgIxN/WAvT3Y1uzlJQQVEIDXg+Cb0e7yZfW
eVDH7LVm/i3idDY1WPVQXd7ZzI7/zB3IHqTotZPPzQtKQi872gCSmylcbVnJwMRFT67Dw+m31awN
p5iugikBsha5yNc5DE+W1271ZW44LPKkHp7av2Nm+XF/EeZD3VDOV0ifwhve4ZHDGcwNY1VLOOzd
+r2/B0LAmWRrrQnGWbqK0D4oQzY0Knsh72pNTApe49wjmZMcObhI2pzU0E+iQSV2P7trpJfVqsvI
MkdmegLQeuz2WY2wqJOx+G0FLFNIo8HJkseMHCEq1eSBJLp8kGYM+lgqVz1uJQzdDCIBdtQq7/5N
34kTbfoMEU5Nn/54mJ0IS9ZOKKz66ar3tEsqp3F/t5Nt2CPbsJ0SP3zMRJKqny1HtlXZZx8fvSx/
+uNzTkPeurA7TtsMyDvo7Xm9sIfQrmcEvRuwG7qWb5DXXQGx/UzRMsVayFVf5Y558staJhyeUrbv
xyV2d8i/tdjbAOcV6cE+r1f0O07JUFSQTOSPdsUCGdpbkJTpMSsLQzoTIybW6vlRw1yGkIZPy96I
u4iuP/7DOHE4jFRvozd07kPr0Wk2aNMwO4AyNFBnVzDISRm0WHcVT6yfjYOpDLoMsmeEjlpXOpzL
0e+zBkmlYnw0oqRmmYERHIW3oTJMckBaWTk7hhOvUudD/g5X2igVsjOZtm+deLosHrMATiEi6ELd
FTjdQMVlvT3YMPwqSexy8bFGixkenTnRsse2nmliR7j/Oxn2vBVUYzoAOfTunq2o2pM66s4I2yg9
ItMf4S3YHExuB3MXqo9k7RT8ry6nbk/PZza5/Y8N5YQhqkgP6dTAwstXdUZM3dzSHTO+3FiyssKa
OI5XYC3/grDUydCdWoG5GlPgZeJ5uml5oE2Xg7eV92VU7zeNKjEQJAsFNsmldAtl1mXcB+oM4x8U
jKwxBO0Ud/A0JhEsjzfE6NGCH5o7JcNxkRarQKjICdEp0k9hJYzpGdmxilASZ5Ns628Gcm0xmd3u
EXQaIchInjP2JoiVkXsvNPjJhP3Tg+TBDbYXH4kD2hjlIh3sS80XZvN4ovLbLWLUaX8OrjkI4oMK
z8TM+DKS/X+xpiQRrZHHqRWRExoikbBTbYGxUpkk9LF15/32wbfgN2mnff+UiuYC5yZ+7sKOLKCV
fW7Tk291ni80tvVBvE3oliQ9zEfr/Jhlj63chAkg16ykmhI8JeuPCZP5xxAmKCJKlHgoQeN9UI05
ysRxgxTfqjZrLjGaN2t8qMawOq9kNAfIAFpNH4N8I3f4Wo2QN1QzKCa9Z2LfvDszXJL+vThtU9Mn
QFpj1fWSlWIen6v4kq/BTbJufv1wzhWzpmPf8n7GWIdBoUJSnQI9hWKBb0y2JQBGLQtWlPCk6zGo
I0l0ycstvIxs8PNQm2t0KtdJJlC+bemgZNRywRYC8caPoiA7eoKw3R+qdToX3pmCBsndnge50JNU
hy9sMys1aL3pzaSl3Yk9TjwmoagK5IN6fGxNEFyWaJ2mi/srSuJ9YuPCQ4fC+WDumvogHiy0VVKs
mXd51O0jtjWpXlPFe46F2R3AB0JPw1wNAF7+tCFP8tILw4e/V/H6brNfJ7+5Z/CH5aDskP+gUZ7X
iBwEmiQ1ch2zCsHZYHqw6pntpn55SSMn5Msmii7dqNU7Y2UrtEK1n/kC5jG0Qw9otqhTKORQcem9
KdwXulhg8zxYVQYaChlinDSLOLP7NAPwtOGS7m8V6l72cGJl/A0dlMwYR86oMEmhywfgHSoYCFpO
4cBJF0rFIL5EdguOaDDjUP+kD4EYZi5yJAuCeIDyGAU1WKj6IhiBELOMWgzaj1/SYLFToIoGLGbx
1+isfC7oK5KWr2N5obhdzwAbg1bF6IaUapQFr592elK7ftGRdgEeQJMzDInUQcs7k+UrZzGkCOCq
l1hXaC7MOv3IWv/LO0jETvCAKPnyvxM+SSMOpLabufuDnJZRw7XHblrR/dwz/rk4rgkFcknNI4Zv
nHB5UeS9QzVSJQ1tJQX6rc56/fol4DKs8pkUcN6t2IBC1KAl2qQdGGKGSGABzwDFxrGRQy+t0bf2
lIldul048apuuNgvWzaLz2Xdkphq4RbwPDPbzqP9cH4/rWztwLKHCR/ELHxBQhhu5nhCzHprQ5JZ
KDA8Zj+pxpKc9+qk1wtYH1CjAMDelqZFtTtCT3FxeEaTf41IegE+MJFBYsIUovQ8N4m1w4HUsiDS
FWnnDcztv7v8Lh/SqTJL/PcjgA61ybAA52EtT+/kavA9mHI2PXc3v4KhejtNOTNPx++CcXBi6t+C
JWxU9/WxUizAG4gg4wsWawLwEq6WYaOBWGa1DOsAjMJwhMusjO9GHgRbz2JgN2P8PpheFq22gF6q
PYeanyYjeV9aE4RCliImGwAdvT7SZmSrRSjOr3aklaDDugtd1xby+Ztb1JikcANSgM76/rPqYkky
k0y/rDCv+Mak3SmZf6N6mcDWrQX2aLIoDc7T8k7wuXqGe4J8z039URb1BTWvE4JJBJjo6lNlvcJ0
8XZh4bH/UcPsmVFTjVTK+oF2fGGP/hK/BF117GFa5p9XISnRLnoWElgfLIYxw+VRKbN7eERBdY62
xmQaljZhqDKCamb7+X5GjjxE3klN0ByOC3gF8Wv+jTzpmVgRlpN+KAGmiIw65RX0pe3qiDuizxgJ
4PXY2zEjchObNV11EXo3lVZTDncCVicLsqEQTSRPHe+crw128fT5aunGZOqVN1zJH9H8elGIoLQf
UA/2E02KKMUmxG8vmHiI+6/t1ukcopO+J0gxwte/J4kAxEaviQPK67dv5RT7WldXaqk+LyHJJ4FD
CtjXHNNFyCtkTB9URGn4Tz6/kNMUdWM4x++5JGrAkJYxLIpmxsMxkOfSMMZx0fhAch0hqC+GUltn
/bzThNrhi7QA94glOCEd8SIhroWmZ+5647QuR3Jx+e8sBFsgQys4AxbHJRZxy9NHD/HoRNS+fH/w
9+JB94OEbCMQTwl/oJrXPYp5vCIBSKOIpqPraEojmzn7LDqW6uYU0zAgMHRbcH2e3kPHh4PFCBEN
p8B31wxZ+XfnxZcrNHWb+GuvxpJihwBWnooFtxjKEZRupHQnHzdvCtIcPosVTT3xOkHG2Ww4rYXn
Dogl36d+r86AUIeZMuZWXvU5UtWHkf+776EdFs9meZdNrczc/qjIBWbGmC+fNrzqwID/p8nboc3Q
arvtMuAb4VARgHOa4QWSZRhUnwrr6MeigWShAxmkxpYgGw8+xOxR1U4sY00piKlD2gQ+jjWnCAuc
9wDVO/MPQ5cAylXh+z7aw/AfazQGwf7oe4MpIBwNLWXmLrCV+6VYoZrimVtnuZWtHSkH1MZmoovj
wt+rpvcbscwIW2gnMuT5L9O6ze6ccu9v1WPxVtE6q1fTSHm4Nebgj8vpOtwfAXfbum9NlsBOUfr8
UBp6VFvkwkLMZD2KShlaewZvJywjktOb6O53t6Bso4LzmFNMQ88k3yqcMeREg0nWK5jusKDhE5N7
9eXgYjbdWgQvpIHy4cszetgNPZy6Ex19U3gOPxybK/Vv5y7GNyMVQtD9T9rXflavSiHGH610PDWb
eDjvwo4a9bdggYGX8pI9ZUj5NMoLn2nWxJI/YWMdG5YtATdqInoiAZ8hkhjK3EP/eujEYIvP35PU
oeboDfSHQlgi8MTyBI4tf3Kn1u4SpBlIYClnJQ2I0Aoa8UzZuIYqx0uNFYXQUNuk9Oz54kUBHSC7
nbPWavuzjaccAWiV7sj5tD3FGQqAHIDee0cWH+zAWbXqcVBWJGs7y4Wj2qcGDI4U8ffxWMtSd7Ao
+72vJKJioBFNWElPdpJNMetu7p6aWHY9iFNl5ot/qpaxZC5xB9WESr54z//lVvJVQwzA7ApC7CMk
obHmhXweKa4sMn62tiq7SEfW/0tuGndPSWlEwdHudd0+0XNG+8oMapVX3mK7IHbcAZ7LrZt9ud0I
xMIqziI1uuFQ8mbW/yTH94jGqL9RU9N4FLhRKPPFwNDva9UtPgFgd3CWA6BxMc0xirIYO/M5+JT9
Ajkz6/UluDYpnP2BpRsduzs/JrzDuS1OtUxdvJjmqkT8XSJllZeTRuKvnebTppd66lkQ2Hpl9e20
IH0ozmmyOLMpR6RhpkAb0S7hqmXgn3JLmqDK5tKht/siXTwu16DmxtBjpPRUS5hkmgMpIc/fc+S6
dH6ZcMst1uG1/3gwaigfqw==
`protect end_protected
