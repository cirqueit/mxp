`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13920)
`protect data_block
iKO7nS0ewjiROkFT60kOVlYxqbP3nHPNr2UpaqtjzmPp2l1TGOmoNyrC8877pqiKPJl7o5ac+9tX
axojgJIBth0Al+mJV+9Zp9Kb1I5aH83o2Z0yPsw5z5i5k+ILzIO19EC4fZJGt4jxZ7KcUVDlEDkx
tnI7zCowxYJUGZy3m09la56XkzzyXO9Grb+aqzZgkCv7MZ0NRC6hbkLWlnqjpgIu6/stexGVgjdc
MBkOS/xDvGp+hXvV6VfZzsGWNIWScESUUn/mdS7PkWSfQ/cnPh50MQa1+UkPBGyEExP1eGOAfoAW
PwGBPIA2B29i/btEo3NdyvdrzKfnDeinfbRoWjjcC2I+P5+NOvAIRW6Fpu8JF6EYlQZxwqtRARyX
8QDujGPvDXcYu7RZeTblq1sr35WSI42gxOdrLYENokE2qaentNDCyvptfTR5SoRgwWGqB0/xw/Cs
T3qgG+Uz1vmb+pGeTn9lPsDVJ9KGe/wKCl58KJE9L3HlWbYauz2QM7G74tchsP6QpFtKKKBadGtj
tWlYWKMfMYrQNg22/z65KE3HCoDIWGvkIK3C4bNt9gEuZYYwNXbIgRqQilF/vr0fCNm8I2gh3UVm
X+App7qZBl7qnHDUbHTGSanwnAfyjyTHcxAtE2Xbdk7qUC8W0NBLtFUTm8xBHxf5YqZqASJvHLpg
rKeqRvTL7mw3B+lTnM3fm4aphTigRC3lAbKDiNtaOQoyzN0vqabgn2iMO1hI+i2iOIPyt7GbRzrh
stsyj9RmGKXQ6Ru2lGdY1cHAvPvfSctAllcIioMVHWdXREaF7ZilnMJgvAnmxJCOb6uckp+R75QV
uE92T4k/7/uVO/BjSynTbdpt01SvS26NUaDjcFMGpwC9v+Q12bpsYvaGu8ZLTR9dmKkPD23tZR0a
SYBwQMX8o+Larch36SF3VFse0VR05Iix4pcZ1xA5s/ibnNetQTly0prmJVMlP5NsWgnYseuYefkB
hptbx+YdqgG5WxGDkHJMBFvfnWda34WHIG7pMO8GPFhz3SspU66N7H9o5Q5UxnCOx+BDNy9sRnot
sd1ll6dt616CLR33HOn40n3g1RFhID1O3S+J5kBETS6DEs5BcNR+atVZJUa+O4fRNzFcALDZvCuU
w01UKHuio+r82nx1dCSdc3n0/4tvj6E7QpmzozxfGEhYozybNCdzZ+q2p4GLeOqgEBqcoq2AWcSJ
VCgT2sSSq3ts/2OB5FH09RDgtHTX3y6kVp2g3MWyyXMMxnjXL/UV/Xy0IcFKj+ljLJ7+gqHNWhsL
CSG824xfuh8C+ne9sfECuz+zjs0WqILvuraLJde8bZ5zz6dON4KCIi0m2uLMGTwdEjM1QOn6WXtq
7rZ2fywtoXgVKX5r+uYSQftOU5ywIb02+osOKix7eaTLdFfY5QEpxriTq0ohc3t5opBMTFjNSVvu
yvyxPXH8w+oTS8tTkq/Itin2mtFPT5vSEPMELnY9DpLybuj1lluMXX7y3v80hhk988S75qHJwQD4
XP8y6haHT8wfwU+DwTT0IdOxutIEGsT3vfOdpPDPCYhHSqgnnKSqwVxJOKy+HvKHtNCiEHf0cqNR
zA2gOsQy36wFh84qgFOTaRSDPSjBj65UiZs3p441xlEKqYUHeIH14no9za95DKHuTz3MHYC02rZ9
De70fWxlEjRhAXa+llKzXsMTL/kPM1PlyJ6J0AcEilr0zBYAUMWUUkarC/0RKBXFy80npYEFZTIy
iLE570uRYtvsyV+snpWqcOTj3AMLxpwy/D1t6Sqp31reRkQFbkrxGlG9l9Tdlyq3+LTQ1gRrHm76
sv2ccbEUHzwEbe9StdeP0rkFwDKOxHz/32eF+ENX9yQ9e8aQk2cmYmWuVQYtA/bRgVtQX6hztR6K
hQTaHZiMkjSv4lH8ZdF2coeqGEu/vZvVW58b41m4LNJCNvxZ24snqa2bi6MQRRTE41WW4Nwxu9Jf
8KHOgA3aTvuTAHupE1I0i9VFlj70BqhtIou2dIljuOMvCjA+BXzt9Kf0qbnbMgn13C3etS9Uwaja
HFzG9bDA3j/TQvYPFUdZgsCUVOrS/5A51LzvZHEPSF3jWlA2zrxKJNZWm1dEK0L21C1wT08qB98t
eKpThV2EmV2s5p6rqswkhSASkzpEsdlGpknVrDpUdZD/zqE+JKcQSkvzMVMyCtuNl1DPElFz8NP/
2JeSwMAHT277yu+5AZh56SqFLJVvLw73ojw64bq753t5yPTUWFuisOdoTyUz8E6j9G8Z6r+axHpw
CGTDp/RFFQXOWzdvBJQDBDBLRYay/QkiKX61QT+R4NvS2YzMgb9f6HtiT/Mm4x/gLYkM4ZycF21v
K3vEo2oC71V+88HJ77LNb/ayfmPJRM39h1PtHmJt14WX1HgCUhsjo/ZbZ/XjasyzsZrTLW8watHu
9y1CEo3hBC5Af4lEW0K0RwOuuyPGQdj5qic6B0RGFrWs6aFebYULcEpbLmdg5kJcUrdOeRcfIX27
OGHo1fiiNSBSkt/LVVWvBqw9OEL0rPbuCpMM9F3XrzDCHzfMaupLGIcDZF+3m/KA0RbWWwyvPMiY
71yFDu7PfXC6JS0QgE+jE1zXvidgPVakc0nhrLz6luifkrApL4tg2/wlRHNHr76RBsjSTMdzdkeE
QL2Bum7q2bmle/QezzKBtfgMOYS8bK03DsYgZ5Ybt06JtY5ibadIVVU1EuNYdcll6OopbRCBayW4
bJ+XHPle8KCoUUdhG2V3kLwWVRrWwfZjBKCW+bNeExAqlcK3kWcQkuIiIewukn++cGH9aX2t6hog
XcPe7/+3bfHdYUwMmvisy62O7wo/RFfA3rvSBzUi0WchUzh40L6ujLL3AfgTMU0whGDQASQ3tCHV
YZKKQaR6yNgjREiLOBmw6pfpjkBoxkKSecym+wKmunMDW9hALajYd9jRqKXYMlSOzyw6owabUT+Q
KB3QMjIHqQZ7Yr9cWt7KXn/NS2MDJWk8G0JcbSQFVC5NPNT1nIfo97LOdXB+791I9Zr/cXkIpyK5
rJh9IsW06+Su5/7FoUBmgnI6ICwGX96alitE4eje7rsq4vUcfViBDGaHF2eYVOk3DpWL+TdLkBx3
2f7974GkJ4mZNyL9kBGfQCpW0KVU9cHI7Z51y6ulNgGSWCS0K4hBZdiFMMacpVfLBwuydXEvX6kQ
TffCeef/xCMCWh3rh6Tt13FWx2m157CJ48BZjgxzDnrNB8u/lLDSsCk2Rbxxgc7DJF4ePa82Iu4/
r2RU5q1WTnU9mmhf4GEV1zs/1CcFmqrWSfElIkTXCTcZPlWlVOm8r7QUSLEMZNmsqKhkxeoC9Qk8
8pTFdKc4j9YozIfBaIB7E1FH7trX3LTEqDV/rQ17DDY4SrkuxT2wfspiNMy3PD0nBPS6VNqjIoMz
BKUxYsH8onSpW8mYE0pjatkqiI3Vkzfadh2/g6RHenvjXkutkfX7zZFO0nu0Db/06nnocU05LfkS
GghiQMczCFMRYYebONjADMVjvqID9kmHDbO1+YuFCudNIvN26wvUtzZ7m0/gW+KSc9LP0kIb0PM1
GUi4jn1qivR/fWymGhv08UVXzr6T5g17O/881yPR1CSx9oUsv5kuKdLBKQi9goYibYgQ+SAIz1jc
gZxzhqQKevdBuJNyn84rABuLJjmRmnPIXNnw5nZL5qgbvRjl8rr1P71imbfo9eJCL1PxgS2FebDj
Rcg3knZr3qX1+xbTVbFHp4wWPCK1KmbcILJHScsTx3leHs9acsXuJSNSkwEVue5KRH15pO02K39T
ifU7bMqjAIFqGMKiiMuE4yF5Ulz07Wi/f3Z34otzLcjy3wFVDC6hELKc51/bXviRHsXMcIQHu++M
uwzZ6NMbMlgXt4sOcKH3qHgMb1EKsOdnkXzofhPYGFxrk7ifsDYXnK46jBScIezxluRJ2Orb8T6S
mxpJQvi3Sgbvsrl6uf1yJRokhAfdCpAPJ7Lp57JYliOewC8lyXJvxEZ9LkNfo9NcQEbhs0RRTCC4
q5zD2RD1j78us2N8+8anmcY4B2L8LwSLIBBPYrBhHqT8/7sK7cubSTfYHqlj8hG03X8zHvO7s4kz
nb/wfygwH9PvThXeAfGH7DcB5nxJfH5XXYlXtrxFtRWHeja6k906oROom3DIvdn4RQm4TE1xw9P3
CMUhKjAWTF/ZBRW9IRY5FImnUWOEKfgz6YCCN5aHe1GXsl0HtLZFr5FQRqK7b7gRzLVywe5S1i/+
ZTGYPta/rRi8MbUi9RwHwARs1fQlNgXNr2Sbgq2j9hxatA6xI65viJ28yvjeevoynj6hDp9vnOFx
pFWTwhkDQQwIWY27Ct0aCOJIDrExSI7G90SAynRqc6Df+aXw2UIw3bdtxV8YOpFebF70qjSKeajv
fkryMIPwzIAVxIhtkkOqFXiuRd7Yea5Hn4nZo248BVQgi1yRFFNFT9Ku+J0SjV7rfVr5IOw2N+y2
4TsfK9r4cHD+0/3bT1xuqHK1vcXWHNNgFiSnmdobEH7zIPG/qacOPBw8V6OCfl2BM+o0QDZzKjTZ
6JkAEbjx7ETxxnrkn+lQCXBkyTwCKJVfoNsqG/zKgO9ykvVexQJiMjETjuX2FN7B/XOPBBgZCHlE
DEXII8T/3USd06h072UZB447S1klu6P3YivaIo/OrCrfFnKdKYWMBb3L6BSLacS35a23wI6MVtg2
c6eVNt2ocoKCtAkRBA+wvkM9WK5qPj0hxzY0BA80mxAb6uou8XsnmNW3kyRbNlQhEHE+6cyu4vnB
GVr7XGoKMKzHstEpFAc3ubqdUJAJa8q0xFJ9ErQwYqBqJKAGUWY3jGckD00fn8ykP+8s+RRIpmEn
96b3uims34qHn8xyyNhP9e7fo25+gbBCMohxD7ya/zCgQersxSFOajVhq5Wj1LWpScHKzjM+QNMJ
gLbb8yQLcwG1Rgwcwy7nZBpDMJ7/LMqzFOUKAGBHiAYjxmb9MWs0H4D5ykgzT3ZHWHoxsUKQtzKR
RRF2dG8cJztv2nAKtOrZaEXqKErcFpHanGebvR2w+PIODVtHPk3/59YOyUSaKP7s29oVGZQDEoaX
PZM8t7xOe0zy2IalDr2M8DLeyVfuVCYyyMqK8IZQJEPS+xQCOfgDvtWpRSXhy0DY7BdkoRB+Quy+
b4KpWTfya/zRxml7ZxtOK6AAt2p0sSPAJ8pp3eAw7iz1QthVYhcwydTta+f+jUwsXFLVDHHG4JsE
O42eUJCyQHDWY4BKP8+yduCICKOwcFhNZmYexBZjiA3p0jEoeu2Gpasa90n/5P8DuLyW/cj5QxiD
cKFFbSfGbA1mjJR4dY3dtUNczzrjP5KBmU1f6z7iF4ySYD4L6fwuiwSn4TW92q3cm6lTjwiMNfus
SaVSaFHiWHq1SfD3bkGJmRIUy21X1X4tv7L5N01E6+qDRGIVX2PHh1RksjPp2qRcp4rz267/7CJc
pQ7vl1Er1PdNRJ8mXAr09D7gUQEq1v+UgeELkCFILKF/klqUwQdtopZEmODQEbh1+dwiHKFCVzJq
9jWIVLifc5WYvpaxxe0Hb2zuAVHFiRRk4Xz5OJ+0+f+AuWcpVcSsCgTRcw8ApxriVswn32KUyFlV
9SEKIoxdTQhHyJLhZr3BwAOAGvgyFS0lVjAZXiu5x5umb1d9Ttym6CX74PEWaQPwrX5r4enDiokr
FnLm5biqBGWLGPQvDSpPyEzxqGCHTYEa1QAxrHOaAcJGrHkqLN06TtiSbm01Dm3JO2JQ0yNOI9WO
PNsO+U5owfLgdnwfVa6pjRtkoES3NpQP7F/GX8pJbEbQ2PzAZ20UtX+yQEcfedH4rdom7KoJMht4
QkHErtrTJHUaROOc9t21hFqUYkzgUMCggQ5U8InVxz5gT9zPiVBOQfuB52YuPRxCVgxMw4fGRUEN
d5u0EmyFnk+LvkmLYEcpAns3ros2ShxZG8ogcJYfrIj6tQMonTGLEgXxpyJ03M5GSzhqJcvMWqOm
q6OzGQmnuXnUs7XpOUw3QVynf/XywTnJVfzyk1xbWn049OTXJlAAHGgxcLL+VgOmSvSfomHeigQI
9FGC5ORywKPrx9ZBtoLOj+J3C68D5vmS5a1s8J0qKNWOuvHSNDj4awodSO2mIJFl69NfJ+pWMKzn
YR2Z3h7ujeI6GhJqamQDkm8xN6mWKu8oL9zyb9RQTzLfc7h56cmPib45p9WpiY6a5xFvlU859W2N
pLCklZa18oKwhPx2JU4aGgCBWjJJ1K/ge+AdYzcu3FHlTeG1gY+umcbtz6bEMLgsdTY8DnoskJq0
RhRI+8Tp2woGB7FlY7SWJmFwZAnrVFU9SDzQymQMmHovpsQ+RArMPYa3hKaYRgaeMKb4bVZB/Gms
rgLmSVufoy6BFFmJS+YSUYe0m6suQ0DEknN5Cef7Ov3KUevlLi77T4C0TQYfSTBcq8Tf20vkliXK
0IWFNVU2Vb7ag2nHqEcOa2VRHAYg2OVV1jN222stJ1txNTAKO8B/xawz/BzLVbxtr5flm/3dzmyZ
WmisCA+0F+s9xS+gGmSdETg/pCWTTPExyzvjc7RHG+965HmDq39AmszqSsatq2gngDoBo3qz6N3E
XFeV/MEEfYAp+1Zaebufgsj+QnQ0uuOfrhvZ5uLBQCF4pa00/vlxDLReg9qWCfcySWYin7H3wQ4i
3bxb4rhmhwk/SMO6hvgXfukMJuWMGn4xFoDY9E7Icu1XEUn+UgVs3co5mVfFBeF52EeTvJxVK6Zb
cQOA6CvHmtaYHdBOJO1xXYdX0xZ+rWP0e+RlsCebj591/IrcuoymbB3b6Jnu6JfpjEdF10e+vCq0
+M0xjA4Mw4cT/yEqlN39HGUGHdcp9Hv+TEXFpB/vQm70FJFaexH77Z1TRVGeCeCERgUu4PHM6MIk
DxLdSPZDOW77cek7IaQnNpSvLtgLhRtIRK820wt2hmA8X+qimWVwhMRJ5LcFakY0AGkd0ZJKu2CO
uhXTeRY0pxBRuhdJiwyQgPvKVK/T/5bwmhAfiq3JQoyRDaRZ5TO62mXe2ZPv518+jUgNFSCdaRQr
tw0OKpUTC546c244KNOfdUy4vI+TQcxNj99UAt0eycQo10WSWdddgSlWdI82ZVw3Xug6YCK+xFM6
tWqAgDIajmYnTXtG1RGwe/jdTLVOKr7ZVtEUmmthxhrGjIDfFXqi2u1nXjjyzefoAB81cp/YTKFC
zjbrJSypGXnXInhZyi37Dm0aFbkHHxDynqFvCGgJ7sVx6/DI1sW2qq1esIpbQ1qnbH7R/+u+bR4c
COmAIIO/jQ/9b8mGxlIkZ7e8k8kBWRP8Lu2/EkDVJHH1yfogBuDtbtdimgG+Hqt0uAvPK2V77wH3
3pKweIC0UEKsohxcjtbNq87jnbUP/sL1o4m6+hIyHIfdLQSN937TDGc5ucUz/v5MMECrIBKoG0IZ
vN+wZEfp2rDo4XysMLEB/wEGT2l6UFPLjVCaNrw2P0ayq8l1AEg5FD+48Y5lS+h6he09mQ1Xwkx2
ZVY0b7vszCjZ8AYm2eZykzX3RleT1huZy/fPFTX6s227BZQ123s2Obmw9aZYMcB9/priybvWxjmF
cm6khFlFGBXYlVjp4R4uig88aDNiZIg7euM50uN3E5Enaa7zfbHRdyzs4l6ISaFs4SD5BbzhFzQc
3C1Ph0rhTOZ1OhL3pX/U9o1tzLO6T+Bo2mihfgj/tovApqjctQo1pX1l26pKbXeDmjXzzacN/OC6
PhOzChxCXGX/Eg3W5HTTcUA8w+QzeG8PKwB/yKZMZeUBIv4XPGUUxglrE6A4qTv1FtJjt+32kDT/
QM+/4SeKngAHfMsO3dQEiooP91hk9QNnx9B5eH7rl0VaK+87vPrwoYWhUJtbD/80ybbtIQCSf95X
MHH6rd+bV7HDICth1wWrJDl666hhHYg7bcfuAruIc8J3UDY9nVupoV5uJ2UkkxabkG2M6WnRwWpv
gNwqnUeO4TPpcyz9aJDCAbL7Tsde1tgTNQ2alcFpDt8AFMNfahKcll/0P077+b5hltbmfIhHP1ot
E4D6TrB2aq3QGBGrnZvQEJQ/cNZ8bYUNyxGqXL8q2HjIT9JdObEsviiASXOQcqfxI51sVjHf2Wgr
5hZ7iooul6/WYASOixrzbjXYRTGo/zIHT3k2ZPpMXEyhhyFiu3T5oCuROGsJRruUGhZb0+1mR4WM
izlVbYFa+iPCZPaVp1QeXUU+3DffeBwp/leKW/gLWVPg9N7llt5MDzwcWCCSr37vs/eiyfH9sCAT
R5Ub4s+DBHt93xwg9NVZprwtU1bxhvyyG8g1Y6UScmv1jJY1WqeZY4ibbKKDUg1HWYuozZ78Qgsy
XFlcMvQBX6WstISuZk28nadRwWDwNcKhnCqI++jIfXv9b9EfP2VKtV79FDXDr89vgKUZTVZN8WH6
+7wKP7VHhjDbt0m7+PtwOXxZyf3fURPiqch6/mUyOPtFNkbG3jrUJ6Dp04U4ml9M/ZVj/wgFks/+
ZE/mrGmdW2pBuBNueFtj0AdC9xDo6w7FBlOlNp/FkTkzC0ilIMDHsJC1n8sSP4o3EhKvZ8faIhJI
nY3kw1ZMPvdXxSbGTc28eaOuZAxTSS65irlaOzgi3sRN5pz7ItQZSyW5ft0WXU4j7JRZf0P4sk37
kx3YjAoqswDDS3K2qZDXNqmpps/R7pfKSSLU4FWtaIN3GuLYApvBLByvBuWYYLuOgOcxo9iLD2mi
QTeo5ndPasXHpYvMvZlmzzAUf91389698gvAmHUP+XAO+mi+Vn1Mqp2yWsWsMotF/niIrYxGmLd9
J5EOn1r0vEUeWRL33ufcajhybp7V4WTPxveaM5/ls2zPzJ7hUz+mF9izUjMjuGDWFW4eBGZlwrUW
HLdV1Khwdt+Q/zHD7Kk4B/G+f8q1rUp9Gq3ALDKuHew64qDSTDgO9TEC3KOtG2aqIVtmidHVywC0
oPwKIsMfbnGNplTKQk0Q/0grD4EkU/5ExStDcMVUUoOcDb4xboRCqwzSEtMI8bkTRBuVgznQs9r8
Rsf2cUMJ4ChdpVnWzqpscz3k6W0cYV5gf/m+a/TmLQy+fmdTB5KGNBCegEc1Udg2aOXDz5eSwHM/
xAQhXM0Q832ZZaVjm2IbadNOfA9OxlMna2QdKhdtB9SF/IqhZkbOp4cY9ACAOZ1n9Lz+BiahM+U0
R6C2vVNQNi2i51uPnZZt2Bt6UBrjYpcplmRicAr8h5uXBTPTq0vnBrfBHMnEo1Rkx+ZsPbPbjvp5
ii3Ujxq5j19cOnjve8/nqXsisPvWl+44rjHg+Lb/ZKT4FwfLw1n7lYqKpMzW6wX5/iehWgo6ACZj
dwImLblDbso5OqcunKU6DVjgC/E2pT587is2JShL3JAIWRnf77C6NwxlOqX2xk6CBpeeojl7QcCm
y3UQsKjZ5s+Ne759xGe9gLTEgQGzZnpoOx0WDKN7M+1dDhHgrJbtT+S05ufi82FFJ9w2vtHHX4u7
Dj8OUTJ+HApDrhaaDhgC7CTH+MPe8WPSLE73BhJzxI31rLK/9Fl+Pz8MjXTLYE12tJuwy01xzBui
nN+HMjmm9TAyAm0Xpfu1lejwqspScsBTztAX3osgFbEtQTiBOYa3IQomauyLdCuKStsJoYmoBU0s
MLBItb3CtbaKnpI1v+EeM7S+D9KCdB1IuUYSFWj4BAKJLkzdpRlF6E81HUh7fA6iRjl86L9EJU1V
cufQ83kLFNasgZi1uwPPVKF3Q1YC3cud/ZbKpcwEl8s4WPNoV2BlV0f8hCOYK68z9UhLiWEZyLBN
GIOHMDxsBlvjpVpehE2Q1kN442cWK8b3yB07rDUnvgk3tpE7YjEI5snxsiIjD2f0Kul7+zeEIuxw
Ls+K/xn5hRbiQEdgs5fdU1j0amJIftFyUcJ2m9K1CTPmCULYBTnShNXV3iRSL70GmKTMqXF248hc
6iP1hlwi8J52kQ5FImohoxjQX9JoWceFgnZFWQ/kzpuoipmj1bUiZqbMLDmjefCkGqR0DRbV7A/X
VwyZAnSTPysQvF5+wqsPGDFutJfQq6uaxBR1bBynTkIg2RNqEpJsw5F+FnXS1CCp0inYN+EjTeYH
ksfrdMs4RYXFoz7XlM91B5kFN/bsRg69kAkFef/RxGJF57RlI9gM3fktamgLSLLf+/2c+fqHOTmX
m+vJIbUZjdqVEedR+zIbxjRe5y2wn/qfJt3/jhhNu1QvY8sHkLQ8HyNd6PTUVvde54NPMbGVnVcT
pdbs55y8fmHXRsJhTnLkqqsN8cvMxAP66WW5FWMIGGdqInWZaFKFszps55j32kHPqTaabCm6xpsw
ZpqhkOWNAWlR9VnrAYnBCwpP4H3jTvS5X/d9CPyKy+Eb8Dw1opywRVGvyjrIacZiXlmYpSjmmOc7
SQGvz9ce2umBmQmgCqqSeKHYcV5pLouvK9nS3iMQvSowBLe5+0In3Uz3FzONDfK4RmRkwSYsqQSg
+XPzYCeEUb86Taa3VyTVbvCi46KhENiUDU+FALMM4dgp8FG8HF9Bnn4XT65pclk+TxxIy0mEK3bg
IgeDIiM1BjhTbSzSc2X6KqeBetnJbfuY/Q5G97TUIYyWENY0JFdF5UC706SF7OjC1/MZv48Libp6
NGCSDdCrBOJTK20HYne5381H69m6YG3Y0rq1bAfFGrHDS9kEY2zZGcJ+2ACGxiLKXRkBfXNiqDR1
+G9VfImehjk6FuJTqnpG+f27vRSVcCOMstN2nLyq4PVRwH70yLkBzdsILEeIs0bZpwRn5gwjYeFn
s7fUmGoDzbMWPAd/UH8Ucdpy9FZ3hPCoiH/srIS/OeaUashPyVk/YzJK6tx3m4xrQL+QZWzfGqLF
qZt+SUkviRgIgIMgr1f644vD+grcoTAgesdZK3BE/iKGiyWYVPiE15WcwU6+qDwOyQAYiPIxgLmr
QN0N0Y5+GInJ0KOXj+Tslp88tgufPghAImV25algupZWgVQSr4BFUyeKLfasPLH9r/xkR80bWwO+
XfSkTT/okYJrGJ+ymE9oNlDPtCa13rG2mqHJ3IL1KRuCiCSPPE2RXsMT5x/6I6o56nIMkktwoRtj
sfmJqB2U9pgCYJFIsjJ8QhoxI0BeNaT8ub2ZBJL5MZdjs/yiTL/KDOAG2gXxOCl1djyOFT9cRp7a
i2C83vLK1VfJ6gwHZGVzXZFEd+eWXzW4OOTddi8sB6rSxgZtl98JFsac8DdRgTEBhnDFVFBQfCz6
NEdUL781o6vSVGXDj+DsD/fEwIpOUkthMNuyQNsMV8hLTscxYAD9in4HvThMaD8iCzhqvreIZKEp
E4mcaVmD625ksp4F+Mk0rXeUwEE9t4xZWgqROOQnLk2q5vlDM1IEQFPje6FUh+1VwFdufdBm5n1o
1Vd+Ht9+a8xfSSb5KPQO7XVSLnITwCtU712hyExj1Kxqu9Zk2hAGmxEOi8nHugbPLjNN0yGLSQ6N
XmVkioKHVK5UB20yxs/EYRgj5BQhehgtgPATd2TqQqd/ITw2okx053wg+PqnHcGaY4WvkaB+JVN9
zqg/lelQjl+MP0q09N3WPwiUI5KYNcancwOEVVu20Oc5bTuH7QtJfJ8YrskaztSSVvRdBc4mWBe4
Nzvz7Inv1tsnmKiNQ27c0ITjBBEgc9op9v2aIO4GfkEGyn67gocpo/UQfNfSS+701GnVRd8CU0jN
oDwvb5AJ0es3yj0HDrjaLAKD+FwjgT+tZRyFud38rKAjFcxDjJp2Jz+cXgvvDjc0+MKesyYjHT7w
zm+/g2OtFx4lm3gw0Ox/YCBKRDXkjM2ePZtRm+FY31WGx+WLp0Hgs+5PHgjOKt81jg+KMk31CLNA
UcgAA2UyPkgh/s31MEoKnCvEI8+DHjlPyI5BNdQ5ENL/3RLOY2t9ZBNe/J3zSNI9tw7hcT0mddL5
MDea1xSUGTTmCa7lfdVvFNn5masDwvpEj5T9zTm54wWADzbGIWEDOTfNZwxdMfATBLNOYZcZEk2j
Vr92S7K8QWSJf4YEbL1/d1WtzMPv3iOCuIzoLweuPdT1h/RyGUl6fdBZGpWFwGKQ6gRrirgBP+vQ
NwhODmLumElkbLjmxaRHJ0Jdslh3UOm+2CvbBZreXYrN/ObCUrtyqsDOJo+tVSau6Cr9TBkr88X2
2wSp8CG7Mko1Bz/+bUdOwBKWdXHdoMx7lwm+ME/CGZskxDhhRjgAINkI5EefOyMnl0+vXAOJHJuz
vt4ajha67lcihC670ByufeYq948Ncvh0oAbwNvnCCvIct7yhGlczowOkwT+cpqF5VOHsfeEY+HaM
IzY2D3alXJVI/TNgOMvD5xD1NafkRYJxOp2o60ConMFj/6vll6KyXMtEN2R7zrhyCq/pscxke2XM
I7MjyxVyeM1QYl3JO+cZmJH6UelKe+pN6v+gFgjdhexaZrs0vuGjxD52O9fjhRK/aR32MUuNQyVp
ItpX321MUtZGkSvJs1aohJeQMbfcN1PqE/+W2lcSPXco4OiKvuKMipdibh+JU0Y/+XE4QK23SNmb
pR3aEaPkQNak0hVakfUG2wL8uVR5ks7KKD441tG5otv8Gtt0FebsU9y74P/jIUERl60MaLZA88wx
QTTzryZ9CIS+ss78YLZEYssN5pOiDjImnj7kYnBHz55kH0WGRa06HVo4iLslifumN6j//ac/Ys/C
OOsHtRBmaEg+isApzQi2gaV5bEata8NpRJ35gZ7Si/MOr+im80LJ0lYwmbKuIN36qsSa4j8PKG9u
u5h7KmsTzR+GY4MENuu8WeUa19prtmvEuIB7SnYsr0UwBQpSsXVvMp5FrUMMQwfNLSKdrlBHEtIz
8mViGSql8oFNWIiwSS/0OwZhbnaRB/P6uyr3UyaM61IfVaKcfFXLg2jup4BtLPZjdRHjBrG7ySAT
nVNmmgbLluwn9RP7+JsCnQlaw0tIk2fZYzB0LrSechVLzdxBdfVa47qGBEoREyfAYEnHboR5lENt
xZM8JhJXP/tJEAC08h3jziknWgB/SvZmEmcEHKNS1dNLucT1mndrSbSeYSey82D28CkHgnDw2Aab
+irgcXzfB4pJXz402vQ9zoSp3P/nepdUJxiwMUKbwW4jzfociYYOLLDHWbZFlWnT17cbyR124K93
N/vEHynMsVNjuh5F3+c3PsHz2Rw0Mxryf1hmu8+5webHvaoX2Ud6QXDlbyyF6RsDvVz7qKTEvyFV
BVV+NZm/WXzUHaQJUpsFxt80xUbZ4irjjwNuxGAVKxTA4gZgX0+r+zv5Kz7d8n8gNhUNsoSqfvsl
T9n9K1NNGUK9QZS687cS5iEdq39yriJoHbO1sBnmVAT/tvVIS1/cwOq83sfV+yybuRkMvkJZKpJL
j2eKrjFaNc0VJUctCF+Z50wAwFCOJt6+m7h5c+TFqAM+xXU8ysFM0xBhN12b6pPEMM0H/nIDpg+f
LsKz3CafsDXd60ljkOyEHAz48nCFmZrES37esknlnG/mfGwUuPq9j3kSguGTpdPjqh5qJE+EXVXA
hgPUdBPk1eq9hxqjSRENuRylwpnGM+gcv+BR8vyFSULg9EmXe1aiGdpAVcYKdxMgk1Zif80SeCOT
TaLF/uEJVwA4oI6mpRIUpCKGn2yqLWLVPzWAHGp7reXOrZ3cjJz8IFZCfZEk3i/mqvJLN5jkmWac
XgQybv24TbH3I7j3TDCOStNaIM43GN6WGi2mlAQlL/Rvi4PwvcABFSV7CzRsKlH203doXqs3dvey
zV7jaHRg8708MWKMlwsrmETsYM+z6PTCTB+5He14JMRkaATMq3jdoKY2bDLJo7TwkdIze3aqiCGC
fuv+YxCuVYizZMo4QVSDTYtEnjJHiGuwEnYYgbz9G2zdFKbXQEnsOXh687eUL0LhqJEZwlHBR5TY
FHhE1g4Pj66J1nSL6RRFRo0ObzcWtr+AdSOYxGIQJYJrWA1KqLoK9FvY1ST9YbYTcCliWCD8OzgP
aPTYLffYLqwJZuVmHgXHJCOUCwbd92F4fwHRsDXVVS5be3N84z1QLNaOBVfO2Dq418vuDSCwC+WD
WXBdJCdMttVL0y6MsHdnji/Q+XWIQL0XIu4c5+Fb77RJ+kffuPqbrk09id0J8ugvwg6Y9UIr+B0R
MAGgOF8YyiZ5AcH3TK5z3GVih5eNaaVtMGH6Z1guZTy4Om10Xp/o/63eHto8MvHB30SjER0C5Y0/
Smxzb1whVfM7uXssHtEywBMCxnI1PoABend/QsL5wSOCMcwSa9oKF+dHImWJs4Ms5MUxxCqADifL
FUjPIeB5cXaicvRK6ZeMLRV1GxyjRf2+/77rypl4M4D8pMzmELzPRk1sjAiHJKeGdW40oPtUwC0o
2LXx1CZEsZh1s1kl15rmKCvtD5SIhS1gAiFl1y+mnrvgMfihmzZIQfYD/EX3z1HG96uM9Cqnr6ks
dGNRQNVuJlh/0rg8S3iDf7B39xoHJAv0808f1GynEPZj7gyIGRxW3lU7GSbTlSEYYLBjhT0DzhSs
xFs8v8zH+VR3nhH7xQd1kYw3GAhRku85dsiszXDMbSgGVePcxS553UtOwKTPH5ZsMc9UWZL/h+yq
IeWpnDVgVMyLqGl0Y4jYnrV/rFutvZYaUpX7YohqfMEqfPMAKg8d22x/sWkKJL0ef4UTGRhnqJdp
mPatynPHwWrv3prkwmSpGuh7w9dWIBBl1qlZAe1a6wxajZRWHFNbpfUz4/W2Z4c0MzJOPhzrfHEO
mNZIN3p1j+QFfsdwPrkS8tTM/3OKNVw1yim/kVF3nRxb6reZ4MVBRLk7yINdij2t2+Drly1+8Ouu
20FrQ99274Q6T/cBhi/R9aHa21wU9rsWHq+sC67vLevc+bRMzZqiyotW7Spkq4gVaf4fPtTd7lP7
sL7BW2CBwi6VRYMflhCeSMMA60vHv4V4n5cKwp9Ybvl+7oUkrIklniWOwS6v4pLr4Dd9tRCzFWjN
xAeoBbkZOr7r/NAFS0PC1tdEIqBtI37npOI9yjDWxickyQzPUsrcCsIGBhayO5ap0vFl7JZ3F1fo
tvzMSF+2Vpa+dNg6aIiE7iRa4Y8ZvXmkpDNqd/IPfb+uHn4+k+jCybaB1o/fl3wBG3uye+vwiZAe
AbRPnAsoHrR1u7Khi2o+8A0M3zhL1W9q4HuvqXDHjJvkAv/297MehcRFZwiNFuvyUZpZl3rno75A
onmywr3YJM3JMj3ZXZ/3paqWmMojfIKlzqHNzjAje/dDJahCM08WU2oIjT6T+VMnmY7ZgYaENhWx
N186biLiEDO38Eh/zSQt38J98Vk/tAFUxx2lfrxhzQr/6G9PTUzXpqrd91sYEZ8E3X6HcmyooIBg
/GFitA7vgCzZt8/dNES1//fyHIYTNW01BVPptdXSYt0YyjASrod7q57YO355PxdjA/ZwyboGQxMg
iCRezFeW1BdaQeSS1Z1f5RYwnKQlCdoTTBf0LLyjRVcm7gKF+fQ2VCSoKKNwgq7tVjv0rtSUajyr
laWszFgO0EdDiFchs//w91CuyKod9gp3U0HWoSKd5eWvnuZbyCXbJ8KO3bBEx+bU6FVIxqcZp82i
u2Zl8aIDghU3V923Ui8EuGn/j7RsiSDyJsQoEzDaPaz1Ks9Z0s5Jsgz5oZJxTrO/Hx26FM+8B3m8
SuiVMmiEqCNC0A2zeUaW4QBkL0zA3eNAdTgq3cHLaJXkbrBjMeJDy78KVNCc3gR4svrjrqKgv1jJ
PRy0AUhHQ7WG7qFXQTOWUWr9DBgpzBVb9fb79jsQ2UWmtA2kiRqsHHi80k58qwEHyGbeOumFOqgj
vjFkOgcBcWvWHB6ApDeaDl4FAiYmbzsQ7si4tyPh2gXKbnLz+C0yuGvzV1aIdmA7LuQqmvzPLafz
tKJfVudKjYvY+UinViKdbfnLUvGc0pGwLZkUPXaDBK6GYyYtosAI0XyTKQEDgJrG5q6xC1mnzdbC
q0VIY4CE1arZwWLCPvmb5HItoZK0eNgU/FrI2sh+icCQ40RER4ym4b2IB48jmUc0t6+4YZskvx3L
me1G5M02ynAlrQ4Y35bgCEgZd9Hf7+kQjJ/bR5TU2dFjGHVkYivwtVmTa4b2gGZp081V6YzcXNx1
B6Q8eVJfAckZAUye2qNafhJsGNqX2jYMAe02Gde+EFs8Z0Fuv7OjP+UFIeqrk7PFkXl712F70DXI
gnCM1eA9+4atdO3AwuXglYlTpVkNYcqhUb3oLIsAvrvtulSgzqK2wdPc1o+y0I34Yltis2eu9SI3
EyG3xqhm5Zhp2w9xEtY0XdfE1bcnAYHNkfRlng+AZqaF0cBbEJyHdi5F+oDd5u1T55rMTmbNSkwj
e6OcqYrsYaULm4TrD+hz6l2MXPw1Lu8sROioB+65dxP8mdePVylsJxT3L+CN/v8yhY2l7nMKXy7c
3ouVkw6pXLlGnWC1rgu1d++3KSi+NrVib92QcHDnMsMIjBL7kQ4xdK2tZ5QDAy/5zY87L409iUc3
ete0iXK6bISX4bgOybCw3NaJHEoM1oJgMfangSn2MAE+vTYwbJpgkK3KoHytjMhMwr5fiw27iZAZ
KebCl+NV0QjazEuYjv4iA5DA6b8tLeAn7R7g4oFss1iTAxWZvDWFeToz78zuJZ2wv5n+k5VM17zw
W0LXZLeKZi+iJvUy9aHhxOQlbIpnETxgV9djBywDVnrOX5kP42XRndHQ4xAcjzHQM7KrM8YRuL0p
IcX4C11mtdDdlsiZr+2sE85U6BwhlOuI8Fm7av7b81r3iBz+ltOWDSMAOf/teJhswk7UyETkWTh6
H8q1Dp2+Ym73P4JbBSrODSL+RBE7Ujz90BqlUJH/dvdqeW6/dyNVqysdg6kgonkjmwXfL3sbbpFm
UgWzhctcnxV2gAk8CzCnmj+RDlw0EN2QmPqgavVa4AJ0FijVAp9/aXzYCUdwkxPuR1DEN5OcGQn/
rv4PJNNlM71xYwt/jK6aLP/OciUbG+b028K5SDDdU9Q6N9tPqmGBTaOsbLwkug9rE2f0xA9B+x1x
lLZHqVLZunncxCkAxjlyTr1FHu1+JjeysnEuOyMlA1jymMEv/UcSJYq6x/lJO5e45c94cCaXW27L
6nik0iMwOSW7HnGa/2aQgMyyQf6v3m75OuCfK78UM5r3F45LgUgANnhkthi0tkuwmu0IKO8J0Ima
Jt8xu4W1WTIuxSFEFW0j/NUmhixjk2hO7r3AbuAbnuKnbstinLExrf8rHE99gPLzYEfLr3TWjRiP
CKYCYrO94na8wheXXy/9GldonXYjgsRNzLnKwNSCvYkBZwB9ccc6cTcDog6ANEBTbVB67PpCxSUS
IlQqHiW5mnykI4S3IiADcCw2Ga5ZITF/nk3JZhGc1H4c9fn+oOjdlSr5DYuIowv27G03it1ImeKW
xjDpKn6zs06DJBAFhtmrbbGyAjXvFgqT+QhDc/4kqFRnzxcARQc7DA+LU9BJV/fxXfQTwGw31bf0
UvYNCydAejkXvRGBo0YducPGwUA2kXEYKARJuOEGcgQhB8Mrrhh5PZoxZZjWt1jiWDq33QrYBxL8
9NjW2rS6/Jz4PjDUtQcx/oG+kBPJAZ7byE+3/QegGB7mr9yy1lUCGbJJkHnISni8r179DUJmkN9j
KMnu2p73QdVrAIGmWRFErulCJVLDaMg0Zb309tpTrI/Q7GlWcBW07mao1VXAq4UjSXkWRX6M//+d
uzLkOLNdkkdDwPMxiT0ThVr3qbF1xSB2ClqChTQeENf1ztR0QPviK7FHtVYPV0H8boIEJIsh/hV7
I7nkCNHdyHioNFJ83jfV12M1BXO2PDuQrWjPEIBQeAVkCSauwCDJLqQwtejwF3p9r/7e7G5dHrG6
LuaEkaZKkkdqCp1L1WF2cMYe4YfP2PJADh4y83S6wMdrWa02121lOjN5ILyW4Lczy7oHzZ+WnExW
aq2ZrHoHw6nHjXaAq7wo/19690eIN6VQYk/iYM4syAO2vTKzniGblDZauQMlKLawS1TWbHV2Lqk5
hp+wb2rDMbJUZXMs6/9QknONcpCfZOgZ5wuEgybNohhZUHFBid7Zd/BepXAw+DSTU3adTCqsdXm8
93S8aGV/X06Auh39B4WmDTOWpHsJfv7Z8LGXtAc8oemcb1Clrwf3pmX91JTF/aCoBTcLf/GRMDEb
sPt6a8TJ/O/ko93lQQyEbpW6lYdg7UfF3kyL0KoKkI1xaj/cKDFMWiCxbakiZL2Nza36UlCNLJdx
QhgQW26DxoMF+MrkWa37rwoUrbXky3/fxuTZFjZhm9jxyW1C24ltrv2BNgLUz0LpM6o/9tcegjok
UINIuO7eDV+M7FB0fisLesHd8A9Ie5g/wMYjwPPsTfw4/YcTlPeDHlbkTpfhzsEydLA28kgf5x9H
dpOstnbgQPwdqY6azJkYgdZs9FOJhJppRWVMBdJbME6KCRaWrS8BUHydzSz9eq+TT1/KOxm1wfNH
5JAjjp771YfStOOT+uwPoraX9wgrHlX1O2zL+CXsEda7yo0aWl+AzI+YNWlGvXIXXY629hgx2EQb
YMLThufVVSyF8tNP
`protect end_protected
