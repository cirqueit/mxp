XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���("%�IMF�dH|T�C��ϫ��c�h���I��D��Z~�!�Үl�n���ٙ�r�݊4i�kG)�{��������"��I��k`Q��qV��MnvI&ȿF�<��M߇= H=� a��g���*9,�L�/Lot�M�џ�!u4v��}�c�d�z��7��#��M��U��2h���	��~�Q4˰\J�S[;�;�Y��ИF�:kg/��?�#���=�7��c ���Z�����JKY��W�q+'�� �5��N��Ǔ��j���i�����d�2���R�C>��K}d^#��o��H[)�?)���wU���-L�H����_CEI��[�� �mN�v��w��	�o#󇏏��ko�	��v�|�
S΀EP̵)�+��4;�M�+�t5��/ӽ�2ڃ���q��|�������Y�T��$���=���G𡏇�2O�<öH���(�����y.[���܃-��~��ja�[�2��h��+���b����cN.�k��J3�q���s����V��5X"��?m�vx�I�tf0����w�T��J�:�C&�~��tu�T��.x��G�о�O�-K��QfiK�@��$[���k�Lŷ7z��L��.o��ir���W�9�b_m�8G:y�'o�t+�g�����S}�9/�Q�N�����C��=́?� 
�m����)��V��,���i�תϵ�[AI���B���	��
�Y
n˜5/Z���Є�,G� yXlxVHYEB     400     190��L��V�~ѶM&��N�`ѧ�TO���!�~bY��I�����s;ӱd|{9�yT�nE� ��Gg�{��ȧ�d��>?�����s��ixf<c��/>���#�l'��Sd��=�ޅjd\�W�K�ƱS�$�?��T� ��ۓ;���(˽d/Wx�6����lxӟě����O�T�?��,W����W~�d<�� ��<j�a�e�v�2Џ��B���$E���z�@�'�^�A����ϊ�ն�]����\�f��Uo�F��47{���B;0��^B�t����kn��0]�1C���v��1�t%��U�^5Fm,A-��÷~U�ɨ^�6E»m�-��Ҏ��PM�1��	�h>�L��Hx,8��TV]�\��`Y��ibXlxVHYEB     400     180wԡf��A�#s���]�"���#�s��L��|7)_�K=\�-Y&����«E�z��#���6�?�qƀO)>%/aa�C��ğ�91F�Ou;h3eU6��ߌ�~MB���/9��4�K��J�.�Tj锆:�8&3ќl�k��_B����0�0��0�|�3~�&�$}��E�|7o�()��]N���Us���%������;ͫ�(�5�<�k�<�0�ᄹ�B��2]ٲ��G�Py<�aC��ϼ�3��q�]w&�Ě� �@ެ���
l�?�{է��r#�l�r�<��)��u�,�Y�Jm��	[T��5~��?�a��	�n$5�`�]?䧓3a�l��[l�XȭYd�o� ��Mr,�o���4z�SnE��1 XlxVHYEB     400      b0��K�>��
��T@ �n�[�9��l�#�\�T6 �S9�I�'�$��C(_8�C�yYyطAD��[I���d��+RG�0/�b�-J���o(qq��ѝQ���� ��Y���
��X�g�c�T7R����9ou��ז�â��TT�^q���t��ߒcF��v8�V�b]%n��XlxVHYEB     400     170�ryIH���u��y�$��"i�P��p���7@/jȜT
+u�R*&�b����ji���=QU�Ȳ�_8���"�Ds��څ�4h����I�&����y��B� B�x�-��Ec�"�s.�G&�d-���Z����?x!�t�Y���O�-�\݉&��Su�%��s�4�n��`�s��=#=��V��z�7'�ja �D���Jf�Ä-{�(Y��x�Ҫ�~��n�k����͟�+���
�:�cܿ�M��c�<7�3���RV_��@XoU�c���@�z�)�F[Ys+]���"`�S贁�)�L7�fw�$E��V�r@Gg�i�E�9��3Ȑ-�X25�ܝ٢+*A�2���4��8�LXlxVHYEB     400      90e�q;�Y0�9�H�p���|6�ˬ�/Z�0�����Qv���
�����Be:�ͺ��_Kڌ������6�5��l��¦ ���X�ta�E�=������"��\�8�YV
����9�L+�iE������n�����ݼ�R�ͭs�=XlxVHYEB     400      90g2���a�m�6ir���(���/B�j��9�r���|a�؛�ǡ\���'�?�ۙ�N�,���{�u�e��EQ��O��MF9�j���o��8k��#�^���g�#��$����C�������uz ���B����9�6�XlxVHYEB     400      90�q�g��+�}�Q׀�Kia����r�J6.;GG.�������q�AD�CCS�
D '�u��9z���G�����^����K%�bb�	���f�8���yp~�"���[��;��-�_� 4�a^ٶ*!a7Ę��.�� �oXlxVHYEB     11d      50�$��9MPT?��z��<�(�I��6,TK���5���Yf�.E�/v)_���2�c�Lt�y��qt@	��7�˂+E���<�