XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C���V��=,	]��T�-r�I�	c� r�,F��a�p*��}K��%�ˢ4ϧh�q�=����i��:H%�0jC�����`��_��w�{�
|�(ƣ"D~kY�
ݪ� wM�1��)|b=��.�-P:�wnU@���PD�DKy$��+�|sɴ��r� �PK����͛$ai]� ��6���@ə�3y1n��48�	1����fW��*R��_-�
t2:f�H7�\`�9���ğ�w[E�Ц��(�m��J��Ku�/��	�ңiyA�i�c�Լ����ط9�2+�]�P��1���Y\�M*,'�����#�>��*׆C�婼���!���U&�y�Ї�@ʺ��#����O!kJ���s�����5Ƞ�eJč����I�^�� rP�S6����\����� K���f�bd~���1m�;m��K��>�Akǀ���PD�:r��+X���]i����3>(�>@�K�����#�j>�D��G��ԟ�].{�N�	������xZ+��b���D�	�#3U)�J�@�:Η�Gy��ي�l�<OH��ޯ�OPT���7��gh�9sFi��Qྒq_��+���Cb�'Bb��m��
�(����?����;~�n���e�C_7�mЦu^ň�R/S�8��3N.n�`C.!�)G�����qe4f��=��ȻXW���b�L�)�z�f��	\^�4k��Z�3p�x�T&"6�JN�w���������44T��XlxVHYEB     400     1b0T�!MZ�N����¨�+�;+=�k�sȎw�6��������̲�lab4�Q�F3�p��S�,L��h�#@��BD��5v��ɿ���8t1M� 	z��E͓��wd?z�/�x�v+LZ!z�U�`*k��|���m� -�9��o+�	�0�-����A7��[��`q��î�9�ѕ8���y`�C�2B���� �&��d����:���V}��v��t�U&�VTW�JO5�J�]f�B�b�.�bc�U�7!z~h0��aj߅<�x�5��@�*!�U������<��F�3�R�y5�wߒ���6{�fU�nA�+ V�h�g/PMM#x34��N��y�f̵�R��P���֠v�nmE8�*\I�^"��A1����Q�J/	��o����<���5=3��sO �UI̴�0v�H�XlxVHYEB     400     160h�>cZP�?"���\��ַ~�wՖE
RP�4�p��D4�=ɍ�RF*	���1m�h�+�
s���6�F)��K:Qh.��7���L�mr��=K'�$%�_�58YE�<|��Q���N-߽o��{��c:�X��h�3`V6H�)Y?���ĝ�1?'�G�^G)J�?_KP�K����_rC��+��v=���U�����2�H���x�,؊ٺQ-�`:���o��=��N��PF&��#BE�?�⨵ͬŝ���^$���8?��� i���S���j����	J�0����	�B��A�JJ��m���*���+���/�><s����DTa�y����d��g�`�jCPMRXlxVHYEB     400     110`�+�#�B	5��]�J����؀N_�]qj}�Q��R�
rs�+�=P�H=Mw�h\�q�ˋ�ս�x���<�{�l��"_{�,�-yT��Ɠr�-�a�X;�1{�%E\�ΜV�Kݰ��5__t������aZQ�)C�P��6S`s!�����)-�X�f#���7�Y*���*��������i��wW���o��6Nߥ>	)"�}f;j�C���D���U�*]8NoG�5��ɒ����ńC�MG��q�o�2룃�/`�Zj�XlxVHYEB      42      50��%�{�?JE���/Lv]��X��=�BVW���%#����>�-���U��;�K�JjX����x�J���p>S����