��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����ϑ�O,#jj:S���f��l<���djf/��'��K����G*�	H���o�

g����.��P<�M�Wv+#�Ql|i�Un�&�7Q�A�	�:e����&ipk�E�wL�y^N?Ưq$��S9q�6�P	��}8�,I�q]���z[�k��o>΀D�(s)��p�l�A�6�v��t�f��� R�l�_d���Z�x��}	�,@����Fn��T����ȰX�yb����L�'���'&~#�o���C�z���)��2\��9��bt��IT��Y8x�Q��u�S�V{ϕ��)~�R2Ҏ>h�3g�S�<Y_��e�׼�ܵ���=�/�N)7���E�ٔ%=CH�2�/���/˻"��0���d��u�B�K�I��F~샷�`���^T6q�
&���^���V&�{���ƿ�[��Wxz�J�Y:��i���~�t���P+;Ck���Q�G����� Y�] ��!��)���}OJ��ހr֦Z(J�>����̈x% �O��B�x�d���h�Z�ޤKMt��;�E�[��az�Z���fA�>+�1��ÍL�%�ѮB�� �,��.�)�n���EZ1�v�D�f �_,/+Lc_aV�u��e�9�i�9Ra���r	7ﭛ3�
n^�N�|؜1�Y�,��-����7���ݩ�?�"��$]Np����&�$�˽�YX�*M����#�������8� P�9��'k�k�|s��x f�1M�Tf�D�!ȩ0��ˌ{�pH����о�*���ޙ�ǒm��.k�ią6�����є�8B$�q�C[T��Y]Y�8җ�@w38 ������I��M��=�/��:�k_��$W���Ѷ�M���/R��`ԝ&v5��,|B�ݡ�A�����Ĥ������4K1�M^b��(.�cux�~q������"n��̩��S��Y�>�o�ύ�g�'o�<s���]cz�N�%�%��u'�p��r*1K8�T6��Z����r��!JEr+u8�b>MaW<)v�k�KĎ�Ã�z�ewN+�8��0��'c0������E�ˀ _���jz��Ǥ
[z �>�:f"��a�O'�[��x*Kg��}[�o6�/���'r�}Dd8
�P�����������t��H
k����\<���k!�P\�Ŀ��\�[�����>���L]���SѠ4z ��Y=(�S(�'�`em��ɟ��ԣ:���ϙ�趃���7�9�JK���"٤h</��u��@�Q�gbo�8���`剺 7�#r��Lg��Wa�YX>'���Cǃ�mLy��� v���'r&��!����E��nǷ7����ޅc-�b��|��{�,������o�7�"?��M%���fAb������1�����G ;M���>�9R�	��c�x��ZL<gq����IJ�I!V2�}�K��7��
{�*��e����Ѕ�I��[1K�Rjm)��Г����^N�.	�މ��H?B=��ݩ��j��5����?�u��Poý���0܄1Lw�"ۆJ����-��E�qH�׶��н]}��O��w�S�ˤM��-�"2�+2Z)j�&��<+����J�΢̀��IM��(1�y \N�Iҩ�2rv���߾}uƺ�LlR��ϯ�B��D�����6d��+���$�80���O�	_*�K�@Q[R �����PY��0���6	).�^%-�@;�6{6sM�{���];}n�*b�B2P\\n�ůo�l�̃W�]��m�7�=�}Ϡ���spl�ſ�)�|��%<��?n���@?1��>��q �IԢ�l=x��I~]�v�h�[#i�ETu��jcvS�b��3�3��]u%;T�턖	�A�#��J�{ށ��]��,�J�͢�]LyFQ&�=VJ��ռU�bP>�L�˂���A,s)�p�q��	\��k:>K��VT�:f�B�p��R��:Sv_T���������?1,��ppd*�j�h&���7�OC$��3�:WC�b��s�y�!�۔�.N�����9�5�a��	�Kl�ۗ��M���7Sw����"��v۾a����Dk�Wq͍RT��JY#�` n����ݝ����u�A~�ݜaa�*�1{����(�$4����!
�)(P�<�?�����{�o;��7v�0���
a[c&����6���Bq��T��B���ئ�#�U�RЪq���֖_O�W6Uv���穉�ѡ�q���#�)*���D�����=�l�	`��jaxA��rJ4 �6�
��9-�3"+�T���<����"�Y��o��ń�s:�Nv����InAAf�F� �1�2t��˷���E��[��ELE�(��px�<^Z܃