XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����m��� ���U�����v;��i������"D��Pr�д��D�e�{�j���x��{� ����X�HP�.fN�_d,jR�����So#ş9DS��Ă��q��0��j���G?����s�o:�(��nY(�M?��l��)��d�61�;U��(�Y�v�5�:�F�I��{��f<���E_�9�b�5��A<lI\͢����9��[s@�=�5�4k���6��'O����r�Ò��3��+A-"�	(�:�Ԯ/��Ը��L>R3��Eh��b~���ۏ�Q��:�6X
�U�e�\�f,0�����s��b8y������}�gY��\"�忉ߨ=�bN���z�BM��ز�{����"�����|`��XiGU�̤:��ԃ7�d���k�=<�����߫l�1\����ý)R�����~����19�؛��\ǌT���BC����0�
�|�
�����N��y�`{���BF���dq3�v��b�sT-&� ՟C'�*��+���Y�X|�I!�_KM�0�.��&����U]_2���4��Fx�:�Kg��A�	{y��4J�(W��"�������Б\�ǳt�j0�}�msn��,3����@�xN'rI�4=a2��d���{K�y�8&��^e<e�b(i��WW
�����(!��9�5��K����Q?
�As����
WR�-c� P�Q�si%]�	�5�|���[��CՉ��9٨)�6VhOXlxVHYEB     400     1c0�>��oVO �1����Zr�M�l��e<!(��_?؆�%�}�.�t�z�
{v�?��F��3K�+ٛ�O6L�����m�\�}��e�Y�M�(��6k7��(`Q��%S�- �r�l������>�щ�G���Ghqg�b��,���qplU�]����7�0��u6&B��u�E�D�UJ�|�Z7�g(A� T�XQNZ)!��l ���%p�-JG8[�{��E�X=4ߍ�� Z ^L���K��c
��@&�2$K�	~w��t��:j����h��<�4�&V�L���b���_��b�O�r]�'�I��52�נ:zp��j���DDZ.-H߱������� x��N�!S�72ܬzh.`�B��������{ De"-�!�~7+�ؘ��_Ey�HPGN(����+��&0�z%�޲�\b�0p��-��FFZ�rfXlxVHYEB     400     180�w���,�9��Y���Ze!cg��񙑇�`�ܧ}&w��l�h_�P(��A�K1#2T�uX�	�i�X�rQs�;2�o瘑ՅT	�Z�&K�8wE�j�y�.W�6���w�b�Nt�/�=[F8L^�� g;-%�G����Ç��7{q�@�����S}��� ���f�y�f�ۂ�2_��8[���>)ڒ��[4�l���t�"7щ������)��i��W_�b��e	f�t�dח��!^�?Mw���I,2�+\���� �/OX�ZsH׳��r��'�-C3�J��f�V?�	�#ur٣e��7��&�� ��(�@���p��d/�O�9�9_���)z�ߍbR4�i��.;�p���D�eB1P��|Bh8�D��,U�XlxVHYEB     400     150-:Q/C���Dk�����}h&{s��Wf�kĮ����k��c�����;a2ڽ���S2��_vg#"�c�$�ORk��7��J�.B�w�+9(��^�!;[U�M�Y�|��~���AP�o�|�������
_�-�ۼE���Y��~es�8_,ڌ^h$�怋�����~��~�����9t�)�/W>/�j��M���/M�zj���%�s/#��%9 7o���$�]c.*y6���|�Bb�b7Kۣ��l��,�uCI������J奔33N/����y�K�y]9e������|G���ٓ�r�N!!@h�R��պXlxVHYEB     400     1b0�����˲�6𩣵1�IKg�7W���{+��i�����}OF���h��w�r"G��G����^]����*��pS�.6޼&���{�V(������u�VD��.���ų=�נ9� �^oO��U�����r���.���Ӄv���Z����4B�D�j���]�Q	�/�X&�r�d��2�^�s�Yq
��r���ju��:��?o�ռ�!ڈ�D�oӸb�<_���|u�@�}��g��a����:�s��o6���qO��2Kd�+>˴+��Ճ��*'�^F��`�N 3l�Ty��l�|�D����B��f�0�qC�ωR�x�N2�3FW��SL�o����9Hހ���M��uڟEI�v�������k	��Ι�d�����VX�v�V�7��X��א�` =E�a��XlxVHYEB     400     100CgJ�`�.Xa}��fu�Kf�]ZX��j~YK��b���h&w�~���P6؟��jb�Gv�;�zpp��0K�,�1i8i�w�L�fmwd��Y�:���J��?B�������tZ�W���.�Ne�U�"y�U+���J�:�̑A����:+G�q3o�Y`�R�ȣ�9%��kՠ����^�����e���X�k�a��U�M1if�S��;��j+��]QȺ!�di�i����pE���To)�\K9�:��i0XlxVHYEB     400     120�:y����3��'�իz�IuX��iW]�k���H�r�K��jb�ڪ(B�7o-�}��q. Oh$&�A��P�:���HGi;���4��'hbc������L=щ��ܓ#��/�	���z/������x|`��<���z��UG�m��)9ͧ@!/���&8�$'8������D�9#}H��1����9��B"i����FE�f�ރ-Áp��nQ�w[�`��1
�����)�m��v�(v�N�~�6�r�z�*M�n����s��-��c1q�vਣ0��FhG�XlxVHYEB     400     160r˹ ������~�x�D"����������^ۿ#�7:�ɝu�vE�o�W�hw?��S�9s�3�
�9<��<��	�d��oD���ƿ���tY��L�,%T��qy�h��.�"�A��A�*���n)H��>���(H�a��kA�w�)րDT��0��廞���Bo\6v���UWi���KA����xa�I�D"d9�6d��lhf#���^��g��[��p�� ?#�j�� m��>����⹿��x�c���*$�#�����c��n7�~.;�V�{tHA�#�������~C�~q�J<�M��\����K۸���	�C�����5��PMR��XlxVHYEB     400     110y-��WH^��m'�Y�a�[u�2��e92@5m��	�DP��@QV��}qm�ҹv�E��lt����n�F���k~����sAv��8b��k���h��H� $0�J����{���|~_Z�EV/��ݿf��D�Q`��m8ٚ���6�;����%�<?��$��A�� &gs����s��<�4yhe?G��ss!7�����a�»],���6l�kC�a�&��'Rxoh�Hcl �����ax�(���Lлބ���L59XlxVHYEB     400     100���q ���y!���(�ZL�E0�&���0-���o0K�.I��?X3����,u�k0�!ċ�U��q����%2��C�F�I�a�������u���tsu�� �9��*��\,�i��Ǹ�9����t��"����ᅫ��0�x�V�E���{Wp"G�`�$l�_(�BPYb���)uu���%KG��z�n��ZM(�7"P<]K���d��s6��ۃ'���`��M;�s��FN��7�y���XlxVHYEB     400      d0�����Rr s�>��ʷ.�mw�%���u�6��gs!n��f�����[��N_+j�e	����}xU��H�(��f�$H�
(e��K��S�^(`+�2'Jڙ�T�́oϙ�Ǟ�>< Ί��L��t虁=�3�DO-|��N ���o�[�;��=/�uI�K�:˪��,P>�0;�R��4�#XQXlxVHYEB     400      d0�]�;6P���O�E�	p (�s�e1��4  ���yd��O���>Kj���;��!�վO��?W�P�-�q�!C���54�
��?H�	uƬ���ao�����\%�ճ�'��ߘ���Xs�.h�U�^�uqO�霆�BŮ�#Dgk%��ʴm#6�:YB�U5�Yv�o	��yn��k�a��]�K�'H!x�>b8�8�~���P�:XlxVHYEB     400     130�Q�Ĉ��뭕�qR�T`��]%�h��
��� �o&�`���4DM^�3P�"I���
Zf\q�v�o�ަ <k�^��p ��z�K�S*��j���T���%�x�З0�9eS��E��~��	k�6���K�u�i��H�x�*�O��*Q~����1%��b�|�i�I�i�'�+'�zI��Z�\�_)�����Ea�"����\pZR8���C ��͋���,��}��C�ǫ
��Z��)X'�a��~t�򡦘�,��!�Mz����h��QKK�ܲ?��^���
!N�[����XlxVHYEB     400     1500��#�B2��o�w�5rrT�.H���J*�4�ׂM+�����?���T�ґ���!ƶ8�E�ј�3���.Oy$ģ(����_ ��/���MVN"��5�SZ��f��fp������eQ�B����bVI�<6� �<Xv�J�=��:y�]S��&�XUr�!��ZZi������+�"��ElCb�F���TgGW�'�g�:�C�[_[���q��1W�#s�s�}8�:Pݴ ��/#ԏ��uTD���^ƽ)PV�?b3ES�������Dat�d`������s�Aa�?����mrl��9�I8��4��!L���t���G��p�XlxVHYEB     400     170`��| !���w��bb���@+lz��� G�4.j�0���;f�4=`g�ċ�y�<�#������?jS���(@t����~���>�Sv�>��~9��������(=<t7���Вm�w7S�2�{�~rʮ#H{�1M���'� �7ZB�*E��yB�G5!�jW�Kr�u<��CmyVd�`�.������2�Wp��%?����6���K�j����JQ����������^J�kc�y�g�!�"g����E���|X�*I������"�HUo��T�3�cʷ?-,=|z�¼W�����:��\!��[)pЪ�g���j��9A���l��W�Q������;�c�M�sS�A8l�%�c
v	XlxVHYEB     400     190�'iL[�Mz��i�����3�qSP�.=^]�^.�)��F�;â��PDAr���ܨ�I��bIӣZ�A��,^��y羣��SmuԹd��c9����R��ck��3���]�ݵu������P��B�>3����?~ke�ywx���.�6}C0�E�%eb�X2d����N'oW)�6Yç=�KV7~��	p���7}X��m��J��*�ӈs�Mއ^��fܦ��H�u4qAj�4Q�\�g����!�	�5�rdw��˔��$q[l������'o$���I&��1� �O<1)z����l���?֩5����÷����s���1gF$�j[�T.��T
$��u�	����|���StL�@��(f���*�0d<<1�%a��E�XlxVHYEB     400     180�C�eO��%?�G|���,bz���C���uԔń o^"c]"���U�H}mj�r��	{���:.�,]X��n�7�6��N4-;���8V#�TĖ~���;Ƀ*V"!��`>�8~��0��:�~�]�!K6���n��ʓ��|����o�lk�k���Wos�'�ydCvd1z-P��涴m���,3�%I��-QR��*'l�Hm�0���8}[m��&���1���^&�s�S�GtN���k�����^P�;���A����ֶ�T���΄*d�u�>�,�N��
�+[1�$�+�mJ��#����m%�1�o��EY�� 
{M�$DDp�1��nMJ݆ܕ�\���(�	*jh����\�|���XlxVHYEB     400     140GEJ�?p6�g�DD�&E�d5�L�]�� gwϓ=t]����-�G����]��
`��@�rWI!>Vz�2]�JK�6�?!��e>��ZI�b��2p�gF�(
�L��)�t;94�/�X�{X\Mɞ�g�
2�$����8DA��4�M�&]u��Z�0{ܗoF+�B���%W�K�M��ra�́��w�0�]1֢u�������ҵ�AD�,��ΡR�aƓX�F���ȼ���Mc���Ag^���u���P�QmB���(��� �dN)�~w ��t�����$;`|�ϵ���B�/}�G�Z,3җ��29�~B�$k\oXlxVHYEB     400     130��w>b�ơ]y{�dN'�םa>4Pg��r�V�T�:���M��G��!q;�1C�F��7u��6m�>f*P|�b���)�f6$�G�;�<r�n�	!��>>�SZo,G���r+r��:��Х�|��&o}����~��Ĉ4 �ٽ��1{��Y�T�Cr�q��'��{廲������vu���~��}�j'Zm�h����kx�u�����%
��\��}jcR��80i��M?��!H�qy��OV��a]jړ���3��V�M��?�s�O�(~?��i➐����%y����>XlxVHYEB     400     170�:�� #
��#Ӽ��qX�a��+�
ɪf��MYP�u�>���0aDҺ��$`�7�k��Aٽ�����7i�C���3λ�K��L���;Hp��|`qݓ�Exv�dM@��U�3��q�VF�?P#b� ���\�H�'���u�@��'F�Ln�٘#"�]��L��-�m�.�(KG��c��ո��`��ѵG����Tx��8��AW�q�?L\�ƽ���S�j3���O�Օ�pِ�p͞�E�]��Gu�Q�X<z������[n��������/P:A�9��`���!ŠE����Vk��־ �}D��,�MsJ~si��s�H<�w�pkA�Io�E�֢�h��u����;�lx�XlxVHYEB     400     120���4b�7�!/T�2(i[	�e�bP�,-��,^��Ys/���_���:[2Q��7~Ir���e��5�
��^O�����w����|�ڔ}����[1C��0��2�J����gۥ�՟�r��U=Â�,��e\�W]O���f�Cy;!v�<{".!86�/\J��� �$���ٙ�0	 �$�i5�g̿c]ޢ̄≔���Dq��9/(��0��dw�~n>|2)�в���}��k?C4%�T1����h�谕p�Xdh�7#��
�1�M��}4i���&;��F�XlxVHYEB     400     130�iJ��?:{�a�2�	#c����o"��tجW�nN�w!w���
[C�4�́��Y"_�M��/ ��y�H���7���4Jц`W�Ix>�MEpd���\��80���wt��:	ƴ��Caa;2[��:��: ��X��,���?�/n��ёA��fcG��+7\߱h~��l��z98���X�oT+�f��
��c��E�Cܫ:,2^~*���[�8����燦���w�B��^�D�T������ 3����0ħ#�hN��z}�$7I�O�3�V��F@�U��;��XlxVHYEB     400     140aܱ�0�f47�c0����S˜Z,+Â�/��m5*��"�4�B$P�����r��S�u[*cgV\��9Pf�
�5T�eb�3r�0Kʹ�v��`v^�7n�ρ^��{2a��]��]�|M������%f�;���b,�EvQ�&+��k���l�V�+(~�+����LIh)��_��x�%7"-Aʎ;����l�����j�k�d"�E�g>��\
�U������o�Ǜ@��ǽ�8�B��&��2B��.$�KDdJTLM��,03��9�'���<���*�MŗM$K�|i�7�1�/�}��Z�-u]Gq�nHbG$��BXlxVHYEB     400     1a0��c�GvNΒ|�V���T���e�*��˒Dگ�M�}��G���]���F��w������d�۳QW��.��ڎ5:͢��AqʟwY	`�3��"��J�o��-�&�G{�4G�:M�ł���w��&�G�Y�U�n�F7�.�/E,����|����K��)*��1��9S{k���8
5G7Q��&�V�.����-��6g_������xG�Z0�bj�ї���9��+-�(�<9i�S����q����.Y�n��AW��]�;}ٔ��=oח�iV�{|�x�m`���4����I�X�VYS���̲���,c,��.(K./x��7Q��b�1w�3���0�D)=�AW�����}��0 �1�S�>1��H�r��b�2!΅x7g�!gG���w�i��$9�f|XlxVHYEB     400     1802�ܾ�\��5�\>�-��x�2���x���N2.'Q�O�~����2��DC���5���ex��$�M�]�Q���k����!�Ҍ��i��:��� -6V8�ˬ��%�/LfȂ��^�s���#Aj�l2�֠l>u�욻ؗ�η�'ي��q�!Fl�� ��j��L-��<�����I'���:�	��*a����T���}6�ԉ�Mgiv_,�.6W<xmÀ�v�B��7�aӞ�X�a[�J��2<(�T��2D�W�g�?�o��]�%�����dkU������*���e��\T\�m�Y;��X-�O��������<�**<�yd��9��2���մ����v��=�:9"����XlxVHYEB     400     170u��R��
�krඍ��i}xl�!�Z�:�^�|�o(�ԙ-Hn1��)G���2R�/t���{��o<��oP��"	���b�������y>�+3���^p�S�a��ei�ϥ�
B�`����MQP�ɮ��>����.�老����L����R�_u
V��_v>�nP���{.p�[yb&�hTb�[fl=\����0���L�d�>�"��Xb�D۔K�W���&�~�3y����f?[n�b�Z�oA���Z0�4�-���W������Um������Y�]������,�I`���W����w8 ��i�tH�e��,�eb�a)�0o���m�'��C� 5���Y�MM�.���^��Z�B�XlxVHYEB     400     1e0��񩀥����m3qE&�+�p�X��M��9�������>��=���77S����B+s����iκ[h$o�6^���.�}.�t�#c�8h��s{dG�M��D�n���}��xy��-L��nk�V��YU���(�&x���N:��b��,�ۑ4[���o�#ڦ��H�a���9���l'�%=w�s1��3��І�8�0�?I�sNC��P�뼭����%q�cu�{h�T�J���9�پ��ĳ�� ��Pc��=R��F=fCϥ�Hzu�4$�4n<��b��I���6��:Avf����7�a#����
��i�&RQ(gƩ��'�R��r��M�BM5K��RN�^���r�(�� 07m�v���N
�@Z��:���u�9wJ|�>�՝��wY�:\i��i	��o��<��x-(������q�&vT������N��yߚ�M*L����H{�{3XlxVHYEB     400     1b0cK)O0#�u���� �^�h6�.Tb��6�Z����!TB�~�
�£o�t�F����Ǆ�:��*�}��	@A&UJ�0 Y��l�K�m����ֺB����Q'_ ��OϫD.WB��:�R����.IvA�춵7�ئO�=�϶�?�IÄ*ּt<��fWDUi�0�	
�4�{�5����������!Q<�����M�7`����ܮ���u�b���7�������f�ʃ-�6�5���_U�ʱ��2�*TH�U������wU��;�D� ~qF(ŪCsx^+��z�l�,�w�~��$�ATabC�v�  �.�m����A-a�`�yc�!ʋr6���7V~��&���Qh�2���l�]��I��߽��O�|��#*ۿw=u��uSn ��m)p�݀0��_�~E6.�(���2��||����;<�mOXlxVHYEB     400     160s���/b�_�{ǭ�/(�پ�)E���8��S�a�M����<�\y�*�W�����G��t��*^ND��:]�<��"�.n�������%O_@�S���fV�(2�?��ج�o9[��0�"��k������O��}��9�Ց��V�Z��OVI�b;x?`-������]�j��!ŗT�nU]Z�#�L���ـrЁ)S��R_#�G�Ǚ@"���(5�Y����v���3^1�n*~6_4�t�����e�y �M�����ʂ/Ǐä��rc#o<�Q4vj��,B�Á���y:JiA���N�Y�Wkk�R�^���R�>�?>��ZUH{JOy8�2�[��XlxVHYEB     400     150�2�a�1Ze�^�����T'�/��3��!ϗ+�`�)`��3��m�Q�@1#1���G>�_w����R^e��|�q��&e�m��*>�w��ݎ��#ǒ�=�S3�#/��*W��5�o<���yB�X���uA%��5�	x"Zظ*w��XT�s��?OA^[���bH�jf"{B��:��C������Uyy.���m.2O���K}������<���aWR�i�~�nP��u&��o�����k©ƕ��%�W7�!7�>�j�NVӞ#�S�0ѻ��)1�5wo'����h��ډqe������%���J<T�ͳߡ��C;��2Q[J˩5kA���;��XlxVHYEB     400     1a09X�U������_�=��2$������B��5+�$�%�2e&`�ߝ��!B��1G���(�2w���jO$7�a�=L�ǚ� K���q����l�_^�MOH�s�F�Uy^��%��s0i��+�Ƶ�P�bɇ�ge���RbҐF�
2���G����u�g"�`��vTw��k_(�U����U��]v;�ӑ��rL�ʪ�u�l3�F�)@������ ���)�US�R���tҮ4�H�.���ȧ�0ux�`A،�~�s�p�v�I|,��#2ǷH�6Ȭv匳��v�KO$�(9h�B�2M���U*B(�_�DF���C����a�����Ԟ�K�)]9��V��
=��emT�� Q�|���o�L��g
�nB,��kv�X�<���s,�٤�`�ދ��!XlxVHYEB     400     150V����񕏩��k��#���/��?��n:6z��.�ds!Q8����tH�"_ީ~k�R�ŝ�����2e���}�:��ݱir���N����&^�z���`8��5�,������y=��a^w�=uϷX��1�t
F��ʜ��ǥ��v��m�G�[ �&6��>!��_%��X�Σi��oAes�a��l�� ;���Zq�kGW(�U��2 ���̬��Or��׸���w�\�y�(&��WVm��'�xy>z��������ί4�D9�t�n@��d�ziDn�aBLWA\n�8_�,��(�V&�ه���9��Ҝ8�XlxVHYEB     400      e0^�w`#B]��u뢕�@�b�X dL7��xxK�S�m.����Q������%� ���2{�Go
{>�����۔�GN*��r�W���Ű��d��y�m-{E��.��^�������@d�1��j���Ws���yR�F����D�/��.gnA��
d����o����h�� �2�i'l�W�x���i�>�Q4�P�n!�&:8���?�XlxVHYEB     400      e0���^����*b5���{N	�̌J�+[a:�����X�fע�<^�6��48�|FQ+2�C-Z<� ���1����]
,\PHRW��P\-^�����F��^f���R�/�&� /@͍���Q���MSBK�������w��(�x���ׄeC�H.DW@���o��-G���.��˛�5[P}��!)[+k�yt�fڼ-����4���Ɵ��ڿ���XlxVHYEB     400      f0��s�4�v"RS~��^�c�ݞ$o��][a�8�@W��u��_s[(�g�p6gR06����-���/��`K��?���c�I8<����=u����ܗ\�M�xΣJ��}<��߳��M��������ټkk94&�Q:̠O�{��P�)�G;��Ruǐp�o�CرZ	�)���O�_�c�ɜ����u��8K��y9��˾���F�a��	_�{5��h�� '��c>X"_��XlxVHYEB     400      f08P)��S�p9p�!D�橅�ZȒdK���_�����!x9F'1Z,�1=�L4����\�ʽ�*E!��Y���l+�)���<b��68$N�zӸ�m�1���Aq�9����ʚ�T<6p� sºq����G9�s�22��R�!�F�}yʂS7�#6�J�pd�ZR�ws�j)�n�1h��a���5b[�h��gM��K�V���D���N�)�i��H"�.��	D����D��Ǩ�fXlxVHYEB     400     110:��(&l�*��҂�M �Wg)�/�r��};�?6�2�9�+�4�y��$�F�&��C�A2 ��Ix�;p�j�k�\�&��O�9\��Zꄝ�6&�f��Z�Z������ԡ�<����JX��*�.n�k|�v9�s���F=9Rp4�v0F��QB�����>laT,��W����U���@{�џ���ĢO>*a�j^�on�c6���r�N��C����ݙZ��V�3��	z�N�4�8A'�ɒ~Qv����}y�8Z����vۋ�ή�zXlxVHYEB     400     1b0������L��� H�1`|�߷��O�M�1�[��E�L?�h&�`h�97㜢DRCZ�)gS���������M��N9P�8&�4�� F�s锱70~��2��D��8{��m��11��g��k{�r��2o�L��C�˵���'�S�Gtc%��a$�����~	���(ڔ��?�S�[���m���ҠJe�U�4�p���4z�c��� u����uQ��ZON��kIS�&��� 5��F6��0?�Yy��t��Iks��fnǭca읚�;���E�k�z�k�0bj��*�ļ��آ|6�{%�����$2wǦc�L��'.4kX�o,��_��9�a�?����;���<���������+�n@�H�������W�>���"�	��|�L3��4I�u��tW�UXlxVHYEB     400     140w�m�p���<�?o��1�:���T�-��=�Eo�f6�$"�����Yn^�"����Ѽ�}��[��"Cb߶a�0�*��d�/>����2�\��G�&�������#�R�"��m�rŔ�_�����0QŹõ��9$ֺ8���f x.�V��p�V̳�;��9d5�� |ť��4N=g�1��֎���G��I�m�����-�����T�	�B�Bx�RnYi��ν� ܴ�m�d�{7{Gv��ξM*�אc��9�@�p[/o�t4�>"��Beئ��-�9�G*b�K�ǽ|ׄ�J��_��s� XlxVHYEB     400     160��t����ك�'V���O��W�L�ǻ���˚�H�#�[5�q%2�� ��q� 9�1�[�=~;�`�חaE�g(s ��*�:3���io����D�ksx���R�!�x<�&;�J��ٺ��%�3MH���z��5 vS��h�)Օ���F������$dK��V�⯒��Q���e���N����SềS,���Q@�R#-��ԥ*�hO�ɻv:�&�XW~.�H�-
�h�(��w�4���5K�rtbV��c�eS��Ε#���u�b�`�-�nf#�i�[d���Ѣe�Ej�U!L��1��u�|5:n�\��᎕��9Me�X*�*��}J��?�XlxVHYEB     400     140��'��H��@2MO�%.�E��e�o`���[�����_x����n�F���_�-��0č�z�c��9p�$��Z<%R���{P?7?�-��i�9>��R�0�#v�Z���:K��թ*��A�iNK2�x0-�b�c�����cZ��o��O�|{������x7��AC�,�[��n	֧r�T�
K�:=|H�Hu�*�9Y�{�1�+�C#�-8�����X�!Ȉ,��k��qR�n$ڮs"O�?Ќ��I5c����܍��2���Do���bQ�:���]8M��s��#��WŰVb�A`�'�S[XlxVHYEB     400     180�������xd_��%�s�o�4֐E�4Mz�V��E{�
/�*?�}(�W��Ao�">��j ��~P�����+K�b�{9#����ފ`�.	�<���z�@�&%��aW)al����"��j.�MsL^�Z��E�~��<E�f�������<�#vYd+g��[Aj~<���af����LwY�Cv�ׅ�I|����L�ڡ����Ibhk �R9ƊY���m�LE�GN����f	��D�����C۞�d0�s�O�$�l�{^���.x�yL���f_ ���|�1�����O*����j[ �zf�����>�y�2M��M"�z��pC��>}@�Y��A��96l�Ӊ��������,�S�~�ҍlUл<lQM�R��XlxVHYEB     400     190���si_}r�ש?J����-���D�ޗz�~b��=j�kIʲWi�J����#�� ��j�Vc�(��<�{��-�a�8��#ȍ���8�����d]ͼpѷ�KӴ�����n'R�����;�|�p�w�^w���0�ph���/F���f�?��(�pc�ͨ��Q�tU*�w�VW�[��?󡫁�G�;��EX]\����]<�A�$Y{AAn�{΁X��1J󟿙����O�&�\��l7*�I�ܤE��X����y1YB���-�bO)϶P>>3k[���{�e���Q�<���bW��r,�e�6w��D+�[��o$��@|:�l�nm���� �B{�=٭�� :�H��୑o�3;"����`�Aݷ<XlxVHYEB     400     150[��Y�/�7H�+[�I}��9��U>�o���-JPà�ԯZ�V�@������ \�i�9SH�׈ �G�aZ95��;��������1ReK d;�%~��ey#�m�Kh�U8Sb %,{$�F�WҨ�t��\� �:O�v)$V�|fk�����¥�)�6������e;����!n��c�b�^+~��H�A��� �QSs�e8�h��%��.����U� �L��C]��1E	����3�Y����6{�=�|�d�����Cq ��q��Ų��ً7#S&�Y��R��\7`dd5��(.
�-��P���X#{�7�XlxVHYEB     400     1a0�VB�y���lĮ�Aj�����	�GM/(M���Q�j~|��Mrpm'x4�ޛ��rte�)��d��9�+�y��(�ʼȾ�&Ah�Lt�b,���Gy.0���=�g};�J��܁6�RĿ�=:�DQ7��ꃄ|��F��츝�Q�̒�� 4��ŀ�d��'M	�<�|JN氍��M_�C�uK�+!S��Q�O�?̋�],���B8�ν���Z�#a����U��W+V'.3�}`r�ur���qtD�m�*1��2�-�2��=�(Ҕt{��}���) s�~�YTݥ	��B��b���_��mi8H}k6���6������oC�݊�O���ƧoV��E�z�8M4P�L���暑ΑF��k\��V*�H�s���T��&�a���[BXlxVHYEB     400      f0ph+R;L`���Io�^p���3���%ue	�y��t���lƤа��䫼����K�z�
�'��N��W���K����,��z��;�<o�و)��5���'˩Ȏ�"�U�ڦ���h(�mm�+W�-��>A���*��V���f>.�xϹl���[4,��,gV��4�\��V��P��#Rn"�?�&��\3⥔��W�<���K؄��������7yܛ�[F0�Xت�XlxVHYEB     400     100PU7��c~�t����np%3�Ƥ5��P��Z�2i	-�U����~��HJ� %����V��O�-D�g�2��=�f@�e�&��k��}�q2�bzC]��]�Gu̯U8�\'h�s����w�{线�"�N���	&x	m'$!��6��u^� �F
YvD;�A�_Ô�7W>����o�,��4��2��`�4SS`߬��eӭ�*2�M���EE1m�Ў�%0�ג�R�,܃l�k���_d�ȦV�XlxVHYEB     400      f0������]���Cپ2�C	��豇7�g9�V1�>o�#$����]Ƚ��֘�sop�H-�����ʯ����Ѵ([|y�NL9N�)��i�f�f�=�������@e-�����,�����=���n����j*}"O�T��y��Mw�}cy�&�0��S��ԠFD�Q+��l�(L��5��[�	��6Fڬ���$�r���.[�;�)�r1��0?}e�ź���p��ЭDXlxVHYEB     400     120Z���]�ʍ�`�d|�'�(��6r��V��*��p>�p�~��
5�:4	,'�?���_b�g,���0��?hC�w���˼/�4�Ǫ�%�*5��'�4{�r�b<�gUy��-��P�%KjFYm�S���{T�n�Ϭ��3$י
�����Y�����}ײ;��Ԃ���#��iY�$M��{�;cδ�����ﾍ�΍����ƶ���Vܙ�iF0'��K?nLrrȣ:|���>��	�(K2A�+s Q3w[��?,'<����_�z4a��H�����l��XlxVHYEB     400      c0�E�#ij�����^�ԓ$���Y�9��Z� �с��5�����z�s�tX����Q'bzQfgee���F_O �GRR'ث��( �_+�7q0Y|��zK{�������u�,դ��sI�#�#���f�[&�8���ר�E�v�@��T7�a�i�a���6���gD�����/�k�}�)��9w�XlxVHYEB     400     150��U�jס+OV���C5�&�8��x��1v�-��S�$��f�)
������5���;�st�@�z��*�F����+@�&�Y#�j�:����וd�5�b���]��^/�:g�%�*v�d����,H�-tQ�96��[|;�M����9��0�d�ǖD�s���G��?��0{�7Lp��ܧ��E��g�������C��WAQ\���f�*r|��?q%�<�lk>��6���҉�Aa��k�I����t"B��QQ˶.��Ǻ�ĉe�7�rЕ;j�[�Y�AH)7��;��Kk��� �r�$��{w��+w�}s��}�_Bk�Q<,S�ZXlxVHYEB     400     130i�媚f�IAA� �7L+M����s�E_$3G�p��%���,�ox�6l&^���$�h"����qԵ:�!"������{6(��t����-�����̧�_p�:��p�i&��qp4m�Q_:gf�c���+lFw����$�۫�/L�98_�P���.�(uvs�	6��;u� e
�����6���.���.�y����J��R��n8�ӱBnW/��<X����YRa�|Mz��5U��S�������I�_Y$����M�"Q�R��;�!��1�z;*C=�_覰���	szqXlxVHYEB     353     160���Wc��N�V�VD�.'+OI�(��4��H�eex��<��Y�MF�I����=84�	����#�$�+SX��}�%��.?���C]��e����%����H&�'p�~�ȺY6F�'#iro��|�܌ڞ�k�<��y�]X����!�#�l�ہ���۠sR F���l?xM��[�PO+f��P\+��xM�F��,�S�*��dt��Y��h{����{���ܑcR��#/��F���)â�N�Mu�8A��b
�Acs���j������\/��|�Nz��(�b����1�+�9�K��IOb���GW� �&2P�U�(co���.<���EXJ�4S�?