-- lut_pkg.vhd
-- Copyright (C) 2014 VectorBlox Computing, Inc.
-- synthesis library vci_lut_lib
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
package lut_pkg is
	type lut_memory is array (0 to 128) of std_logic_vector(255 downto 0);
	type byte_memory is array (0 to 128) of std_logic_vector(7 downto 0);
	constant lut : lut_memory := (
		0 => x"ffcfffef_424182bf_8daeca81_d184a3ef_fbc5539b_00042087_ff458d83_c044f0d4",
		1 => x"fbefabab_d20b12ab_eb4aa00a_cb47b8af_e1d78007_22010000_f1d1c06f_f1c7aa8a",
		2 => x"a0cae8ae_da26dbee_eb9fe009_eccbb0fe_801ce01a_5082089f_f8fc0099_fed6fdff",
		3 => x"ffe3e2cf_8345b9ab_128a008a_102900fd_db7f509b_0010508f_d313c283_60da62f7",
		4 => x"ff275020_d7816075_89415299_f885faff_dfafc187_d105956f_f78b8385_fd5fdbf7",
		5 => x"ffcffa9f_bbd3cbab_bbb882ab_c303f1fb_b9873513_5943914f_33113113_3197b333",
		6 => x"dddfceff_eb47e313_134b8082_e302f053_c24ec70a_00112002_a6bec1ad_e6dfea82",
		7 => x"f048bffa_bbebedfa_d28082ac_f5b3cd9f_fe2ec58a_1800fae6_505c029e_e0ccefce",
		8 => x"6eef42ff_450501cd_05190980_2044604c_ac0f698d_9101a37f_4f1bc713_f5e9f1dd",
		9 => x"e20bf8a3_d313d9ee_7a40812b_f3c7d74e_a00aca42_c009c2df_e4cd481b_f45bf3ef",
		10 => x"3f3bdbcf_e95befdf_792f280d_eb53c8cf_0b838245_d543e91b_0a83ae6b_dbebfbff",
		11 => x"f79f7aab_75d907bf_f048098a_706300ff_df8bd1db_f881814f_f1d3f4bf_faff657f",
		12 => x"f52ffea7_c4c0c174_51c36809_dec3fb04_fb179b25_81d55194_5ff9818f_fddff7f7",
		13 => x"45510044_e3319b1b_54010100_c016d1fd_df034b22_4001d001_db75d146_fb7fd5ff",
		14 => x"a8feaaeb_ea22ceaa_bc818813_9a0988bd_dcc63597_9040d94d_e758de31_d77ffbdf",
		15 => x"f34a7267_c002c322_de60c2fd_d52f61bf_d286e0c2_510146c9_d718f382_fbd7def7",
		16 => x"b70ee306_e347da6f_b38681d2_b021e233_c7459014_c004418d_db39511b_d24bbf24",
		17 => x"ffefe29f_e3812289_9a81588b_6349e0af_d79140a7_8103240c_31f9d51b_31917500",
		18 => x"ffffc200_f987f100_f1dad0d3_f48be9ff_dfd1138e_d101416f_db4df1ef_f503ffad",
		19 => x"fbcffbfb_d893b18e_fb82a09a_f98bb8ae_f72f604f_1103d4f7_75d7c3df_04c0c98e",
		20 => x"fffb79bb_f7adff8b_e1e490c6_b9c7999f_30c50b83_0040bb13_d25f6ddf_d0d8faba",
		21 => x"b8fbfc1f_9a331430_ecfdff36_ff7e2c00_fbbfffbf_bdffde5b_7bfffffe_fefffc5f",
		22 => x"dfcf0bcb_da030a1f_c2029080_d289a923_c0c7c1bd_48422102_889ec6df_ebdfe9ab",
		23 => x"fd2fc25b_ce2b8a42_7a3b8009_f90dc057_d2c288ca_150182ec_9cc2927f_d137d4ff",
		24 => x"ab3b820b_a24b8acb_fb83d081_abc5a081_edb10197_d3fa0a5d_50909990_fe407f54",
		25 => x"cfbd208f_70cc00c0_e78889a9_c18270fc_dbd18955_e019865f_d1e988d6_eb71a1e5",
		26 => x"b7dbf9d9_e9089cbd_9f41ca84_d040f09e_3391d15b_dc0c55f9_33515995_b989d9af",
		27 => x"7147fbee_d841e2bb_70400043_01024047_51cf91d5_48018246_f00fcb0b_f2dfeaef",
		28 => x"fbbb9883_6384388b_fbeb2043_3040a1e0_fd4f9172_cf01b1bf_fdfa139f_c024dbec",
		29 => x"d593e582_11628000_8900230b_cb8b938f_f5079212_1141a0c0_c1eb9191_f173f3f7",
		30 => x"babafeff_fffeffff_fffcffee_fffffdff_99f8fff7_ffffffff_9ddffff7_faeecff7",
		31 => x"2d2f2c3f_cb11d2fb_f3000010_fc01f771_ff059009_0540c0df_f5100014_f97abd74",
		32 => x"e25b7821_ed09b0e0_0013802b_638bd313_6052d019_53104052_440b81c7_f357d1bf",
		33 => x"0f6b636f_1a23ea8f_aa03c002_024cb3b3_8d89043f_39028127_ff0f2213_7717c62b",
		34 => x"e29fcb8a_f921834f_ab018063_2981c1ab_081a404e_45c589c7_ef5153df_605489ef",
		35 => x"fee2e234_b0afba94_ea5b8033_ca23a08b_6ebcb042_910f10cd_e8ca0113_e47ffbfb",
		36 => x"8ab8b988_f2a89abe_f90980aa_e392f89d_d74c82d2_d10b88a1_d396b31f_faeef7df",
		37 => x"ffffebd5_ff099250_cb8ba18b_f30bd295_f906b273_801992df_f21ed28d_f96ffb57",
		38 => x"0dbff5fb_a8ff8ccf_8aac3f75_3db7dfae_1b7dfff9_bffeaeaf_20a0377c_1032ea94",
		39 => x"4def5a9b_7b411d5b_09aad088_584b5546_ff09d180_9001dad7_3a92d82f_5d3fd7ff",
		40 => x"f072d8ef_080818aa_e8038c0a_648be1fa_5a10d296_0006c856_c21f000d_d2dfecff",
		41 => x"f5cfb3cb_fb81e8a5_f0808080_7311f4ef_424a1542_c2018c0a_04cba0d7_e0d7ab22",
		42 => x"aa02fa26_a9a7e863_9ebb8412_d18bdcfa_ec27101a_87006100_fa032903_d101f77f",
		43 => x"ab0c008d_82412f8d_81009880_d80091ad_1f41915d_dc014455_55600083_209c08dc",
		44 => x"ff0f79ab_fb4979bb_f320c201_7b0e4c57_fda90159_73835893_ff51c511_087f0e73",
		45 => x"d5bf44ff_e7feffff_0dc6fe63_2773ffdb_c6e2a6a0_bfff7e78_e662eee2_fbafeffb",
		46 => x"7313c203_a343631f_52230023_b3421345_fb0724c6_000080af_fd71921f_f3cb662f",
		47 => x"eefbeccb_a40020f6_da804c80_6730a1a7_dd05ca8d_e01d82de_db45d919_60e480f4",
		48 => x"0f87400f_1c525cff_48884c05_aa90ccb9_5fb70453_990d939f_57cb86df_7e03c9bb",
		49 => x"f202e312_f01830c0_f84a4880_d009b872_e218a204_0048517a_c850c1de_fa43db6f",
		50 => x"d38dc921_d2899080_cb012154_b90cb8b3_95839103_10839810_1a115152_c367a733",
		51 => x"a8dee07f_2a9a083e_88cac889_f8c5a8b1_84e58443_0504c017_3893bb95_d0d518dd",
		52 => x"8f1d7465_4809e9ff_faa3008f_b300b0bd_fb57314b_9100407f_fb91829a_f307f3d7",
		53 => x"f6fbffdf_edffffff_eefbff7f_fefff74f_f062ffee_efeffefb_d2f7ffef_ffffffff",
		54 => x"d59fe4b6_51ab4150_410780c0_dbd3e3e3_d5c5d052_91411110_cc4a612b_ff7ff3e3",
		55 => x"fbce41cb_fb0a5adb_d0880cac_42c80aef_ff8198b1_55c09437_d543e583_51d30bff",
		56 => x"fbcfdaaa_e581c240_4848c108_f201d023_f643f154_b111c3e6_f091d2df_eb5eeb0e",
		57 => x"8888deab_f182998b_ff024202_b40a8b83_dd04d191_d013b011_dc07131c_f910811f",
		58 => x"ebef336f_139c79d9_a638220f_106000c4_55c70031_35851085_dd47c10f_e4840254",
		59 => x"e4feead4_6137a000_c88e80a9_f983e343_c00388c0_0501014a_c1039800_e94fffdf",
		60 => x"9007d90b_930300ab_a3241014_e08981ae_0032c00c_44101013_f2530051_fb5ff3db",
		61 => x"45d5914d_81049284_29018093_724cc3b1_d5575187_80d7194e_715045d5_fb11eda0",
		62 => x"bf9c4434_aa3c4bfc_bfcb8028_f84b88f5_ff5c409f_8002981b_f7d2d227_f38cfb75",
		63 => x"e7bbfb9f_c342bf8b_9b426800_e2a18d8f_c0308103_500e41ba_e8934285_eeffc6ff",
		64 => x"dbcbe0c1_1b035484_1a01000a_3a279087_3b4bd480_d0418191_1d891008_f34fd7b1",
		65 => x"002bb28a_2b8122ab_32020084_c01f88ff_3c905004_4041201a_590b90c5_d95ffcff",
		66 => x"d78ba2c6_4309002e_051a0002_600ba0ba_f741990f_d2000a12_0293934b_f54ba9a7",
		67 => x"28efc99f_2e01a298_008a8088_b883a2b0_39d3301d_11018017_a33c5100_d107d2b9",
		68 => x"dd2b88fd_c3010001_e880c080_f089c480_f5c511ad_06019116_f429c1d8_9211f131",
		69 => x"d9cfc14b_e308ba00_53008088_6003d131_ce53c00b_c004000e_a3519183_63efaa0e",
		70 => x"8abbaadf_c4228088_a8839181_c009c9ba_1b55c441_810041cb_1ccf0111_0683a1bd",
		71 => x"f5fffff3_f7bff770_fdfffffd_f6fff777_fdff5f7f_f7fffe34_6ee7efe7_ffffff57",
		72 => x"bbc8ba1f_de059bab_dd0091fc_8d088a3b_23911589_1d093691_9b5115d7_f918fbbf",
		73 => x"ff60aa8b_f014c3dd_db89a203_f181d124_2202488f_a088810f_5ad7c1a3_40b644de",
		74 => x"afaba80a_ef9a8b9f_81080000_18238a9b_ff0fc00b_00000053_ff01d005_d094caf0",
		75 => x"fb7f6063_628a88bf_a8aa08c2_a209f3e7_a7842200_808850d7_e0c690c8_d83a99b7",
		76 => x"1f2b0838_aa0b09fd_d902020a_5bc3f0af_9dddd4d9_a2118913_d7d5319e_75c8bbdc",
		77 => x"5052cb7a_4402c048_f20a8800_f9593304_0282b01a_08085010_f109c1f8_fdd5d36e",
		78 => x"0ffb239b_3a00001b_ab71c21b_712a0040_0f05030f_d511513b_0252d515_03640972",
		79 => x"fb834a8e_e701a243_8001a080_80008087_c20c8885_65054d04_46ddc247_ef8bcfaf",
		80 => x"ffdfefce_fffff7aa_ffffbfef_fffdffff_efffffee_fffdefef_fffffefe_ffdfffff",
		81 => x"d0b5f0e1_510244d0_c11b8497_ec01c1ba_279b54f0_cb33d1c0_02a38013_f69ff9d3",
		82 => x"5e5b424c_d2081680_5a948019_481ac99e_5104004a_1106649a_dd134333_f3cfd2fb",
		83 => x"f101ab23_d390aa8b_fb000221_f903a3ed_40401805_00011107_fa078007_f28280db",
		84 => x"afe79bab_9d81329b_e500208a_33403080_37dd2181_84004153_b0ee42c5_62040274",
		85 => x"c2cf88a3_e3009601_498b0082_f10fb137_c40f535a_9400a384_ead28085_e377f6df",
		86 => x"2b88288b_6000c098_e8018088_d063da95_5dc852c1_5100009b_d0140015_d0449854",
		87 => x"efd96af7_f8831b42_4a008004_0a0050a1_d5920000_80018107_c1440c00_cd0d422f",
		88 => x"9633efbf_79baad20_fe7fef7d_fffe1c34_bfbfbf7f_beeef9fd_fff7bffd_9dfbfdfd",
		89 => x"44c5c5ff_5755d445_6de4fff6_ed76f7f7_dcedffff_feeec5f5_d6e4ffff_f3fbf7f3",
		90 => x"5b2d005c_1080388b_d0800008_119808ca_59111041_0004401d_51539190_11501232",
		91 => x"f2da44a7_801042ce_db0b0088_80050088_70184012_80001052_d5837190_e298e2fe",
		92 => x"c10f524f_5a402145_c0800880_13c04099_c011c001_80000951_91004081_d181ffef",
		93 => x"bb33e1af_400590ba_10840880_f2888b56_f580d100_10000044_e0844844_51518652",
		94 => x"af3b242f_7fff6f5f_fc752d7f_3b7ff5f5_ed6f25af_effe64bf_fd309c95_fe7efef5",
		95 => x"0a8b0849_0281280a_e9808080_48009029_04001147_01003101_52572213_4808b59a",
		96 => x"3203dc2b_b8015208_62882082_c202b208_49110018_49048104_53038081_f309984d",
		97 => x"d5a7a0cc_80818101_d08a2000_1312aa90_c7010041_9104408f_93808081_0307b110",
		98 => x"c0bcdf75_eeff77de_457fff7f_e5ffff46_b2c2effe_f6efdefe_d875fefe_eedfdee3",
		99 => x"48ac0141_000002c9_20000080_4a004088_d1052040_00004015_510600d8_5300c0d0",
		100 => x"2d89ebcf_763f4f3f_1f2dff30_9b1eeba9_1babb678_efefffb3_12a00b00_5d00e203",
		101 => x"6231f75b_fc7df497_85355f75_86cfa644_162c7f67_eeffae6e_d7afae2a_c7fef64a",
		102 => x"453fc567_ba7cf6af_ccdeec6c_ccaec447_0fffceff_7efefecb_5eccfeff_491e84f3",
		103 => x"f3d33e7b_5e773955_55777f7f_77fdfd50_9212ffef_f2fffee7_66eefe7e_5ffd0fab",
		104 => x"6bcf460b_80400009_12000000_00008388_a900d003_00000010_d0008105_5080055c",
		105 => x"0a9b800a_01830822_81008003_02020080_10070085_05008808_d0004000_814200a5",
		others => x"00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000");
	constant plut : byte_memory := (
		0 => x"01",
		1 => x"00",
		2 => x"01",
		3 => x"01",
		4 => x"00",
		5 => x"03",
		6 => x"03",
		7 => x"00",
		8 => x"00",
		9 => x"02",
		10 => x"00",
		11 => x"03",
		12 => x"04",
		13 => x"05",
		14 => x"05",
		15 => x"00",
		16 => x"04",
		17 => x"00",
		18 => x"00",
		19 => x"03",
		20 => x"03",
		21 => x"03",
		22 => x"00",
		23 => x"02",
		24 => x"00",
		25 => x"03",
		26 => x"00",
		27 => x"01",
		28 => x"00",
		29 => x"01",
		30 => x"01",
		31 => x"00",
		32 => x"00",
		33 => x"01",
		34 => x"01",
		35 => x"00",
		36 => x"01",
		37 => x"00",
		38 => x"01",
		39 => x"01",
		40 => x"00",
		41 => x"00",
		42 => x"01",
		43 => x"00",
		44 => x"00",
		45 => x"01",
		46 => x"00",
		47 => x"01",
		48 => x"01",
		49 => x"00",
		50 => x"00",
		51 => x"01",
		52 => x"01",
		53 => x"00",
		54 => x"01",
		55 => x"00",
		56 => x"01",
		57 => x"01",
		58 => x"00",
		59 => x"00",
		60 => x"01",
		61 => x"01",
		62 => x"00",
		63 => x"01",
		64 => x"00",
		65 => x"01",
		66 => x"01",
		67 => x"00",
		68 => x"00",
		69 => x"01",
		70 => x"00",
		71 => x"00",
		72 => x"01",
		73 => x"00",
		74 => x"01",
		75 => x"01",
		76 => x"00",
		77 => x"00",
		78 => x"01",
		79 => x"00",
		80 => x"00",
		81 => x"01",
		82 => x"00",
		83 => x"01",
		84 => x"01",
		85 => x"00",
		86 => x"00",
		87 => x"01",
		88 => x"01",
		89 => x"00",
		90 => x"01",
		91 => x"00",
		92 => x"01",
		93 => x"01",
		94 => x"00",
		95 => x"00",
		96 => x"01",
		97 => x"01",
		98 => x"00",
		99 => x"04",
		100 => x"04",
		101 => x"04",
		102 => x"00",
		103 => x"05",
		104 => x"01",
		105 => x"03",
		others => x"00");
	constant flut : byte_memory := (
		0 => x"ff",
		1 => x"ff",
		2 => x"00",
		3 => x"00",
		4 => x"fd",
		5 => x"00",
		6 => x"00",
		7 => x"fe",
		8 => x"fe",
		9 => x"00",
		10 => x"fa",
		11 => x"fd",
		12 => x"00",
		13 => x"00",
		14 => x"00",
		15 => x"fc",
		16 => x"00",
		17 => x"fb",
		18 => x"fc",
		19 => x"00",
		20 => x"00",
		21 => x"ff",
		22 => x"fc",
		23 => x"00",
		24 => x"fc",
		25 => x"00",
		26 => x"ff",
		27 => x"00",
		28 => x"ff",
		29 => x"00",
		30 => x"00",
		31 => x"ff",
		32 => x"ff",
		33 => x"00",
		34 => x"00",
		35 => x"ff",
		36 => x"00",
		37 => x"ff",
		38 => x"00",
		39 => x"00",
		40 => x"ff",
		41 => x"ff",
		42 => x"00",
		43 => x"ff",
		44 => x"ff",
		45 => x"00",
		46 => x"ff",
		47 => x"00",
		48 => x"00",
		49 => x"ff",
		50 => x"ff",
		51 => x"00",
		52 => x"00",
		53 => x"ff",
		54 => x"00",
		55 => x"ff",
		56 => x"00",
		57 => x"00",
		58 => x"ff",
		59 => x"ff",
		60 => x"00",
		61 => x"00",
		62 => x"ff",
		63 => x"00",
		64 => x"ff",
		65 => x"00",
		66 => x"00",
		67 => x"ff",
		68 => x"ff",
		69 => x"00",
		70 => x"ff",
		71 => x"ff",
		72 => x"00",
		73 => x"ff",
		74 => x"00",
		75 => x"00",
		76 => x"ff",
		77 => x"ff",
		78 => x"00",
		79 => x"ff",
		80 => x"ff",
		81 => x"00",
		82 => x"ff",
		83 => x"00",
		84 => x"00",
		85 => x"ff",
		86 => x"ff",
		87 => x"00",
		88 => x"00",
		89 => x"ff",
		90 => x"00",
		91 => x"ff",
		92 => x"00",
		93 => x"00",
		94 => x"ff",
		95 => x"ff",
		96 => x"00",
		97 => x"00",
		98 => x"fd",
		99 => x"00",
		100 => x"00",
		101 => x"00",
		102 => x"fc",
		103 => x"00",
		104 => x"fc",
		105 => x"00",
		others => x"00");
end lut_pkg;
