XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���`:��w�#2"Lܓr��m�f�"=���^�D'��UgQ���67	�B\�O�ϐ��_(ǜB��,��2B���Kݎt��&\�7�(r�L�a%�Z��G
c�k͝�;8\�Z���"�ꭁ���m�P��_ʧZuG�o�����(�c��H�+�c����z�l$�v��c�F�b�C�q�Jb鼷�)��t�=�J��nc��+����R���� WHt�vA �ζO��$�H@@�~*L�^�/Qg)�����V���I�Y���Wźˬk-Z�&^����x���m��s`2Q>��~���@�RѣZpL�.�"�^/�t	o��}�0�xa�l�<���m���wl�miY>�.�I��;�v���9ە�[�KJ��~��wޞu�P.�#�e�lԵx��=����Z�;,M��Z���)w�l�Bh�����8M�K���NDa�J�( U��4�\�xO��	�r�m��������AN���: �s}$��n��b�iĦ+���%�V�>R�Q��ZW�m��wm��ɓS�:�0ƼsI���e�-��*�[O*���;���%����G�V��]���r5+X��a�+�ȧW �L�%m	g�?_ɖ�G��FNL� �K1�Ff����r���߫=�Yl�+s��he�~c
J��E�	D[x����}4uP�ύ>iJ	*)|��y�m-��u&iIn�bk��?�"[؋��k�_џ��U��#�W�ֵl�(���D�H��R!T�w;��N��*o�XlxVHYEB     400     190e/����Q�-�BK%�X_:(��=|��g�i,�c����=�`"#���{x��y��$�m���o~�|�"Cr���i�$ۭ%���a��f����?��w�i��@b�m�4tq��˜�^��ш��Ha�Z����Dnc\[S7T�@����Lj�[V��(�[�P�y�BJ���uh�����Y��?�M�D#.�0��M7�ޥV��>c`˳�#p[?Feu݇.����`X`��|M��.�HeE�?����۪�-�l�Y@kn���PӒd��q�0�n�V G���ԗ��n�\���.;�����f�=}��$����c���q=��1U�vr�̛�B��ߢ�lJ��V%K9�o��7��y�%�Rϲ�zm�&�C]0M������a׋g���ZXlxVHYEB      3f      50��%kgU�?W4%O�B���OͰW�ux�X!UH&O�R>]_C�
�����-xf�RĀNRoٞ�[5%���j�)�g�F<�