`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45824)
`protect data_block
/zVlpVR+6hNk5sBKmCovvrX9WjUO2VSec3heVjxkrys/pbiRYdIkYgTgROagiuHA1r6wjR5AO4FR
+IxWVjkly7hdT8LBuC3WtoKG0/EwVMnOZLkNs9D1+24IGqRNpYZm8nL5EU3oib3XRgWiuG+zjXZK
30w50CHA4+kRXJrZ/A3RRYb4plrxB+b4rP+9pZhA89E9w13OlNFY9zgbJfN/1AXVBUq8MZBczI/V
rhTK2QkBvjAJ2++AIZxfq39JgQ5Nm7Qwy28OCJWuampXF5MPYvsaRQDdTNAEfbis3prS7XjSSpKo
lOdRenU6Y9O/mUuGjUjQ68gS/EhILdh9WM2ueAcE6HAgiNjzuSPkoV94Wr+SIEeY75pIbafsTPKA
x04Moa5fRQz8/gW88Y3+NrzalDFagCv1JxQ1+jOXz6M4UkrxrWAEbKdve1LUtBFF0IgGVwYW8hqS
KHMvwFr+An4u97y8QvDa3KUp+nSFUN5t2rnwIpnpIPzaN0g/kOZWJHxSg/a4R/5S6zGC1bcZotQX
V5vfvQOBnuE94hMN9orqSHZ3ikz/m6FJA2gV6D5PiKV32zIrj1d9IrWE7Z+k7P3jgKZ34udMi+J2
DDX0ID2eBwQ9n6thfS0BaHOCjAqSPdL+pksm+coJB8xbEIZjE3uU9VDPo0mqEAEQvucGku0Uxtn0
84EW/WhIKPD6eFY8WtOWMHslxIznKE3PDxq8HBp4yOdA+DuQ1W5ZxElyzVSQ6u75SRheoiErNdTf
4sbDxMiV3lhINu23A2ntYsnTgD1ENygolP746GXEReZM12ERNX2nHCqsrBTcbTgdiYV33t2iG7+A
0seidVs6X3QGLbxID9t/OOpe8Ys5APQHjGoj0eQq728NFyM23hEnmGMkLaOTL7LSlsJELHcIaNgU
R8Fge0kVRv8Ckqi0PkgHjsCi4OKfUFw/T9ZXopOy8+PS/xA8ruyXNWTVHEkyCKgRVHNRhtptwam1
0wTdW53S3RMI3SpKW8b7Z+L8mrDRLDLKpoP2hBteo4EAukbj7dSjdy7Mep1l+TS0CA0CkZJPttlW
UrlfTsaHE3S+P9gaGz/6xzZmcwm5VI8RBFGuHDDjrdYVuzB0Z04OLwibL6RPjJHGqKwBT/bX/etO
dv/cE0C+v4lQQkRj6AnpGmWZTnHbIeq95ehlfwfGDtD8DT7dOF4tUlV9vuvCflNeNj0HC6GYgweU
1kcfYeWu36dZQ0Ehx6QhQggPlrdP7iA7gUT+BbZ6jDez87tjvgYE9fL+n9bOh0n3KRinPqeJZy5a
+tCLVO4t3QiHu5Vtk8nvGkpeLQL0ELGxXOK6LTXsseUNIz+JT349vL7b3SPIxmciTaQaw6wTdKuO
dWTwc37VyUg50HWx/PH0apyVQWucYcP1+73zN1VVqPUEDi/R/kGAiSwRifFzcXq+ljKv8nQY92Z5
U2tyDUkZSw8+KLVadaTbgVJ2wVa9t8dQLq6nyvmvuruCqSX17+1fLWzxdpXCq7iYLLgwBFNgklaK
/EoOZWTi5yWoi0qp4PSZH5cND3aXQXx+oTntK2NvHy9njX4eDJoyaK2nHnUlq5gQ7f2AWKSLk2Ca
vQUXsErv2Buipwq2T3hjO0Gzm0rELyC+4QNVGuTpfS72hsq4B+MgRXWWpYo0iJBhszhV6+vz+Jfi
E5c7IdGtPCraL/J+0xRCffM23dhawghYE7/kckda520OMz7K2f7PoVQsw/aGN76+sJpKx9IPNOvQ
LUjpXJ08wXiJwuEJOScZ2nobHYX6XSvdkuorbRwzmabnyxmCqaN1Y/spvMCBl00UY3dHq1emENsv
tHQb8TapI50YaEQ+yKyJcPyL8qedFA9ICoGeBKrMNqrHQFuD17xrf3ysIY0DaMVq1ZLsbKrFD4Ke
F707oaxB+QtMgnilVKMPs6ih2Udc016RrcPpav/dEeKjqcmOB7n3hM8dKKrwV08ieYa04ZFXsiI+
jx/LWOh9oNbhRM1C+41jtenp/LUHNBdwZEoKI0v9kG5r0aPQBAzlae8vc5qcJekGZTPVKoyE6QSf
8wbAWLKHkCnzDkQsoBSqiyuiVjIk8fXTW6aILIPollMHItjgcMKcOUKbPSAxv4sSZ58mj7PGX5Vd
jgKbpFHRiFFfwgGAwvIYefBsAM3mQkqQgdZotUcGxAoPlJRVjj4Pp6hAyJlrq/ZHgHfvODPlv5KR
s8MDpolgYlkGcw9SxG2i8/+04U5/sJ7AOlOpOBaqoh7bjKk+6FMDfztJmg9a/ouw31HKR4RpDE0D
/QoQA1tqwhHzjNQOk1BWP9snU0ZimWHj9oXQzW4ieJSNpS3bnF3HLZuSysPhuQJXD7d5THfrzT1y
9sCK4v4SKcLYlOa53/R0VrQOKnvnJzR0mBd35cRTp/J3Z/I7Px9UX44w31NkyJwiEE9xOrjylPxW
K8BjrZ8GHoLwYLYuU4oMvsfHFAt6A6zEFADULPkXqLbUHO1fKDbtB+4cunpJ06MkonfV+rFgIBo8
oQmPIOqTNzxd+Sq2/iRtOQETa/aIUbo50AeLW8N9RBFWA0T5/vVG+PhQFivEJsEVY7DMR3KQLcMa
rP20I5IxZOkjF69Q6GE7hvJ7yKtjEU1RwOdUWY6uoHqSa47vfCxWhNOjmep300OBdC3zYIXmUYMS
3Sn56IeMPDXHmFgw22O1Ltrda1V4sVxC3dukDJFaC7ZO4UcxHPQTMsetLJqfvpEVSBlWYh/qNAFk
9pNovY8DZlPQrBlbxidC3q82sAfO+/BMt81ZluLydMAkDfDKZL8hikKz5Mmlq2+OTNu0jKoXZT3f
wOYPhGAsZ+GJcYTO1XtYPIvtMLdTFjq3CU0roUZAkZa1EO9LQgiJIdz8DAisIfaVPYM9gFJPzYsI
Fu8H0Jw3rGz3l5GOMLGYTWtJNbDrbPCIeIy6n4w1zVUyT3LuWLA8Z4/ArvVVe/z/qXrSaNVsKHhB
6zGUX1RucYaPFImVJXnKK/9hrjbjorn8e0ldAMaY4Ub1wynnbNWrAjIfWGvJfD5KJBXZS89uRFPd
mkQPaiz8s16NH/gbuTNgqDdWuOd4FybhE8OPmSYzqpOoBT/zFAZLFGfnCjmoP/8pU1aSZWnxlNYb
AWpPdOafWuGzPXR8PTpwKthxgh4tpFMMiEO+OCrG6VlKZD8dhsOFkDUk/OHG+w8hUmJeEsRxz0mP
yHUQz/oEoEWvAykhxHuPbu7wqtm9iO4n46RsoXK48GYvimyUGjPGy/aI9r5d5JkQANsVtquEAvjp
iKDhjQi5DKUbMunRcEKTho21H4IQRANHOfu4VDr1VjmBysosUfeZ1fA84HuMZK/JKxspbxurWUm/
howBsEUZccaNzj+Wn6VLcHQqrY/96SwiD8t+0hJgHeVbosThT6ob/PrOrOONvXNkWFmuufst8RNS
7NQZezRYvnYKUeYX8ZR0K5HVgEM1g4H4Iz1zKB8sCkp/CkPgOrVpg2DSxMaMn6D3NmLQlVnaGiBJ
7yjqc/+P0iTfDXzIJbVtkj7iEvIbFsKLjR2JPH66N71IuN/oRiok8XaGab282wPO+NsVGwqn3oTq
B+p4cPbTecd69z4yCLuCasXn5q5gOAHkAZXPuE/WsQjve63DB/ZKhzHyiAbCHO0pXDiUvvF2JjDW
9Cc8xbyKX50WLd6JfZxC5rf90wzF0GJqA/Mg1EdGBRUw6H7Nlf2J5dXDjpHBoaw7AzYAmmFaXoyk
f6K5sOdn8ZorsTOwAFIb6KVkiEIQQmUgvIgFPbJPdZov7S3XX9I0TYqkm1iPpYE7A9Tm5Tu/haeZ
vvc3xauoDg5fcv60FrpoFJLNAG8ZP77gP+6BCjjB0NJI+qdhhL9VSHY+uLMrp1OdjQsLqNOrAhdF
j+MdauQooHE02r9By3P3vlF+GF0cZrG2j8vaBY14vV8yKOM6LaG0lw1ktGwrE94305/zrEI59ish
DMJ9UKeyCQkinirAfK6aqrPmOzY0Fw0sinxwY9vm2sbjw+bG9G8SfaGracOec0yBOaW/3SJ0c711
GQLPt7wsxj2nO9lPNsJOGcb9RWKUUVl3ahJryEEt0mGQHyJ1ycwdvzMpFi5G5TZqY3zSE3s+JiFT
j/qGL0kciCogIzuQfwH9nctwwcmHwmyZJUSbVuUwjYFn2MWImXWyM3UeucweFWMfJcNrURqxzH8p
ZYyRY85BSQvZJWu9J2kuF/lc/sX4wV34CmwTbjpcoBJ/kxGDxIyMGh3d9gCov0uu13YGuLOp454N
cQ9R6MV17Yr1U8hcVdrXVwXR+sp15pzjLO3FpbkPhKRkgK6ipn8vYFEKMY/0IcOPPabUUxIyCn/g
S/md3H8qoqzychc8K2MBlOciRnT+iej5ViJoQupBBTmS8MDF8BoiLXHR7gda1KP6dcoE2tDZy/h1
+IJazOpaXhE/64M0h7zOgVoCNMnnA/YBmkZrm8Py+1/qSEkXd+j9bqa5lcLHJHclUuZ6BsmRhFo2
vlU2gzDvJGJsuD64YoLllCvjxS+ZWrE2CUBbx3QegSm/QbFRDqswxpDmEwEPtSoZqUbnowda/wWd
CNZ0w162rph4KBG4+zM1zEuALqnWfxY7mHNuFrOOl8dkrrao//2ANJ2ZngXErulym+fDAVzVSOgK
BKyvNS6rdVaZ5simrAWqtRNUZkZH/3DMHUesHzJcnT07HGXNWZGr1Vq80qB63qyKBehBgV7ZUT7L
hRQXaSTMEPdup1df13JdV9Lkzfn0O0DNSgQt8/5Ch3U9bO/MlzC9XypzGwy5X/PpyK2WP3wsB0Ep
HOIjKrp5iToRhlxvHQrmYT1siUWypyg/yCSQ2GtPsA2ah3eUf/xVJ5Yk/4PDeUOkbij9v300gSqg
5MdXE/Kgy9JO65FRMkV+mMkEmT0aSI3qDpRsBX6IVKLg0u10iFBn+FhHyC1q9mlkJhS0Dx8faxjw
uP7bIJCDalnjC+GZWWSMAuGONrZrI0mGOeOHOhjj4UQ0CPhYhyi9Nyl2FzuJ51vjkQiS8YjTC00X
irSqbVQMyPKNWI55v7QqEvHD4i3uHppxUqRqhJ/XtDW3mlnvU2uRQNCuyPS3q4bEat+fmTuJNQBe
PIsUmXgaODFdhZnOnlFrMFbS5W7wclgtpoDzcN22GIUcpqU83iNGZoz0xcuWdNIFdQaXA1CaIf12
JqYmLil1/KywkNlr/jpbB/OSR66MATMWrkjp/I0khchrkAKO4PRAaNJCJMzWclQgioMrCHxj89ob
yYPFAGMUWVUFbH+qRQ5Ko+6rMzTHqiSLZXVPEXV+KrlM5gcs/geuucA4/3YIbU4nrr0mlgyA+bZd
QyTspMa9fA9I5th93/UiRERSMuDMjpsJphA/S53qfpH+Nm5ekEGXRRKhyZ62jVpWBwYlAfRhHtbf
poO57vQEtfn6S/oRMZ2TaDC3urg0HRkwOqRC0zCXqsprS5hxd3xxyOyGaJupJDiJ8EJCkUF1HVeg
4HiSSF2MH61Jth2k2cY9axgP9ifTwx0v3OnlHDwp6csuKFlQqTTrO9uZ0kc9PsVYkAKICBajXoIa
aIiij2cdAkcpjmg4x8dS/JFeQlp+p0zSbsPRUnpY0DToAIE2mR+mTzfzlKCB2dYO5ZMu5YoXtH5s
jRamKItDBekiTKsiWBORN6APJEaYtFFk7KqhRif120edHpTddS0sZ/mmWmIYa24XJjXszwV764T6
JVWn5MqOdD97aOCAiT3bHVmGrZsGj74lKFKXavpeWV/uPEN2/dTmU3VlHI9p8yfi9voX51/hon5d
luCWdMu4HqmEfDK3VT19vnSFEjUgPsiB6y0FaxvzGXpkxusvQpeORlr6cb7oFoJsPTGcJz9bR3Cs
lkrl8jzguBtgAUoipyJCuN1u2pqXrGyIlhmNfrENimcGW3Ur8kp+hsE4l2VVUFubBgbPL2Zgw8Gh
OogEbIy8sPKz8s78/DWtOx1jv6YUT0WTw8KeYPJsMe6K7rdOPGb9bHD/EZhxlgbl/CoSVLD3AcpU
mBKq8tIdMWiFDNXb8l0Dh+05A8cbfElep83rbjrb+869yNYDZjIvtJ+qjhqeiWV5uVNU2QlbSZI9
+JiYO8DbRXo2a16IGefTppCfq6SevxQZX2mXpUzYeq5alJQHiWvaf94Gp8zyj4Uauu+XoC2CxWkj
ei0zE14auPyH5S0q9I6Q/Vf5KwfMIGsPR2zGUuml8I8uqXaVZq+lWxioXBFGyQC3EeJ7R5d6kRgT
nDKo0le7fJsIYefr8ejjGbOuApBPpV8wdVCrbafVRuUxzJegg9drmdb7ejSJuYjyg2BHAacbyPtA
ipq+b+omPWWg1O7eMbvnIuIg5z3hHCPoGMHpvtGpE7Zr6bcmT2pi3WVnKf8os8K272+BHvH9VkC7
9emdi2oxxv/Rjf6huVRHkweZq+NO1qiaLGE3eS8uxp3dahCsspDT3V9KSWWuL+JQMGS6ehDYqNA7
2bR2ODMDo3PLu3+ZepTr7fVc0S4lLHtu4Ak8O/E9hwhafa5dFN/nt6KAGLK0hi1ZzxarUBdPJ5Ev
SyS+O6JZoJWd/d85dbZ6W18s6NvBlIBVb3ZVE+y0tWMu/jrPvV2ogx2iP9aF1QqDQsC+1ld1LuOy
TGtfnzdtLROAz8Q3r1EJSMFuJlk5QqjfE0+L8RYvsVCJDpwrowvKEm6Zxrs1goOaY68RNzSiiZbg
bs59VDriYTm6VD6Im+jZp5K5iPyaln4CxzcrlgHDnFQ8traVIr9RPm5BOkp9AQ/UKzia/U5wZwat
zfteBiLBoNDGjBEPGy+UFwSsNKYZeL1bHvGHbaA6uuzoLeLl72J4yY2CpfP1kaBZn19bqQe0fkIq
LljNaUfmcXkvnB9Yykt++7b+h4rINmuC4HgwDVRVSy7VzwRgIjBm1wXkOBbI1GThXpTodIVRtp/w
qZR23+D2rRS2q91k5ZfjAak/h9MYkL4ghzrKdGhECZDdBrUf4RYoHRxm5kTIrDPNEXAtOHXa83hz
Za0Ycf4rI8M+VNM6jAZEXFXyvc2ZOvBwUMFl/JViVk7xk/ZD0pEa9kQQKPgl+NqIFOtA68rOfh5D
JG9lDtQnNaN6zg8BgId+djsquPKZJcO39EV+JJzAMqqfpQjE1VyW3S7tnUaWN+JKXTJK1Kd9wETR
jlDEi+HrPc/2AsGhxjGFVlvcjDCrF16uTTIXa+M9knP/fixaPSxQKdsJQLQZhVqStg0L1oe3OYVj
psiTD1tnv4cE9AVkpoQpfGNpCh1l10dUPvXp6Am18ABAnXIpFNtMSLFj6dUpGayzBa8omMcg6wf4
OQaSK28lvVj5AjRwW4riQVd8rhBaBXyqwvkv+oCFs1uR/Qtw78Ouak7diHcCxgflYCMPG7TFy/nf
0M3p0BvENfvu7QUxdtY1mbpeZj9Dabkb3SNLtxTlwY/lUMyL0tpQC/wa2Oko4l9rZQhhO5/bZaWH
p+wI5IYvmE5+UEr1OelrzPL3GSqUUWY5wY+RLKO2hPfGYWSJSbEOfJY2bYVaGPpDjLoqx0LED3Um
qvPgU09i75/jzXBP3dCbueNL/Q8eCZLFAZ/2evayH/lfGUT4xvP8Hjkgbmp8eXugCFWpV9EXceL8
yTTMw6kWuGrHMh/5IbEbSM8tSMfWRxbaw0nvIGqkAxP4mcW6QQ21Q/uNtUDMV9X6Sxa+Ixaqx1QV
RIomVHsMQp74fXl9AY6W3+B4V07bjEX+cbFIeo0Erhl/IHYv7tw1aIghgexGT1JpVhaWWWSeYYBx
Ptx1RD6NthXRCDhYr/hBEqDSGt/p7hNiOpr8vmkz6n9itnEA6/8vASClQs71ZLbd0beN2+Stn8Ca
lne1DNIlluamnGn9zav1g9zsVQTM89hQKcCneMEYqOYDQ9+OhdA0aul1zYUlt1NnhqLizM4ZZouS
RibK+Bxvb/axbYS+Zw91de6Y9mR8HOM0fmLdBRTL7fUXbCnT8uf7ATcYw9RbraxHl+nMne3+AT4O
POkP7wNBx+VpuAwHI6Y59zadBByTHZ0iey/pavTmVvdW1762QwXcHAEymlv8FcbFrvcnktGVd9Vf
oRrYq8XdqTK/ZVlVhVzrierVxSpWCHXsMIoY1yHSWec/s5b+zHHDivi333lOsi1+omcRAhjIKi3y
IXVy/ifOJErldRYu5cAX2EQW4oOMyUExK5jN+aVYIaJ/Gwwl+1rrcC4j+vTnYZB9x8fnghv8/REq
TSVN9ca7O7m/Ndn7nTiT9CuMqb5/NsFM9mLXtjfStvEusG9L9z95NVY0BxGgultBFJLgLhyn60M2
B5fCCTL/pLHxM7uZqI79pgzZTBdzI4lYtyulPDRIuYOW8mbJf6rrDMY9MCwUKlG/oa1qpW9QEi7B
oxVf7sH5fZcXpKWVq2Tp2Zar1vTfYNruwDBcrTRU8xh9PcWo8apfl/RPRgYCfhKVbSB3fBEcXFq+
3Vb43iA5wZZn+qE2jBfoqQfZv+/UA5/zcUtB+m/w0J6QLCcb0cW6uvCXXacxVwCP+nf9Yyusj+ze
VwwHYSSp8ixxZdODM6m4tgIhDImZkNBY9sBlT+wxHVhKVic88blsdg837Te6xApZtXIGo5C66Xmb
/vs6tM/XA9UpuBTKWwgATcQgKz8fzpvdNRqSYKSsTmqCIfas6yLQLuge0Fet+VD/I9tDpmgyAPN4
bByJ2zk6GWA0cVGhg6zZdA+G4HrlWyhKBUClQN24Rb6KGK7nDFDStNmqElZCr1jCZhe3/1tJQQuE
krI4jovXamDciR/9p8HC7c6jgWjm0x7jKcWS9ep11FBhnFiClMjDhj2UGJ9TIPE8SICbCcBLhMAm
DeHkQHoTewpxtrsvY0g85VRqbFPDs5L8us1N/ev+SarGHBPna9PzrGrMNf70fWpV+jFI/qNF/mPT
EKghyRwIKe3I9JD+u9QnZNJ3nrp44nVt/pwBKJw7i8WQpyFLZcXN11HFLzyXMRMfBvG2HGnCFcOE
llvaQpgIU1aC7IkyGUIgz4ky6DcayfxEPQS8lflf26B48PbwxCwKDd845f26Lc0zi1dflZb9fV/t
QTvBv2AXRDqnBQDysIDSuhBHwPXuHssxOoyBAudfDRi7E7aDlvaKpk2VueQD5TeuSZrOaJ64bV5X
QDYPw+CJYUXM2CJe2OQsNNLjBfTtEeC5STmqcH3U81kPjmDZsQWKpncq5ZpCJQX/Ea6DcWf0sjDB
lRozzKokU5IjUN5WKC2zegC2tK2gQbR46T/3VFu/17P/tNH2Z2VIjyQHjGiqSs4w1TUiSpfgmajw
mxsoOwaTTumjuZv3hqdqt53jD1GHlzVoD238cSqXq/DRuVWGsCSNwq47SngtP9wW9yH5eisjgafF
DbA+zx5zOUju3zVApxMT8QQd/F0p9roBm7+8ONn4LKAW6OUOuaEGofr+ofeAnT7oZieAjAgJYT4h
1S+3sMVAiI0+MXoZVwCta705G699TL4r6hgNvjY0l/blDdpv2QFRdjw/HhCcjtFcRFjcpge+ju6C
OVL8rC45rTXGxRcd7RJDgu2oTXANrsaT8iwnidAmGemBBywYfE0hWc5oMLrly/lfVfFIJScWejH1
rekAP8k3oRSkZlzGC3gtvxdXyY5Vu562LT3i3QRcVGmp82JHFmfKS7pF1MJ40+j3z0ZQtKY/dSwW
6iMc+MH0+LQRhEfXU5UpCE94G6i7mUJyv8ge1NncobqscDTlXWCkhDfVyMLJRneRY93zal7aL5po
55zP7RYrkb2nTxYC95EnC1O5GnDp6+TU9tkDB6y7DCapEljVVYbzxhwUWfXrQxQLpN6hbz8M7DNj
/r/C9wvVa12Ahgq8w4+u6JT3SoVA2tG5SzaZKsf0VC7s/hzW2y+apoBueqqzV8bOF3Aimydoe5mt
xUMWVsKlXOnwToo56SDojfflAlq0bkkogVzWmjKfvzNWDiMVYIGWLmJwLdIbVuYFsRxneTO7OqC9
8CNM/Zifsmsj+80hgu29XGTfsz821HK8iw9jCAYEClt8/peHYX/xeq0rqhcKYEvYc8qu8d1TS6Ei
9spAG+xAX7v3/jAhJ85zLmvr7jt/wTLvJ0S5hD2DYnTG46JtkYE4DktcOXEUaOvTymE5a6vvorHR
/j6bMbCc0TZ6Jn52Pk7xCIgM5KD9MPSYXm3gKpWYovo/uFoM7ukiXxnX9EVRPaxMbayS5F7mdSbZ
jHPFt4VLqh3sDV8xraycTn0ECAmWqtzKsCsLx6VBdveSSrbqDPIPIz5F79fCGCtOGE1IVB1heGZJ
U1YejA+AAwo5mvSn4rZxr+XTxV/2y55B3LSPzmnXd+n6zxAJM++8TIe244s7nVSuCG0tspfGdZ3u
m/FJcXT6MLj2KoIvWK03dU06N64DEBSu47VRzyiwRHdFR2jdFWtheeFYAWwJKtssyFdfdpmbCkyA
vt/kFH7BS5iu5fZ2OHRxu/LFbLdVCSwDqiP9oZ3J4kmoDu3shB3ieGnXPWPhQup++1UzmHjxL3Pi
LYkVjhHJGhAo9UKcEOa6Gp20A5tJOvBLxpX8r2X7mkS00fmcucm3l4mhzpujpQtY9hGIZfU5IV6x
k2CDNaOC7fi/JlYandmBg8Yuu+nyIkfYj4tNzjlCqnaeuR8y8rLrH5L3YnPL5NtTe37Mjsaic5MS
1+/Q1j1ps6UhFYVgR3S7CL1N+n9blBAOji0Bs7RccuqaYV7BZvOgRWc9WUG1k4/CQr7bJLxnytbw
r2AqDIqiXYEcNYIMWrF7fdyiDhqUN5re0Q6FgF14z2Eedg1SH3r9wFhJlddvd3gTdKeZkGRHZWaH
OMVcpd0YJ9V0biQ+cErOKljhSp2Qa/aq5NUE5P3lFiaP86yFBfiU2HYmn67ldoFHrRQlqKaT3vET
bbm6cGyQGuXokucho/+jPyqgJ/IRxgVPTSCHn0QYiN30R3KOn7t8K0o8g+jw6SrbzS6hZQoJDjop
KKFsQrpJ1NxjygPeFtTKhtmZXVA2T5Pw/zF269ktjm3lhLsd9P5+0dwAzq+DjXIx2/1xjz1mvNVV
mJaR/3dJ9qLyigjjwepNAT1QKlz5pVGjvwlFO/uy5rsNWevim5AMt365NbjOQdRakURXZwdN/BjJ
mTfK7md2is3X1Lj10N5aQ8w4EB5CJ5wWKU8U2KdCdiqLWBLmLyaw8NZ41GkgfgSobIWuGeSSYO5I
gIXqp007jhDl0XWJMGV6tNDb7DdfkQttEusR0272OSknc+G9hL1SnWqp0XOEPmR7hhekinPXXT2b
qcnGrv76e6G9/8HmCslYBkFUTS3hOYsnI+6DmZ24+uo0I6LUgnETVAC9Xs/F4RZ+tTU5biX/u3Yg
i4uue5pDx2jRG7g9nXF5XuvNSEsxLa6uYJNSMWHUMU8q9aTviPAqToGL4ERdCTY++xhy+DoiWnTE
0qNyaWhFx3NmSikShSj9+SzXPngQpNl+Vulrc/PaVTnRUtra2IZWXjRDRQFm3F9KIJiJao9lcW+b
SXLShX+ygSK7IoCWyYSyhVPD/PWBu26FjARkmoWIb/2Temm2c3Oq8mYwICq/feVGkkBYsgBK9tDX
lmwkQV7Kyb+KTFBVikOd21knipH3pFCiu9BaSbyGN7sNJwnE9OgND2BszBPVII263X2e72b7iQ0r
M6rXMFip8/5Of4THua3CBUbIWJpyct1ieRgn2/R6lyrkmnDQ1NLiiJje7zJAOkhVEo0Ilsmy5oEt
Zb25kJIyIZ4QNliNTrnm3+TLYbkYZKQW0GGBymB15cOdI6FDrokTmZ+5/umEFxvhrCZzHCv7x1nw
fbYAr9xEjIXVXxHGAhUGH9vLAufUhS92XK8PcXbkuy5vdzRGdVvkJ5i8dPy/w5Gywubn3/llfejD
zsLTBg5oniQjuWDwtalObBXjgEOPMty1zmvn0+qXuSGCty/QE7QTY8ljqgelJVboZrRq9MHJTT5d
yTTWqURArvZ6Eng+dmTBcxYpKboETX/iI+DSp7SaLkBlBM8Rgtww6jLIFOcuZiI26UkBTzV/9L2h
zzEVZP+cbSAIrXxtqNbjrXYD5oY+g4hX/pEb5y1923Fy0/z1z9Gv6rIDIrLd63HdWHXQ9OsNlwGO
UpudzdbtfqdWFWW1tgZoPz6iOBNKOIGCSOMm+IJqjZJZOIhvtlWFD3Q8hq8Aa6zZMVuLCwkm13qg
0WNheMVtezaE76VUb7bcom5c9Ft0vVlAZLBomFbYzjIf+fKDhh/KjiaJo5TVwnNRecasY9WkQbdI
vUyuqw2Kik+oCI8zmI5olAXqmBVeaGFK2LFewIRr7EQYuxpt9JZ3r+bLO1IuJkrgi5hU3363Ei7b
BsF2KnktHAmi+fQ188BR5RClnanwZz6bu+FwY7E7qM9/6Cc/r4F0jeleodvHVUbp9+L+ZntTSch2
XGW3wEKVZ8Yx68N+hbJfiQnpDDmSLSXiOG2tDCDw6V4vZcPlzJ+B4c0l3NDcWVNWXfVGQUwJicVh
k8xQ3N71XJUiBzvqQdKgQdYhiCs7oX2JXiX6duNzNoaqktu7s1KNFm3d0SgxohiHZxJnL8v5AobF
xPEKdejchiCSnWbENfMD2gUQs6G+I8rf966OEeHHgBolVUXlXcVuOTW5oN5tYWRCblwcnsS89i79
ftNmDyNpjW6ivd3mIcn2amAPny4FzgYadIY5wSKfNUqR3kxnNv5/4+pSZ4tB0bHbmi4gYGGOXgIL
PmZj7HdqBF8s+o3T7yD5Bql6nKqtLpu1Jpfkytzj4g9U76hGReWCo0NMlleGMKG03HtLCPqdBial
Rj7tjXt6YVqsnKN24EHiCQwH5u2vSls4JLBxLfK5YI+mpnjF6saw0wQeBtU8B1nziNsdprP57oHj
FG7N5iC02WJsOHQ6VYvpvdMtllLjXd7PnGnnA08wqw2Nl8gOonbd8x+xE8p1xxBmcuM8pzYMxInn
QFUDD76TmcGJf5pHzs7Fezlh0I2VLnGwOYzLVz8Sk73hW84kJLD7rNIRFT1qJRJSGsVL84mzv1n8
7kAjcWwCWDDpmdMV3y75yRJslIt3fBYiC92SggR8WN4wmZNaii38kb+PHg+iLeYnAWi3P1U0Gs4j
vWbnzIkeeLM+3AAwJBzYpRHqmbBEEPy4nuoqxp90xAxPhfejiminMBJTCH8DEdFQ/o285Gfdyu+U
ZLMmk8v+czQxDyqLPHms89un0NFWlF1TowwE/5PwniV9o1Rws/hMxv9yzIduwd84f2OagxqjK46V
aPCTXPar0oXDBDBKl9PdwSYJBe0FL6LeQ9+VjUizKllXux+flGSmvkajx+eXicCDI3E/hGqL2kqa
B9HYnjtIljSoM5nOFoVZM3UgLnYG9fBVI5N+IQJ+NgP9fnImKiAxMrF2KlKbrMzbc8/LWNyrfvV5
aMCcBwMCIbaFJPNshddE3agee8d4flEcdigeG8WHHqietDZfvN9PuVCOWs01Ll14+Uvk/X68Y9TS
+Aj5KEHORBWPLUo+VDbNgsggqfw3vqNQoQoDFRRZkgckSlHg0cOaz7ZOSdknYYgiBCrwCbAjE3ic
gZnqyEx5sp1g3+QxcujLUYnRB/Bfk70iBEdaZS9cVuwRTl2Z3R0U/MQq6C0o9WqtGD0ShwmPwWsw
vB/qSX/a+F7FA+lAmkhSOmrRq0zayN4ARipf/A0pH8FzToH9TFFjVbnNoswunOBoFYeDHZxzZn3E
3MfxA83Ib+y+b1ELWV+nQM7ms1kgb2WM7WoeZdHNdrdrdkKGhNV0IxffLR61ZXYpUsWxiJQDADz3
EzHttxHcidnZqvgzlnUH43coiFbwy1kWOwlPHKYjig0hqyO+i1gKbhoG2euvShlNpRZQoOM6/1Lj
IIMdjsiFu8pBULeSRzR1xPXhkOf768VP3Z8hxN1USnfwB/tg8Kr1v5XEduseP0FV+BL0wkPhmeau
krhUL47iyb0FcZd0BZ6yrfn/bg0SyjDuaAFHErwCIhhtfSLjFfTUJILeWGsH8+/JwAgkBHUCctLO
XMFLchhWgUqxcjkr0mpG8sO0JocP53G9mqCUKqwdG9F5NgyMhUFvPHZJY95WMu92VGojNdloSXeE
SaRcqy/GDtAXXcyRkWuo8Dnmux8qRzxn+P6yH0D+PN5ouzgSRgkwVN212OcW9aIGDjRPV1BW/tVM
8vdAgsKDvvhPHv3Sn/+EDoO+s7XbcjsVGeXDc/BCEgs4P7YDx/nNHQZCsRUp4nb7UYR3c/3i9mi1
eQA/CYTZ3A7A0tFkg5qSIxB1octWi2aeRTgS0o/mPk/U/+2mEzh0TNSUFOr+BiGy5StYwTbJJsZo
d+dpkeZnNkgJMYgWXE7BgEVpOG7fN7uz31r4SyLuxCwzAT0f9K9/nZ8DNl1jheQm/Ba+m52eYK7u
BZiwWn5Ria3Fjdsez8OPvESB5vUHwG9XExWoBiLRVg6MSB95E10eZFe0TVZHoYqDX+BQ806iKp+r
jwVUjB3TQyACrkYK+nyBZDmFGECnB9vryurAaVZP+ibxYOPGyH10kVUx50TccgBFGOg7vbP2xP2s
nCHcXK6b5WqxIud2oSUblBOwKR6zRQCegTVex5vlDCNlp8EgyhUqZVyrY7c8lZmWYq7Tit2IXdPH
51yLaSs724ddzJuCvbq/d5KhIMmL4u0GA6WAhF452oq0RoHCPhXTCS1V8w0NZqid7GRehb/lcAch
1vrgeXc3oblRx/xuQKxpZdkB62pHNYHiOR8a1YQ5T4uwVAyWLzn4qUnS4ZJwQs3HMD8xuaUPQoJX
CIeYa9+4kVypKpfsugsscq2lzOloK0JlMgWQXHC/xBXeVXU+0rexFFXMB5vKSEPvVNw6syh29b/g
PcpdY3KxauZGeKXeY5GTzE9SkuGUAWejo3lZ9IB3mef9fpBqBxxYKors5K3aIMbUp1BkIci2EUaT
Y0Pn3X1y7LHvs8hrSqwh+IeHCp+5HeMeCb/PlYiN2viAkYuNnv7rzlvJSYUBqZ8Cj8pRQzYlBUFy
N8u3XE/ZJ4JSvbP9uPboh7Qflj+ujp0Q6ii2ya+Gk6/BmbC6PI4CZOxd/uhGnUSaDCR37XV+gxwk
P8ujQvvRqHUxFmWEdfY6R3sKkQhgQrQowSsGqiqKtOo312R+Stubc6gueX8kHfhKA0L0+pG2M1Wv
dMsLvqNBl1WFHF85wqrY2NKpPFbWPq/XTP1HtgfKWUjC42iE+T2pVTw7Y8dAZWZph5n33Sx+GEuz
wl0LtcvAH+ORxKXp3cpyRM0P0mPhwBk5h85cjjGZ/DiU74/rMfeWGu25wGOluN/OMGfzNfAl9Bvx
MtxS2NEA/zzwPpsWmXUH/Xsm1LVlVv7IsqK0Qrw1nedOXfyjSthh3kpdPI9HMA5M+E+4DjOhPpjA
YzrLOHwDT3NIuKuWFSX26YsNJOx2L1x9FVLo3RjR7qn3t02MmfF8/gh4VTQD9oVFaMxZf0uiFkSe
VRNRgMUvlzsq7T2a3mz8gFQLMtGJas3qfe5b6FEWNf3XgC0/CWdSILWbYMMf3oXYzDB9cQ36eSQP
gFDt7eon4c3dBXSe0nmIhkAi/MN7B7mQUvIyq5RcVaJsHwSnMF2KKBUpMEGFxqi3hoiUKJHcoCUU
VGgdC+KUdCibY1oguFFvhq+JcCHQ/LOb4mXQKRyKy1FoslCQflMbVNQvHdOYQ9SKSOIDe7nvDw7i
1WPpbUgUKW/DL+DwQ8OWH7c06E0Y8PrljDas046WMm0u+yrgtaDGbSRoWcPSm6u4Nn8urRRVH6Dj
oC0CCTN/OEgHiLFA71Gb8oSf5GYuIcIcAt0IbSmavucln+5SxM7i6faxgWyBN3sjEGGKLupmOiie
n0xD20uIZN+S8ApVm+fxw+JngvSRJfF466owBKeKoF+n3d8//Phmg2sj1sboATw4+K/WAqCj07Nb
fwBvi7ebLG6VmBETCqyMGjansGVopj9pF2sOT/rHShhqWO8vKjOdfbziFypGyk3itGn9+8jCpmD2
k02yyC1/JmNAVJ/8GDPDdBYsr9caHdNzm1WJEI9vUnwwlbnS18roebeWwDAs11njaaICt1ggDjPm
g1z+DARPqcx2F4qjq1Z60JH1nldSzzygSthr6CDUFBG0e+pX77nRum0KhWY0l+Bknew5I+wClK77
mvuGme3KsWvqbdpUZDjTHK9OjVireAWa9mcKJ0aaJ47HJroPgi9kVISVBnWfonrNpOKQtv9OKKqM
a0dDB4gpg8ogyCAX8wF3wwsHLWpdnbCbvjQWr2TiQkW5dcgySH4uH1l2GPfZCq80WYJI5IgfrX0f
1Tb7/SR8HZsZCN0Iam+tmlMTEtRakDjTfAH5NUQvszgT97NY2L5a4Z8QYoJivLBPf1cMGEPKptC4
wnxniwFgmbIN6bQoMieL1UC3tnfDPzGMYuSGP/0Tl6yBuYEstyoyLqtDDFXWy8VJbUqngFUho7lG
TY4VbAZFfwKzeHCJ1kvA1JFQHnzj9brlG7Fj5GMuIZn3df4L3vPxgdIaKkrqEywyIPPGbSv9067g
9TOr2nHrG7ZDWX2ta+/ianbg6oqRBc3WNoFqdYRKJqHwhvnKTKx0VAcixwxMhhsxPQt+k3ifubSv
ZaxdUnB7V6x0lLwR64vDXQUyUziK3E+hHTdxq+47UkRfRBOcPhBOHCgH6jUV56C3pVrPe6Fbm3lW
VpgR8pZnmM034m+kx+OB2xJ6NVGL368e4iqqMnDK7NPQV8bidxBKSHO0cVm0Y/e4YlUnvbooRQRI
F03xvFyOcScHkBhNrslXPZTusk4zvW3OygxfPjOMSaPSTPrf5f2ESVNrXN0YL/XCORqirBhbU94x
tGNHg0sVzlsSDAsnnCFS0/0dAOned55WONVrudqLyO/zTISZJonV13llsw92D1400aQIzCByYyB6
1TbGfq5FmAD8INF0azUBuSKLRcYLrjvxlVOzYoe1gX38q0cC45/GX1zfrzulfxUWi+eARSN9WyN+
zdp+40USCe7LS92HGlMeP+J/+q1ZnvbtdZ3muPXDImKGYStF0WVc4QqbIuchB+5ww5+HgSslSHBh
Q4HNJlGKTBuBSNGdpyQe2Q+hyo5Ma61FYu7UXOgvoP79Lgnb/5FO2/T8V36VP4E3MDW/Xxu5wjq7
F7SqDCXY58QiTG1DeJRdqWzxwbWqOqTWHiTsUaPsxrQZMD0OSHMS9+3tavlKvnpAq6FOSAae00v/
3+8I46ZCR7tOabQ7hoGe7IdFsYAAZ8OAz9jZ585D4dvFtxNnrCmcP4BsG2BhjxxZZXWIyIrX2mcq
KuKJtAy9DH8rFYp0iFg3vAX6IVJYD/NiCeso64k/Irzm1MYHmWJYDWkh8R8ywCpr/r5AcnYrQO45
h1HRSa2jkjSTPnU4xpjOqZepmgBGQIJyfduxG5T8Xx22R4yXvvUJaslycSsC0S9eFM1ufH+ozAXk
fmwsFIyOAPzVFzzayWGMo7XCWKzFexmQRhvnxXGdDEj/MEGnWpFah8RB5IQedoTgX5nYRfgPduiQ
NENuYp686TRTWfbAF04ElcHdxBGzBW+ZzkQLX1BPhUbEn6Wo04rx7qzWbZnVnXHWOC3NB5M0SamQ
Nd0fvJP337EpNPCcHTsrMKrORl7JktGvRWM3wnKLXwSAmo/w1tCfOlREWaLnPIiQHCFfCjp7e+di
TleKs7+w/PhZfGiUOq9MT2aZbl7x2tXTNvUy/WvSk/bCm/7qp8ELgs/HXO6umnSmWAYNairxgLtv
WwAFmtWwD/hIbAu44DL1DdNXpcp5SlD6jp1ZGrEgzFApbl27+xoBs8+LnOjLDaHxhTS2Px2ceX/X
fQ1zLVKU8+NcCB9K8YD07tBM9byLIcoQA4JnxWkqb//b1zIgJjT3lC9vBNcnLXXcOxklKxpX2h2y
Wih9NvC4iVXKbDZQUCfC9oo6KcsAdIgiidQq4DzTjD3FRQAPkFORwLU6MOfr6V2WzFMKb8DVGUID
8YwGnISQPG6jA6F1B54vfK8+BURKwnBL4XZyoQ5kjZcvpgf1C6ZImrzreBbWcbCcnD/sp1waZqx1
kasW1/qtiVe3eikpqzmM70eaDp5EPBPbgG1ANcWxYYEHSgEijsmE4lqRFCFDvStWZq5JR5aGSFF6
YkcnSby4FzW54jlxrWF9wuDLIO7SyGWhtk2HHTiqgcxlNrLDz2NHimJWTmA537dRapStmRgUkkJh
0kzQwZEN+1uL4VqTfB4Qdl06hPGz388QtWcaAzNVx1YknT1cz6y6UiDcdItP7TBO73l9pYZZ3f7h
d5dI7OFfFExLj8Mmnmi4nc2tRlfJiNV/8vlBoNn/FyRyM5LwAuNc6EZ3gmWumwPdO8BCf0rw6/gd
qrDLwV02+Y/u2U+US1Go1C1K/rCnsbcYKSUq4RlgrtElb6HG00MUXMoa2xP3WVswvPu/nsHNglIs
dr4f6IS5nPx8uTNREY1Spwkvj16EGF/D3Ze1s7fA+oyfcQ5yIQ3s32cdyzuOca0rTkq3bWzb9Rby
4DYtckqMphWq/0ivBHv8phcS3T5RUtS+JkmUiyiTgxDWyxm869eD7aO0acc18nZj4QTsSqRg8QN7
z84XJxLmxCCLXEEMX5mDoxxjnQrqA3E3cYkl89zYT8x2XC9xjvrF9v8MVugfiDlNcDJM4h1So6JJ
ybnOowJEAK+odUD6r++ijlghPHhv25MhOJlHkhCsRa4ShyoEyppM6pbTBtt9IWiupQC+lgVdkrMN
lYmO/xHFL+TgMJdiq+1WAtIq/q/QxXL8ZFs8EjMDiQfELocnbfhRqS20Fz4cwRzEKsImBnvuxZVZ
FlUcsL+GDOl4k4lUgUA0tiV2D315Q5X091iUcoGyypiOco3qNj0DS7B55kG8AdzHliA7J4euPfKI
JsIhRNHhbQ7fwtti+/AOPNssZRFgcW0AUslgD5N5xM3ZvuB4SpDA4GdPxZl202slkiCApin8bnaZ
uxyxyv5pYrDMtQc6tPdkziXjUhag4DVYPrmfYiV3cab/kTcpuK0+bHQcVoJ8pLdL36rfr6nQ6QH6
qhEVAm28W/1ZauqX9c96Kr2Z5hahWNeh64Qp9EjzHnpNmkwLxel85hHRm/drGZoL4TXUnRM1ZHq7
3fgRG1SFsPR0Z0Egb1UgE8ldxSUhKVmZ2cnsjQiOw4ydNSwgSuya/gwfwhphkDxodZ+E58RaS5bC
NBUYVWmwNNYafAkDEPqn59kYvIs9NwiLhPIryAIO2zy9HMnt+Qj2OAypWdoXnkVF3VNJ53lWr2dY
zUlrjgyXS1mMHlg8Ag6cN0kYnDECQUXrU0ZwZK5EtsMTIAx5uWLFl/oRJv+OrIOWFRrKWGKa5dgo
mhuwdtbI09qoNPVJBtiDhG/IeYIxSi49JZPrr+f7X8/2xSKDqg/3hDIHvywDCSrszKIGq/GK1XJf
YdF9o67GyWMgmN0JLf/dm9vnsM/xjhJ6gefeAccXz++HQygXEaEkBF16WV54dRmEIe2Eabih9+Em
DDzqMXS2p+fAkFfn52/PU0YalZSO7pPsxHh9nXfk+z9nblj3jdyoaElNH88KVyOHyQrJPcXddQNd
+Lj3NrUItZPfjKVivNsMHW4KrzM1dRTxSiicYxEJyVE2MZZxo9+1h7gtl+Cmr+IXMmN+XvnzbRhf
+pr94ZEQEXoFk5FlVKVUYQxyjwtiWlXINyCAmmsq2HijOPCctF/IFgkuRdL/gdWdbfgcZQF1dEAn
Sp37ZPcjuFP74pbYREMm0ZDTecsUBwGoAmfxJl6MJt1o8lYyinbe8rnL+I1tFPyhCxNd+Vu3lCoQ
xGYjoTD+V+m8xeLX58JxMdH29W0cUeqO9VgnatUnF4SmDrW1PNMH4RPhIdOm3eIrq7dSyuAUITzg
hghMvPq+RKu2/0dRMhIt1tab+BtDX1O8W++BBdbjEVHDcgAmwaC6dyXtliKAs4nu5CxJpJQC8ZUo
YEIsRDkBBVGfvDpSWt4Fp+GuaotHmm3CkUKzJRJ42X+uqqPDY8jVqtI794sbH8e6vwAmZ7SM6/c4
Y8YOaSAxBJA9VjjdCWkU817ieO9z/JxAOZ/3AoXiX4/NZbrsFg189YORBnooHEoO0VMp6QwN6Zrm
cTgX7Kn4qrnHcG6Hx+qun3anPbODNIxUdIP78Aur6HakdkWoHj98VXmQIr7XL7jjBcqCM2nZVjxA
WKgUBOhFQVXLiD/M7RyhwNFlrPmwKP3mYtSL8SVh6gMoDUNPGCxRUi1y6EV/nGWR7jDJlITMbcn7
aae7XfkuHnQNzuVU0RYpQYl39pOz3F+/Fw0G1vfx0nxmd0IDn1/mNfR+w9xZ6pdmsZsa+Mwv3b+5
s2dys6pgXtOz9knBJpfUxmNrPbrFzK0G32+elfDOZTNxsi4y41n9hfgWSHGKWXjY9IMx+GNnPNKZ
4FjzHhM6PmOnk6W4KPEW3uXj13+ogFEUvjQgwDg64LsZpNKKdDFLYrgu5/xC5rQWlj0nmKcbZrL9
bPwIES0lV6o39eJFfQTipmF2F80r+/4WRp1bCrSCGnz/CSoOBiK08wFJD2VMMh3xkWLp5MLDwHbq
ewl5ILctXVDXyXLxLIjD7ASXZ1PB8RIXY+AxQeSQfJVnQcmj3FtjtCogzmziWLxW30L0VWC/3Hcg
V0egONyl2zUxt30M94YsxbM+PxcrO5fDg9guqS3IfTe2UQV14DAb5ocaOo8HaPRr9d/Cbsl5iUS/
TrDqHhhz51gRc4djqNAR/MlRtRZz9mocu/Rizinuxokya4WcjA/WlReJYzf6RGLhn4HDgoTHmAqs
gssTnWQOCIR5KPwMmuZHDd+cxgnAX4pPIB8BTsYWFCo6M4lCeSAgGafcAJTRmoPCc5UMGtVtycmK
h73FwEba4T2iLV7VvuMKFD0N6hYTT2OO8UwWlgAa/EdtKLOjROvJPe+69gUHsL5y76dHGyU+GerL
6p+qC5h0GJREqpHUqsf12nbGaatYIpGBOU3on6R7JYxCSAZfRYhdyR+vM2Weho2oUI7qhrzkXjSF
ht7qe+lW6+h+IR4zUdV44w1gYfr3/VeJ+OVEKmCdxk1hGJ2+mDmr3sgiMwjMnJVJ/X8P7uweulg5
qE+4bMAK5tU3Fx0y98G3JTTWK86S1+lIRLnq6iurVKuGl/Lq+uvrltEv5al+TQxjHDEexW8+6SHR
1qkeWHpB+h1770odMZhmZG5rpova9tev5SZm5c/TxrtAlXLQdCfQqz4ilA8LQJJXwI+3Fhtb+59A
wjYnbjXBn+/6Tu9nXzK3xv/Z2qjX4BKcCTepG+Qera6iLqoNDafcD8Mz/3P8dd8JxXHRb9kVttwW
47TmMX42TOXQ5WK3JJlKxzH4yXmpB5rQLahyb4C4wMGK21K6RPneQ7hVE2vfZd9p2WBKmnQuzaka
Ej6Z8lvuMCZL8v0vmzBbHtuD18f1+rEkv1kU4kOaY3EtO65XX211a0G9S8Un+b5wXUS7h2usdPlP
aFVoopo1w3ctOuOO20bUQc9A8fbhFuvGVsox6eYGpNy+WeA5Zox7UqJ325yAdkahQyghB+9t0fEm
5rkshlLVtijqzCr/OmHhndnyO/tP4GFaUQxd14CeyXrWu1gzkvt8V+Ej9+LddDCPhmvCH0y0KXTI
zHOU3NRb6sLQkZRH12NQshaYnSVViNRuryj5bKS7zI5S4Di6JLm36qpoHNH5w77N9lbG80rd+VGv
RcdibFAW8CuGWsZOCstALzxq3EEE0jpdinfLYQDlSi+ac+/h3o/BzSsStJ5Pz2WNKu1IwHkLdAFe
wS4/NjfHsbqgSlz6lfdnF4bPC5IMsUxUeyYbKBVFQsONVLZPAGfO7KPwmhl00QkkbJvUjicFb/tX
hz6603MoslZU1AapiBsd3Neig9kvpEdcGHjxvU5x70N+VC9GP1Hsdp+55QWkbi+SBH3FGwnp9DqQ
OxgckMLQoeNUmC6ObQFtR2Uq5HFcrB80DTdEnMc+KqnQ1g4TJXnNXx7jPMb5GmhyyWM3T0K1EyPZ
1Q9nhrKhZTh19abGYn7WjqeVFWS2z9X0HOv1dcs5/z19e1hGtaV/VVf0+f0fkzOPwpLa2KqIb4UN
FiJV0cwe40C426Eo6hXeJe+9gHlmxO/9ooSHPcwRSCv1EnOia/MTxWctjkQAUFvB9r4pZiWt8apY
FOGt/dahv7ROCwmJfhfU3/IgBhTMSWjj/yK806udYYkA3w7+xIlSbvvFp7XGlhlkw8RUX3m9JTqu
foo1NKuFaq9AWuEvZKcBv28mTQz816Z9KRb0XydHegxBp2gSflD4V0GUG8GTRHzasgLuq/JJDRsY
ZXUZi6bsn5RiJgtxXK9b5LkZbQlWV9g2noekXC+Fre2LvEYo6FgCgbGXUgy5WKuY3VxljJDklIOG
jhcBsENhru30El5yTp4oKE2sd7l1eMXMV5sdRf/bK1mNO6H4d/jHSRzxfgBqZC5Gxj4E5lX6PzBL
47UwXFUml37fdXV59yV+yUvlccC0BrjkoAVqApSZHXazZcaC8CKcHR0s878cnT/XQxZDOO/+Ua1C
rq/HRyr30VS79F2asO8vo0oBP8DHd9L2g/8YoShx45VnfsbCF777Y2Celh0yq4lkhP8DtM0JqCiY
oKKGUfDyOem8uaX0WELD+7CbkBZlkcZ6XjheS+DHFuSdPtUdTEz+RUXVmFSbuErCsB26CCZHy1VO
GIEcg/OjxzodQHwFQC/q/UOUAlnivZCtytFEqq/8pFqSVXjmUQH/SBoTkHAd59DlJSHukQ1K40nQ
1rHF4vfV5loYolE72J1CaHL8UmYJrgJzhbiR2985tEgiolneOrU3iozrv+1ch1t2OEAKdB4Ib2cN
FqhiXL0tBrLiEkF8nqIsEyf0IOlz6hGxjeAJhq+7qCXMjL4EA/+GIKBgvcqjdjvFOxFtbtU+/8TN
ziiyx29KH1u/b5GcS0lFYVP/PLsEhBb+ivVWq7yfBk/QnXXZk82cFAwRj+fgP6ozvapmpRYAHHZn
l32l7pqKd8LdvNrat3HigeR46efM4UFZoUFL47TlSpzx+6d5ZZwia6Hu0JekLYXjBSelU3EzSJPp
dk6NoPC8ua8aix+UfqJItTJgLILZzN2fENrRrt/SwmeA2jztr0zflSvrsTK11pxwLPEbPpucNkRQ
YYx7GFEnqeaquNAo0HdmvpAny/suopYM3wSGfWLb/2LmYRhf5xAoYX8NsXEMt/WxTsw9if1ZYFxx
wLtYbF4gj2o/UiknUeDnoidB5ynorcILuLZs2I1KmVgmnsfZeOaFFk7NhtVJDnPOXe5+tkrpICcj
3Al7QyDe3LB2mUi3ErVUo6DPqco90Cz37wstIVa6SyrzbQ2yTVwjimGugViGlmqiLZdTnmb4dMAX
CIbkyA66fSHV1FQlAZnSJETM2eIf2+rPwnThhQQj5wYzj85D1ZVzeqrst8IHVpZKBPP4Dbf61uoG
HOhoqySNoO36QExms28ft9MTfYF2ZgvJ1SmfIv2IU/cYQjxOIh3UdvWdeErzcVCvqiH4O/pICNRW
pMwJlSr+RQd22g1F8CQUFhSNacA/B+n9o1fmQWbc8UQx6J6nSXfs6X2U8leT7zU6XmOziTH478dJ
I+SPTa7h4/8xy74WMptTejEVtinh4l+rZ+gQkTNJtaVdbLuVelPMFKLpyHkQZdl70QWlWw2WhAbZ
kQrVuqpDasKmeZHLysbvJSGrZ1i8LikDB1foWmKZfzraH63k5fTNNAJwtL9S7YOTpiHSMiBLh/M1
ik2bZpNQZMzZQ63G/dLAvdNLo93w79EDzojvVPOlZ26B11H2gx8tmqdO7/P6kAMLFaq4D7R+OVXA
Ee8ElTX78C/zsCtTjW+5XIfGViamjCIX6INhnuoPDNIF992loCbAluxzipES5wZYHTVJPGPNhJc+
coBMgr9no3DNNFN7d9Y6AEJACf5bpA5C+vX9QwUnVa/ITjnarLjjIQ1wDpwRg+YyTPP4uuo5K+BI
3+iXJCAHpZ5mofyDWcgWqE5JxR1Zv/w4puPk2BKgYh+xs9iU5+yFdXloYh+2wZP0GFmsJyriQgRZ
99OF8B8NDs98Q3/KWuR270MFTUtwZQs3hV1UMqcIvwSEprbbP6gfD/4m/9ymOuAJuC5xU/Ufy6ex
ByR2DNZBrmDTcOMy7U8dkatqfSblCVxppQsVggxsu+ugww56Q1vpQJ/zV/pmAu5LQ62j3mnGn8EW
xtq9b+oCU3Bva4Co+0KZj79MFwoLkEOh/q3Th/dSen3QTEqKXkoBDsfYrRyuPidC5MqmeiLlTjNI
8Um77XcVZK/jRa/n4/kPrfjxFvSKpb4jglc2tFGnxmGwtLoHYSZdmjHCYmOWGxQtWxUC86Otv165
fEKeyukqdetb4A1RT5x44h25C7wQX1mRc1AHLS0qvkDgoQ1YrDZyJdHr3xAyWnonIskpQRiHVEA4
qYDlnRlNtzc823p0lQkw/sCM6CByNtaFDjnVWcSk8+tgZrMp+RyXahD/IXNk/mG79DGd70Gh61v1
SumYiv1aiWsLjLYbuW7xuqLP+p2byEeDxIciga5rADJgF6g6Q/MswnOG5MtiviN9FTyjFydT5yIu
Fl9T+lKVOjC/MBANtt7Fw+wtflZwMXMxw7xIMFdjXE5E/CDABzfxzkVp+FTMW7pWAAx+qJNUHD7k
SRX81z2pkKG/chi+r9VCmaBNHFWq+xjchjanNIKd+tKzd74Ph175yTtt8xukGVw7QQrCaeWCG+zr
VvmaS8km/kYzJP2jetd9PzQfETLxuyD3mkPnaw6t8A/Msb4tMsRsH6ujgqDuFnnCgawLE0sWLDp2
vD6VRvz89mI5wx+rNC557OkhdPK222CIU8I/1CIpuuEbfYppIazOLB7Q/O6ozTaZuWrDgRj8gVfq
jkg2UNmq6iWzSqCsrhSf+qMHeWaFaUaWV3b4gEgketp+7ypVSB0csrqZ8EAIqInwmxkYecei3Ftv
/xGFe3lXxgzN47x2yZH+0jIENn7tLgbhonHj7hKEBJ2nT2Cpymw7T53KZAMkX3VFcddAeBeVVfRL
M1GZRijM0pFXs8i6IvOJMKcf1lmw4ysOv5dfytCLBU00j946uZ4koaf+v4cwvC4dHszLKFJvN8Tv
f/ifdNdjq+LGDV8Yx9IqFJ3RxQ5SjYFJRDqEs4dWQ+5tFxvRd3EHF5SkWbjtPwInK3mSQGwh7lw1
16aoWOfojzNTHVTmbBrL6Z215NEQ618pkX3oHG/oWbUYyV+A7bRmBKZdGMt1YUNJzt882YiC8ifX
m1Y0Z5HQXHaYGeSXSXPJ46E+TU1EiSeIoGmC66NhaJuUGpXi76kMZyDaj6GXdXaPWgNUfE1g96AF
ZlK3HF33YsNnRoEKjAWWV7oBvOyWRtkpk+AdJCJBMRbONhCAPKYIzk+SCJ1UTjMYpXlwPo4TdWW4
Bxan2aRUy+/xk+8/MSMYYpvMi15R7/Lgo5Te2FpPlmR8BHznP+L+idWyOAZ5rzhnSzSvFtj+1e6+
GeKCAEJq9ktjR4dUTY5xevQ7Jk9jro0+7zpmiy6J4AJMu4QedUVgSDq++BgWEIFTV/IW5xiiQmNb
L3w28lnfkrf1201ojCTRAc6AWi1TJ9iSsAT9W7ce+bvF3xv/qO0wRbnfRy0Mhhe3medUsR9XubfW
o+iHf9KdeTyY5fYYTGX+RAjEa8Mvlntt7e5OGHKUfUIDeEKPc9nIFeMrx+qbTQeW8TMds5Zy5dm7
OhQqMM8kq6ULLXCr9ByaFePHsmcOYhP9PTX72yVX7VnvTS55rMNeaQS29vE0DgKcSva4dJAXedjP
FbH8yPj8FBD7l0/17NFb/QSXQlEf2H73glXdj93ReDmqRBuKDsyVrjXvYSM8kOOJ+PEtwVHGQWnl
uAv0GBi+L5IQ1kzneuUxJt41fXxN4HtGNJl6hRQ3fkYjy6NybEAnCf3+ue3JWW8jseGfOTPsX0z/
bH/7KMQP3Ew07Ie5HWhhp9AuU/EarEqX+zraBicDHVo/xSrUsmGeHQQE9OAKl5KKaTI6RGmF9bro
GDtte+6HnLX6E9RtnPPOmizPD2woqxjlObq197DYIj+PslBv6eBPkRY9U1dLdWRKAMmIAco+6MAl
Pwi+ksQ56aFt4Lzx6rw0hEbDO7G5N+MaiCd4Ca3U5x++RjJlBGKrCmWUO3PvwhZkqbjEDnbuMvPn
KwF7CUH0CKT6rqrF+iupwzqOVnJUNFJao4zXCfZ03h4e9gYVXZNuy5NIH6jKodBDoZG8kqB/I3NL
tqnvdAIhKczTSIhiJbO8I94ntw8i5eD7tdE5R0ABHn2YQ/PmyakkZjYDE9Bau/FuM3b7O+QzaJJo
9qmfotlWcqnUtDTytSDqpZQKc5Tfc3HyFkPwc9THt3zHHz/fSPukXPucCo2PHfZUcneVoYLpje2P
Ze4L7tPjwHCZ93k6go7FmVHWZgvAIVo4/5rHQDHwNp30+sjThuQsRJ5aYQ+Wm4PHmj/EMw1t7ZuI
NO72lATwUTAonJ0mLbpuBAo0dYn5OGcyP/UOXx/JEVJmS8Q3/nD1n76XpXbclgDPeRELxkvCdf3F
dDVaAkyQCUmvYF1XMin48jb3g21K45G55CGc4ry7+3ZgUKfNYT9Bb4ZnbvzohpyFfWeE0GWAx2eI
4ipr08TE/YPaITcBp6MzgxsuUUgoRuWDZ2IuA3UtSTgxjba9PZStcMSDctDjJ8IqqjIegXVZ1Nd5
6XRMHV4U/iDwiGeWQQFQGcR9up+OHEYhaW2JlinuPbTbaVrVDU+CLOZH0l3JlbLR5Z2Ssjl2BE1n
y/0PMpyFKFHyg2Z7yTcX1Q2ywNbZqqd7Kb3bD2s37zV1S4PWBP+uMM33j1zcYjdiRX3E+TJXdPqb
GqDProTRQ6HhBlwJ8CxsC2e1BakhX8rVd8+V5OepYdKCxz8DEaY8jHiEG8Mgb8sPVEbk1guqynhg
Xf9oBzimxv6JYq02lRGHxZy0iEUceAAXl8XhFsleVjdMoXIJvRkTugxbVOjKjV9pfk5qbfVHXSNv
YtqwpYuIIUC79+09BpOk0HSAdzzD2njPVxlH/wEsDxL+7ZH8uEZlLLzEvqA1kdwhJ7ABtGfEEv5x
5lpThUxcN0P/JNE7yjkZoJ4xpZiLjMFouMtgNsCGEuKzqpfn2w+foI58jHTRE0q6B0gO4+W5NwLu
5gTJ1qdvwLViITLhsna+W8gB2El9hvav4QiKI33xfqGp0AcHXpp9wk3C7N9RvIoAWVijQF/FTRbi
rLqJLqCgPIr0JLDiRZqWGWoNyAGW1GkseCdBYzK/qvCdClbKFZ5xTGjj/Lcq9eL8meNwSqYlRmAk
J2FK8NPU7LIr224WdXvdsXcYQtRdxLPtkxzGkC0aEVgMx2r4g09sdLJvSb2LT56//8KkDKVd3dcg
DRDyqyC0VHTUsiSCybieiJ/yitqME7OfH8LBwvPZHGg9PYqDzjcxYqdsBc4Lur8w9Y7JL+BpjIDo
bPcKyMTYGI9AeTygmrwGcZNNw2oqA4jvnIaGhUbHqTKD5TB1EiXMvnZlMBHiA/Ba07/idD4lrguh
YYZVwoRKhFg6aL7+5GN2iyLPAmJANmTPylUupRvqhXxE1YZ9Aft4bZWTBe+4BRs5MChJ5nlUDJnt
PSS1j6GBV56rMKW9pQtHZYAPVTGOME/gnZGTx0mX2mQ6RC7IzBmKMH7O1rk9Huhl0sqaxDcXHZ75
NU6GbLzuinEMwbBFJiL1ClTIx4kDMbS9PpgOo5Kd1kQ2JCziQjl6nReWk7ZsiVz8sP/FWfGG1VIv
Rx/Qj/YP9d/NMkY5eA9HK1YSS4XG735kqBzQLU2yQMRqnmNKCJPISzXr8wy9VMba3tqM3AdiGX+V
saKyIE8RlKov+C0hnbooMo+LImQEdhIiX9VbZXxXjVosVBiSeekUGZlhyuIf/oBAT1q834Sooh+R
jzvZqRmsAkEbE8mF9JMRkBnJ2/KIrAK8o8KBtts3+P2dxot/gbIhuiM3X2Bd8r3Yg9gQJrdtg7uS
C5a3nv2yz4+s5DPIaAncWramcywcljdEVBm2Ekb7Eh39p5MmlDXoC8R+jZNeA3xG+hfS2/XEGBIb
USfItBXgF9VoP5J0qgkkkMzYYNBOUnRtOjE2Ql9th5IYW33Ti3aPmCxXRdoU3GapMoVRowKeB4/A
8wP/4p3CKpVInv0NxjzPRFZltyLOAR8Y6b9KHm6kM2LqoXuF8bILwBUeEfTbkPDy2qCbGk9aK2m7
K5vJySMn5LyxlG+fBS1KP6XPDkerV5gPZTkNRq/9wBr8k4jSLiC3ctoQqsfFglSJRqF59onK5xBj
51RpOC1YAZZ1hHU6t9BPXEzpCpVwCAtevwbTY8fA74sbT7TH/KqOT1qui76WIZFkCkk7idW6F3hx
cElWM3Hl1CpCsPrNzx+bEisWRkVJ31AN2N/CbutpFOMU8tZU2lWTthhYTrvWuvS70bBqXoGUaclk
/d1AgjQ3If3buFazRFl3m1+mJ5rbrBgIfDSd1Dk3YfHK/833dlMX14qYQYqCKPCS6NZmu0Lj5mrM
8SoLjdN4nPioUo+W+PjlV0Vie2K0itRX9ZfBFy8wOiwLVihC+wtEkYkqo1qWThIJ5D2TvSi8EaY7
KeiHife/cZlDdWjJb+s41mR3RTtukGRFLmLwkowjUkSm6D8JtvAdRW3LPJs/+j2T54MTMo7jXgaK
Minf/e/2O9SqFDOMDrcCMdrdk9G81znfwyYpJv4HDmduFUinmgj/6pADsbwxBQDf5X8fFwTqfDs/
hPWHV3YbR7yFOl0MJnrt0E5n0wkjK4kA8tEPtJiFORvKNM2P2/BksCyyl9BP1Q+iWNfzw8xlnsoS
mdc5ehpSGd3ptQmkYhR5sjU8rW+omM939zb9msrE4qRG6yn9AiYWAlcuGLFfXXW+fIKuvjV+NTSa
o3oCntdh7l9W0lTqn+S/AnI5z+1Zq3wl+unIn3ooV1i7mkG75Qa9SHYICtm0nPlI13nk1ctNiqf0
7Oo5goLMOg1EVlz8a7blSocrAuw0PziJhY+5S+5KkPljNhdQtdPOUdh/CieXKv3r+U334321u6WY
uYq3FaKJpfi5InAE62Xcb3Ws2S1f8zWW77bNFTyOgdpyUPFOHLghx/XcvVWDsZSd5x9kwUSEYEZB
tPohsD9qvyzz8tZ+Ax97fg+MsuiQcprTeGoodLClLrKLjdZNYGJxNw/8Rv5oZClCZRR4Mg+TvJ7H
a8eXK7qRVI+dCzCnnK+a79kl4JzaqZzKHb/3mm+OKTEHejVK/IU1KCSrIAdEVShM+/WbF4Ts7rto
w+dzz52ZBMDPNJpePwqQ5UymawofpT6u7yxXn8jRZIxDarz2prsoFRK1wQnDiwEixIKLG6Oi2sJc
3kdFlR0VPuY9LUyn0CDwl5dFeHFlwj1xewSFXgOekDy36Ux0MNLeydlMVMBHueMfBgQM/8PsIM+V
6rmDHpur4WB1jSZypGwVJRkfPxtWgr0tejkeh+zF+vKee7f8tiJ93fWpz9quYrZAvM0cpHXW40v3
lZ22j167dFcI0U/wnDFpahDMYoJLobAHcvEgjLxnrprCpellRcP2FQCOiNguaFCpJvi9/UWqgAk7
4ppWMB/BlM39JNHFskuqmVBXgkpQaLtJNJUPpIx7/D5lD0ALQSMDBIhAi1aeUD7nV4UvoHsehuiV
hPe7/JG4iIX4GOw30hWUFfLqimIlJP8lfVd5TmPDLRYvjIQNAFt/swUCNwiQtcEh+XaGIPGT/eYO
0nUK7s7F2JJluo/+gbzEEnbMKC10yonfd1TiLVj4HV5wJ9G2rWKAFWngoj6Hm7PSNAvWAkC1NAtm
BM7CYUAWuEqhT9Tl0DA6VFzesPsmlhkrGXYND6bW5FMYjDTxah1ta6axayKNtToXeZzCfEKuLbYn
X6f+aGaBg23lwzvtZyjX7a1gHZqjp2Aw++I5aehRKzZXAS+nlaCvnx5vMNWSiKz2dtT+iqVbpGWe
nPZyMf48oQHyUvRKL4xpeaxNpkHRNjEWEgAGiq+IEjOk+IPh9IkbG6VOz0ADv78SQZ//H3M45mLm
eA1ldptuq39vvvq8ul34koIzr4P2w4yOYBDy+aDaKfGsQdj3hwQo09N8DCrFUQudF8BllEjyzJi4
2sCAHithZ55iyafELyluZehHsU47BoKs4ZhgRYu2nfR510YBJS8g+i7bzNED+TAv5pYdUc3yNdtZ
p840SyXsMbkgopkL5G/CZt76XL0eRmD/4v9eIhVric5hCDZQNlMCsURrI/mdPzP5isADdhAH694h
VbSH7zaL7fspswmcOo7EEDnBaJ5PHU8524ObOKP2O8iMPMmGCYB8ZPr2EagbSVSpzh2CdB0SM8zM
fnRStBb7nPDHkpEKprz+rb+jEzRh+RL79GtlghkNfqm+Qi9Tlwhg6g8tthvJcinZR7JDVn3LubxN
MII+Ks/JNJEmmwFcqXFCdeemSKaoCaA2XRl9VXOr2a92EmK8SQ/10A/f5H4bwhNy90EwDpExTlnc
UDpX26BEfdDmdkKhEvcZWa4f4xdgnJjgHfCvLAlcLn8de0CB6VbzpTuiM9t271hsebD0wtYrcyhu
I4KbhpUATmrQtjMpFq0KSCqvuo7FPlRrpcWr1Jpo0aHs+jofy3PDWd0KsV9DLeBwp3h9Nw91RXkp
Ox7JY0exujfWhyz9FWmXarnPbzI7ew3CpsZX1wI8exaTRnLcsiCEB9rCJmtUsz406VYM5QDEaMdw
7+xFyhQpPAWLgWmuZzwieGrune4JNNkzYBMWKhc+M9k6nG7RqPyAeDYaxeHPcJHPoY61pUTqiTsZ
Ek0Sxl/8AmotXwoaRRThAGN/GeQsLvN7o6cG4uxCt85yssSUycK6dMsXIk7wtQ93Tt4WWN76Ehej
1WQOBjNHpbTkdjO8R2317nnZyhZJ1zUjZ0bAG+1uXCX/CJCvOfgJybvhSwqMhGcfhpeMUZ+MSRbI
tlqZ6PsDuKmutVXa6BpULaVzHIKScFY1W6HrGrrVMrgKMzOcEz+Xj1ClPDlUbIoYoZNPUUS3c5iJ
rTNZhy56wpHXnhzBee6FffobTFYDwmjS4InoNxl8Uwd2o6JwtOQIzkTLtYHfCUhJ+iG3IxlCEuQH
J8EXbu9q5UMdY9bgAY/w+kzLj5mvLjeWWmdDplv8oImN72AP08ILFM1Ti3oqeZdDX4jsTxR4KoST
7bx89IdjoaL+PsO2W/pCKLeCJ9N354adnH13ICDK3XeOk4IwUrGD6kDb0g7V7xqoaFjvdwFmjRK7
d8sjVDD52+AFbPLjnTMBTBCOGSfvJgTEWm9s6ncMle+wAMCHNEXTVPumRxeHYaEYm2d2rq0b73PI
RSpa1bjhDk+Nmd4LXF9M7KiUKfebfEojJ7XnMTwvvL/9+Grr/T63gXL9hSRGGq/eE8z/iZ+6bFTq
BxU3Pr6uiatE6/icsEhH5n3dHzWJg3w7oir3lihgEWswRT+zqgyTy+QwbmjK3Xz/Wq/KTfDIoB+h
ALBou3+WAaiUdbFDRvn1k5B4SS5hUJDpC1FcEPJFF6w/LFIIZTi6g5rl5mhUY77U9IzG/SBnTMcP
IFcazkH+JbuMRmyhM7cK1vhTGBJukW+KObSyrou7gIR+PKWLPYM+ejISOEq46iB0ZhqXDwWL1HVW
qOBAnCeyspk/v/5wxH3LAy/IPjRl+unV8s2Ts9/AKhWTDkf3eRDxmbmofLhkkHsu7/h15BFl9dq6
ObPJLFva/0GGkwWMZQqODq6Nonq9yiwurN3DhIkYjTlEfgzXRnvTNumRPTLNkacl3+bVUXh2v/ku
Gd00fjA5bGxyeYVU6Au93uSAleWiCXcAR8Ejh+Uv8KgQArOqNCQSGXmfwY/ALU9SU5D7hl0Bj1tu
FFuePHGSYBgu9ciTOic4DnO0kwUu0omzUvkzGi8YCXRJV3WgDhgE8nb4KXli4XGtGyTwxFxYNj/g
wCSYSWPCdV1zQM9WXHUEDf1k9tHhtJt18fqdctBOYfhA4Ggacky+adVlmUqMJxltLXsSQNJ9L3II
aEKH98Gcx1nuP+5jSimaOrRHFWQ2PLyvANM87T9EI8lQeBK6vUGp8K0bAmzB3Y56vdnwwqEt1VFw
OwjXPSqZaBXezpkFbG0VrOpmdHnzJPIX968uwByQ77i7L7/Vg+XoANjiSyNTqfKiQlQP2sEWoqIC
WvBDhlPvlIfsGUWTrTHRp1sBlou+goxsxoDZuef9XPRXgua1642kz6YVRtxjHPaMPJylPKLfBYPO
m+MFodm4cU+MoF1vw79EfR62KyEpfrtkdfXMZtK89gDIK3uBuWCS46jtnvB7X8yn70SOR50dadzQ
EE5g04RQDOhYGbG1B1+MKeyJfZUdO06nqMsv7xG0nh2XpYtAMrQ41xySkH71Y8zTb/+UCPRFawUW
wiW1K1KO4/A6iAmpwYA6h4V+y97vE738RJC6/Fe1/Vhjs1lj+AlY/BkoIOSwILiWIcYT493xtAsj
73odQePH5GrKSaDoP+ZxtcbAgbx2JEeX0IeClbf9cwrDkMcRIac4uDwa/BrmP6amHPzplPdfoSFV
t2A949d0CthYKdcJPU9uoexHbRar65RByvM3F27SWQU46r1fKHvxT5nGJvda0Gdlnp/HNhi5lkfs
iNEzFUYS7TiJZRKoDuuKdt5LupRtNg28jpxLRVbnIYbLVwLQz1vLsUT0SMWVyErdhh7T2iBb2inA
2TycpW2bck87usnqr31qWBAD23YgI5/ao5JCgqlS4dv5WyZsgtLKqVzszWhCB8WzWK6emm0G8r0F
wnD+bGSAF+7X5yeinJJbzDU37G2q47b9K/s273POb4sL2L/6Unb7AWRtyymfnl+yrNfo8eUGHtku
giwUWiQmEnN07TObo9mg8nd37IlPBCif3lKCbI075bDhHy5yfoxnm1ZS6EXRS41sMq3EAiL81WI0
+1eGyFrAL8n07CHX3L0q0De6Any5mBZ6udXCDDwSZTcp7r3+CSKMF2Yx5zlhyiRNFAa9DiUenRY4
EesBn6eyzahAoEv8cgPIffI1AnjPQ/pTYJNMz8vJSuR/zQw9vgEMoeN6jDyI/slRphT6oSb6MIBB
6hEFtMJh/548m35CCkJT5ZFBbm+mw9+OsnyeboztleteB0RIYLwt+gxYJr0PcfuuRB/78TZ6jN1l
VpY27OYTh+Ym2wfzGWjUn8/it4lIIsDBVjaOWbOEdqNJdbawxsDX56VDVp1QIebYyvOzmu+j+VTB
xqJQ3Jejdxie/RVtWVWHPW7SLBLry8yrg4MesAA6/D1Jm/3kPIjtC712dzd59AxHwaOtbFZ0mi/R
Qx47B3ncg04QUV4c9pJ0soolXOd0mfJXgYscFtp63D5P/SPEA3mTLe8czORiwlrKLcOKsOT26mVF
4Gh89Jny7v8ZxeUo6pvpJTLEdNm8QeG1Jd6C+7DnkiXJcuX/Cvnsq4bBA1mzkwxJGCIEZRguw4pg
xrvQG1XVJ6tJm/kjvDWjOZ1J+J5aoC6RQLhlWjAbH0mL/d5rQ18b9FGfaUick9Zbfu6ySWRqxcQj
JJV2R+55+B+nuYlqnNlJVvZ7TTxULZMD1a0y5eaUDAx1fs/8JGxQmcx4s49nNYAOwiJNdhbFt9v6
OS75dWhjpC53okEZyV0zlHujsSwuI6Ft+cn/ricMXp3xoT+GlMdhEQCB5pk/25BlnKS/uMYFFIXd
R9yw6S8jMISRPuJFlbb/nZCkt7IrmjZMRx1NcPMcIjIMiBiZqbuQ5PbCg899yr8KdRYDgkHpwdbt
epFy2emaHTaV6ASgNH4AsFyfJL+dmcaqWSDoc2ct+PeGukHVSzDn96gbeUbepf6El4Prl+s7ndLp
E5IbU55i+UubKurr/G59JcKmLqeB5wTnXBjqSPj8REASHr2H9rxSpcW24p2ok8FuKmEC16UTe5N+
UsRwbn4JMiuPKjCSNw3ryh8f9uRJXR7z2HU1K1+f7jz2HXXtSc8zD0+NvfvLV2eLVtL+Z0h2ww0z
dEToeQsiYxGEMs5+Nv+x4ls88YlMJRU54rbHs4oC9H2sDQyDpd+mfAhoPxmrZ/uRvOLXq4Q5Y7pP
1rx3MUVUPCr8hJNwicOw8288Wga2n8Wc6IqWDo/WTngTTaiIMnXGfE2nAi/EVMoRFrgMuegwgC7P
RXja+7e27ZedzMis9ErJYXnJjHqO6776iiFoCTH1VPSRB2v2hNCEAJ9Ccy2FzPLoRnpdfb8dd4FC
nrDDZuhGCR6W7avSQsMoamS4JeP8z+XuZbCHl/0Mi3Qh90oPN4yZdklH9IJkQGP6PBUrJSV53RHb
B2XJ1Kr7GmtvUbs4Mv74qYVZm7wK3K2vd4z195+Lv+cPvRONVUT0aOEVW+iBN6p2ouLIcW+so5RK
CvGnHZIoLCKoopxVXDS3npSE+4HqTfS9YVj2G1oRjsIWyVmrCZoUVwJqNt0IhA24jZXR3LRxPs0m
gYZiGYrhatqpFfpVmCs5ldCt9fce3w8ohLHPXn2TfIsdT/Npc/ab1vOf1M62M0kfCCAz/sWVqtwe
O36si83yKKPX6Ns7GiosVNTPn7Q/nz8gRp6sjmHFItuc2kxa/+HY5rFggRu3ofhQat0rb+089Rlf
1FTZQcpQRm0mRRKBe9Al1Kpv6XB4RgmcXn9j6bcFdATOxXt1fDGJIyHeU3Lw/WM6mLoIHt2Qj9bQ
1AF/1r8wa06JDJJ1hcRQmbs3yU3hDqgCqmJvi2KIBSKjYhPYy4tdzbIxaykiFHYhUEei2Jo+fIWx
M9THkh5gXu0NjRO1Gdjm/0Z/HDj5JlRLOAK0pJo2Trrw03dCKcUJfShkbWSU7GBqeGopvmsnUAjj
S84SHy25xq6rBGLMOXk8C7MJ129Da4a6yWf99dxwzRs7ZoZtca76GuDAQzURphsx8SRYKNF3VGxC
VnWuIoJD+jikFG6HvnduOmU8Phgp3eNNLaRhBFf8nh0NvOPfwD0CkHB5FPm3Po5ERAoDZLpmyjg0
qaQr2AX/pxa4Jfm2dL00vOUkEv1BA4wdr9jWv6Y0UAYPZGmZVdNVcj4gBwz1KJZ+mM/uj49betHu
xvvlJyt1CpbCgn9tFwV5rNggJJ/5cG0vtG7cw2fK5YNjs/XJiIs86AmlJB5fxVkbWno2UoYjpzhv
RY0in+EIlvge7ffWH8hfb0RIWXyWTGOGxA4wxT0CqSyYoks6TG9/oXv1+yjsRyMXcok1Ee9DfzY0
Ydj50Ut2E1a7XXXnitXTM5Ddsrc1AqPmLEglMri5oTdITOcGQ1ZJP1U0PzFP0YnLFHH3ytTprZdm
NKKOK6ig6DXJZMC4H2s6vrczqHkWT3FL1GuBpu56htQ8UrkealMhNdQ7Hm+6ufKB2anx5WJ8s2/G
qiYPrzBNjFuODWeUIGHw+SNYVoBdQFqhgkOMjHOWTUmp/jyGXPNIxeQGfAor+/C/Ww0SCsX07wPF
NWVa+BbiHK/hDuVHxNoDpC0ydxw4QrIngfI9lmGJ5RSe2/fEd/7QDDSTFEoiQVtrZQ6FjKr7ml8R
yUG+tP8NuG19zEmvgN3EETNsqjQjbnKStRSPkGJVBR4lmIRAq9UG8+eNnadXNKL/8tGRas+g+c+N
0aolcfrZ0rmThs+H1ZmW1cGPgU4LpdmzfJ7sxgF/iJ2ig3ZM5MEgStEN3M3xZzf1QRX/ZjBFJCdH
TitAUI6izPf+vXidojQAOtKF+MIE4+CkIhtiZwI3sDaHIdnEaI6H2bpOCSLx4ZYqQh/tbHhifhFK
hWFNF4rrxOQgiiKDAnJudfdP8GK4OEbdWS+dpeck222d7bNu0u3gmwZ/qPK1YcD1ftNI32Y0YIJq
xdiLryMP+aubLQljdKkJuvu4ON/k1xp8HAA5wWSUp+k7F8uEknXeeCRr/50zNFVsvRlokt/LL7jV
rFnSpeUVQAPTkofOQrJNgkD32UBlLW00ATI5Nr15LYHU76Bx4p3BTqX2y+ujVKpFF8+wYVbjxV6/
DlIpz6r7bAxm/+yl4tw+aJwJZKpQd8YHbqK8M1IVJZfMyh427pU+Wn5VsRb9t2Qvf6azGmZu4lHB
9P6KhKWC69AlKDedG27PLOQzBqk+itox6wkOdige+RqLu3UtCO7aj5lwD65kUfxWKQWVScMxDB53
gtj2NoNs+9PGZQxbaKnSC3CAwiWvq8dSNtkVklbISWNJfy0jNAv9DXwkBP4lAuN4+H3qVSaMvqte
q8o3YvrFgxeSr6ZWlGrMK4Lm2tClkSODCOH57QPGfcdfFuwboeKcUkeGlfqKXy2ovnnKAHq25lUw
f/mM4YLaK0QzKaDcJ4UzF82cNLD6GkMN2Mi64bI9olgCIL3qlBmdKFBZQbwu1Kw2pFKh79tTItWW
FHUuUd1a0fxqFazGH/t8YvjcoQE8W3QpP1pEj8mlNzTnxrlAZ2rM/LAXLKEQBN84hMwVko9knLXh
Hynkm2OgOd1Cpe4qo77yn2nu3DIu0cSJXccdtGOI8KIBGnUMSdjAnwmxHvulIQkq2XdVvF4Mlzp+
2tLYfBFMkuXYgEafXjbZG/3oBpbT9cwmZlwKpWVXiin+J7cUhAtVATzv89ztxYeNwyMDh+TU0ECZ
CO4K0F/srlBDDvNRqPe3jKCqqZBp4nal/2W/wNQN4yElYeA3p6APXgvUBbEHyyxsE2n1aNu0DUYX
PTx1WCLKN4znBR/X/jjKMpu7OAxtNDi8bH/w8sn4EY7vXFXfAzBM+q2kno4p+BmcN6J0ijHhVbOE
4o9klL+Rl8GATQsuTBiMqiXMAc6tKhxVq4V+BVfFi9GVv2/p8iPq1Dmlumto86JW+6BR1fDFozr1
yt9rwdUpwFU5xxsg24mlbSvKgzE/zyZer0gR71PrZfczWBFENRm4r7UbINDcLh4m/xuqMMHBdteA
ffA1Sk+/VKhvwVd4syNukZg47SKbg4ESBcCktp16EUYdNDZzZNzl8fpHTroSuLYlUlqolkbdGYRz
k1AeHustvaaIZPhX2ji8uVYvnOYBB7AqitIid+Y9eTaBsnYbl+6I6N+K/jWAjm7wuCumNX5ThyiM
azGSYQVniMg5/FMughdys49xigOcqfaN+cq5cIJwqFpfLrtaT0XzEtPDZPXaaRYwXOVWAOvkI352
JnHrHLoFsjrP7flUocuPeBuK76S1htrjN6PQelQ1n0UTah9+DRoJEp1hZHTffAo4kdarPZtF1NiL
ywlTIPdPFAp+3FuxUX7qiMLD7Cis3bBwbuZ2zhwuyrPV+sou+OvHDlpmmjK9w2DHNp9ppLUh4XMa
tk1wsCzwawyvFzVwWkAJJAuOTbUcS3812JUVZ5haNJmqnTAxDQGZMEBU06NIvBiB3irOT62TmF92
Y67L19FT4LfAK+RhO39h4RUD410oWnSUuk0G5ms39gp1fWuec7XMbRThnVEUJULjkGXeNn8SWQKv
ldqrLtgsR5jCqf3Vasuh3uLTZhf++1Q53k5OlS5Hknfx1X9fu2R1pNQgYPMZo+q3BrILfglI8ri0
Pcy5EYK5GA+3fQ4+3ddUssoO5TWhfCYb5d5mBtumilkKnRheYPaYxlKIDB+jskyoTfUQYr8M8ufh
Cdvcru2rFxmWV4YNU7evRhpiQK0Xjw2yium1lQE/dIXNqPYFEjucKJAV3iKx/0Rxn3vlFM5lrHXw
06yzbqKlllT1F8einKvr9+mwLTDehbqXB5RtqPktxaz2IozsH1KZpsBrNOR1juLXsfKRUIYWvCw+
ABD99G7FZlQwgzTRj8DfRNlxuOM0pTceuPKFRDf34csOG1au/QvEhOqvc5WWbjzBWYQLTBenebt4
eoZv394GRCLQS6zRbsIjTFs7zLzzzp6q6o1ER/FliP+eoSFhNu87fDYP9NBqzbGtv26waWzk8IlQ
L7o9aEXATFbvbV94Cv83jQd1obPPIZBGukmVxwMH0/ySsKRaU9X0ktm7KZKJy9wMYfkLQtZFh36r
UckKsd+spcc2fdPTgxW/t6RQQ7v25bEilYlCov3QJdfJLkRvzwJtOoIVjZwxDV/pEtWxrCOK8myw
MnEgRh5ebzLT8CdIc1WRHYKuAYJ22LYpGlBR6jNPuzxN2qtUd37CoyQxPb0LRp8os+JIM7dX0c/J
KcpZMA0aIiZmEs0DfNEBoJcUwSKd2YkvMjRIgq255Xzck9ud7s2tJ/8ygdiHkCv/icv8PYTndGkT
7aTtPGeTyzIRAL+N2BqUudLrYO5TS7oP/ppfwv3GoIa5NqIRv/uIeBaypALyPdjvZAtSLhhS9FMy
6pVtNV0nyzjpFlUjU9nF6lwVICc+EB40Owd2Jb2UALcRmyJoyrNvS/XsO1KDtPAHap/kSrNGt0xw
VN904dhK+9wcTtlgL/GQJQCmdVkQ5URdq7oq4gDCTFsWLZGr+4UPH3or3MsIQAthE+WAUTHmuS79
WYMuT2bjbtzIeHyUUrBeK3lS9CMHvea30S2XRwDBF6EiLeBka7yPjcAPe0yFzUdFTJwq02Js9rFS
xdVhD65xWAXVB6+NvAG8brLymH9mkBHZlWa3s0UsvsbJPJjZUjOwrUoKuptFdaV+FDDAonMmLDsR
sTvTvbHKQ+jfseIWM7ii8MPQJFvJGhRsSFRsLsHoG9XMhaPl4++GKVMbhqrIld6+AAbzFM8txw21
CrMrwABz6B6xxEV2YRvJAt0kW0QcYy2joHa2iOJqT+LZGAUmdGEJS/emtmYfzXMhOVKDXisU/Pry
X6M8aT/suk7iZnsL72EXWtn7ePEI8AE/CoZLbxiHgo64cb21io2EgDGz+8D5ZGZRsKQ3Wb9vS8Ju
wFm6qn5pk+MtC11oJk/LAy9uGVwruqqddQciPJvZOQqGizkFp/oLwX7p6XFZf0Bnr/jIfB8qVwSw
2hYt6214qAvIVKtLKaoH0aRfkaFuoPDdnFOuclHDV0hCHryoSGAOSDtNxlGYxCH7QKX6ElUBhW5v
CWBvjRDuatcPMWxUgLIrDDYtoW94G1cLk4v1WMPCz+0c7VKh9JrRJ00Fbz6Vp3//o9Y84Y4vhMFY
QkO1z53XniF8cZgMq2FRppZlIrgoKtSllaO2Dt6iAlVP37Bxbt17gLFh9FLPgWA+qyuXPFYZOq4/
SeaGfo6ILDI8kMva3cGPQy93ACso+/ySyVJWbC+Yqd142IE/5N0kjW2d+jjFfpz1UiX86tv5t4Oz
ppDCb1vJm7wTi+De7rVeajDryfd9PSWvRLdnhpaEZpWkLHGrExgQTumSGh1wYdZPPAVhN81GD7UI
pvyTIVFdw2fwzCEuNUyBmFaxbe8QgujJ22Bx4DSLBlHXICLBDqvJ0pC25Pqy0BNN2thwoaI8dzhq
8UiRK0TYgTvCB36ipaW2UVWgywn7sDDs69jV6JTRZSD/WAcdpuncCRUBMFxHz0zRJqYaTgoQT6Ne
DhY+UyLuubRDHM4FzedBDQlJcjtdrNmn8pkvLKUC0fBIjnw6FYMKcemFjMvESpst3E1U7g/AOoVr
28RVVSFOoE45Pa3ml5apx+E7MexlfIMmOnqPc5q2AHztodL/fsUDfLIUDJf7553pI3541UafopxS
t7aRqriSVN2YeEmB3schVhgWts9IoiF741px7U2mP0AuNZZbvwfpndxfko1wEDv7j8w6eoFR6TUU
uVzTCFqRElqg1SfkDpMQM08edK0nSLmTbzVEa3FMZ+9YIcA7iJEk7Pa645RZc9I6FPmHkVSANrX4
3v5qM4/uR81lI2zeTnY+g4JPvbFMbirDvlzlMmeaezcCPBI6pXQla4IOHkXVoAZmdNS+Dbm2xz6F
eVjkWY1PkWamsatMYS46M+PGtKqPc1DS6Fl2w/SY2VJ14zrs4mFiVQCr8FjJODd6t+po1V2fMpb6
fzXIeRg1lnKCiv95fmvZ2EXFpsIVurbDgr7R+A9iJmeokaOrdH3AZha2unH0Mxdo8MiKSGrE7oaA
nXEJXBrmoRXrsbBCkJHVKEOQd/TCWzN23818M7+jP8LW3AlEilNfFT0DAOr8CmAobhudIeHOiJsq
n0uUoyFlFiM7a+RlZhG0pGTDtjF9eES1kRwU4zEBRVIRdYXKc4W6wSUaqAXwC5JC2/aDoBer1Xyd
NS8v1hSVF0eMCSd6wLHCLwcAccRFC5WzP3Ep7l0G5iNedG0XH6uQauvyW7xr8ScKyrdebzyo/7zZ
vpv5M8J44V4EN3zp3LVHoMhHi1M4d9X5hs1R2vzsPsSIwJBDdPW24bdFUB1OIAqQbQFcGIdZ3K/T
DRvdHHIYp4I2xjAoTihzaulKFeOtP7pdIQiRZqMRsOvtgYYl80IsDaCQJ+FIH9kjT3JrBQdiCHNO
776GtxfSirxb4IeeCeZ9vRWRDr7UXWQLBGFCWCij/dumbQCKiKs27/KLLGDbJYCY9HCw/ZpRBepY
uYjXHnJ3Z1wv3hz4nuGXN0a9sDkFfeaswsxxwYwyzIuNtHp7AVDMh/CY0jf7mOVEDsknHZNaC3Sw
40ACyqpQj5wGN83SkITzPVwZcttP/lmkrk40EAS/BM7YZsG49lS+JS3ioz4YX9vDZ2v4V0GVUD0c
E+wKI8tBGNpxOI+2cVdfJP3EV621uUz4gebNZIu1x4YkRVS3p/w/0f72aYFqwAsSmQRCeNCP3BQ/
xtSjfM3+sFDhjMraWrYc0khtVzF2h91ZKz/SDRmv9ltMw34307z5KdkkIbuGkZdhaewEzVIxkxtJ
rSYx1PKMqPCHf6pdGrqe7Glb2Xlcq3ikAU2pJv4gjoqvnyRsUsM3mdaitfbwWYs741uuKtY6FUlp
hWlhJvB1Sw87QjsphGx+G8TKWgQpDQrXtUybRon4Kp3UBQro6OEiNkFzbvZeDe5QffdyK47g66Rw
zY3L3OZhAYRbs8dZd+rkmA6u5RMNiFDQ9zilOMtuHhtGRUYKkGFj/QAocBddDrzUqfrl9nd1oaF5
/hdxQwkRyI1CgxVE8b9jBPumXdZ1JpoDO1Z6ST47dD+kQmmLqwBWWuay8bTunhDb0pDk4vQRquxD
ndY29OZ5PDGyOAYxmCyMistTs1/Nx2NVY1n9bwgmyCNIAeMBe2mv+Hr8pw7rvrhzZJ734CWr58IO
Wwz8pRB6tO3I0WkvLpMjZjDLtRotlIWL/i34+dSQ9eDVHmNtX0OBHW1Tgceu7VkGY1hnOVBfJeRC
o0D+LYeGOy7jG4o34UKPlHGhsjN0ES3pu/s+ABjpx2QP5LTeJsQmj8ZxHXZ5wKrkk1MnkHzsT0pF
N1OJ3OMXTRwYEswLSc61iP3dpruDK1Fr2ZKf5KslVEZ8Zj6wKrAJXtfq9aHhI9dOfjZIoB9f3bF0
Nim7pn1oY3DTGa+pdIZ9PwKcvb2gViKct6W3ksGMAA+r/ryGb7A02yiIThDz8iGxQXPAcbdRE8HW
lN6VDIBLhbjNPDM9XcGYUL54OPYSJRJdsJqTDCqV3wQQKgOdRPmWCEMw7KpSKPoeuepk/NURbGOr
L+3b5z5JmoHNEW/1x3NizMfWDUmRZsTYbDMOaTl/2U/kNVqUYs/K2drsJsApiAIGXEi1G9HUCI+l
CxrmFTpvSSQOCNPGYuAeVfojI63XCagjkEYM4ydzN6YK2Ze3DCOXWvdJ4n9mzyFdlzxfesUmhvv3
m5eD+9TjCLRiPGoYFF++PyzzMvTH5VKw6wL2tNEQCE+cZT2hLY+xQL29RM2Z7YNFPwvjQ84nK5h4
EaVSdCsGmFR8kj0ITP39zUG8pHiWNwRWlRq6LJiaRbEHlKMiKsubXLjXtn0KR+VFoUpmzsx7fHgl
Y4I4/ZbDQ+eFLpnInwDuI8hAKHQhpaIsMe+aqgTsF3J2zizRXaNZuC2d/eh31z6fbRYvn23jJRqj
sIlz/aPUzc9PrNV7JQHVbNtLEB8E6xUvC0Usrik4Vy1G/dFang09ggLD/sxNu+0zOZPuhDY2C/kR
burBaNFDOBM1WvDDg5RvhtKBtAfvlgFjvmwj3rP+iUA272gLOWoXhBIfJ04dstFJudRbuulm1NVj
uXEsgvY/+w65m6Ez/u9X/1pzRo8XgORysu0P7z0fQsfUnuurtYTbgAFo5xHmxnfo+qPXqgB9KSka
PvLSTOtj72bOLmJp1LnkKKN6ijK5pwN6VOw+VoS+pqw0Ea+c5bqBe+96Zdo5ddHypyjKF3xXXqHO
q379GXRoHdmzqrzZpUil48DkW/Q/dDOktcCH78A8CgPvKja2Qjc6NNGJMT5ecFqseEqRSF1eraHu
zbTErT8tSyPhCkW3PQ80bxCWrCjNPIfOqyXfR6nqglNej+aQuq2elEMgGQ+WG+fb3LDPBEFAgECZ
us1I9QZHQRI0aB4PkTM9vwTGk5cbNmmoGpSvmzbPr4DW71rqGCL3VFM2+FIwOUmqns4GcN/ABevH
Q/Bw5VWuSgXegVelhnxXWzUbMJ2xLlHGpE+c6YrkFeLHpLbgFxeZ1KJ2gamjiNxRwwP2V13gQmJn
1gk1jNPfUrWfqj44IO7o0eBMUiiWGFGVB5zlwZMwDT7o7KybsobhW4xkUctWPdN4S5yZKQ9Q0Euo
P/0WlqCqVLqARVCW8mM+4KL6zR7vollWj5zPDG7EEIQLPhhdjRLqNhhWEPV6OTRCPNfVfGtLUmWq
76SFHQMJjbBI//GiBie5Xuf1Md1MwmacUVjN2tRRNBZL7rsPQxk8e4eZPFuhTJi0u1KeqLFeMwo+
eg/jinUP5ypmMr6W1Jm/TMVi/Oc9oheBl3y41JNgn70Kyxu1mVc+S51Jt8WQLcpHRzYvc6TmKILX
dnRdrBpONygabhGfF+UeEiP5LNm66V6hREHvgeMRrzAFf3FGCcOUi0DhcnD0b9RC4ds7WN4PUCDs
PLVGt46BoPgV7R8b7gh7Q29DKlxrzMhtt1kag90bPv1tNJw8cG0ijTWE7+zipKbbwMhqil4uoYnU
bzMxS1pw3b2fXPCU9HDi1Z3YIodcGddCQt2zZL6YgjL+M4ZZiXgxshUdlw7Mel/vbVJjcM4Z8XzC
+HG7IINJUpjKWZmtHCG4oSAWkKPmngO7rnjxN2TMxulKNbYQGPMIyT5gikYy6y6T/rrQ6PmM40tM
t+Wa9StA9ao4ciYqif6xXWNXpwx5ccgfCRm+LdD4N0L8z0XtQWwjiWus3IROHTMT6knNocxtUEk0
dK3lEvhTNRV1LaO4brvoQ1MXSKM7O9pp9ea6jibuvr1m+1iPAywRAsYKswGeiRYk5HtlhAUKI9Rh
SxE09ei82W+FLNTewbwgob3O55OlnIbDJLhzaOTwYU3b19Va96806bti7SJyXOYiWiE9HFYwdTuc
JmGKcuEWXNUWEm0Tr7lCq25P3ZuG6BE4lax8mFL6n8tktNKDnnhBN7svr5/WiAxokzPLKPSuLYE+
v2w2qQ7pDIehnUNKIm/PJAH5w5nqBNdDOoXukiNX4LonBK3yHl4qMZ2lEcjPYvUzJxCjWCrI85/w
8/KQizPAjWsoB7c/6UlSEoQ/WejSM/ytzi9bXBC5iHiw3OyjE8nDyEsjNWQG1HFckbLhOxVzKXVg
HHY2IHJxpbvH9GGdVDAUUhNHZDpu7LUc4IlYCeRwqpRgInPo9Sa51LiD4pXiBqnGnWy1zfvuP/g4
AjjDH2ypzGinFVGadhBLDkaGDNLqMKWGzEVODXYkVnuFgMTcgVLW+ovAGtkWBp0phtkbYhgyQFNN
Sxo96pOkFo1VEfR8DgARGKNZMWjR2DtExtcxjMGl8rR5ZgsK/78GcM8FKfTFqsq99Q1+MIGtAEyt
yEBliMUw/yhTRk4+XLsQ7oYj5heFbC737DkYMV0oQIkfhJnxAx5IxNhd4E08gicEdgjME7Ou6I6H
x8OJwHDtOKRFsotl4/fHvaBNZXoK4VR+X+UBybnqRXuqLmij/u3OQFS2xCXvxFvGGEVvvKtQ/HYE
v/KQ8nuhvLPaPQwmj7iw2oGe364q4nuWhDURTUmjbOUpx4qogMF2lX4W9AGXoWvvTSwt6uVRZJM0
1Q/vqG+2UdW7x33Qc/CNTEpwcF3PkI1RuUJrYFRXLcb8n97PfDL6RWJEdOvqNoA70eBM9nx727Vw
OuS+CGxKhIZCVMpNLOfUn3yfioan5yLSQ/VmrvYEixoVGlVD1SthKhPB6Xo0SB2d9beCoY0MtegF
CJbW4ad8UYvP6lzGw7CRtuR4WFgEoOsVxScsijFxLMCheiOYGFvwwTPomkxt3vtgfL1Xq4NVfM/G
aA+huznGDLVfIgRSwl8093BCtjwf1Nc/8XVfBcMnSOHavCKYepgZwB3vdJQW1rrGqjCJySyNcgzW
fgoJ4v5j7j7fXXevp8t0fAqg0Y6mq/IDaDFs/WFJlZY0J8THJQ/j3nM/oGxXgspFx1SanSP4FtDC
ZB0xUp+nWEpk1C9FVX1JdYspfrmlNZfQ6QXQOs5phgKlMlWz89wtCKmODhSB2G1JfXHGkbiqiLxg
qAaXm1YkFATg4rwQYdPX6b5NiRiEQS2rmSYap4KzWIt4q94FfkwbL54Nedqc7DZOUH+B0PCiswhg
gYiPokSe3MdfmmmkW2StIc12yGW/u4okZmquT2arjGIJ2xlOEm5Joxb3nPxi6aEoRMJrcf1pMFQt
vdevEmUyLOZx/ulC7PwK8FdWAt6dhStrmryf7i94IrGlrl3nsK55cCYF2ogYagIUq5SStnNp6pgo
ZRSInDJhJfRgpCOwaCVG1nWRB67jYZtEH/20yIFQh/UYHcaUmWGOBcny3dzN31M6vqWnsue0MmTk
TBa32ngzKcmmRPyGK9+fNBwJdHwpfC1s261zqR+70eu1sryLx3OCzHxo3xGm/S9Ftw+VP665DeFh
eCLA7xqW3OiiR4NWNwAhFoH9jMDeyBU6ZNI/L16Lh1cWI1koToZk+t6L/TQOxN65Sw4eEv9UYCqM
iA1UGZYW13lm2XD4G1ohSiV9FDAimL2MfIAm5twOC+ltwyy3uavfxxuP/FKjQOwo06HIdVRE0Cuv
CDvslzDEozEpv14hW1IDFMfq/Zf6aYXToK/bXrtuH4ue8k8er+bqkUwJwQi96RZEp/6fnYHfb1w8
+GeCQNmxUvUwuKmnn/cZAfXYipXFpWWjK5IBHJQLdRzV5XP0eYeV2xvisrIsWcJePxn8IC0Sew82
hk9IlV92rC6hV2E4jA4rLl3wtYI5KEXxSZllX/wY1SKFBRehnbVovbZxdhwim7nmCAtNRU9H1N+T
zi79Kb+nbckffTSDfhZ0PKyXMcsI6tYpee6BdAqIzzVCCjL6w2VTmhiwJydPBhnhQnzlmWTmOcsw
Q3MKBtI1R1id4lpix6C96yeZCXYSYmMAiavXMkRwqZgSXTGFXbKioLlM+uNRnntOCGKOo7tS9edP
3DJqUmKWfWUCW3KXnMTytwb6xlkEAJ1khivQiHH2pZp0p0o0MKZE+g6E5U2r9XkUr9zcW9FCLcp5
CaGN9amm59xYwyQOIbbPrKPJs/0XcFeIl+zbxos7VgEqg6TX6bQksvA0vvtVGTQ7lECPn98Lzt1M
UkMeiApNNp7zm9vsinkrptRUvf05ybsykuwjAyxWQjyjaS4Lxlh6RvGG5qDdD/38ycGw+mcheNqj
k5b0SuWQ6AeeSyHtgmDwvClymZo9i1UUGAq7WEVoYQthaX3r6HcCBq90ksEb1SFyTxGczFUHBEIS
RdxGcJYHEsxRpAvDTN8btg0EkjnnOA1F6SdTRHa3w7vcHmWmUV4I7cNzUJmZiePOyj3JYliPuqH/
v73ELKMRb0xRFgL36M8uWh5+oduG5dMMPtTKeSRGQ78w2cz93vHa03XkYFwAfeolywiNqpGXdnD4
tRhJMw5Ylsaqxy+mduGHqRy7crNGsVcM3Mgi+AIfbL2lgrQmkXOm0mOMQchchZ83ODH8/h9n+Z3Z
BeK3QzeEfBR7CgBorOF0z6gH4c8fo4S52FP4YhGFIUPAEGVQbORrSBu9Z6j44S8KkyKzy2ANRHq4
Of9GNtYs5Zv2kLa2jc3ehGuBoc9g1cXMk45m+NNWesaXJVePVGNg4N22p4nD0I5Dvk89eLX6hRz0
yEXUUcpqyLJ+sh9rVO7Q99njP/vJnJBJgRnZt9QtibqscOt49AhjLztUTDP9oVcSQAaT0sU0Pv/T
Zpg8BFsKfzlKYMgGAsunU0sR/+KLUMhtibGhbca8KSs649CD9GwEcZQDwqkrpxYB/Jle+16VoyJi
+/smw3Ci87dzdFY5AqvDpP/9nFOWdeYJywnAMKPS9QKZX8tpxI0hxEGzvz+a5JuwSvV01hbW+SkT
BUfoMu4NSSM9g9frkIGtAJKUCmoSbBkWvG/Ax0ZpAXyjrDCBPFKOqL8KjCq/0MW6BTmV1w+PTjlk
ixmOjsUkZbjwqHyKJ3H62q1Ol47Zqxx3ezbo8tO5wYA2gYnZOn3jxf67JvRrri3bQzs/pWoqasqn
AIGJUgDn+NZkG45gbk5hwzhJWIWXYlnHu1z1G/uRq1K1CoNTZIbS1I+MZ8iNSp/6n83dtLTPTfOh
iJej0D2s27pTnZRu9UplcE2Lx2UTK7qvJkXwJoYWP3BsPAaWLQMHz6JP2BQBUQ3eKheB9DC60HaR
G64AfE+da6s64yMqhCTxog8x+sptajmEohqvNxpFYjVvtexhq8OoOUGcesm5kmV+/IU/aRLQzdMt
0sDn4k0PIMNbPPJpNd6g9KF2nmWee+WjkQUPnQSaN9c5R2TBUlLE458Im5mIUr3Bo452E38fT5N+
NXtrlTDdGJnPp2ARNsLOWENLI4/wYRHEmwxMhD0T7PsLVqYsxBSycEEyGykcn3oVAxyjTExQf3NN
4zeKlQrVHQdsbSYcuhOsVo11ClMqEmoiEzGLwEf+waVFs61Z6Sz1IUWYE3XQT3M5vE0BF8pkvIEk
xYkvTfI+3piaIkMlNni17g7tOXlVZnp38QGCIRWkiKXr7lWhNCfqTefP/nciTuixwwSdk5eEYJih
ksfx4gSXRG6bAAZCWxxIRgPHyZ5QMmR5vHbBrjbM7kUmgpwwQMe3dagVHox6Yyc4PG0vXekPibVy
aUjnm19d+wp/Fq+OtSMcZy4g1H0Bzcin8Fh+oNh0pAsfZDA2GMeKUT7t/VsRpaKGbaba5cINuijq
kHf4zPNNqANQygQEIWglXaTwxAFq/NNN71Yw8q9UWk9L5FbgMZ2iUZGuuU4iunz1KbVc1IGxUNmU
rUzcyPiBjNvp4wQcJ8EGUSqfCo79J7EbpzXaW7m3QKf9qzHKkbgzkF5LsCO9nVr3ZK+ZJn+HtrtS
IOQZyoINithaiecUwUXFm0Yd6fBRsGy3LFen1D6RSIJky0lAskU7Unj7UVEFKYxw5zoW9Cn2694J
oelK2O9NYPsWyEx1XSjR5QrENC2+zZ8H0XZJKweEy517agoQwNSvGxSSnUO1ijJTA8fnIoWboTcf
yS1mbbnZ2qXIiK6X4VmLP+ftxNqoH4lXqYTq434GX9jiBhPeNF8VCZRMhWQIMVVYyELx4hg2rIAA
iWdd/umVTYNMKpWZ6i0/0HwcwujXFCmlXoSE2W+2fFAGW+jMe6gi8ShxaVYFe7jp69VFwxl7ovNt
0cB1pjpK2Tkz2uU811wRJWSaTPdUaEs7h+fSTwwh4Ad7QB8dnCbvFp5W3vumx/mkDyQiaunNtfiA
G9vTDadH4G47G06WrMuHucnsXZj3ZOfMO3JQpsm7UUIIn2njaLB0b0eJuyk6Na2sYYMXhoeMPpFV
RejvG0PEM0m9xSMIU9JqIJRC3gBypIqG6dFZmuOWpzJ3kMUociDbnWXRvgR0YCj/znRnovZVPoDw
+dvVxpKUqzdodkAhXKQx2sxcJB1GDqOU84Cz/Uy6qYqrUSu34i37GE64KjsSkZ4xVRX6CpWWr5J1
xaJsQVj3gBycDnKCrMzAeqeUMcoUkeMguGgHX/hgCyVTV1DjuuXRILw6+RrvlqWl5DLD7zC4pBtT
iSwfs7ISqSM2leKs6vGgmcA3LL9jJWzZAT6FP3YvG2wDzBY/dieK2Q54cncoalEq3Xtruh2rajNc
aEXIVsOvz8Lfkv0238EgCKko3E49h6LPS2tgolEN0UhB+VLr34fOIY4NYGwuHPbT4o6NEtkPjp+g
ZTm94rhRkswfKhtJ9qmELmGnZBRCeTrKyb1qgqdehtWE8Um15jlW+S1u7rq6qYA0RsxvgM8WF6oR
vXBflahhbtHiriLQKZWlwVufeZ+RkrgI4qEPSfzOVHQFcfT4WWF+EKcEFFzUFqNLi7FA92QzjN0i
UIzeXCK0ChwxRb3w0rRvaVVBe3SCBnLBDRjqJFyktYs/NZ7zvSYrOBbgWts0bmC10JDafTnwZZuZ
G5FDV18gRlk/OqP7SDjFkIMOI9mRwF+KjClJ6eTDQUQrLAduHp9BGPgw29MjmGorNijTxwcalGFi
rbKCZmty3LpkjgXc7fynvjkT+ffw1XivskgEnbls1d4OJVFuXI/eUjZ3SX0USaodXylSlQK3cT38
aEHpzlsBjGQAaFDEyj8DYl4skHSVDXYjWb4sz6DvvovBQm2IfNgR1eM/21OSDGtaZeKYtT4FNxDG
7G6MNyBVL5BTxtn/sUPNYHpQOrrGosX1I9zLDGdXFnvrdzl7AvXUFkamJ/D1UUbaHx5qXrybh6xG
aRaQE6Alry/myqQR5tt6Af94kFOMLiRxCZkutyAwQZtpwv7MbRkkDBhnuVdDAWFEI55IdVJlpwlJ
0hwW4yeQWeOCsWMqDqZjC3oaIPJY+Re3+Xce+xynq/+Gto01RjFom5yIPVstCH0KBUa7UAGG5Yd5
sUdkgO3m6A5rBmbsGOR/WIYnzhiQWWsql1xMQLr2WAW4NGbnUfKShfzSgW27EBbArnNzIfjXMRJm
t1EFZg/f9RC56th53RRQw0TWMKyb8wNfUb6xAnlmFJV/7pSGIeXjKEJAlhOLi7sod42Bk1MvBMzf
SgPGwHSNpiGEcUUx4WQMl/i+PZL4pq/1XW4vOexJJQxq2C5svc378oX2bfsfbfInRyubZT0C5MTn
MWiv0HxCd+3xrbuMhF5DInnvghGoPP7ZOhVI5JmWevpuPDZZ4dfEdTN2a7l2nF5A2JTQun9A35kG
4ZNdGWN/U1fw8bs4ei+g1D8d9d1B6RU6HfRZgc3o++rmWfJwGtMRm3wMy1ax70SEGW6ok53MGHuY
1MjN0IKMD5hH4WzMW/GOdJcL3d9yN09K04N/q4tmV7FgKqRX9kHdTYjATDMb2PqJQtpeeaSEcYAu
8CX47/n/fMxB57pljs+zhKAxJ9INbbXMjLy7tDZYPgsBZMvgDeIKI6EAdWmnLVT4QJtYOlVLtU+a
LP45V9y4NHzDJQFWmFHaeiWgrVcBs/WJ0PjvASbmaEnG1gcK3I+wX8RGDsU1KIxXbtA12d2hO0kx
Ah48LGczmS8PszmKPBf2Ywi6G8xBpcF4RL3A+cndcSLJ3TMKo1L+yD4Eg/qnrF/K1JmsGF5xQ/oY
s7w5lyBnL7CbvijHpwSK9FGoQq0MVn0W80f6+hO06VnSE9cNQK+W8aB9cxSvXQeiU3LWsTzgkypb
8UaBUQ7NGlMmf1cJei2/HnC4OMqjN92qci9MiRle32oHRS2l+TqiTTCTLIBUBUUZZng7yTRz7HaL
A7xTzn7nlNGIwnmb5sVA67Kjo/l4Vtt01P3lnlPr2RROuOFmAJ7X7+E+9DmInsXkmiG/l0NUFYsY
bZFrtnWOn2wxlkYCIowUEoMuu+cUuQsqMmeQjmTYEJWNsOhyucwSJDwLYEh3L6f+eSBO/G498lNs
xq54fal3NY/Xs1THAvdXgFIbmP4fnmjekl3Zox/IffKT3LExB23+IHe1cvHDAt58owhSx5yMehHz
pSn5JLDzzShblW6MvxnPY0Q13w6INQLTt11ZwdknfyymrbEe+uxkUgTavHCHbCuOtx1C9GlB916f
vkzxMmbpqZI8IUbgco8Wdb2QmlFyZ1AnTP4BC5/oXRQWAAwzsndIa7ZuFpMg4CqwDcDS9+kpNaJR
RhQe74WeyCI9s1R4wm47mKOYru3+bmEBDaO06RrHZ22TDP3f4pqqIu9L76aNUmeAR5NAILo+IA4G
hkidPmcIFOVHMPudyY3xOmJdRxWElRyk/ne5D0cyTj7RyoSrAgThIFLLFIOOVRmguCwTsrV/D4jR
0WWYK9bnmTwgF6FeTj4/tp2L66l8QMkZ1w6GnIPFi5zoq95OmFOABZfN8CWOTwPYWXEOsornyhzK
Xm3d5yul1jFIZwBmIhe8BRqS7xQkW+o5ZN3uGnBG5WEvbCyp/vpWHajjLN9FG5EHaXZ8zRqAEA0n
d8w0PR0d7CLIw4URZPk3qYwdNojXpU6VegKmYTh8lk0zeTqp78Bk9kRaj/IvGKeZrJz535Op/TG9
KEenCnWbDxwB1K64av9cWC175xOvA5LtqTcOt0cnNiT5XH9n0tZq55NsUwm6PFHu4uejOUF/rxtS
1F/j/VKvVApvxLeTDvfGeGJzZSBoiQJKYPareVM9BIDXKLeTLXWKEwmZIwhdB3Vpn42ckgQhndgP
N6c61IihkEsI6JdJeRR4q04bW3Vvqp+Vs+SggXaZ2J4w/g6aAk1oYM1ZLncBCtUMDP/ebE3iySzk
D8FSmYq7Izyqwuhu8FP+LK35CWAEgpx52nM8DtCkjDblgv2pFJPl7lCWBA3+R2Co0VtLHH/dcLD2
dWMHAKMPpqwFkzvEpaWz7HbCDYsG7vRIf2Nni+M9raCX2IfSfpgC5R9qSaSfHtraxRKT7pJ2UtBV
sv5dxqgJlWjBERegmEsWLKL609V593OtH07OCAdpG9H5vTkEuHwu2IgnKLbkXNvkG6hjU/k5gXL7
+lfg3xrmC30Unr+3FrExx/p92500zNkg5/rdc+xRNSVaI4eQtC2H61fOv/2T+yQw2k++RCbf7G9E
S/b1uHXZrM2GbMTYKzoyISpdSok+dQY5FSAN+uZsvChP1nBhlGM0ck1/V+LGhZ9QYomLar4M6efl
ElzrQz7YuxD+OnMjhj/yLA63hvJ7aDAzSjO+H883nbL5S5W3neOQQGLOZ5qVtQssBXQihq37jHrn
cj3EHQhojNI4M7HhYbx+RhdWePx0DQvEDwTvnKDxQclDYoxvI3OUvfmTZzYmKTgOS6SKI1mNhJ+W
TIHupxCsb8Yob7S2uRXGsuLp8qeakO+3l+EKjMhIKp/KBXE12MiiuXb8wnM8USh5mPuRuS41noWD
IbVCWoYicXBzErsSp0BdCc8Z01QNoaHYxYMmUxxY3WJwVcSdAnyPNB/w5MdjiB2DBKzqjQy3FYm2
+iyDGEsk+z6a1xrMkw4/wHBnaz3vgYRL4KTRmUIPQV6DHNo5hc2U6qsyj5VPtLlf0wAtHnPpthO4
X8xLkVX61UFhoKL9EvCQABpcBc6WBr4PjxsguHrktP04mJVI0uAWJVHktQTcSxE+ga5u+uzfaG95
+o4VSztY0zTdop3e/7o448O0Ehe/VCnkytyK1MrGa7R/XrBe0qCd7iYquYz0dbQzhKG7MjfYoKX3
b/zVCYLR3oCFS1mD1WJGj+N/S2wflBoEBgYczBkvyg3OrADFBf5ZhDiUbUyt8QPBm+XGs0cGhEJH
xdm1R19YYp4h1wDmfcDsQ5Qscp6t2p4PWlzjEB/7rCgGmQZqdXQQ6ln4O5EZQTWe0ydUxNrjrfdN
FwXdVHa7XWRGo21Mp7DyWNPbcrPGXhw+ECR4tMK2byQpxxLv5mV69iNxwYfVCQ7FRkSpoUvF+FwU
VPdFy6yERsjgG0PdHPi8VxOaSRNTeDv8XKC4xRcShdV5zxpxkZ6pl4CvFHIW4fr4TsnLMAd7rySG
JCvRQCW+edxboj42IgAm7bWwJ74v3CAstdVDHHC+P1366T9XCiPkXmaN+R0GTr/Y68C+s6r6Yb2N
glLgeZwAA0S62qkLVacL6soMzUvEBXtEb7m9Dv0siuRnzJ3oCu1gb7LgbpuY8NRGWIbUcQMpRY9j
DDQftoAdEFsycJnrXNjMR9Yqi6wJyNi8rAN65mVe5lobQdXIDypMPjboRiEre0ycn8GBIFSXuZU1
SZUyvg3dZiA8fIePxg3w42E12RduGNEs2VidNkc3FDoV5I/PsIGKhHeNE1o11xMxpH0mQjfdM9w5
pYJbDiiDgH76J+DTK1t21Ceqh5xnu1CgYPRgh96/5uKDm5mXyWs//qaQDuF4Oi6LiBqDVkKV8qfm
LIe8qRRxrWWc3nRhhjyqmsiFQxzRwFIy39dxsyuzRdYKRTFSVRWm4Kyf3Z3/RaOFbr/xWyB7kEaZ
k3s7C+Ay9Uee3AUtRcnamEImDNMKl2WZlaQe12fNFs3iVe97e/liyMK3773yvn1lprOeZkgMxfys
p6+RUZt6maRLg3/ptK4BROPnDvcpEk11fmTjRRe/c2Caes1Yh/InGomNfwa5Snx7HygZp0eqYx1B
l2WJNvKbPpqcR35vFd+P7OrruJR47S7n82WaXv9Re7hjWdx6jDKHnr/a4FyOsO4AP654jBUYtmtN
IDRA1VsUCfQRb9juvhFi+WCLL4fL9P0YAN2tyYH5UOfaYZ9wvsk1f2TJpXMSv/CSTeIQtlzyxLxH
3lHl3PAbCyu4zmkCZFREhkQKgNfB2lbyorTMRXFIr52A39nvvcKfVawXVClteo4SqMtq89nfGEfQ
lBcw0IoLzfkFhlr4rJyR4Xq2caL+urVqNhwogbpD/XD2zMyAiMqLQLCkQDtCrotv10J0JNlAwuvf
e/Dhmzt2OPmPNt/SOfew3b/dIzqBiLKZ5A3EPsC9xUWV0x1zRvebsSyzgsPvR1vMSKvcDZil8LKU
qw/3WTnWnbEBewZUioCLX505twR4EAYJKP7/FhUHDRdrctuNf1RdwKe1wFAuASY4EIYHn0QU0m0K
PyGyTLBNTr0c9xznNnDO00oW5fVcZWkb5odVLnAcI761qiVumo+V8SSL1oLEDDOWB2futGPHOBlu
l1xRyRWbDdjmjdWM1YiZBED+94H/zRn0+1BASJIPODNy+zdaHPSbPKSz4JLz+WBnajLc/morC7KP
KG2WDfXHfPjiugRkL6xLG/iflV65JyaYzkAwI0eBd0FR+ERPQmOM99mkzR7JlXIdUnxMaAtT+k7n
fNCAPd9+D7ahl2Gm2/VZ1YWMGZKavY7aLDYv0wjrcekGYRVShJQAio2AxgpoKBlgxM9Has4p5XkT
TFr/Ac6Im9csIvUwKeaZSaNmrS8wGCoKteidusvjPzOE1VUr9N8R2Zkhp0aK7fk5flxwQ03sWWLw
O6wnSLdF20KuuinM7fkKK9cWsfGYRGEo/6wlYkBa7aoVA/WwIyo7XLMGEKZaois0Cv3pxLFWEnJG
5iNphGxGRAs2fGF3c3vzMIXJ+KZ1I2mf60/IR46ypDQQyQStlWirmxNTMdwSfbGOqE+GN6gwxvpk
aPczz1pAUfKr9zROGcopr9fGn/2eGAiOogy05POxjWvQP7qsmYf1TdQUEuTEe/sAFw4EZ3fK8eia
6KZmMlqdExZuuUMSzZpPjpkFFolzA2hSoPUNXZh7qkYBm2KQ4/cnn14dCrWKiE9XLKAsEyQXxwSE
PN3WdUe31bvwTMngZb5OLMqyp3r0ZyuDmfPE3KHdmf/lFTHEfhWHCJfpvzSMiw9Jx9BCV/+wQgd/
5ttu2YfyIzJXpw5Vq4rF3bk57GdO9Ow+8b28etbPbe4T/7AnKflqb6fexBPapj64fCNtGtWmnYyW
q80CDTL2mEcnesllzyk/GKHsTRfSu3iOvr+v7EdzmKUOesNe7iHUuTXLF6SoDEIpUT4KYn90LJZo
jpHQWl35Ivg/C8m4o2HuDZByHDh/653oFXGcqSUcvrxq48a06OfHT5mIglnUtK5n/rlgPu6G9r3t
LV35XhxpzcNRYWBh8/vy+cWEEVlHXX3+aq6s9euqkl3JNuDTT2ukr0JlGQsvO2Prlph7uUNwgwj+
OlX2iCNQ+OUkY2FK3HJp9lojQivZ+uVx73CTXUen36hHTTTlrQVkt0k7rHLa7Svhrf11MskG5Ya/
2HY0XVqdL2WcJuhkazQEQzWMcgqZhXXP96ghBera12bKokOXwOPdQZFW5stZdPVsWgNiw1ArCZvo
cWfrcCdP4Ko2hAt3BNP8VrnrshQbxa4CvSiR7ESNjCgGOmBu7pfdhEBztt5BKeDPSe3yYWXfeL5G
nfwPWYzELto/TYcuUGnLRQBYpNrw3iMB72T8Ch4RIpOUJRtbNDAcUFWfAGQqFVm/TRseEmh63Jls
QdG6rjb5JZ+cYyfQLUyyTWHo0drfMnko0TGO1LXc03tbIRb8wABws8yNk9rS2NRqAk1EVtiEaV/G
PIHwFyrcndJ7QHjb0jst+ByHXubpdhlDXetDkYSkXJToFnWSw3gMBKeTmVk9Xs/SZ/CFrvP68IZl
QkYtjyGcWRe6gcWjsYLdyGiXK3eha4z/5qihsopU1//op82O3UGjBP9dMiHvGZQYzOUDQ7uhWkno
x2RzAKrrTd86sKJly5CQwi3qTlABQq7T5FiT0+LkPfrTacfDxvrVRsFMd1iHy+VLvsUQ04qutQoD
1hlvzZIwQkaE4KI3YRDYFLXj+qlkchcsFITwQOATKzvrrjlFEy7FlAJSMg+r1ghW1m6hmbqfJQGm
cYaBFjDrTzflg1DZNlwRqY7UbTgHMYiA3uM6gdNxmc2oJnP+lxlzwWKY6kXC65Nntk/EIqSTip8b
TVgdVlGSUuAyCj8w02bYxEXjS1hPCchpEVlRyG1bXnJrbpwEwst6bX9TY8cfKWPf5eAgys9HGqKH
GmPsvofpgYJy9jmmP60PhEYKQe5prdJk1FT5sNMi8E254c4RqXsX9+Cf7xP6ChiZdAQ1Y0eOEX6h
YghQGqmA0UCbcpotwXki+DroCyWbBvny/YlGt5hDML7rYNZG1SlbCJgLiAQDqWJCe+uBz2/l0e/t
mzZaxRjfB+1ygznH8pJLZ6mRjqJW6vd1vmgIlO0EcK6+M10E0EWZ694ufclEzzE+0jLDikMqoEfW
lk5At8rkKwFpHYITJTW1K3VgccEcMlNP5seWi1yHQwR+rD+7U27XU0Jjh6qTGd1K3aEH3nBF4/ip
nVPmqFXkJDUWpWFoa7RjBNXFvI79yoDI7EipVb8wkS9trrRZ9MkuslBXBidcPUfnUSOV3DiRHhxW
JwRAJORAUAQ937JrOfsWz54AVjM1+y7RX4BaZ/X+xVEehR97S7Fp918ym7JFolfc+zwr0XrBP2TE
dH/RGukEgAawsNjeILv/Npxe/QKFYLsBivFfkj0quH5hOCdcvpbZoOz/e8XpAlP4mhuM+Yyd0lU9
Hic9EMYyOkrda8iLvSa7IddlJdg/AI8AEzRgK/A/cIwPHJZ0J+zQNKsAhM9Vl01vn2d/9l6yHxAU
DlDLrSSOiiAQiaYgzpa/jMOqoVK3v6ezFHueoLFVRlHDh/43VFHuclj5SlfM0HDWDD9rAURRXkYy
cef5yy+vCY8IstT3fbeMhsxMFktBLS56oISn7++Uk7ELu5oKonPlmcn4wSdRBxU5pKsLFiw8ZVaG
Mc/pPA80j8UhZoAXKYClZawes2mBUIOm1xHqufrmBpyKAbwc8luVd5Yhv8wV7ni4F8xRyFVaTLiO
12dfvCHIvqBohaxTCc3i6tmbu3l+8irjuYZCMuRPYOTCeyZq63xW35ibuumgsZsT0J+85wGivP6Y
TYOuzwBw7FfxM4kmXywA8h4/k8Wa31Y1hUs60z8S3MUPlmFbahWuwYKw20FTDxtKvY9sXlUQQsYs
+UJ+feWbVESA1hbZ+HoKMPbFIia3gRKNW8neOC1DHSNnoJXcC29HrPKAyeMnezQ2IQUmbDxoc+hN
RABEKtNgULnp9nQS/aWv0HcW2SLeOSobHMBlmM7lyF/UbcOD/HmcQ5Gifw88+aFWasppNA63wKKC
wrdwn0XWz0PkmFX5hv5LSf1ApVn/VJRQle95Vg1TKKYWPSBEhSJwjBuKo22+BNJBNR+/SN4RRHtY
ZQqZxvWzQhLxgm0dHNeDBqovNF89xkhSp6NX3q3SEKx9iiuEBWL1yAKPvHklF79rT+yX49RupQJo
3PbNYKi/Tnt5rhx5mAsVxLc+RGipihipC5YcC6/6Q6b03mWUKP8opJCqRXegtB0CUS4HddCX2vjz
ZucsQ5vX64uO8w/oQZ49a54q5ZVdmOJ+zWf2YfYKTLd5wwmi4uCMlpP5S3npN1gSA6oJnLhyctKK
Dbzs2dVkDc9jiRi8N81JqP7OKbZo96XbvP6Mgb4Et0+r2050Pj6/CK4wbl48K745ft6sivZ3PEjN
DdtIiCsZkopYYgpZrjxiOO8VgvZJDjm1t9azAuWqd/GlwYLlJcqtG5gUlwYDeuWDVDY1nEcyB1zV
2EwRRXVnbLUpJnziM678NWGYpR8zsP18ZuITIWcBRKQdxOe0sPywMZpDTiB1QmtNfcHaIAW3XwRm
7dM6jFOjq9Y8E9uU2jmLjypmg/f+o6nqOtcg2dw88/O4FPPhoj/PyCNeBAGe6PMG5p7JqYxcA2eg
oxgIr+2FuA/r+7if4kb9FCGlHBB50ZbvpqeKoeO/JVEbebt8JDYEscPv3lvH2+kXF5IYvZ6oiZRr
BMc1JuZ5zbL9Mwyr0GRplCas2TAzz1Wn5KbQQVGqnia+EremABxp5wAi8h4E4XtYtJb0BJSEJQQV
/p5tKuyIUOINIZKt62mg9X4HZYA2dmfvB4hzaWMFLL5ZAld7Ak/tnAcjbYomYuBsfuP+vS7zDOvt
ouP3eVwtVJlZbvqqwTgWXgH+Io0dphu8Xwvw7x2eQcJ2spfqClK/oUk7s91be9vZ4YxSO1prIXT3
2IzSyeeVl3K7AWowE17dOj4Bv/5ufY2LOiKSL607jvRCM3gVWubLmWJiWwIh0Jk4rbNIM4LTGWvE
3aey6oO3iK2aWDnuncuePlQUVGh2uMJjFXAqVXHCaxw0XE8rlrXRd2kf0fdeYLpU6/9IPmFnTVI8
EK4428uHqd0sytUkEM/Qe03Oi6HZofeeAsn9T6fQh7UUkUSJwxvGYT3ZsFIubRf1IUFx5GnYqHwX
84CwUo7u1lVpCLgI9esPnvko77PxBFVXZ8Jmd2ofN483POI0+3TEVHtr5J6NtL4MM/TcjAKQNVJO
rzX1Xs+1u4pLYt8xty4+UxOkMEZJVm8m2oPSskMYbCmHP08VZFU06euMI/qChjEHXONgQPiztIJw
LVnKkI+bR75i5XTifTh5d0ZZLPDuzx2Cy9yZMcSXQGGwQ8VvVfy42Rpxyad34xvv6uIMwWQrF7G7
b76k6Vo4DOG0VToPbWQKY/NvguYH2bs+lQENSmkcHpJaUJe2XljW8sUhNI19sQHmjCjzomr/vZR2
nb7iYDVSh/IW17UHsj+DRBg379ntkeynWaoVdl1Wu0OIDeTdF2pvts9hLhOWEDhvjVvTs5n0bUZI
4JBk/1JL3tdQtb98ylM8hTAjQmrlG2uMUChtekiMPfZ6AnETSeut0KMsTT3AyjLah4PAeDAUaVNy
q2ZKKsHmcOJKQL03yqSGG47pFfkpZymvnCSWHgvXyPwOZb2tSW2DmAhXmCi+eP0SX5YkNc+Bz/xb
K0wUdXN82H7bfQBIlbW7dtpHmn9TGBbmtwOEUhloG/i8QmxrCkUSC5d7rMmWXcHApvDazi+t+4cQ
NvuiwmAnVL0MAT8X5cIlc1rz8brkz54BtxwyxEk/aspigfi+RTx781OX68T88C++ZkCm0tUGn08N
kIl/z/OwgXWrGjDuVaexNhccsjgw9VRPxh7agS8lmoV5LBIOlvKfZ8JltgEWBVI/e4LXX7fmBTkj
kEgugIMgIX7ybCL4enhaZbG5fEsgb/Rh1Z8FSLLV7Ym84/vWriLzHkxdNQGSRSY6o+G2WTH9lFfR
vsd2QS2icVnwMnW69gH2/WlDYHM+As+27D6uECYnN9safEpI5LtZjXFk3JyBHmF7ZKJ6Y98Z4eN/
id0HntIiYxY69zdLYW/f64awcSfqeCljpud/um9FoXdZ3Cd+/STEkhGwvyIsZhwGpsDyxes3BGVo
PwfwFOvpTQmozvn2bd2ripxrT40GF8FgKDos7bNtFvgxXvawOQdgke/HL3SrpoNsvNnIXRggXF/r
JVYiIN9QHNkx13sSjWuw+pXLUwDn3sAI5y0O1gZsk7Q/gPehzKqFSWfOJZHU4ljQ5lDOtT/11Pxs
4oVlkI0OGmp33Iz3MhbTqLdakE2A1vCVyMCzxtMLjAkPPr5iG8w8/xYWA2Xic7nxsM/SwmRC0121
WEE8V0X/5VBzRSfdFN2S8yD9rQEIVWD/gwPTRhAhTR9+U5wcdPPXQc2o0x22KgtUMRKJbYNb0VLB
tkRvIL5oSwGTKwjFwK0wKYoKdf4XrVx7zKyUgnb8YDJEXlwsNO7z8rnu9nT18zdbRfvok6T3mal7
5uSs4RnWobjnfZqhBlKL4I+1WhWnMWWhtQTJdjIXT9VZW/G2QECW6hLwy9WyWGoMnyaYn/L73ZvL
dgrCzZQcY9d863pO5X1OeQ80UOpaJtOSdY4ee1uihy67sucV2g3PFb/js6ojEJQEgsTqVQFk3RJO
Stm+IyDVwCEW2ZqZRDNnMJJZYrUIQdV/kJmghMuULs81oVWZRBbQwXH4Q0RlsRv4Izp6eMhAadL2
kJp/UHPPevaGWf0KT3scbrY34AhRkkmjKz32Z9NAO7t2sDYiYeWAyzBpUNLASXRCSqlsoOLz90tY
uQf5bX0tW8zGUGU/FXzVqbVgXX706yZSvPmd7X3aF99UGm8eTLcQCKL2QSSe+Y4UAW2rssFYjQNC
iEoMB8CUHpAUTL1LBnCW3Ja05+itTX4kPNxb+lnUrDjpWtAJy+bDO6tS6yvPlEvZWM1lB/Auv2cR
Wq+rbflPDh5ncbYY8/NZkhwAy+lizcMm7ChnxReAueU5U3eqga94n5QY817dzTUbp34uzLnQAf6a
bGxZzE40+JeHqnkqkzhMSYeKnS3Gnvd17SqqPU4DbjA1P0RJAoXCBz1kTguzZN07Z/vvsvwectXY
9I12lyS6Ies1VKYrDRpXd+TE2diBf889egeFed5YIMjvs5vgEKv/vlcqxiiwrbyWTgdlrnpac3Bm
lTLpn00GBFaephe7t+IelcM4Ht/tbmMttB0wuCwSU31vKvxmvJ5ygk2e2HA5MYSvl7SZZcsdhVUb
1FxpmjR5WbxGuiRJlt7qRKaNOYROYLWJiRTV6QcK9XYVBB+JWU6M77u+/P2apC3JD7vq2WcLjSzd
GkNuLSSZgV3f+KZr4yDPHs2Owu0OD0zBE948amabvfAb00r7eK2Ct0Ag5Hwt/0w8p3XfvxoCzQjf
1vFeaMgMZoCOLeIIkukDEcBooYSHfTx29Ua60Lt61v0BYM+LWiW7rZUNDhW0f9hGfiIg66HUoIKu
ujyuJgaHRoA8zldwvlm44FpWCOhWL3WdXys6DTvztT/+Xo++m2d0JwPHAnCJ86XOPYm0Ukm0yLRi
IMIuzQUckYWePKFILBg5jOH+44wZDOIvPsPEjFnRtbpWwix8W7pWvOAyyC3BlwLHP6i2zSkaglgk
p/Lc7Thh6tMcbeYFFU2Fg3MtDR5QwPHpgW9sP15uETOmOPXP0JM6+Nf1g7taB0LyuXf/7JiksI1k
4oAS15f9PDIqbnuWUx25Wu9x8+wfQhh/xjjWJCdbbI3ux/2OzGtLtWK8r6Xu+eNG8l3DJmHjwdYA
E/E/zyHaCxK8t+ENPLXJ+0P2qfq4FCRrIL3RhkStRfnO3RFONGfxYo9tXjvwntKBdV3+TptVrpHl
xEn5fsOpswUM16Xyx6ZESFA8QtJRRRnYsRAJcAUVXfcdmGmRq9ELKgrtcuhW40wwAx/AJIm4hbF6
WE/kxEAWkN+zGJHEx8oF020KdjY3gNzj9nHQh/orqdXTT2BMeokupoyztG3NUBXFBpOjSFTejOmD
FhZo4fL3XZ+Z3p8JYRXlWf+FVGXplYd4PSwNaFx0oKszxkLwT0X4/HDg778ZJu1u7L+uoDYj+694
34t5cbg3rE9jy9EqAR1Ga22sJl6fisayyPItsQMUsyz9DvF9rc7SRxtlDgWsoVJwiNyjszCjUXhi
xYd0wRVXTvEtLQxfsldMs1KPLcZ6q9Uf1qm3FUa2XBBetxTNwwtelOGQjGZ4RS1kx/PVFwn0n29v
qcmccGSVUPqZsgvfVGPHhmvF37gjPY2e/8NJLDrF6rI0Ndfx8ryl29dTTcoi7zOnpSZsBuaZUngs
UhxOnx4U+vJhs0aQ1YjNRHWbb+LjA49BDwt4YGhK4Gn0ipfcot0xtxaDlVQiXSFWjt8n8sOiUKJ6
fG2S7grS0ihDM61M43hGipUZsb89x8xCE/39wzyqnrjtaFwEADM2vHBv0TBkKCuaa39oXKOD6yZw
PBYLtRp/JQ7Pi8M/q3Y3qZ7ui1o5CsOpLFJ3aPjqaJV1WzdcwA7zTOcm74sB/1SGZr2c0bOWj1Aw
UivDn8zaei4jnZ6YGn9g/lRKNO93qQ+f2AOWxWyT4lUjGhN0sOhWW/CkJzInuTOtWL9YpGPzDhys
E7uJ8dMFzwa/mrHpKTDVgGrH6fNsuMFsY0pKM+i2O4XcwEGGoZ8VVXfxNTXFkBIRBr20weCckD8q
/C1mv99yBArhvWcuASj4OnOg8vU6Htrra5Tq0rObXcalot28m5LEubR6h8RnWugrpajpkyRH0i5R
K22NQ2Qp3GgpyVhkWW+CwYsShFwaWGyut8veuAn6cdoWZbQEKjgiGPZuZblh10YcGcnlceVaA9CN
j3n/2wMb+FcIHiDSU9uYgANKyYXJ0i1v5kcpQhmVayi09frgmIshQbpKsesvnEfyeArAmt3Fm2/Q
+7kISngHoDI4OVJRaJ19USC8UBa3s0kq4Wohcr0Q0vfNX4Rrt1TyE3+7g9oJ7TAeU5sWvU0ZfXAf
1a6CCQKgASdo96agjzrWxug/3+T2OmKnFo2W5HpcPxG8I2eHaUY2NFW6XKHiI9A04g8QndPnz8DO
n5QXBPE6uyLtOjYcdLJ9rfUHeZdWgybkNhyb3FvlkYEXEr4atsp+p/CDIHbHjBYw9DGJvWRGy2+9
1DalQ2zW62YXpUF+7MHTgeDnoVMjMbMTGv4TlvSTpMP6TwCy5iwpsP6jypYXRqmzb72I3a0=
`protect end_protected
