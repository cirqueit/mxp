`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
bPoNnd/Fm3bnYjHESr8+8e0Il6+4aaMb3i2VJOf4+0Aj5cV0+RKTm6ggxsNKPC56a8V/TtC71fAh
+ZVsZewLnR12KqLBqdlEu4psgaXlVPnjV0OiLWQE40rQfGfwhiwNNNNhdHUyaR2IMy4UKJFFtsmm
+hkI5Wkn6kOCvEqQkf2RqsoM7FtmRuCeGN40fJfQzYEHf4qAlfm+yAuAHZYrwOkNCj2GLHMq7+aQ
DJu/AYSb8LC70/IxtnYkX4yk3G/2qHmv/gu/KEgrSq5UMv8YVS9pXvZxrVd4UwYY84y/JXhU3OxD
28nxewLj9AG2jdg82EV+df29+ruCn+2jSCGTdwL9QGiD/31vrk0CABMfT/sTl0rwLgIA8GBT6lIZ
0Pf8o4HeLeVn7Ha3b8pH/fcOjr9s0H1uQuOj3YKZrcKFgvn3bFU1m6dygXlWLZhjhhjRTM2XBBBO
4acQ8gyRIZp9gTzpwEnnsda47CsjvNEKHlaUW10m0cnT8akFjhAuUDAzMFROmdINx7JAiyC2tpAa
M5K4CpTjv6BVMUMZuC5FEdfOsXIKraEaLNhVhyNCty9KjBtXU5Bw/Aye0yu3rAHA1bLb8iEVWKZC
PeLxBMLVzI7+xKz4CZsWYZ/+ezEx7Y0RDoqITEzSZsFacULy6ONnsxspHbxgRmAgX2xOAzsdVEHL
z/5TREmNkbAcmVkJrMM+Vdst4vTGaPSjPSZE9dgq8a/0bNTcZ6PDGUS4mC/CwVoHbcMNY/dpJTZJ
JWOu0Kar2NgWAvT0Mu1ihxcICsosp6yvbhFzzZI/V+1Kd4RXJHpdgE75qNmGkC/vjG66u0KPcfDT
sQxQz8TKzog+29xuJ2NJ0v2sRwsHuM0nsPySkmeFs0maaFaKj1hvALVQYnFg3BSs0JHjLCdAnagn
OdWqJQY8ZBr4tfR3bqEL0i47NWApF/WZFHyG8nCkm3r6HsLzYBpJ2Rt0b2/R1LGo/UBf55Td2vKi
4CPuSo5rgSY3LICrnvoFlLer9Oc3v8OsISWbAw1QjevG8Qq6G2VUO5Av5hcNxzCMJIpvv0xEmc2X
RowRVb70lL0jA8WH1ILQxKSFXQOJ6bq6fbKiim4fjif2lZ/X2Xt02hIa+y5+dR4zbUz7j1dxAD22
2EGHTAb8bgmj6qNrwCAIa4eOB1u0hG7cxBv6gaE1nM/RE/2Dr8VQ5ww9IJ991aELXp8RBnDf7nZA
jG074yNskTCUihtnkxwsrg==
`protect end_protected
