`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12192)
`protect data_block
s48oGk+4Pw7aMISNDAfylVqWqd/v1uj5OTa2X8dtLe3Ss6Ib/AwqSGjr9reZI2R+OlmYXpJFd4J9
9Hj+uBjBZbyKaSexEN5VTbfHQjnezYhEITNX5RxOuHwf65uC9m6RsU/mJSP01VyUVs56Z0pTzWO+
VbZydyXLvzVinnwsfvYF+MjjQTZcvyj1SV0aZp+76Jk+CqJqXWPIAzrgRrfP06G26d13JXl0ciPH
TjEDjmuKAuZuBCfH8Ek9GgEZmNJT/1mcqqf5KVyzPsJtFW0mmeoPodUtLFFi3qp+WArctTihgtUu
Brq2GTM5etawqnN0BfvPRppWp2SHwYXHu1dXwxDhx1XH4KkcLtQfPuI5qbBx7lRg4D3InKdNzf24
rXCVxYLk5w5ul/cnmfkk76Y6Vt2y5QLykm7uyabT2AoeBsUW7atj7Adu64BwgsdD/7SxKXcNlkMz
AtRWNxJ6AVU0i8JCkfJYvDGKeDaEmABNspcWldxJ84rVegKhrwziA29U1XG8ma17tRyc1GWPyyMH
flsawcgRVEpABlFhAhdIL5yxLtnUn52oZw7VrerhZixJsz7Xde8gvF7lQQXH1MJ1jWUJANKqIoR0
2xKujllSE4jc+eWewvxGasBCBVmpCj9QEOr6M6L9lAffKolFG/dsosfAAc76jAu7cWP8nxikjiQx
5//bnwU3WFbJjzwN/xLWjcclsX87Q7bRGcNxK4M11bDqGNeQoMkZJE0OZhkwN/pbbImWBOAyc7+K
bEOFdB0GT7nqaWhi4zbS9pXuBnpjAGgsaLo7/R3eQTjI5mnVMhBDfDwtNkLChEv5w+UJqIkOuMSr
508xLvtr6AkfiZ+pvTps7Bcw2Y46ve9WgGo0AX3a8G+lAWe6FX5+zJl1eTN1bLnVC5cPRk8kmaBt
QrG47b67sRirmkxBWl3ysyLr3TPCA3hndQ6bm2Wu+x0VraLHfHBQy6+dRfpQJ7BIEVhZwJY8j4Uq
LAIjWcKFHOr0uPWzFjwCqXsnlGuV3Pl/eSpjUYEGOCstDYZMHCIbJw0wRMvB+zywOZagmD0LOGsA
uximmDCXm2/y1/dVa+2+lHIf5x86I6ExwsNlvl1NlyIPxlo6W/vxeohbomkHYunJcmjIvASgkQZ9
OlWGsbshEieQUgiAEAHxglwDFzWihqSAxMJOId35Uo+SYJ0e6GpUHn0A3oRDlabxPbG0tnsJqdJb
bYQ73txrEkrcud8s2unxaoUFBH+97iHX64bGfbd9NUzWbN85671rIuaeKYCq+m7kBQqQtN52WARC
C2/jW6n93Fyv6x9YNYn1+EtjYzNs11BV4ReWRnLJ3xEOdNAgDgbqlNkQMs/OGaQfeumqAIUS2KD5
4UdQr8oAZe/Tm8idz3ecftOrBiI1S8P+rDrsZRPkRQ2RiFBM/0evsPRhhANVr+CAeSuNCVpx5CRT
RYj2LZylEdCuWrR3CeXWFySCdkibbEJfm4hIcLQlBDtwqnMcBxMbjlSlzgwhrojC7b9HhADO+tO4
iXCLnaRmk0fkOC9wuWtOISTQzAzahDghlwktRbS5W2G+TlddmWes6U9PQX6QWdseF/Co7zCml0dD
psh0Y9EJydLAxAgYmIIV79F+3WKvrzp75VzYnARfLT+hF6sx8UoKcf5IELC8/7jg/Zckhs5ltFgV
nsz+T9Vb1sgIAHvf5SpE1Q3ccGzSt/932kf5EbOaI72zPEjnLtiFxXDOSf/Hm55C7XhmXaTwvLwF
FicZDvs76G7phtd4PlPhZNdSjW+FhkearCxfM/JZkiJWyd7v9LDsqyu0+M3gusRiyrtX7ehKiGSx
Lvyr2+8kzZeoKVv2h396XNxUWhJVoRS61xmf1DNY6h47KdRdGaIHNGbp1nXUlJEX7f4W8pg1SDNp
NEPoiq64Y/1Vlf2pP9mz75HCDUEOGBs8ZI/KdE+K0v+AYYak+57F7ds8jqtizRueNvWA6E8dYmRj
Hu7Bm/Xt/xTznjorZrVWNuDvYmf4kkU+8XsPdxrY1tUg4rlnHzMM4SYI6I4rewdsP7I5BxuQMoRE
tx+/cFWBX8s4Mqj77TQyn1TNfLIQn2Uo/CSBoteRc4Mz7EdAzxfr1yqsZ26rvCmhtr3pW9LfFGXU
jfhpZi8BrUVSAgXs1EGAJv7apH4bg3cM+9XXevaRxJIszv0UFXy3wcUJi44S7yQY2td3sEMcnqa/
Im9LoStsiCS66a3jeGwYX5HGAqU+s1QkUL//TCiNgnaVxZiyMvibJ4Blo1aAuVD5p840FsLj1t2n
8ndMlWjb/24+zslgKezT4cMYEep9RbJhO/ISCy4JYLobQvDhCHTZe7X/ylD/fMHBCO+VxIfY0JX5
zZUS3sJpdjTFGGvDc0UPZaiigTnkL/HtyHYfNrKdg+ZNa/kwDhX+CHKUMpMkrE8P+RW73LhhJq79
qUsLxLAhpYbmrTSwDbzqCkx/ra5JoC9AQd5lowkg3QVpXKLOL7fsfpI8MWrg5C/ESx0CskEtnJnN
H/fk22gQuOwIMGDxJNyfm6HTcUFbocS7ChNuQ5TBuziMv4fNANE8wqsTJt7s0CuDgmIVqMkSlE4w
TvA8GUWHAbYUthLjCZ/S85cx/yd/AS3y26qyUqbEDQM0TkzLydSEWA8FE5/++CFCt6RWgodc7t4j
3dXm270JxEYvAjO50dXJH3uUF3+tKK7mHdV6Zmwmm3bUqEpYYjPmv/PM85YuhZDLXibNxru+8Wso
ePXaarCeLQWsEiQXQb8wzpMwjgtLvtMH6dELEdb7L0Twqom2ZWobbfNyiKgy6REEC3ZDSZcUE85N
admmx2S5c+wTI+gmtYmsj9zBZfZ1RqP4jx3Au3946bGTLQCWzzlsh1fFpRLuWVe57CoXcTblOQPK
EsDBP8FbH3HCO0+MiP42TM0gTJZYt1dR4kyMVC4Izz/gf/m7bLXgndlMmUMUp/8bU51F/2eLXvSv
Cxp0uHesGQeW30SbHUQtvV2I6mLz5fwKIVVG47jF19yxgfnmwNeRdxXTXfBNAkutOB5hpvUe7GeZ
Pwm8Be8uLUSaYdcMrjxivDXue1cNEgsnq9nR/0s0QmHdqSCQ/XUdRbmaPe3tPFcrXOiNNr6523+G
+DcOe9RSIlF9CPdjP1HRc9ujeAtmxTU46RxZVFcGWboOU5HLjt4IrLBX05VJdE+9xRjRg01D1Yko
PWbZrN0gn0qIifSnXWwUizh8xTD86OozJNizVgioC9U2VfiCSM1mTmNXAg4x8YwziKSTWir08Aqo
aU/REXZ2YWL87Px0wnB711YvVGuUPS2REEuBtq//HBJPjZF3M5+meDqAWYmvflR26+OCuNDnRReK
JysmsLgpUyEUjvS0u7vDxzdpi6hjy4GFx929/EcbXcreyTm45015eDH8bhKSY5dved2Vc6cfhC7I
TQz7ZgFGV2/bjofzXCXQBWRxFUQqHlNGvg1hG980OPRgn5ECDaqJmFAIyKMqftYLjv1NuEcjj9b1
E7mHy0VtsKAs7BBmccu0K1Z7V0r4OFFhTumVoz30ODTbWyb+HHfDeg/Rh5OtoNnkQBEozQqFIAIu
UvXkQvamvLenYYtqsVmfPtG8vvvbqgjN5ZZ8eLCN/3xhW7Z8r/eI+hlbkm3KnH2o1y66r87A5RqS
It6WGu+KTXnDlxGXM4G/673jAehUhzJiXQK3Sx+GIRNQn8IiNWgQ0q3UulEV8ukyu0EkRI1PJAXv
73Io1TJ8J3IDmzxG6atdiPxRfacdeomC1/QWdXgHVOm3HOqLrOMTcx4+yXumnkt+q46JZx35NKH3
hGrbAM1s4bSQWw9GxTXRJpveFhx14nOU1kSXtCLDCOYcYdGDjGKF9Rh9NfLtAtnpjowLMx11fuXK
LxGYPtUZjC97LsFp21F2HVUATbdrvgM/z8bUysvGyxmqybMvbH/qjyKFbwRSNqYFj7PCQpWQfp7a
HVdqKePxk/URC9eHf61lrYbiYgrqpE+kASyEZYoS5W98xlw1Bgsb2PIl0qjITjtVZXTEhDIbuYMJ
jH9LkMBgWJC2rrbNbJDkAadadrwipYPyadzYWUykB4MzrP/8gqw0lm9KAk+t2H2xHmpgJhZ086FA
5UM/1Sc+lFwNez0CIJyRKGaRpiZz8a0gAOvg9w3W+MyMmBQxVuozZ3XVdIna6vXpYroiVCR3Vjrw
V/MjVeiMsqVQJ8dAWUJ8dd4n+qAdOOjSuvAklgg10d3LFSJWFooyLPFDovyNtkUjlO6vJkdQE/lQ
lxtW2E94fcCWG2Gw4l/wa5kO3aWv4ohWuQ6fXd+zRsfNZ1THjSA1N4u0z6N6zbip/hsXAiT5h5mB
H1zczdLkhAJRbXTT6kUHPTEBHVZQBlrKGF3ajzlWSP0Q2vgUaFk6BiETYxJg6lHgfWuTcXwLzTaH
Li6Ok+Jjxf4/b+IXd31P7IuhQrzM5HqI4qe5/rHC6lj4Ppf/rWCnhEP3ktfVmkLSQco1y+wwC2/s
lMiAeUA8kkKgZt3vDLZo15ETLciBv/YG5Qy6UThB7qK9uU3roPjDFjd9j+rrWMnDOMqGsWwMrifl
ADoMvSiwXI3dz5JhxnDhUWXUCq0GlCc8LVJ30346bB7ojdoMXorSTyklOalGNHTFwT2PFugYZMHh
MxfiJhVBX5fv8r6HjZJNs8ePBKQnF5dRFwItS3vmHndxMe/H9yPtBmJT4ffNfA0IJV1b7Xaa87eB
YrL+k2xYw8Plh9kjVxpYfwzR4JtULpJRxrjZqMXd4n+zJKL3H4+dxR3VoGMlS7KkJZ+Pqgy410nr
ZXsTg8CnvCkW9aH9+Zb/iV6rhgnMCEGXwWvjMCj/GMI76UAuRpYjhgfY+ntq7MKBNcXSGyZGCwI5
PG4WKeKCDL2XWBGgMMhOfiI+uN/m+yv/E0e68pv5NnmBh64q0nCFJiReq0AFXSzOJuFHkLWZcieK
CBu2sgI3R+Iuwy9yKEdCOXuXTZ1oHemWlGMiihTDvpNpKEE+5PjF3NnfcZ0PKGm7vnS2+8GYvEQY
/2h+clAwGi7NptsZmwJZGgAUQrTZTuQD7fZY7BqGm3rNvccHV/rOxEukqrJYDqWkUfensLxGnTs3
Rr4YaF48WUqBNDyo93hMQwVZrRZz+azw4rWi5bOGEhZqefuOsUpINsC68vh2acqona9i8R94CFFF
Wa9IekILyNduvbFUJNgqfjFEhSJQDTEvTfYxICeMNd4aGr5YEJ0Sl9lExbws90t/GJ6l2D5tXJWN
kYJm5hxF3RUOUMnBXdMJXpMistJgkkG6Jveze5HrU7xwM/Z5H4Cktmr6l8CCN8eWpDynYiRLt7Lr
folbJ7byCxPiSEbj2E+RDHQfDSxfxLXZSdmosXN8yEFCPle/IoCT9VFojCkdVbZDgNPjJYyCZvE+
8BH9PbERM3FmTCEzdOEU6L0LF/8iQ5As2C9pG7pOiXPHwk3UekumDWWBQL7/Q93O4jroRI6RBIwt
1fbSIfdCX9ajU8GUFAB/Cp2ekEbBLZ3EBIB8XQRw4hix3nYzXeDA6sbxzjWQdhkVogh0qkPsi40Y
wxHVj/jXc5OHRifyNySEkfOu3QFif/v0IyGTTHHY8RGP5GuY0sEHvILbZ7lznHKRFy87tdeeQrdt
53XPAIYgJ2ml01ejTtxY5GU3eZrL3lytfGycwhG6ELgYeBBOFAt8DFKlz5drjfsGBzYEbSeUyzyk
EKMzGWLG5mJ25NhsJt5nUtS1Y9Ry4Hf13c661cIaDMuCvsLNeS7nToseHbCXYBi34+IAtSnMd4oP
WZWUHWoQFGqEB8PiupEI1vDUCov61OOp8e/WH5fcpX4MIj3fyCmNAdivP4lu13XT02SWLHRFf8qh
07pYd6skmKPDIMrOUFxXWnguPFFOBnpYSRNrr/Wm3SUnCJFC//3RVgY0BDUERrc9CZKh4AYZYVvd
y7H4gglXchtw5jqmQDeVswydlRZISAiuj2P51hv9BvlhURVnxxTqceLRIEtJxe0JBEm3ORc+IAPl
HJSAQayCCxiP4ngGhP423UJjMtA62sntDUHGGlcjQS3CswPi1A/UrpAWpP05VP/rdxQpw1abju+O
+YuS8Xti1RG9B3A7cokG35tga7nUOqry79bGay2LSZyiWcVpBF/AoYs3Os6UA2ZZdiHgG12E6A/F
qRVeWgaX7yAaEMd+Ga+ZzTWryk90JHYTLKITuvLMWyQhpn4TMCT1A+MUvB4GUUjB7FeM7I2ZVAlE
TOwQGYXU//n/B0L3ReupUipJ4Ec2s/ZnleT9V9bPDmKC9i2tIckRJeuG7K/ZC2jRtlbPWDD/mUtE
Ba4RlUy+wvXE+Mw05BoRQEWve8FCer25cN5eWweLKOd2Q7OD9vTVnq0m0sxukI7Qwhu22OfFlUgL
ftAZ2irJdIAcRDvAL3XOjZ72TQAqqhe6BoINza40wmyA8C0aMfY/Ysm9ufOfJn3BTEOzbq4erMZE
SrmzT7h6glH/gvVHZ++7fnvAzqBR0Tqw+URRuoibQeNRXDmQYaYdznEYWmYKOPoGwKqFZpLMskqF
8/Ml9DQYPACucvCps4DfSOnSh8F1h3Ckt3u7Mh/5gJxnDk08qR8bmvm7tnDVJCeZuU5hMdxq6VGK
ghI9HIGcx9NkuaVbTDkxBky/R9vEpFAM1hzMXDGV03NuK4pEiU2bvYLxdKjuZqwUfMh+HzVbCaK+
gWzCgsp96/L4jcmDKhCfGJa4xETOqpyV2nXduO3UgwPq747EYuosA3dzlIBp5cIA1Qtt5jYiFG3q
JGlW4SyUW8YspJC6O5Le6tJHUptKq44lPQs0EDsPq5N9U7DKGpWwvU5FH6C+4sPp228/jPjhfmgw
L4x75juBxzg6TOJ7RKtnd+mersLQ/VVuwem/GvVvUVke31cvno/O9xNsGtWYYwrBr27FDUKDhc5Z
0ds7jCAs8uyRzXAg+jjtNqSmFLH9FqONykPXgJXzfWdCBASpY2yzSiP//GTQ2n3GoyzEAJU856ge
LBzvVQ1PyLNbKm7dBo/ocv5RAv/yTKrIqSsvxZFec/1wzQm6/78RrScsGC9vyAYHUOpx93xriHZd
FQj9gofDgw2CX5F3Jd2gGS7G86IB58B+dlXmrXyU8dvuysldvP3SJAE1ID6R6iH09Woitjf1xu3s
nN4QUFsJbOSWZaWCVKPE+mqK8NTKsNa5gnLhQf53GLQofMBBIpeAbOh4qeJ6B0iB4cPP8FKdJ+SK
Why9byIeEQ7Kzv1B0KX8cWHqyigowi+s93qg9La0RtIVyvEQvrYtHzwM2bWd0kLQuTyy4r6qRSeI
eRzr44p7eqTXoMZtZQv8/PRslijTL3pVNXHq6LwjC4w6nw6KWfiopyofXRnTtyKRL7CzRmWi2MGV
KzyWYCCvKK2cXXoSD64Y7NcQesaLTAZA5cwXYrs00zw7TCNwePQ9CjQLvr6ebNnpNOUjvRX1l0XW
VN/sCvqVUqWOqlpjadNToD9qqgmt0GsAltM6FuumT4zqXnKBq7ENaYDXIH8TrQK2CJO4O+s23+o6
34XKtFELUOLeXNjkEuX3hps9frUyHlJCsQZ+YAKlYDpHdQD5nLXn3HhEnUD2XFMCSf9BDSsx+QBn
ZaBoJgWED+DcpPaut7U1F7SbQHmdqEwLaTw85rC5VkprZEaR4RkOUj3B3s8x2KxlalJUvZXd8Nd3
eGDhwXpbfj9OOzWkmNzbNnDWNh7hRZVTcWcTtH6PpJawAHyJ6g37CQ/5styrUKfj4GB9fTM92F/x
qoMFwsV1/jA5M9RFzMsi8rsPA1Zsypsp03oLM55jG8wicTFjf9GmBpfpmTkTqNsXqIXx0yZro8JA
fzLxZoos2JIsnk3bmzMcqYqC4pK+HQzMhe7yEjwscL8KoGeUpxPXo/3jzXqL8Nob9eK4wSMizen/
sFVxQayJe9UYOs6bcx+QVyCDoFLWtCP39q+qr13FfjR52AdZsMbdqVGGVMzfgvgz5vdfOny1bjLP
b4eng649XnAU1aoH+3w4if1WVSVajrTMeiDv/eDCbKJEBC1m792Z41yaVF5VU7aGPRSIE8+wJtNE
MrlkH6kNO231yZigv9CfAHcclZabyFnJpDRDBMCxtXzSMRXz6RVEMQTls67hhOLJB8OWIFYDPQQM
Q4M/sip/Pu7QWCTMFsjm2R4gVidajMQ6jbBpYb23DrUVqgQLm1gJHp/24zTRQWPGFSuibGzoZv8X
uwRyjmQ5aygn5zUSjMOyt4Z+bJ7qKl5Opd15iBtjdWoa8T1O6mZOz1J7AXv4Om14955gxqE92jfe
iOZ3FKTiDGVcZgJhyd7AOARNCfWv+JKLd5QhIlQAAKotIbIdJP24ZNUeOrpc2rzv2dfvjuIapTDW
3lcC37uKbnRuYlkUIPDlMjCMHS3JZHeME32/UIiXmsbbUi+gKtzvqbLyUGVwNMlZWfWCINLljTZ8
UGIfBpYK+yqDjEyd4bz7TV6RSw4rM7YpuxVv+pB5NDCd/oHBdPwPcnD546aXSRJ+9bfq/aZ+nIk7
0mqdunOvWFack3OV/rMNoHXm8kWFpTKXt40Jq7Qypz+Uhs64HrtGlRbX7UNvvGflxLrgxQrt2rQB
ZI+emaVmDmc5O/JoXIrz6RTeCUagd36lKH3ICKTN3eO6nr14LBqo1ZwXkUHsuxrXVadnbVbKXSBY
EzTsfV5tN0N+D3FeUT3TtZiE39j3b0Z0cq8Wp9/L5K5di1fnMA1KbJDvlxzf8sgLGapKZJCc6Isy
psMnb5WLzJqRrQs9BTkInufOsQ7QQ5rYf3gsjMfCHtI8IEBupEM8H7E1UsA95zPnY/VXQoXSbPB7
GDZgsOttTWBH+nDzwDO+APk7nPPJ7+Nav2bGoSi98IZqIgNFuxfPLufN7JMQ39yhcw9MjMOredOb
dEiYzskGpIJ69BIjqI/CPeJHNkTerz0cJ5GfxQUSZCvK20JYHICmim2T37Ajbm/t2PxRZVHv2yW6
8GxEbjr9wg70ncMbPRXGxOjKQLFSXneKVxMkyo4chvP7O6moanb2KV/Gd2x5Ix+jhKj9EtnHq8Qs
cGcNiDWrH5jX/uBcAbPVryMKwaLhXX1Dcs5VELnOHpyaLqXJWu4wJL28yKS5xAJCzTTk4IDims1+
wR7VT8cM4b3O6BT4Kd/Jp4TmhoMqb9cs0ZKaCgJsYlTzS3eWUhyZadpBXFLKZHjDtOIl1RqxJxi/
GZkYIociFEqR0eqkmCPEYUKFuTXAOvOfIkpzCRyBkgNMIu8X3DiqZ7iJ4yAXhi8TzWD366bjZ09Z
kc6SPH8oRnNB1ciT4uCSpdQRxfk30NBwdgJj9gcC3nYSTEU731qXd6rgN9wBga09FaJ/V7uYNVzH
pjvVVMFIqR8EMHv+UBHtOpnOyNOW2JTWzbousszJ3yhWPAqZ4JDWSSZ3ajsWCkEJ2ws7VNf03BEz
VpUF1nY3+7chh+wVTtqQp5eDX3VYHmlRkkBfkS1NUEn14rLJpjIauz1e0m0hQwlIwMp21rRDq9DF
V36NWsn+uc8iuuq5AaIaDHVjdCaUZjV515lrzmnjnWzK0IHtxeYoeGym5ijvXALcl6JqdvKyA+yO
lwXTMM2z2IQkqUnbz5YFcUdMEU+TFYYvhkV8IVGKm908kYnmX1iJnlcxyr3GYt0iN/M6NsDe4FmQ
PwoRikvzdFXgAjc/E4kd5v8kDplo+n7Ww8ll1tIAd5Rx8UUhiJZA1xFaJ74M9IY0oG9BsShDZlAy
r1JBmEdK4iMeWNgf+8BB1mj8S+gC04SmZxTQgucuBh+dcmFu05uNOtrIWedx3Fd4Xvchgdfz6XF1
JB+mKiC/DlIfEhbsExcYiIbs6q5YxHpPmKWfEEzZeLrWNgbxjTBVZ3yiIi4VRaaZwrgABawtLK6Y
bxbM71/iUje2Q1PoubZ4LbfYnI7C8QImiGZB+s7hJDxKuv0p0Q9UisCMrE3HpnXUve6NzRGVgPSx
GWi8zvJW/PsEOmmhCOsM6eyG5gkUALvrWE47lf9lzMydecKLeAtBVpyTRjWmPxllH9h1xtfFs2WO
eWAurSiASqbPkhOuvbe/cXZMqUXfJbuiRne8fK+1iNT2h6UT1Dnwh1ZqrHxc5Rhhum2+hMDyabRi
nPrVRmctw1G6TZ3m5i8HqaF4b57dpwno34J+wG+h9QFWV3MOFh+49jCXwBl3ZDRrZrEddy2sYBsf
wKeaDIAuT8Ryp4w9LSy2v+IfSe0wXPheHb9/xYUJiNj/rfFMTEWChnRqUZ//Z0ct/QIPwfpM3lk5
FW/mTz9fCN+8M23omBd3lYDO/+6rI8BjVOlkGjkr2fkbb1se38HJVuZu1/mUz/eZCCEFMd1jypNh
Bh66jL8pQgXLUPCXW8u/anfiW48GKTw7kWy1Jm8u2IbCWra0TTTHtd0kWaXXUsRQXoQ/39N35smw
5E+WqtcJ1mnTQdNbekhfXX6sLq1LEHqfpIaohftjoi5Wu1NO6tAh78OWRkjZlWhIbSg+POj9UG4s
V3VkETZLhbBowldVy01DsfN9/KJUdNetjFP2HcoBm6iRsDv6Jldbg1PD1afijX5C/5praAO8NkrA
O6FtU8JXocWkq+GRAj+jU7glot1zt5L9oWBZzWVbmgYliOQzfr+Yk+MQ6JpNF23l2FUyPSLgmI35
Qj3DRIlrRmmAEsRblNF29V6TaZdjVfdNqIOmqaAaQWhKbd9IuJZoyCrK6oONA0S5tsgFT2maVbxk
itA26C985WBAFRQO76Wm1a/JGHgCgSs5ipQ9A6nHeUkCJO3krcS+LKDl9J6eO2gi5tSIuv/4+fQw
nRHPbn9oyhrQ952eGDRW56mvhgIxaFuXid/hzDxPfnaoA2A4KPoCSGxXbqfwjCnIEVZzMjsCBVeo
kR1sC4jgymW4cCJzuy6wtFh3613IfPPGiE4S11ovTH4og+cvBm7QGX3SrTvfAO7B9ClWFY8o3rYW
2+fdgiR7qA86LznfIOWugsu6b7T43ut0GGKscG6oPIqDDnU98JZGHX85Dr8UGYUGRjbwZamyerMu
RGzxZP8+DTh4CgoJEeLytBwC2UIswdCDcxa161ldXCXpnw8gtvSDyYgVN45ioh/+aXlBkGfXJpdA
ed/V+0Sm41UZtod9uyNW+lDu54OCipV6c4NVFtKjCGhhvniUDHYG2GUJ4EjuTBBNoFdsfS28Qks8
/xJNkLyH9zb6k+Su2XoZocfg1HBr3oGjI34ofkmMkOxMoy5rxl75bDJKKifLU+kRpilw2ZFyKNEm
Y++LxSKDgz94VXyk/ZlaV+1umf5Y600OFORY2kw3+UV9T+sPAN1jeghQWM4nhUnQA6H8s4NUlKnG
qIRxMq4kkldcN6dp6+a45NBLmHBVJn/q73eeqMzpmJiIp7tilYDk+Pi0/nTeOUCK/KKXPRvaBQzV
4rlicUZ25VmXpCFb3Nc+uYbL2m3aCTW3xSOj4sKAwN7mPlV6im2Wbhwf6CbaCkoiMUK8MDsALbEL
rGOT6KRfv5VNpvqQri0WojhIaa1eJNETgBEMcyC6wnv3lK3BwfTtovHr/0DTXdhT6YHP6aNlYiLN
+0rgbuQIeKj68R+4a77rzIrA21HvBcEw6cMDBuacT4TdO+NK7pQIxl8kdxBDKalDL8OrVYWNnVBy
dAaQ8xVoayA/i4hd1dRO0FCRcU0yXP1FYgqSBG5LiHS+V92uGpeOg0xoRZL9fqMif4gTP9tj3xgt
fN9x0EKStIYfd9N4wBLyL/M29tBFxQASrM/6qEvdS0rGoWUYVzDUj3ojKliRryAuJvSLGb6jhA7K
9bJscGrMFElWvAGycWANqWTJUXmRoqWG+cVXmYvQIHQ5PiW+BKCn4vstgfxab1K4Ti7df2V22Ecj
z0sLfOo2eryid6J6UQdyumt+piMp+iCDv66e4f/e7Z/dBXqTyBccQAzucHIQ0qY9TaTrFt/fl9fr
rVrcsrisNJAc+OROB+r9khIZ1ia1MYFfMYS80mWM44eEXm+diNOPeruUiZUUT9Xw77Ahhf3+qXnW
/ENoshhZcfA/1OZDa0U5IJEwNoO6nmH0E47jsV62vpRQyp7kFmRos92JSD1zUtXcPpwGQ1Klnpdn
Hvr4V2BcLh2+SCVMQ24r5pJpHFpg+Ezi2mHwn3hH5UDfYFf/Yh5BLxpSpqjmKsPl1fyEtiH6CHmR
N6A5PTh3SP7Y9gPFORabZ5UHIGrKKIAOjIGiMa29qk2A3VLJRhDxwDoJ4GmK4fSjwKBSvQLkZeOq
LOD6F3upF3UuK7qVfJATWZKNyQPXSbjzUKldmQ1xx3+izfWEO52+3sGOy+dWDAKIIkIrY0Iuskjo
Bhm0ZbSYqH+lYJDOPzNDTr+6WMTYN9CsAL+eQJkXeV0lQFD+MKtHSQxLG5IWFpTzhxiFN3foMlQ2
/dtbnNnD3h1LQ8X2C247Axn6ziRiXkgozDIkxdohEsSkhIgqSLZ17pF4U5I5zJp4M07jKuWU/nZ0
yBZ9mHSkprHgqFOBWv8RzgT51YoPLqnapjFwJBTaZd+REWZnrIYIiEEi6Fb5hzmuvKoyAyNv2/pp
EhATtD+Z3cLXTt5IXurxQzP1xruZiIbAOzzjY7VmvIRqpGuPDiOiyWqE6DiSkumzteNBjtlDhSs2
LwdBItncmjgmST4QI0OinhvPxAx7opjVVH2OLkaV0ARPfdNqUM9PRcRQl0hqXylhDTPcZtdjokQH
175UcFYWU95BaPHUr8wwqiEDLtMJlCYtNpKTDoF+0CiTUJtpE7Jbb5vLvDe78nlkdStz3b1bWjLH
AfWRKGgGfHnbKVlN259oH8Pqg7VB4WHo8aSW7KWy5OYQkjglchdizdfwKzxtrxmR3+XMBr5ygSbV
3rmsPi2cj6W8hqZRRX/XyZ6Qx9tvJAzys9Gp81rRkZsvmDdtwqATp4Wx9sm4GZS1BIHziRTlqXvd
SvEwT3oNr1rzVU/PXOCItUD4cluah+d/Lf/qtasV5TVEto3vFyRuhsGZwTvDvweVyYsoFA8Cz6jR
AU9i6KLGywCCy0xHVtBoPhvvMMIfh+ovH/FfPyN5MB9ER4uLf2FvX1g9MQ4fQUH+LIw5Q8i3I4z3
JCsBsaGTBaESRXJnlprZSqbhtapdAsfg2a3kLyL3A0OjmzcvSbhgPn+JSPqfsOiMCIvfI6l17thX
15koZ3kcxecjqQsLdSDcWiYN95CSB/PQUyvOIoud1Ls/zffajY9rxoqklqr+evhx6gGMhX/Uygx+
ggVdKMyNlDhEMQsHqhkAm9hfEsAE+WGbtqSRc+Q+LZHnaYHBQY+xlh2Yta3ddKmQE/yQrDiDSrCO
40Rp/7G7LLwhD5bhxYt5JYSFc6tUIrHAHHA9TVeS2ROcawDtKtTQzBLEASOIqwwGdBEa+K4VcSIq
HI7Q5XH4bNIXgOYk7sDTzJ0MajyvOE6ajvfO7i8Luhb3afqTbiii2Uq5SZ1VVASApWqjaCc2YX9D
YZMf6taDEKsfOML0qz2kJrU/zimlS9i0Pz2nNgmwujZ0t/OgReLqSrPsyoUz0n2V1ycx4f0AQjjv
DXAM8m6K84CcCJ1HoqqK1ESIbmXnSuHQyqmc4NJGPx0oFn0uetlGVXfMrZPUOI9yZCIGHrsFlHK9
G0EQbxAPJmOidgIhQZ44426lrswn4rOJ0PACznR25S+EWrD3UbD+fMF/54iBcr5XyHmAtTvtmxOC
//XZARDsEOmyBXoI0jXNJ5pOgmSD7eNXcA95VSAnCfZSjBYsCzNAtTheQYpyK0+9ItWn9wuI3FML
9rBLOIMG2wOW1kdoe3uPXwKlqIcV7vJTE1HtF3racY0EbjpE+Zdhx86T4mz23SlBkQQU142cBMSy
Xsvvfc2wkujdCG9D246QW1CQB6uA5FB2oVTDLXZ+UYmaO/RajhRWMPsP67m7CaI8dfb6/50Lsx1x
/IgNRKzZAtf3ktQxxh69K4/hEVqPYnXCFW5JY8JzF6rCBWTsJ/1e0ZfQh0XJxqdWpQQ7Z/f6D8uw
44U6YGojcxL9E/QfuLP5NrZ4mHC6AbEhj13EzixiSMqutpXQETJxZtEB6rp9ho9w0Sc49pQv7lkh
Ds6ufllJeICElplIWOHKSHqMaSuShZ5sgFR9bBkdOjSGKZ+Qo/3ExPbzuORUgO0tXJzKKdM2iXKa
YCZf12ogOrjquSfDbZP4fG+7AM5SawDo3FsLwESKFXHXODfdlzG1GEkbcbqgAx+ZIu5OTSPe4oIJ
hS7hsrcaDwWhUQN3E0Vk03NOXPoWSLcfxQ3LV4BDojudnPV0l41Y2OmOuWQudwyTBuQyF+TBaf9z
KVTD38us75HtHjYE6FMZDbw6XVTh+2b00kSu+YgrlUpkVtdRY2i73+HZ3Jxo2pCUGSfGdx5JPUAY
7FCvMrNSb1meQUdeRO89pJVYnd54CG3HLz68p+m0Uezoxt6IWqU6D1JXfBbIXJ2F9myKcPixplTf
9Gvckd6FuDgu+4AwdG+FtT1Ir6AttXY/7Qlj6ndQRYXoR81i5Opz3iLrsnTvGIBgyub/fz14XRjg
mrbpI3r6XQLvkUmh8UmnUXVMdQqhaijyiZpnzR6rJEixHyJkHwyyJ+PWZSxUtCG5SkkyXIGHwZ3n
RqoB+GPCFJtDid6zKQPlb5Qg94DwKF3+OSB5qIpoUMjeFOoOYzEq4L7rAmIxGL/oZG9km8ZU7rZf
57H2HNEGNc5JTmANwpARu9YYc91hTuY+NX6+50ghBc73NST9w8e9wy5gtpWB9VrpHd7mrlsSLnjw
DfCpJtvtHJdHFfwrjq/yibwy0ZekWj6Wen+VSoEcyrwDqnPyQ/iA3wfVU0FFx1hiDjj0daTk4EJc
BinsA1Gfz/Mzk1o2XWZdALFzPdVYuKU1TYWQgtqTnt6ZCKwAIpVSFIKPMhAELy4PvfpQVF1zdTKc
kp1MvH0VyyMqrAs8Yjv+pxgdHmtk7mgU0dGULyH87KYle89PUM1Rt7LK2TfoR1am3i7WjvsosVb6
e0OOgRgd/FgawLpVZVAW1CWCZARBYjUuIgdxTDpFW82X1Nn1D1rbbfTBb/ZCPkFs4axxcR6z+qkZ
udfLWkzEbl20H691oUFPOc+gnac0qcW1VXaS9EttH+hy6GK/vogHaNY4L62sE9mSSPmcyY+Jzvr5
jt1yRqVKWFMrrgLXko11tOjjPBTLtW1ZKpEquTkQ/ZBDgH5R484DfZeQTncMmVfteTO9aw3qyF+3
Z2FmqKpKr6orz2PHFYFbWCK6805m6wVD7l4LPKVGWVnFvWwu8OBfeE9T8VBnS5zSeAW8TFEZQU21
I2zluKxQ/iBN0+JEs9aEG96K0jtfHKAUcdBmgeIKkpek8U17KTytNPi9o1BjV+QiSV/+MvWoUE+y
kCveFK2Qrm0GIjuARN+BhLC1RB3rUdc6V3uj84Rx/sacwP1dOZff9YSRHhcw/Dc5ClJdVVv62cv3
2UgnSoLbfPvNIM/yJwL4ZyDQjoTfgc5+ffF4g+zrIGNSTFUB7AKnHkryP7hgZA6Vquld6Aj5FJ4I
wkJVAZumNhhsSvzrV6MCwasQ5Y746CZW6q/ElcIJpg87FVIbAg02YNAcNVoodiNUpVjIawFxmVu/
n7ebhHpqhjZiLfWM+ELDwA/7+Dy9LRdwKmoJdgq55HuPOPQf9zRQC8FbUo0hsm4HTtXnUTcEPugT
nDr9e7X7m+vcyr24j/nwE863p+vsfoOnFiFQIjZ1qzGqaZTwH+L62gOXdeMBB0ccElDrtjJfcaBd
WowLzm5cpCpoveib7qcXmibrl+ZkwR601AdwX8ORik81bDNh6Bal7R+45hAxw5pjWD6XBDVT9dQK
InTM3clhc3iBlmXf1Qp40XIKIUewLrzmgTUvrP8u1tVbgiTGfWD7kLSGAdZdiJcG3u30XoWqD/34
SbZRFjBbBHnqwyI4DW0ZcRGeDUlciCa8guBvAjxs+TY/X9D+U4IcCBnmQCYjg8fziFKgYl+DTr+U
pWbV+J5OVQ/hCBopLq6rqQvw/MrnNvc3qvP+Icuqj/oovlGiSpsnuyGadjFb0Hqbki5gTECd8Z2t
0qNHbFic921w867ZcE8uZ+SjF0upMcTo5jCR25vTdFa0NKd4K1PLBISI+OKUpQnIWijEyiIHzM7O
W00I7r4Wtjt2wtY8BxdUTGcMA0p22rcHBWtFLyj5twpb2G0LIibG/8nKhnsZa70JV6F2RpbtuqRy
L5gGuzkZVDD6leObeWOnhUw8A+HWsnjvGAiQqwbFQLB5PI6pnZR2s4IhYQ/3zHnxCrQI
`protect end_protected
