XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���W��R��0��Qu�ny�Ji�U��V�b|es�_�~H��[�7��T���%`�k��n�(��$37�6'�aq�_�n�זm�����K��-�c�M�bS���q��gW4e�5���s���8��4=$)D��+��vo�;1|�t�[�����x*6�=�u�������v��zw��N^�IV����A�� �����vg(��
�]������ ���	֐±����ҟ��ƽ�B�<�[�P)�3L:-�<��r'
s�g���q�a�\ ����c>	��oZ��
�����mI�ʢN���K�S@�{����B���,!�,X#��qS�+O�����Zȧ�� ��T��P�<�����%�	���v(^Z"��)�Ư_���:�w�<5`e�2r�A����X�O6�#n˸���
vi��A"�cf��O>y�6���ʛ��S�0�"�	s�V�d�%�#8?=l��>񬄆��D��SR^�El����?��1͂t�h�
~��~�c����e$v�Ca}��8}��q��z��T���(�$Ӂfݠ.����`"�����rE�/D�����
~��Zu(r������,Z�RZ�1��K��p�y9Îm��
��O�m�ٕ��ŉ�~��_2z�='�њ�-&jw�bd�V�X>�P�Y�-�+1Ҭ�1�H�B��f��w�	�����9<5"_���I��Q�J�h�g�>uꩲ�����a'��RZg���Z�o,b)̑������i��ؒ|��e�7�XlxVHYEB     400     1c0�D+�=t���C^2]�n�^q~(|a
�g8�Cz@_�P��9K'�W��+ �z�\�����w�+`�&�����rsh��$M��WR�����j)��37�l���%�Q�t�c���}�DO���q�1��sK.~Oixe�� ���]�;�V��,)�5pf7yD87������H��/�����Ij#��n]S�A^DѶ3F[���g��Ή�������+
'#F�XA�_� l����x���g�����my�e1h��$N
("_ܣ�>�1{_����@��u+T�Q����}�b���3���G�8t5i�dwG���䁻��{�ހf���q������}00k qE�?���S�J3��M
i,��%BURY�D,n|4W{J��H�	DE�3'��,���%����Nq~���S_-��p�n���%��0+�H��'v�XlxVHYEB     400     160lX|$t�-]i��h��AUF�%[z&����!��L�l>�6�����d9�#��rbỤ
Nz�rE�U���|O��n'�3s�	��h{X�D�C�&���q��Ke���[���GS�Bbn�qN�W6�1�rZ��� �f��e�ǋXT�i~���QU��W-dO�Zr������B���ɗ������[�GG�3dd��O��+����dѿ8D�ݘ:4I'8��K$=�'�vo��)�>3�o9�[m8��W��j랿����/��Q:�/D_ 8�~ktR�I 4R~1�K*�#܁{l^��'a�1QJ��=��' ��l��˳��2�"{�����ߖa���XlxVHYEB     400     160Qu�K��c�Ҹn�^�q1�6�lk�jܿu�z����B!�>n����sWgY�1�N./��tG9�c��V���8���b�Z��F���5��L�����,��l�M(��
[,�O9X,��q����!�I�*�2�C=)��ANw��/���m�=����hLq#��"u���<z5A&��%D5�������Ѿ������1m
��;/7�P]�����9�\���T*��aE.����(>���w��zOY�
%m�[G	/����P*2�c>��G��	CY��5y�C�+��t:�Ԏ�Ĳh���_�,�m.�;�̫��?L�� ���f�W|<؞��ȚՅؠa
�)O=�8T'_$XlxVHYEB     400     100�]�sD�?�ƾ�����AM�,)�?�;GS������&M�wƧ�I:�w+�6�!�!~�����K&^N���%}��ZH�Ɠ߯fp+$�)I4	���툀C�6.�!�7r�ќ����1y�3��.쒡��ע䕌1�m@>ȿ�[m (K����:����2��Y�naځӮ�=� �5�'�����'����~�j�bN�,��$,ƞŔ?8~hh�T�OC��f�G3r�͙̐�ITF)['��"�d�`dXlxVHYEB     400     1a0VM�ԨP�K��k���m�Jq
d1="�g.�4�-D5Nͅ �c`����Vz|�x��.3R�$�#�<f�t��'>xߞ�O���( u��zw�����[&�@�Կ�pB�s�� ؼ�R٧�1���H_���ml_��.�k�4�2�R�/�0�u�5�D���F�$�gh8�nQ�� ���F�j�k��I�J�I�9ye�$�8�϶����\�c���{�JV�H�J���V��� G3�{�=E�2Bs�|�s�C9RT�(�3I%f��C�3�L[Ϭxi����x����G����+O�|��uǵ�T͛�,U���drc�~
E�#|ۑ���/18'ǌ�h�ʸk�6`����w���j�p�.���kī �.I���#O��B����o�Z�XlxVHYEB     400     140W�Ǒ��hN�=J$yK�>��b� }�fv��#����5�v�	�c.vO/�'!.��~4o%��� ���=���Y�[Ic�"��q0���:n�ݵ[��FGdk�0p������ȣ
��@�E"A����'�z3��5���ט��jL�.�c���&WQ���	d>x�|��9��c"$	wQ���tg��K�D#�u��?�L@�y}��>�$��I����s�?rVs{�M��� ]q�ྺa�_�S�+7���g@��K޽���!� pj7V���s�9>*�:@"�T� �&�Gk��w���E������XlxVHYEB     400     120��e:��!I)��$��6�.�o6+G�Ad~(�c�<_� [
���6x���ǉ��Au�P�H6��RL��9�[��q.-�z�=�b1�$�Q��gM��TbHy�w�2��{m�Y�b�*�^D��ad��=Uꉗ}sLS+�����N]4�~I�"�zU��i������;M֍KX�z[l� 2�Q+����׻�ПGNx��(J+uw� ����;��2���}Z����e����)�ݓg��3��h����n�$�s<W��:Rk�g��VEv����|��~�j�XlxVHYEB     400     130>��u)�F^9�QK�CG��6PƄ�B�����i�Hr���ݗ�E�S^r7}.s���uNR
�X���\r�3z:����Q4v0Gm�05��P��*����lӪ'o.6���P��<y�ɷ�dg"	fYn�7B���r�6m�3�r��֔ 6*yu����G�$����A��U5��A���yoY%0-c
�ȓ
�M����@p#	U�,k\���^����,�lK^./g�e�q�������C���
���
!fJ{���dʦ�ܵx_�k��WZ��KIx�:��Ln^�4錸����m�5��XlxVHYEB     400     1c0=��p��SI�Ь�n�t[���d�b5ck�j����\9��^%��[~�?O�%�ޓ��S�b��׻�%|������c'�vȳ��Do�X�]��O���H<6}Z�k&�ÕJ=����+^���u�VJ=n݋3�;5� �_"����[s��2!�fp�쫵��@]2�/ė�&��-�gj�9[t�j��"�q���4�a���G!ߟ�z-�c���g����{wS"&7Jid��,�{��Ϳ�~-@�[�~#Y`b)Q�����h��Z�7!K�+�����o��F�E��(���3&J�H����b~��:�����n�c�Rkbd�}ta(��ȋT�Kt������ѝWr=Px���!z����V�:ʰ�u<�7���[�����|:?v�'��r�];����ʥ������w��Iߎ�_X��L����/��ỽ�Ly�RUV�#������@�XlxVHYEB     400     1a0C�;�1�/z+���;��-CԸ�o^���j�H
I2�!/��2��@���]�<�B9��4��C�pvˁ(C�XX�i	>�HL��Q�d��'i�%M
g��N7k�����B��$�������~Ne�N�<#��Jʁ��}~EG6�4�lc�l�\;n��@�%d�ڗ�ܸ�]��?��&����q\�L߾���0����Sy+*��I��9�$-�~�q{*�d�׆�?�w0.C���=��=kx��s�Z�O@k�|Tܴ�xa�Je!�����*+Ό?�{~�T��iN%[���}y[>;��u�A$�����T�E��u�[L����"·��//�8���o@ݥ�v�$m�&�Z��o��?��b���B��%�ǋ�<�u�`��X���o�GR�1#XlxVHYEB     400     1a0yv���}> ���lp�9�Ou��|jsP�������L�qq�����8��S=�5�=����f"�"���{X�z&��sY5�����c��v_N�?�*aC�?�~�@���Y.׉��:J�O�!v$�zz�y)+��;>\���E6�Tp���Ue��Z:Y��g�˝�P6qc���.�BV�}Oω���	��y�x�OQ�ؼ��n4W\���ma�������w@���ޚ�C�Cl13�dQ�q8���%`Σig���U��}F��2p?Y%)H���
��%��d0Q��7�Z�N�еZ�	���3U}3�,A<˔ѱ,B�4�,o��l7�{��U���D���:?�����ɐ�la�b*3|��A�=��(��`bs���!f)򉈸p��XlxVHYEB     2d9      e01X�#�;)�$�;��u�
�~8�sؚ�?�7���'%�HA�O�ȵQ����Ⓝa6���(e?_�`X��o�Օ�$�H	 �؉↰��a�'�=p����p�/:�.|f�4�e���\�93+ϰ�ӧw5��R�Ȗ�eJ�������Wg�S�-\C�YJ6�P���_�F�8@�Ib,�[Ok,��Ț�N� O����u�̰Mp*k�{ql"Qu/����