XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���g��r��T,�����[k[����!����'H<KA��(��{ /[t�Vi�?�Q:�uF�v����֋^I�����5��p��,��B��`�(��W�ZŜ���gk��Ĺ�o���+�Ԕ�͓�Ǵ�z8����'g����?�M`L�]T������̓��h�)"������ l�AR�Q��:��K^�k�N��'/�$�.!������"f������=o9���bǽ���c�� ^ \q'Fw��B-��f$���(��<#h��PHB��
���e˗��FFǋ��O_�I���Ϗ�r�~ ���?� �T���2	�X�~ٌ��L�N/ވi�ω�����lXfrϤ;J�dgmg��3H��
�Rv�CC�,�J�P�c$����"E)��M���-����*����B}����[ ��ɥ-[Xβg�&�Oyu�S���T�/XN˦t\���J��`��\a2e�u���*��4��������"�{�i\^]�8,���bZ����5�a_�n������BR�gƹq�K2�%�F�>��|5=:l� ���(�儿�>��FeQ7��
�/]�H��Y�jT�v<3�$�3搜~���CJ�����o�L6}<% ���~�f��k,K���Ƞ�w���Iw��0�"N�(,�B<ڷ�|�?��`<��?��H� ��G�gݓ���V��d��Փ��J����3`0���_��%n}�0܎��m��!����x�b�h@���Y�7�)}�\Mkz�XlxVHYEB     400     220��/�D�]�S�D����*�K�bه���������J���c��$�u���=���Rq�M �h�;ݾ\Um��K>Ñ�h:y\��ݕicĔTt&}����6F����2�oɵ��a:q;����_�(R8$���q��[>�00~,$�Ҡkl;���X^����z�ˉ���z�~������RJ������B���*R\(��+���ק�l����T�c�� �F��8qk��F�X$��VnPd'("�:'�9�S�.�<���q�f�$1D&��oj�:�X~����$�t(#�2�L�.��_sPg���G&a�Q��R
���7Ū[	��V����b+00_�Щ���c؁�A�s�r4��}ԇ����2�w�L5B\�
(���m$���_oG(�4�Hf�8��J�E����.�����>�VXT��ت����]�./I��d��c���H���1Nں5d����P��4�Ÿ뤋}L��J����#ć� h��m�S��)�z�D�yb74���uWߓ����h�f�tr�S�=��XlxVHYEB     400     220JUG1t���`�Jb��GC��BZ�|U�JL�b�tk�����G��M��>�D�mTW��k��(�ڪ/5L�bynH`�6L����[�7e:����T��ѮhWZr|mjNU7�MmX������Uy0h)æ5����nGy����N��,�t^H/+�՛[r��yը�w���&G��M{���V@��O2��N��7+f
)o>�[�q� 4�}=���\���k#�iʫ*��&M!�Pu�C� ���S��m�������s���ݻ��A��v�mI�Q�O�M��N�A�t]���{#��elC�8ʻ���8^P�uW �����&o�h1����5��ͧ��~=;�U��}@��_�^����}!�#3�����L%
V�..�S���͈�x?�	�|5�!����OІ�Շ�ds��_Yt��1��
ԫ�ّt��sF��à"!�c�6�62e��[vA��g�z��(wз@��l6n�(��W>3)6��.��.U�BB�%ZD+�cp��u�We?`Z�TFF)*��|XlxVHYEB     400     1a0��9� zE���XUGܩ�g�����Z�wQj7�hU�T��j
A��X̾V�s:�å螚{�������`��KG!4T�xȒF2���A�YYդ�s+�YPIG�Ĝ��K�|z@W���E��p0Y�X�8�Vr�!M��,������&$����4��3m���7�&1<5?K+���Z������GM"���d>p�s03U ���y�Z��؊˪a��i�"
�3����=>o��_����M�P�y�� �.ږ ��I���#�M��I�n����Q]jF�l�i}v1ZUD��t�⤬M��i
�f���&=87r1^?7��~�����:t����1�W�)�J� ���RC��^k��B�
���cƲ��Xo����1JbE"�� ��"O�1.����o�/�XlxVHYEB     400     130X�RH,�_P! �H�K%Y'��M�D>�P�;x��Ss�ƖK�u�X���z	V�y��,�;v��T�S`d�q{�?�/ �m���~{��Z�x�F����:޷��d��t����K]&�E����~'��4��	��=<N�ʉ�,/��D�����7�Jvq��C��و�#PE�y3᝿8�,n���|#��A/� ���7��Vee�e���`s��U�zD߸>1��} ~o#�l���(J�6	��7�B^F	<!1���������~C�o_˹�����Ue��l��c����!bgXlxVHYEB     400     140;�r5al�����-��̐7��]0Fn�s� e�� ���=	�k�m�S�����5[V}�/��&�d��p���]ľ�{�'������LS��UyVY$������ϊC�e\�T� B�q�o,	��ۇ N�I�>�������5P���FeK�ED� ��̙.�~����	:�й����_��e,�	ڕ5'���A�QV�n��M���)��Uy��mɇR/|h{'%�R���I�=h�v��q����;�;0!?g��B��8�O�7���=	u��K�ydL���{��m���L.ѓK����;�uֹ�N:��s]��,S�A���ye���F�XlxVHYEB     400     1c0��Ǝk��8�{~�ه�2,�{i�=C}ű]=���A��`�d`�0L��rq"�ޞ�r�ǞʹĆ
���K��k��
��M�Tg|��&Sa+Rc�Ӑ_8���fVq���`��9GU?��˩ǣ�o�[���#�?7���h�M��i�I?�r�Ҙ$p�5O��CC�t]���$1�)L���V�#I�+EfB68Ѥ,ݕC�4J�A���n�E%���3����+�*�~�C���J\��TU��{����m��$R�� �� ��5f��2G���✂��k������!����X)!8� 1W��8�i&�3+6�R��#5	ʢ�h7B<� �C0�ɒ�*Ҳn�nK�"�z�A�kx]�ԩ��琰�-t���i%}:"x�A��w߫`�H8���wH�.�t�6M25d|U��<2B�a9o�q`��A)���XlxVHYEB     400     200�O�Y��SG�ꏁ�z�D�S��Z���yW~���tp?P1���%��%�޴��o=�������;��C���j �+`j/�ۊTpZ�|�33
w�1Ћ[��=��Vj:ɓ��%/r`͠�M.M����	�֫n�4�,�yD�*B�w�x]�Ǟ릨A9ca@9.����)��K�F+�pA+��9��/��XR�%�����b�b���͛�{(?���2��z+������1�)_�<ihЃ���l`��ޫ��U���=��cX���@���g!u$NY_���(�i�ַ\��� �d�����=���_xЌd�p��\����/�T�V�����C<�,P��*��[���!��ny��NWqҍ��g�"���v�k�};{�g����,�r�h�����4U&����6��ⳝ�R��c~�X����e�2	&���s�ʉ��>��TBp6��ò�a�u໳V��1#��Ƅ2�.��67u @7b�0�J�z�Z�e�G�#��v<�AXlxVHYEB     400     1f0l�)�z��j�F�r�Bi�8�4���ءUR��џbÆ��_�)�&��<2t��@U�x-�#�vU��N���N6�-n�Z��-D��e�5�'�sœ��x�0�5�����1;����_�b���=���|�ͽ�$r*k�[1�UM˯�%��zbq-��<��d46��L�O����h4G3F����O�!J���)�i�)�ڀ��y2��;�Y
6�Hd�w�pp��*�r�ׁ:8|�UC·�K�)rr��<E�8�E��U_^����a\�%�0י�jPJ���8��Jl�
�/�iɡ��qT��i�<
����
�k�>�bbƵ���0=��	c�s�� �w��5����W�y��մ�����¶v��C���D����{�<�R��TJ�+9_n��w�zZ�/����Ri��Uav
u�E�����å:��J��H#�O�},��re-b ���Ѿ�8�!&�Y3�����s>��*��٘XlxVHYEB     400     1e0�sC�f�}���[�*��'+�^��׺Qi�>4�od�m9K�}��dy��Ga](��#�X�4M���8�ޣ�lW �lxؿx ����lS�ǒJ0�N�#��v[��,��cД���W��c�ѧ+P��$[��G�(bc`8�'���u4\���PQ|���E]}rq?k����\��!L`[m�JM#q���̨dܵ`~����,t�4�t�[91��˿���T'�<��v�,��� �f$��gP��X�9�n�y��r�q��}�J�X�(\�a�~�����]�D��'S�c_ �5�"x�A��t���f�j�Zs�D�;!�2\T���s�s��lMxV�*	�yQ�E��w<��S��9@�X��BC��H���jO�vњk,[�W��Dg�0m#�o��PL�|w�X{M��lK��@�1�,�_���,N����1��p��S���х�8�'p �t$�ٿ1XlxVHYEB     400     1c0�j���!�4>c�(�O9�7p�����`k?��y�<X���r��%�$Z+pB���j49��Ui�;�e��et�V�#��:2����6)zu��=����~4��fg�E^h�q��ex�BCY��%j�����e�یzc�7M�U��_OK��a�9���tǵ~�Rtz,
�����l7E�U�B/�<�E!p̦ՠ�c��E�#�� .t5�&d���M��aL��lb��%�*���[ϋɰ����P��+w�ka,�-&O�z��y�	�H���a����KVޔ��3�Ʃ�{���23��ި｀��m��0hܞ+����-�ȟ��)�S*}N�����0c���G�mJ)ˠ��5�O�63�nlJl܅@ᒯ~8>��������bQA}<� �2���[~g��S��[��5!T�	�:�B�lv���8���JN:��#XlxVHYEB     400     130eS�K���f��'��ߩ"��e���������z�kYy��_�l�n��j�Gۺ�&ڳ+�������z�e;8�ąD�S�0�D 'u���@؄V�ڎeq�<�]c���H'*��"��ܶߌ� ���a;ө3�	����u��ND��qՓy�#��d� ��z�:��QJI1�΢<�9ů&n=�O��>��F=
��Z�6b��}�`{�|��fB�>,��膨�S��N�L\D�]�Ɵ��o�xx�t&�KK�I�P�c4��i��Z��Ֆ�sO���hn����0Ǉ#N36+�XlxVHYEB     400     170n��z=~�@<AJ��?I��|��+���h�zo���|���ޖ\�����Ɔ�n��8)�M"U�R�h汉z@�g��$��޾9��R��+�����&
���yO%�Iȓ!��N�?mB��x��VV[kq�2�u�����ʗǃQ�t���~J�\z\&=͘�;JpY�A:wc��ebx�čN���SԚ��o�����'�O6W�KG�L7�s�SިY�,�5û@��� ���`Q��J���kS��@L�99�%��p&�����`ㅾ#N�d9UŴK@�m�cg
<�Tʉ=Q�ӊ8�+��򯒃&��S�+gz��Ӵo" �o�)U���í���Y�"(�]xR=���yƸE�XlxVHYEB     400     110�*�J�����Y�
�`,R��7����~}���~��VHC'%(����u\��u�tn�E��>~�kQ���luB7h=���;֋n��:u���]�`�[zw��%[ȤVĒ�{~t�$���+�7����[�S��1�7)�|�u����5�o���ԍv��2R�L�G�C ZW �
{A�5?�v���$���Q7GJ��N�.���y�E��'a؈d�8���_��E+ʷ۝%��YK;�{8ρŻ����/��Ϗ�lX9�D�XlxVHYEB     400     1401Sǋ���y{&�^��s�b=�p�ؐ� ��T�$�t��#w��xZ����kΠ؞"3쉛�\g,P�6�d>��or�rp��w�"�]a��8���n!�ٟ�u>G�7M1J������~�3�� .
Z��O��m��{����G�z�ׅp���GӀ���lc��2�9LS�G��*����!��-E�b�E�<&Ԧ�-�S�m�c��w��w��ShŪ�{�+�%��c�wBS_�b�̗]��)M��>xe؈����&��m�E�"%ך/�j̹�Ca#������,6�����P��ly{uXlxVHYEB     400     130��~���h�^���Z�CI�|S ��w7{H׫�܉<��7Z���=��4�G7��5%?�	<�N��0l�ne��,>�LF�_"D�tr����� :�j�Q�SNK�KD}M'5��Y�`Y��pKX�񷶛����<�X<���ڵv�[��$���H�!Wr�9���;�g�@ɶ��)U-:�����#�"�Q�	+�Ro������旀%�^e�1ɝ*.ϡ��7}WK�u��AW�1�?�:�t)��E@�85E��h�l8MEꮷ�PvvsEm��N�}�3��A���VV�4SXlxVHYEB     400     130�M��V�D{{��W�ٜ��������^ϔ	L�U�	��-z��v����3|�|m	�ߧlK�mu�2�ITS�.�Qz�7��hS��#g���#O�l�!�L�����|��)+ ��Z�
?\K��"��ͥ/����x� ����6�l�M�w���]Bm�xi!��C�&�3RV�)�V�m,p �zq#�y{c��~K���"���fW��b2&i��N(�F� ��  �m�dD��$Ө<�ul���D��9N0+�d⮁Gsq��'�]��k`ݫ�khڪ�^�i��I��s��d����XlxVHYEB     400     150��ve�v'7��|���2_��E�`�SY/��D�@��m�*e-�ۮ6��D�JV0
�Ee�RNs�,�׉�q�fN��dy��-`�N�p4y �X�E�lv���^fg?�	���]���(/|�C����[�������~����Ըx�g�=s�Y�"��6ա�ͺ�!�躠��X�/����=�A�p{1w�	��(��.����l�}C�"�9}����������\���)�h��9�׫$
&����fť���\���#"h�����&Q�5��;'*�>X\`���Q���i��,%@�E+u7͚����k0�lv˖M�A��駔XlxVHYEB     400     180����ۋ��%p��I�fk?��S*9��4<­�/@O���C�����i)�[�!����J$EJ�*�kMΗ�@A���.��~y��0�(���i�3Q!t��AtNuG���uR�ep����;Na	=�͡������sRR�߽_�)����(P�ՙ� ���N�Wva��"^������/V����<[�W���!��k�s����!�І�~�'g�IS+������>��r!�?���b[Ĕu�!�Q�:��!x�����^ e����{_+��n���tFë�n�\8�_ؼvp_�٣@qh�ѝ�-�lR�@�����L{Zd��R�_C���yS���h]%9�KD�1��Ll4cl�+J!XlxVHYEB     400     1d0@V�6�.I����0��
�&9�OYy79��r ]o!(�ݵmzod���?��?y���sWB��&Ь�ε���fm'1�)���(Q�Z�,��'{����x�K��=K?9�2�g�C�iO��~�> D���ٌ\)�ʩL}Ϟ5�Ő�%,yp��Ͽ���E��|A����Y8%�FǙ��+Q��o�~ϑ<��FB~]~���c +�<]�+��i�~^���aǖ$5���m��<��9�!D&���VL�C*c���$n@�}�p���ñQ��u���[�-1���/�.���?��'��DY0��zK2��:Wb�o�4K=#8cOHk1�0�3�<���tTDS�G��Hk��P�YV?��C	q`�Z���8�K��5L��x؎�'Z�������/�0�N�Bt�z�My��&!PID3���o��2]?���?8$��2��.����dE4�cg0�XlxVHYEB     400     180��� ���Ɯ�Ffg_��)������h��2�1�RC��:d�)�Q�2�B���5���hi��a��R`��t$r�������#��cJW��љJ��UHf�\�l�-�#e��[���3���;FW��?�j��HJ�9N�B�Dܳ�;B�W�U���5�H�.ȏ���6�^%Τѻ�E���}�(��G(Eб]��}c����eóue�U�;g��vԝ���?���!�FW��=�ۀP����^�����&�*����b�����n��p*���c��_������GG^� ����{M���������v{�u
k�@D�6i��e����&C�M]b��^�2Ce5 �j��{j���f��I�o��pk7XlxVHYEB     400     150�+=�V9�0ũ�4��K���5DoP��s?�h���j��?�j�ʸ�����Q����$�� |��t�z�P�uq]('k�A ��mΝ&�@?��'�F鵔%���2(�w��j��
�hjn�B9]C�?tH]r��M�}���l}�A�Z�`��׵���bW�m��a���CnA��PS�ʒԅ�:P�OD�qQ1[����҄𸸎W��'�xô��������yF�!�$]�qG�p���NJE����)ȴ:o��$9�,��1f�ՍW�����J�	��=�hs��/U�c%����5�D���x��{1���������̴��XlxVHYEB     400     1f0"L��6f�C���xY�(�>n��sov�.B,�i��m[|CVe�g��#ܓs��W�eI�i�_
h޻�'�I=�=��er�fn�W�X5Op'.~�>�Ҫq�r֡X#���8Gh`��9�*CW�̊�y���T��[d�E�����N�.(���N�8�)�����hP�X���z=aI۵�4����	%�}��&Һ�*/����Z�����0۴-��[b��U--Z`P��$���H�#I��=v�g��P��ҕ�QPO�s�	R��Mf��+�0l_Dw^
H�nV AďjU{}`�U�q���˥�$}�lE���AH��9w=�#����%}�N%=+��E󡈥����xOH?(��}36�( ��t��_Ӣn�g��N��O����R�q̀�u�@��S��&m�t�Űъ�Z�^v0a��V$�9�G�G��	a�0���e�#�RU�OR�Pك�*	O/"(=2��R[}�'�jXlxVHYEB     400     190�޿��Ц�?5e�"q��A�����$��98#c���X@�~�}ĕ��K��Wt~9�^t<����\�9-P�ߵr��z�������O
��C�^���%,rx(���Zdj������(^�5�{�TE�NW�/b|�G���~�M��0H���_t3��K����?"��o?��Q��)uGh��SrJ�И��6D�c��l�׽NT�N���� ����L ���H��������nV�'�_�/ �Z�ԌRR��,6h=��/��=���+H_���J��4��aZ�	;�l�Ֆ/�y�j��B�#(grv}���F�3g� ��jfN�����/�B(`����[ba��2e��M�3�<� ,��%h�]W�a�8�,H�W��技GG��ɦ |��XlxVHYEB     400     170��
���G���_7�r}*����D�GrV���=o'9�ȓ�h.K�R�t��3{�Vo
����h�(�/��7��1�+�6 ,K�;w2��������sn&���: ��s��i�"�&��>���]Ew�W��n/��.�&K��%�����`R"���^�tM����ǹC�^>D��G���G�䉬x����jR�z���Մ�,�ȭ�ڗ<�J������&���G��6f2���#�X��|���~Qݨ��6��g �~��nc�R���x�(�,�_��Ȁ
���zN���TmMD����J[�i�Bٍo���do��E�m��(څ�0�2�=��&�-/g���{L�GXH�XlxVHYEB     400     170�a�϶�!e���"�h�X��c!���_��BO=���Z�@�zn���t���4x`\ЁT}�c��(��.�È���â����p���Y	��9�e�,a��v�!�z�X]Z����:п�vH�v���f�>م)�ҽ:�ܣ4�%Ue�O��^ʴ���_��d2>��6�l.�{�����'�X��z�F�
�H^�H2�����zMZ��)&�jm�6��j��G�����%��'H���y�`����޳^�4����^���3��x�B|��ݴ�,7!�dA�z��?��)���(t�a&�~q�D=��a'r����=�O��*��a6�4���TB{Z8��Gf9�IS ��XlxVHYEB     400     110y΅��3TL�}��1��9��K!o�ǫmF��%^�\�c��ׄσ���tF$�a)�qŧt#V6��T8Z)�Y^�>�o��;V���Z�Q���=���C�;t��߈ͥ�X��j��C���P���0>"��� y��1u�%�W�vȭ��>?�dV����FLXN��!4���%~7��p��5�\(�������Ǿz��3�a�G��|D���Ӓ���{҈-�g��$.��5��o)=�	��Dm�:������L"FXlxVHYEB     400     120�s d��.h�?p	p{�֖G�M���@pe��;0���%�d�s��t��{�@�U?�8����{�����;�sʓ/@�Ty���>�$���D�[�p��bd��-T�����~��8G�5���`��G�A��� ,�[�	�8YgZ ��t����X�'�ĭ�`AL��8�V?�"�>�6�hA�'��R&y⹫ۜbj�߿.���W��*6���CT��2�(R�'g4�()�_~^�0so���D7�#��u�1�/���\���5ɂA��л��Fs����;�XlxVHYEB     400      d0��?�<?�S��g¹hD�-�����nNk L�.�D4�����BF$(hc����-@yR8�lU]�F�*�[�<v�"���D��n��Y�j�\gY1����mW]X���Ld�_B�Oy�\��
�?�q��$Q7<*bS|`X���k jU>��좀�/x�bg�R� �*�H�G��ک��Bj'3�$�I;�J��~XlxVHYEB     400     140?�ۍ����0Ul��~�`����[/����f|�θ�q�O��ZP�u[YӐ~����|PGJ���_o|C�>��¬N��5BA�m����@ l�\�~@ܽ'����
�ɥ�&�}68&k�@E�	�S{�V���p6_%ͪ�i2}W�dmu).}�tkP�}��3בT�hj�� ��ůK�TpL���(q֊q㭚z�y ����}�񾼣��L���vH"�h���n�~�������&�����kde��W�[�'4#hZd��6c��G��vϝ��lO��JW<x:-y��.H���s���K�Jf�WXlxVHYEB     400     140��M˺�T�������q24����B�'%��4_Hq�X���&��
��8R�~d���uVQ�����`l$
f��W��oR�흞�[��>|�֨�X�o�����;�iE��]�3�c�Ac���Y4�q.��F����Dv櫙��+K��qkZX�"���=t���;��5i+��w.k�QJ���Y3����!	s�s��umzV5���xLa�r�U��%�/�S��vW���`��l4b��bz$#b�Պr�1�/��"qͮ���چ��e~~����+XQ���<:x�++a�*��u�[�'zH{�EI��ڡ��XlxVHYEB     400     120���qN���
ѝW�O��8i�A�_�Kg�TX�I4_z��ȣ�S�:��6Z"����)�j�hJ��{�H>�*f�q`��N9�xJ���,"���2c���㰕�]g�7go���o��ʂ}�����*��G�\�=����B�o���(Rz��^#EE�����7AI�ۜ�}�F���b�v�IM8<D-;�ŋ� �ǉ*�ħ��U��p�u��id(�P�� �+�	��X�ٹ,��@'ܟ^jx�t�C6�R���Rv��m?�b�����y���b(XlxVHYEB     400     1a0�'̸��UR�]p����i4����`@l�t8���:͆ZJisU:�������"ɺ-���!����z3T�yJ^?p	c7��p�6S�5McA�A���=qG�3e&R
Z��MLt�Ɍ��d෮�y��K��[Z@]�Ľp,_봏�T�q�h�M�J�}{�c��ZH��@��8��rz��&"5|��$�;ƯN��z���m� G��X�$�N�Fɟexw�e���{}�62�T�y�\������.Pzo:�r6�h7^1�E�5d%���2�f��ifz���ѼCN�o�Q�!#'t�~�0�:�^=��#�Z���e����yC㜆�	)`/y��;�=Nm�x�{���ֆE��&1�D��F9?߇���<���ܷ67�D��H�]��R¡�'T/F@�^�ٿq���g�XlxVHYEB     400     120�E�ӊD�
=ΝdG��=�F�z��n^Ɋ�7�����?m�{!��-�-B}�ҡ���f��q|F��.�j��)��!zp����Z���z��Y_��v#L:Xe͒N���縲�1�5sj��V����Y�s�zF�1.vE�x$�H��"d�)�6W� ��&&"��@Z|�V�h/�k�m6:˭b��Z��U�&����ebS�>��'E-E`sx?��4l1��j�����w�����B
15N�x�ÿ�,�Ɇ՚l��R�ާ���U�D3�J3ǻn�JuiXlxVHYEB     400     180:�Mc��I�Q���E)w�9y�ܚ�S�ՔL_o7���#�	35��8������%�\�����"D�D+�"le�i��26���B�׉�N����n5+*<ٯ���˻�����x$AR��������ra��DW�>w8�1>$�oE_s�� �[���Vo����_��yh�Su6uu�8�{��7��ܴJA���T������ϐb@1��T�h�\�h�������@"6�X�M�ѯ}�H�?[l���:xr(��ܐ���+x����J$���5�y~k���>w������.��C0}�hI"+���~6+�^�q���n2�t�L���)�PU�92(��c��'yŗ�y��<��қ�ᣢk-���1ږ��XlxVHYEB     400     170�S�F�'X�2�������C��p��2�E'#� x�҉��*l��z�Q��D(m�Ƅ�g�\s�sЬ% �HU'󹹶�n?@�Z�g��.v�����9ܳ���D;[�I�'8��ސ���	R~�hȈbq�����G1-,�j!�p޿Ǥr*/2���p10�	(w��$I����J��(f�= ���Αys3F�hF=��ֽdI\�J�k>�-owm�����)�oD����5ǗΧ%�Cd�c9��4X#�WQ",��w���x�GD&_y�
�$���b��д��	�r�E��Ҵ���1ԑ��g�Y�.Aw�n��U����C��`{nS�@q�j).���z�"�	� �XlxVHYEB     400     1c0���I����~e�j)�=�G�H�s�����z$�觲��$���>I����񋞠z>la���h8QȧT�Eżd��T�mg��Z���69���v%���mHէ(�fq�ݎ,�Sm!�?a��!}����x��:;����)�� �ue^_����
�L����G��6.�����IeCT�'�c�{V�"��n���	��}`+�G���.S�Mlw(o.��#���2;F�V[��[�5�*ZIR1\��yJ&������5�""���������6�tL�+��t�>$&}��!)�K�N���2O���/n�b�SY���wH��ӔmAQn7��u�łw�����~���C�FGc4ڼ�d�����;�g���wAY,����j��p3)�oKo̔7���	�\,��c���^��a����U��ޣ�i�xXlxVHYEB     400     110�S[3�X2m��fp�J�P�9��ñ�fh�����] ����=��e���e:�H{�Қ���cŽ�&�K�j�mՐH��sj`�}���ED��h<��9)���r�S��_�S�<���KR|����$QH˶#��Ư��߲YC0x���~ ]�b���m0���֩ۃ9�q����2)V��=��K6�\���2�V�؍N�$�a�N�$�H �p�j�%>��tO��2Y�
�)ⴴ�������Ww�jH���6A�ԟ�XlxVHYEB     400     170`� �p�H��)�T�����B�[9h�9����E$4�	M� ��rVE^������X	���C�4#��YNE	�Ib8�	�a� F�#�#�d'�9e�h߲!�M'�,�H�9�Q�ʨ��:f��oh�>����d+���~�]|��v���"���'�$��cQH�1�<�%UJj�y]����%D�L���]q�'�H\`77;}Ɩ�n7�3��.O�T�QBx4dd���Glw?-�0�b�-]���X�
/���ǥ1�#E�<�@͙��IY��	��N��6-g�؎�9c!`�4B$A �^E�?�j�'���MO��N�-ڶr.�E<$�W�;�@)�nuRG�笆X���Q��,z����*�xP~XlxVHYEB     400     170�/���jM�^o�{6��H�tvZ� �Q���� B��~�R�tB����V�u�kz�J���yg����-Gy%5�1'���v��[z?�,��"���}H��I�f�Q86. ����`d���3z��q���&�D��,�/�jP�A�$�e3Y���=,��|����iSi�_~�e�-!�l�����Ƽ=���ME��ݛP1A~�8vy���]/�v��:��ˤꉊ.ߥ�*���L�dk�{����t�:\U�Yi=�>�t��W'�2"���c%��V�28�/�]��<�q\E#Q�ʢB��3S.Q���^��� -��Ğ�p��Lt�ދ��+��:����o�3CSmeY]��SXlxVHYEB     400     190�tM�8�N����9j�9�c��|M��)��'�n1�I;�H��b��a��:��n)h�:�J �����}q�
K����+��c�(�����a����&"��{J����7.jIu�vYE��/��Z�C��|̋[Kr�)�2Yw��H:3w���.˄�Z���bF���y�MI �p���]FQ��ol�Q�?���a�����u���������(���Q�"���uh�Y���{)�R�G�wM;[1�Q��3B�Bp0nQ�aI������F��x�`I��!�#P��&����.*q<��9q}_Wa�[O�@`Fx�����-zl���>�s0U�z�(����!������J��+���wM'H�YV3,��N)�h�˃s�9%��	XlxVHYEB     400     1b0�-��2���֨%�}<q`1����
H�D��z�c��6~��(����y	5�;���#�j8��􉿱�^1��7-9 ,hM���3E��jEJ���8��<A~C̈N�g�7).3��U��4�8�7l\�u���ѐ!#&��w�3�Y�@�}�>ú0�Ǟ;�v�$���y���D�mq���y˧[�k�����;=��!
!�?]�l���>^ < ���4s��tF�.�aDؑ��p��!5�.>��+q�`͓����Y��A��1yD���%�C�\u�Fw!u�׋i��$��;L�^�3����@Ʌ}��p{��o��Z{��D3�NԲ��u�5���S�š�5�2X�ȩ�G�����e����L�x��>�u����$��T��� 6�
��tx���"MbU1XlxVHYEB     400     1b0,Z��^�:�?h[���|N�jJ^nZT���u�%u���Y�n�z3�˽Z�i~� ����;�b5��ӭ-o+'ɘ�ٱ)��.30J_�+�ѳ �3\�3aq���{�a;��c��&F���F�3�[9=��Cu�%�g'ͫm��ń$��Ǖ\��4ηJ���+���rɭ��q�Cu:�bL��0�u�� =3�m��'s�qJ�`��:"�j�͸y����Ӆ6��&�u�^��)�L)b0M�f��~k4^��$�ϼ���e ���~k���-�~�� P2s�x8���K.S��k)<������6-�za�1[pcѻ��_w�xC/��uA����qt?^qT<��d+�u���WK��ԉ����#���lA<��[^��퇘�ZVV�{E�q������ilhXlxVHYEB     400     1c0W%�
�e�x��(��."�!\{��f\6YȢ�f����9���R,�K��H?�<a@�ˤ���W9渣2"kJ	.���}o�Ǆ%!w0����@")��D�m;��}ݥ�ԼY�]߀�"�7ҁ&���%����>��ÂͶ��`�Qc�x��oYy�W��{�.����-��w�����/��7�e�s�����i�rǏ�tbz�.����C�ez�5�Ѓ���CA�x(���+��d�7D��J���>Hj�{�e�z"i#3�R��	��9d�E���,hi�|n�Mxn<%:Y����_9�:Jv��#�e�71����#���х2�B;��]b��P^���i��x�D:\�ޣQ��TL`.4"'�p1^�B�ԶGE��L���~"�S|ik�pըeQ�f{�X_�^���(ٍ�[/�b��J�i%�
�N	՜ [�n�C.�XlxVHYEB     400     140_�(Q���c�	��O�$T(N�9�#�,|�Q"�:&9��P< ���p��h�o�G�>2-�����͚�@(%�=��wܗ��}�+B%M�x�_�T��^��D�<��:���c�B�q���O���͉q��������k\?)e==~$1��̰�K��{���Ag�Z��~�O:,;*VҀ��<�Q��Z�꿯��f|0�O�� �C�@�{Ww#��b��6X�G�/�qT��	l�r��u� *�R���J�7���1�W��"1L�����'�d��ɤ°O]�����Ǝ���ߛ�g�Q���YyhXlxVHYEB     400     190{�>"����7�R�ʻW&���x��7;q�+q�IF��q7�QҴ�v�
�_�JE��v!5o<j�굙DL�rx�1f�ˮ  ��Y�`��= ��k���1�IȲr��v�"Q�˷�J>��Q �ąD@GB\b��;=q=�X���eA7��w���
*��|���z��Sn��w;E�R' ҟ$`HO��~�l���8�(����Ы�\F�2��8��B�5H!��i8�gn;wབྷߢ�̅,�v D���_k��˿"B`�d[V��ֆ��e�f�,�����<����P�q�\�X�\�<
���X��g�1L��(�)ɫ�]��%&���6"�x�JfݍdI�t���b���W���m�\�p�}w��"f�p&:h�$Z�D|�@��ǏXlxVHYEB     400     130ءq���40��<�4��+w�;4�S��I�pa���p�R����U�/��")�8��ӏpR�ʑ�g+��� �X�(����[#$Ν&��K���`����k���=����5w�������H�|�뾪:�'��t�#f�(m4E��Z���M�֗)�Uj�Y@����+^(�}�RO��Z)|zV5��͵���G;�b�&��V"G�R%n���Y�D����l3_�F2!�޺����c��gWQ&a�&���s�C�B���:���M�N����!T�I���5AP���,�XlxVHYEB     400     150?�u�]�M$o܄Iu�c7��=�� �������tr���Ծ�K�G��'�L��J�T��K7�:OIԪ�Q1"����csS�ً���\ԥ�˳��	J��2�А)?/�(��1n3�2>����:rW��ǱJł��/�^��-һ���s����<Rf���B�{���I�e����/���+�g5�B��E���ы��Έ��FF��M0ô�"Z��a�-�ה�Y�F����.�{[�;�M�y�(��eR6$5W�/���զđ���.`�"RNa�Q�g���_��7��d5V/��s��ƒ��$�(N�8��詞�)Z||XlxVHYEB     400     190tiP�_���)4��D��AS'���iݺ{X���x�ng�t�2P����w
K�I�H���qʬ�'�h	g!o��\К/�������UQ_���z"�h������3���s��E�d����߉K���ʪ	0O��:v�?�rF�v�l�0�G�==I� 89���04�������a�r�?vJ�"�\JxY��j�>A�Y/k8R��W:��a:�ٕ5�IA�jr(4	�:Ao��x!�c�=U6�Xd�n_�&_ʑ�tk��t�?h&�v������#����d�HL,+���U'��*"�pLv麯7����u�Y���f	��X!�Aæ���E^G���V�y�pS��<�Z9đ��\��2�{�Z0,��6-���i	zs����g��#�FŏS��XlxVHYEB     400     130�<ȏ���K�D�Rz�[[�kb�ز� 8hU�H�nv���wf�Ft<����as�T��\ҵ�$���p4�g�$K��Q9�W]�N�܍�	�<��\�D}�O��	Ӫ�n��A��=��0�k�-���F�~]"h���E��%����)���P��k�ZTI#��̓M�3�!:^wd�>ZC��]7N���a-t\m<�2f\�m&�zw���9nڑ�<���»rF���rR��������m��f-�>���©�Jʜ��ϡE�ƽ�n��g��v�@�P�i�XlxVHYEB     400     150���<.Q���>�a�����R��Pc�����F�-�����|�C�s�&c)�}`�l�,�i��$�[��"L"w��t�i�8��۶����S;�w+��y� pAr�՘#z�*l��k������3Ş�=~����}1���*ZO�<▾r���+BO�x��O�/'�82�Y"�r��,�İ�m��>0bb۝�A��Va�� �bo2�a��`%m,�01��r(/�ܺ�)�c�}<�8X�5�_��I�� )ΒE"1���������=6���z撚K��[� V�~!�⦝�RP�:E�C��Y[մ�LH�~9���o
XlxVHYEB     400     1b0���B�fט/�!�n>��k��IC���[<�dV�N� */͜�v��|�/lR�O�[�ck�u�9�ǈ�E	[�FؘW˟�CD�� ;�E�;O�}�Vx8(��-��̗��޺�U�L7&���������a��|�$�Mls��NE�߿ܺT2��6S�}\�,��)K����A3� 4KpR�ktajeۄdz��Ɣ͐Sy|ٯ�YMI��u(IHR��Ǜ	��P3��w O^2�)�<U|}"�Ut��,¶�bV�-����f�{Ă'u����beBlF�J�7��x����h?�C���B+�m-��6�f"eɣo�J��|oW=��֨>g�ߚ�t�
�O��+��O�'h�>$�x%q=C��Y\kMD>�@t��nJ�N.�=�O`���N��#ճf�-*Y�Xf�^�WF�oH�-����WE�{�A�XlxVHYEB     400     1b0�˳�� �S)�-ˁߨN��+)d��@"TI=���k?ӧ0��b�o���Z�'�Y�0��͠�T�]>m��;�đ3v�}k鳢�`01���1 ���L铭[y��&���;���u��ze�֨;��}�̤""���ф�ǓCL	��$�@������O!�C�\��a=�#g�H�ZOC"�N�!���D���ņƖn��C%���!��ȿ��p(a"@C'�����i�)�
�X��i2o��]2��3�`��_q��'�EKu1�]P��X�`�}>��1εga_@@�m��Z������QQ�����* Y�d8�2$�%����2�������u�������`�rO_z����s�S�b-^���d��ڸS�BS"����{�����e��z�ܰ1����7��������:?�C��ظKXlxVHYEB     400     170����X�,C��a���_�?���ɤ6d���)�-������՚�ݭi�ȯa���͇��蝄gP"G��,����Ĺ��'��:{��F�m����)���v�����1k���WO�+�$�������gG~"ݺi\��n��!��8n*W��wtl��������̧�K��\%���a�r�Tv.wTKi]G�5\?ĉaK��M����ӹ������~���#�:�bA���<KD� Q��lٳ޽��ІJ��kѣ�1n6aRi�Q��O��4�?��۪���$�νg"9IXu0�+I���c�i�yW$�A�b`X������G�&�s����Й����A���M�?��XlxVHYEB     400     1f0&>��qP�{$�B���\Rv�G����y�!��f��
<xPZ���T�ژ���Pr=�S��������>❑����![F�7����M
�rg��0k&��di����,�p����8r�0t��.�Q�F��T�0��3�}AE�BW1�Yt��X�%j�Rh��^�P[O�36oP[g�q,*?%�kU ��k��Z8�N������5��1�;�_`y�Z�C//\xM�,v��z3����VT���[4�/��6�W�z�4'�O�������O��1��8FsiY�(�3��쀜7$H�λ(Q9DW��o_W��␹�K�T�,�m�`�P���w��8wv�R�O���y�!�;�@)X�
gS#n@#�����rg�P�a�\�G������ߢ����S
�-4�	6fh!Ŏ��ے\§����ª�� be��
�a%)��SAxQ8&�x�;�^�
̉�;����8=ptz(�D�nfb'��@;N@ +����XlxVHYEB     400     130��z�ͪ'��Z[̛�;_8
�	-����wz6RH�{����QÄok&ɲ� Ⲗ���D{:��rrzE:�_�+��A%�\|D�d��Od���^��;���7m�?��R�d�8���)��%��*��xW��N�9��p���6���f��T:�����EAu|U�}�1�����b�C��^s�� {fn@,ƕR�E-��]�g�s�}�2%үu�n�!K�^J��1�|ӑ�%fWY�8t��0q�5���sw/��$i�dl��{���_��J	|/��V]5��l�K�x|�����Y�.Z��pXlxVHYEB     400     190,�n�p3�R(7>���H{*��</vē(p���V!�-�rX���u(���~{CL��/�&]2Z7B��7�k��{8��R�YC��_}�h7��y�Ϯ��j)�~A�I�D�U�/_��Am��%�M��9�!zWB��.��]�K�����M�'�`O�>Ə����\�ѻ�W�!^|�J*GU*���7|�*��湌Ʋ0P*;�D��#�?���]�j��W����b`�h7Gc�	�V3�PSk��K0�-=\��:��+�GM�I{�g���y���A`el=���\��S�{��T.�QOp%�{A��4���+�@�QYE�s�=K�d0��i{.٨��rΪ]Pf395EW��Y�?��7��Z1�8����+�T%A��.̎E4�6*��ݞ�KXlxVHYEB     400     190R}\�����a��ߒ$�.�
�0����m·uJR��կ�FR��u���B��(�B�֖�5+OG��>^mY9*����A�8�1ܱ�����+�V2~Eh��w�l U%�g�Я�I�a��3� Dd�����qɊ����V�J���)�[)�w'�6�sU�d��76Iz��e����h~�8ң��Ĝ�.�D�o)i�*��۽��7e��������Od���WC����T������W��sf1�a�	Q��SY�m��� ����=�@l�Kf�"s�I���Z��k�~>��[+sO,����?�1���?��z�����8�.oz�%S���U��: �U#�hi4	���!�^qŌ�>���B�ε���U�)XlxVHYEB     400     120`n��
&��m����(�7�����$��M�|ѱi�Fb�k��=���=�����W�Z�L��/�U(q[�Az��~��p��#�{�]�R��İQ��	��0�ڮ��?oύ�򹓪�� y5�\eD�z���� (��8��q�Z����{Lvq[woJ�3UyrD��V����O�|�[��HL�I�J���y��SU��:';���o���/i��xsN�A$/M�'ueNY�,����K��=G�����W@�6��°3�?��
��s����~�XlxVHYEB     400     170��.X��XC�t=�n�C�UcS��.&<�݄&���1$��74"x6�CBO�
|n�{rb.M��:b��| l�!"���s�v�R}�o��_`�t2y�hW	�]�&Qw�sMD@�� �d��Sx5]$'��N"�>����&8GJ%��$b������X�l�(;<��GLv�lD��Rh9��xӮ��&'
�#������@�<I���Wz���|��.P`{����'��6l�x�P�<w��0z�=��o�5�dJ��c5FX|a=��U聽U(,��
6Fʠ�Q��M���!��n��}�*��{9*���}��f��)��;컲ܾ	q�Z!<lw8b��j�mi�sA���w�G�AT�Cy"�(��"�XlxVHYEB     400     170�,�樒72��;�{'^#t �1ZB�����GmYU�& =Fͫ�C�p_���N���)�lx z�5��=ᖉ��慒�'#��K�x����Z]ws8�6Nf�+>q�y�$Vu�	�Y;b���0��^�z6�O���A�:�|�޲�Jⲳ�b��Q-���³/V�|�"��I�����Z�=�!"�x�; ��V�lX�/x�z�a����>2騨�����\b��D�qKwt�p�L�tG�����^.o��BM��o[H�$(oh{pc�D@u�}��a}��=� /bP���L)�����H���=�I!?��(oFz�;T��%�k��qߎ>�s��t�C��FJ3WA�zXlxVHYEB     400     180�N��N_�]��\n�e�8���S�?���A=�A��ٌ�wB��k����~��D=��xkF
��� _y�y̡�,V�-�%�ҋn1���b�l)�[0�7���JR����ЖV}��8�ݙ��q%3Ǵ�DJ���cx9�a,�&���YZv���/C;"̘��qt�S�5����f<Տ��Ba�S���
�1����P\Z+��H�Vg��^h��E�	���f����"�&v�d�!���(��씩��]6�N�ִ3�l�Em�c0$ڲ��y��<�-��q��%�}m��<pռ���-��$UT�Q$CV��	����/]�Q+�9���y'ϳġ�q�
���ST0� �f�K<p��Xp}"0?7XlxVHYEB     400     100��L��+��ߋU��R��{� �:�niE۬��Z?B$����� �Y�s!���N���N�&:tU�5�ĉ�]��/N�^�K�hEy�kb�����ei����Y����d=��jV��oM�ҋSQۧeN��}��P�8�3Ou��WX�iU�K�k#�	�J�������ZO���R5�{ }�~9�����75+pԎ��|���22ZA�`���&8g���	_=e;�A�c�"<�1f�[-o;%�XlxVHYEB     400     150��)�(�A�⺱ǽ���K:����1�J]Ɉ&y&��E]���i����x�F�ԯ<�v2��A%�%�h�\�΃JP�OZ=ȀQtW�]D�II����c�`�s��q�.����U�т�=�C���{�ly𒖻��� ���yQ��rK��3����+��V9�9=��J�/$:V���C8)L�k:'1��"�&h�D�S{d������ƦM���,v���x䥹��vYv	/@p!�g�͗Ĝ"G����71�5/��T�����$��GO4�����,Z���_p�J���
pk�$l��u�@e��O��*��VpA/�V0Q�.���=�AXlxVHYEB     400     150��Eu�K_�?����n��g��
T'��1��S�F������ڑ��tW��L�T���j+���le6	�����#���P?�Yr����H?JH�z�\Hx-�E^���������jkP�CF�P���n*YY�Ww�}���3V��_S���,3��^�A�2l?�)Ҙ�(�u�]m��.�9��eo�O(�+�}�aJ1�	IqP����c�ȏ��s����ߟ��dMh��	�������?n��Q��!E��� D�LH;�^�l���Q�K#H�M�D%\�Ȣ׫d�&8f(�QHUދ�M�;t��?E�G+LL�0�XlxVHYEB     400     150��!=3s���C���E܃	�?v���Q��,�g9FI[��0t�!�3���B_���7N�*d,��-VS��c�B�k40*>Q�Lˉq��8F���/�{-�a�����?6��H7���ڷG{�I��1�.���2I��A��������/�������������j��,�W&�im�煴h�{��#�"�U���s�@xF��b�^�p�����nOVY���BýA���18T�~�D���։ u�Ne��Y鍪C��7�'�_��T�[~T���'6���-/8�_[�!�4�N�� ��þM���*;�-�!��vu�.cקr�p1���XlxVHYEB     400     180p���h�7kC�W�>l!�6�2�a�n������5�R4�	���y2��G��ﮊ�fqz�Z�k�Y{�zZy7_ �s��Ku�)�5;[��j=Cݬ��ԥ��v,����ت��J|T(Ĵ�x1��Ԣ�E�<�Ѷ�H��i�]���q�TP�~�j˻��w[�!f�y�93��Y����.l�E�}4IL��w�#�-��W�hΟ��<��cr-␩ �٩w���E������!��V���[��8��\4z��S�L��&�|Vv����JW�3�/9�G����s���U����h` �^��1�@�Q�KF��[X.lݜ�`�#ȵӦ�H���B{���g�G��K�h�CcB9)ՙ���߫#�~)|����ɰXlxVHYEB     400     160$/;[���2 3Lk5�&N�9 ��oA7��۵�J*�Y�+�֖�$�"ؔd�s%�F�@�z��J:��5��h3rv�8Q���y^�*��Qϣ�#�[���_�V�n :Ź���'�πZ�K*�MX�� �( EB)J�6��"�f��m���Ǟ��������,��˭X��YbzB��! ͱi�ӣ���tũZφS����|UQ>䆹%�`@�#9�Sf�븜�W��A�M}u�uu<� � �(��	� י��L~_^R4����Z�!
Rʜ����n[C�����)ؼ�=B��uc�@�oF!h�=;he*�֬��c1"ڿ��Q�*�^[$�~����XlxVHYEB     400     1a0��w�T��!�XJ�}qǿg��"�Q��.]��u#6ￋ�5W��уK4��1���(���-d��=�u�o=�}�����0Z�t?Ȳ�*vҭY��+�+Dm8��o/�c'1��X�~��Z��k�o3f0��=L�p�`U�v�tJ7
@�T(�����N��.u���BL�	�/c{ʣ���W-���v8+��|���Ķ���J��S����O�y���5���o\#�dE��*�" *�:_�Nk|p�aըD�/��Gr�?V�m�p�D�k�5+���ݴ?U'�F�U1EY�.x
3n)�C�#b���R*��QZ���,-��UL��� ��K�9([���?���������}U�HS�^_��Gg����G0��h;�u�5~����Bo��ɧ:%���)�\XlxVHYEB     400     1f0S@g�&�xo���P�k�.&v���ErPܜ�;�ٚQ�8�������b�B�7|$��W�,���WQK:�!�ͰK�.�L����[��L�3u��m^��?^ u��U��G����	R}������ޠ���%t�}H̔ �p]�N�F�#0�n�����*�S�@����&�1j9'wbć|n���������Xq$���k��w�t�S��qz]�" d�$�Kf��-6B��s�]�a�b_�Q�Q�=�w��X�հ�JnpE��ׅY������������� ��ͪ�����,�.� ���&�/�3��XlND�!}���q�$Q�>޵oo9_;��@u��KԳǰ���A��_O��14��ܬS�N���:Et�}�����p�O�-�(@�#M0�/F��71��M�%X	��ljd,H��s��A��yv�/_�q �2�^�������޽���7F��W�(�һ��=(4��LA���YQ��M����ΦXlxVHYEB     400     140������m�gOw�>�f?�����y����G��C�-[���{��؍fBT�5㥯�b�nY �t,o�n�CDt�K�u�d�mA�3Z�X��E�3���)_��(�:2z��]'�,���Jo:�Z ��/<;�d�QH��#��\���B�_d��G�^QR���/Բ�\�6��9���_n��V�~XmwS-\a|>�8 L)�4�	�o0R��|�>�4l�k��Jj�B����X#5'�
����@rS`�F��x�&�O(p�lǿ^a�Q�M�-�����e`[blo�4��T�|0�_����ȰHd��XlxVHYEB     400     140��d������ډ�	Rݿ��1���I���D?����JN�`���//�vF~s����@�����N�@r��k�2>Z ���"�T�f]�7��b�N>B��v��΍h���	!� o�'����}Xs="�bKN'�v�#���bcT�5�W~�MaX��3�ɉ�c�V�c&&"�3+U<��썆/���S�)[��ug���`�[�1�����ނR]Dr�\��ʜm�7��w���K�s��^���K�#>H|�����}�p|n�7.F`},~fr�c��T.w4��9�D��\S�VTʯcj|�XlxVHYEB     400     1e0��}��Y��SvGGKx{=u?�γ�FGXfu���FC�c�;����_���_��ݦ�̣BB�U��j���m;����B�e��r,�e|�n���D��ޓ��R������r�5v���=:�����{�KX�*]�p�Ia����Ɂ�)�H̾:	��q�����	,չ����_1l�����1n�{Vq̀J.��L8�LL収��␙�����;H����!�Z�x�v�~~�g���9��3h؉��vM��e&S3ֆ_E#v��@��g��`\�������1��<�Q^�)L(a
Y�0�C1Ŷ�5DH���w�7�N�<kK�(��	��P�dW��ˠII�T@�E�?����&��۱���'5�;�Ū��+����0��������z���5U�RT����uy��g\6s����Y���q�Ӂ�1�c_�Xv��P�����V9�`ZNkQ�BH�U�{Δ�
XlxVHYEB      90      90�&~@�j��F=�0��M��ٶ�Sя\�����W,��K�H�6.`K��2��A�e����ԫ��2u�S,�K��i��s+Ǻ��Lo�#�:�N���>�֎{V�u���+1E�֊X���T�]Ӷnv �B��R����