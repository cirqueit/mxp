��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���;��ڄ���>�]2�L���.�ښ�8;����u�f~U��� $����J�K(�з[Ad��5����i�I�(��*�3�o�%dU@�Y)�%y�����}�bCX�=<�A{�[�;i�?��ZUVӐ#��7���L_3@�_:��]a�F�@]��(��2����y�AZ�Ia#'	�6���\��K��s�Y%�͍&L����+�k����k���j[s���]u>�Tu���]��ˀ��m� =�S��se�����iS�C}��V�z?]J���W%�&f��~��qA҅�Z����
��W~��m�IlD�ǖ0��|��j�L4@Ż�_�ºF%VQ���wo��/NBW�D��A���wh��,=��.�|�����va���}�:�,��s�R�a&��s����O����mg7�{�%Ȏ�:��WQ��Įսn�0I�Z���~3;&�z��O�Y�>�ڜN�`�Λ�.��PJ@������0md�x�����2����T�)P��;�V<8�ȭ�c ?C�~�������U}���o���8.�ڤ�>�����B	?R��ǒm���&��S]ٲ�0][����v�|9��9��TV5� پekOg��qo��&]�����DJ@7Y/��.G���ECE�`e�����(mOJY��Y0�«�/�b�$�a�S$y�׺M[����<%�1�D7��<"Rݟ��-�)cw�qMnE�R^f=���/P�$Lܼ�d���$[�i�i�A�?���5��X�-i+�뼫��nۨ�{90��+Bà�P����_+#�]r�zX�)���&�`"6f�<��������`�[
�)�uit#��"�E���3"��O	��" y�W���$ֆ��U�H�a�AqŨ�v�7*9lv0�	�N���KN��Uz�`����jA���V��0	��r�qP��m��>�����>0x�'t��K�G|����<L-��1kT;�Uj����Q�T�R��� )t[�'�%�p-�ɬ0��f@���1X^F4p���1/�`X��ˆXg�J��5��Q.ܡt�l���I�uR�{��3$"�@a�$d!�t�`���~+1�NݍB́>^�Z�W�-+���yA�'�A�G�<�#��6�os�vuv�5L��l��~�牴��m&��1��|�ݿ�]�.��oRG�$=@�V��>��N��&,�ǐ�~���bh]v|Y� i�M��\�О�O�Xk!O�):�i�� ɤ.���4���o)Ar�#��s
+ ��j��ܯʓ���i��W��D�Ʋ��/�afd�9����~� �G�ޞ��OpB�r�GBS&��dN;㽤��#����΅�����\����嚢���t$��,p�����-w#6�0�)8Ӷ�����TLɉ��<��v<��CiT� �t�U�6�V(�'ř�<����)bw�Ս"&������/ZF��|JZH~��z�Q�^�ή��}߯V�(�p0a�	�P_az�{܈1IDb@D��I�����p�h�H�����AI;1�S���C�Y������_%��ʟ��O��Z[��q˨�1q`��j�s���9`����.�u2 >�@�/UP���w�uCO���(���d���[�A�����}���=�qS��g[�^ "�^�8I�:'U�Q��3�Z,0cC��j�#è�í�����s��}M&���� c<���F���hO�����jQ.ʵ]b[�4�N'�R�k�c����T�'�($�zr��%(�K���HxXr�{�r�w��������@��PEq�%	�� .`�!��v��\�R�r^�+Ɖ��"Q���PK�G0���F�#_RR�XK98��^����lm��*Úf�@�Ec��k�cc�7L�=y������Ϫq����2�,�N��c�1���-;���5���$��:�g�h�]Z� /�UV�b�*��L԰s'�t�'�`T38�U+Zx�Rz&��]U+�H�?o���I�i��_|�˪?�#Rw_���6P����?.P~~aA�Fs���O4����,���ށ�"�0�Gt��]��,�Z�)ۜ����z�~���i�ow>l���������@1��&�q?�p��BH�����V��;�i��$"�xq������^���� ��>���^96�Da'yqL�[y�KK��4yD�m2z'��-�G%}s}ZG/Uj���=���/�{���5@�����RЯA���B�F�Z!��ٳ��̞D}J�;C��|��$S���x$r�I��gYc�93��m��?���IɆ[�{��U�����LXw��.A�������,�������m��8�E-9;�jmP��j�q�TuX.��Qa��L��0i=���{�0~��!;N��
8�r�@�t���d[wz8�Ν���o��!D?)b�$���Gr����G�`��c��a�L���{��`o�Ž�)I���L���F9:!��9�2��~�N�y������m����O&�������>���z��a�����IOm35h�_�7�`��b� ݕs�%��{�L�����	�@�l�Ň%�r�|�~����ǨP��Axϝ3����`�,�'RmU����ٳL���֟��Q�
Y�@k0��l�B�aU!d.W*)�]c�7������Y�C]��fX�Xj��wl=�	����9���+�P�j�����z��W�߯՛D���uK*�7 ;���GN�4$�2^�\5�A�9l�L������h6��i���!T�h�m:N���2�����^��zC)�:$߇׳~a0	�D\��e�֓1�v�%�Q�	�o�qb����fy��h���v�\Al?��m �K	Y���v�u� �J#k���xϞ�Ь�K4�#�?�mw:�LKq����D�:�"	�!^d�WK�x��Jي	z��;�4���':�}#�V`�����'�o]�HV�о�K56%jiB	�x+�D�yq��\�>��Wz`ίr~�?ݬ	�����Lq�@9EK����N��;뢘)*q+7��6��_e�򝢭A�Ъ�U�U�O;߬��`�C�6,4��2KG9Ψ�۶`9޳�e�t���H&���r���B�N�G���"ljP+ў��~^�qI"j���e�~B3	�y*�8h��?�Sy?C�&kF�^��������1�% <�
Sg^���p�tb�I��H�d8v+��li(��s�7�R�&|J�����X�$:��sI��m�0�4l�FՉ5xi��oƨ���q��J��p��i�%=��K��W�b9�ҥ"�'���֍5_����$���k��3�Sğ3��W��W�ƾ�}fŰj*��i^u�}������[�S>?M4��uZE��9�>0���2���F��������͋�B�XT�jM�W,�n�k�������%h�\Ġ+�' E]6b9�4�f�n9��|d��~�՗���$s��Vj�>��aV8�z3�4\a��RۻI:G>h\�S�I&�o���|`'g�F�Yt��j�C��L�Q��71c�%����J`�׳�@�!��]H�:. =΁��hA|����8�P�5���7T�������������2��,Y^���y�U���i��a8��9��$���{��N^~	�����Hq6Ʊ���M]�B���]t1�ь��FK�@%��Px)���1Uo'�0L$�8b����AzN�9x�c��� ���mYMX3�fR�!�_��I�|GZF�V)��ۭ��=��c�6$}�tP��%���+�7��3�Sl��c!�w�Ң�J�B���ц�p���aEM"do!oWh.H��e�xO�O*v��M���qf�V���`@��N�pr��7�x:_ga�Q�8ШcC��`��54P��i�{�}�Ƅ;u���5���dëv�MA>Zd��ר�)/@���Pt�<�{��o܇0s����:1ڑ[��F<�t����Z��}(�J��VՀQ��b�<��!^�W�J��A��f��i)�ɧX ވ�Ѷ`�\��'���2��h�=	l����ĿC�:��bN��W$�Ԡ�G��,��4� �x��`� �'�8�3��t�jm֒�M�9~�����q�^v����U���y��Pq7��kF��F�96M () �M���e:�q��r��9�L��[nϛeVտlW����V���C�C�pQoMV���T���Y@������x*23Nb��ۜ�S�&Rp�>�d�_�!�3��q�Zȷ�
�	�7	"��`�bB�X�;�y+K:�����&��� +L��\��ZA�6ơ��-�26�b�zS��)	��!s��ިq2�ZÅVն��`��LO��6��#��/��R3���R���m7ݶ���2b
��Wl��2�=�w]m���j>�R].@:X�����7��/�IX�9TK���R�~����b���J�}��P�REK���*Lll���>- �f5'Jб=4h5(��X-��g��e�Faa�x(�ݨ�����b�8-h�:���\�
'�ނ����t����.S�2����*��U��a���ڌ�X�F��4���IE �Gn����|�s{���;��01.�	?s������%n���y7P
%ǖ 'C�Śo [r~��K�4r� ���}�/oO'5d#A�ȵ�f�&����r�o�H(�׶�2�^˻�M��/���o ;/�XFYވ�����_G������;�KB�|#y�B��}���󣸵�Nq#��r%LK)6�.�6�0ɘy1o6lC���3�ؗ0_*�ܘ�+Jq):��~��f�'|e��C�s�������������nm�Z1���n�%�ْQ3~f`�|W*
�yՉ � ��'�FA`�Uٳ��T�⾥>^�I�FC'h/�;l��nZ!#w��q;� A]F���xr�!n�_^e�� �M>�:�	C,h��p��%)&�e�ml��@�@ɓ�fD/��̳̏\-�cW5�P4�L ����j��߰OM��;���n(�=�1	L�=B�>XD,��Y*�p��+����4o2m����fG  T����/n�d����
�X�����N/n8�vߣ����/J�p_����}�f7(���̸�'�P^P;=�P��d�/���p�W>t�;2�PO�e�]�X'q�e!�r�NJ	���W�$O��L6F�����W����D�2s��v�C�O�73��ɀ9�t&tp��+P~�Hs[-{Aaad�m����E�1�IE:�{�4�F���)�4��{�q�_*��Ѩ����{O��W�u.�Cy����~&<��6�伫�#.Q4����m̊���Xz�)}��!����q�}Ǝ29���8E	1FE� _�2.��nSx�F�����@V��C*y�ݑ0�����<fï^�Ao'��c,��[o˳q1��� �e��Cw��O �$8��ϳ��:�!A۾���-�?3�V��ă9>�*���da�s�r�⠹�k���$��.P����o�i�sW�p�o�N|��T׮n�®C�M�c�"vsX���N��?��'OƂ��v� �{=ե���2R1pS���d�n���7"�����[4kI&�2:�6��< B�G[�4��g�N<�ѩ�#�Y�3Gp�W��8��;�Ҿ:u�GN��������{I�
�^���WZU�j	3 zQ����5k�̽>�-�\��޼�Ybj���א���	�33�=��v��U���m'�q�2xĢZ,g��(Al�\�E��(]��p�m�U�7�I�v]O��s �رĸSSy��A~8ZV�'��r)��A��I~k��@�+����)<*2L�Gr���!� �gKH�����} a�ޥ��Ɖh��b��^JLM;<r��Oh2��0(��[�vD���;��|�N�i%^�$W��Y1\� �������d����{n����o�4�t���_������l���[�9x7i6��+������Y�;w��4<+�����+s�^�����h)��AC�sL�Yg�tݢ��߷�$)��ȑ=>u�� ;����`���S#]��q���|\���ʠ��?�Xhe�-%�d8z^+����C���v�]ɫ��@GK���j�P�_���|TQ�dQFKi���i�u$0�������XG
����`�lH������S��w����q2�&k���N����ì�h�҂O�ܑ���d�l���%����.kt/:bTSH��F������[$�?�0�����q�_Z��g�f���eh.�|�@���Һf鑳����U����p��i~�[WU���e�`��h�� ��'����_�3���X���S����X�����zq_[m�3�" R�lIs H7��ǂ��'�ᵛLX,�L_��0���G�����J�\�5�c}[X�a}����/������߹/3�a�K�U��mE��iC]k���>!ֹ(^����k �Mb/z뿅�]��v�ئ��n\8J�g�:���E7o�բ�<=ꨵ�K�$[�Wg�Sb����7���h��F���х1��Wٟ2<�L�Dx�=��ݴ��;�ظx�jnu�K�i�L��)�=J~W��%��Z��$�W�S�t>@�W=����P�U��"Z�@��CA]ho��x@�����N߽�h:Ќ��R�`
z}�ʕ���صa�X��zټ{M.\0��a�J�,�o7�r�i��7��"x��HL�-T�86�I���>;. dU6GD>��P�֧t��C�����̧��{��1E�� �A�S��G�g�Z8@��$5S�J��Y�2n�m[�y⛱��1�ɷ��n#��6�8ڽ�``��3���>�%�<��X�q�r���gdD��w�`�@���hP=�yEMN#���8M�+qu��}o��ԥ��� �+j��%��p�][��$����W�'����8%}q�(�G(|=�.�|w���x�e�����<s:�L\?O��]z�F�ش���Ub?Y��a2��}齐�!��ET�%�����<:��?��^7�L�6�:����7!	.0z�6YxpP��↽��K���$�|�%;�V�_e�b�%�fV���1�p���,Zs��G�j��w��B�G�9�H&M�yQɡ<Ђڗ��c�^7rZǉ}���c:��|�r�VA4��._
���4[e^���ہ�<UD��-+<����Ba���1?X��0�q~�|�9��R��wj�@����!���}�kTōvy���#J�ApB٣:�,A1tpA%"��=S0��Q�Y� ��
we�	�0�s���"�U8}�r����R�3�bK�(R�P�7/�x7�&Rm�_$��-p�p�y�c$Ǫ��<�pܒj�R�e����!Ǣz�F��_�Ә�x/�^%V��'[��!��am��`��Ip�ٝ���q��%�ÿ��X��+��rޜ%�����������p���>�8�Y;�įH���zX��S���e�9��%9[�m�#������_B$IoB�f��j$�$�TX%���q[�+�Ef����ر7�E�4Hd��A�a!`�=��ƻf�,�����,��ٷ|�-�6N���w�(�DU�_��\i�G����~Ikd��.����;�!���X�	(�$��="-�����
�1����|�+��(K2�i�k%�ߘ�.5��L�M��3n��.�BB���8�������.��,��G@_$m���\`Wc�o��xq ɑ�G_����@�D�y�)b�67˾H���9ޙa�X��u�\4�d�;q���j.��-dD>K:��/�Â�����������.Ujp�g+k�ds����1A�y�`�}�L|�g0;dbg��S����6��=:�&�#��0H~h�0�ߡk17.DAM�@�1�����k��/�!L�S5}��V62��{w�%w
%;���-G;��K���f��P�"	w��e��laG0�nzڛ>��0�r�Ď��- ��+�jG�E�a�"�Po��ZV�	�g����=�Iɪ������xS���N];^tql=����ss^����
l����}�(�t%/4A:t��Q�n���)wI7�#]�N,[��8Q��q7"�ƵʵB�X
�0uBT�0�]r�+	Ƀ�MM�Gy����G��:y�;v��/�'�����aLl� �5>4�"J9^E��X7�H��=��S⶘�Ɯs�=��K5��W�ܹxf<{�mb��,@y�:��*O�����j��6 ����-�0��F6yve���o�S����>$���ȑ��ĕq&2�l|���|-B�6@?�{B�޸�J�>��������gx����7d�Wr+�7p�l��G���[����k�D(%��P�xü?�|%���e$��5���>�#q��1��9�6p�n>�ޣ���|�x)'*��%��ė2=M�g򶬷?X���M5��(�i�����8�'O����8�F��U��VFzV�E�G�+ok��D���R�5#ϴљ���Q��j��w���-�/�qA�4��mO������MOfHe+#�[�I�i�.-E4kDW�f�3��´���.��t�8�� ��-�h`����,|��х����E�/S>���z˞�rd���0�e�C*�Re�
ݭJ�h��^���jǕl�ժ�-_�檬�����1f�rSTJ�������ʁ;J{�pz�����|�(yc���r9�V>��lXcj�\�35*v��Kk�U���$��̲ǙɊ�M�r�:\p b�P�[  y\\H��?B����A�,D582��> ��&�c�ͤD��<u���Y��`�Y�;v���vkq�6��l�g�)t��ӧ�����6ܖ"�|��]����C-�&wi�,'�M0�8&^R�'�c��k̘c�I�]1�_G�Lc��!�/���}�19��w��J*kf_y��H��ϕD&��~���GM���C�����X�	ԬO[`;�@�} ���9�� �3�+%�<a��C9��f3��Դ���P����8
f_�6?Q��g��g�g��Q�nI�ى~�1PцT��)���&�|��N�=�=��AC�y������L@�}�<0�����@���}w�#�z�吊�d�@��h��Ā�;di��ߚ)5�W����Jr��m咚�ˤ'z�0�hٲ�L�|Ku(j5�&H}��؝��[t����ls�-�C7gl7�
.e~B�=�$M��O�	~����� ��ҏ���]5z6�	��@�Md[Y�v�N{�sΆq����7ܢ��$��Վ��g1�-:�S>����N×2�@�и�ޔ�I�y�k�"�s���!Vvh��Z3e-J����A4���=��?��� qJ�Z��"�z��?�ӵ�Y���M�l�͏	���V�]��0/P����?qi�ۥd6��k���{u� c�w^���n��(ˉϨU�#b뢩����Ȑ_J+�q��i+�������>X�h�2��!�C(>R �h�SP2$vs-�l6��Qt�$R(
u�w�0fIڭc���'ԙ1xn�u�j�IUt��w�L��ȶ���k�p�?�L���.��#��Z�ÞC/������Rx�CRnX�8����Sn�b�\0�^Q2;x�>�ؖ�a�}��oR���<�3�������ih�!=-������;"X�&�'�lÉ�:�IA�iSܐ�Ձ�}�������3� ��HN���gk�E�Ō���k/��y=e�E���e�i���Y*��:�t-�2����W_Jnx~�e�ϓyIY������x��G�n�	D�7(_b�AB��bU����w�i;�=B��3�`Gxfp����8��?5��h<���Z�/���g�%���ڿ�l���	�r�g�ti*5\]��������빲	�${ ����*t����~�Fs|�նt���Z�k`�N2�U�b���>4!��z�&�5��^j UX�{��1�F�޲K>�Dk,6�忂P҄���"�BRn�$�҄��Is���e��?<V?�z�bL�:��S\���5õ�>�z��*>�;3'�Z��WLd�,?;�D��4k%�%���< U(N�zc��I2��cGn�%(�8?eoHG'���	��r���`��2lȗ+�o�İ�xV��B��Q`���E�A�
���iw��ވM��+�J�DV����V�7}g�_�#�6��ሲ�w�,���`��>��3�I<�^fѻ�(��z�'��Q�,>V����rP�a(��������,h,��6"����Q�3#�Vj��0�[Ho�4��VJ��LZ���X�P>���_dX�wܻ%9��~*���i�����/�%3��v��j��v5��i{ ^
X�'p0O�O�B� �|��v���?��q�%��|�ķ7z*����c�g�E}��%�_��w��VBu���s+�A�����%�����5�����4(;�*��{;\&{Ө�Y������o�8��������"��&O/�ndg��ArY����z�cH����\�l !N?����~ހgz����\��Kڕ�˵s1����`�6͈�啦����)�1�Hj�w�a������Vn)uI��������d4�ZXFF�r#U<������$%�tT���.^Ï~'��d�[��73�<�K�]�W7�A^�
���yp�aZS(��.�.�&9�!�m��ɛ�#n�R[��f�7pV@�j"=.��ֆ�A�������u����D���f: &��tc&�ڢ��n�<�{�Ćb�!�X=2��@\�W���NdM9�!�^����'$͟�{�vw�4MA0��`~�+�^�z�I�J"��e��� ��D��b0s����ڋe=7�7����B��9��B�����kR�O�i��ǡ�����t\��_r�U�Z���w�o��Cұ�nd����!-�����0fB^l[�8��qEs�n&��n�3A|����j�d���ژ�h���6S���N��>�P�7v�����.榍^�,6�m�_��ϼ�N�A΀��61k"
�����K�0�<}r�liz�ղ}��l�n�����a���.�F��h��B���c &K��<�gT~��O˹ɈC�����Q� �H�'8���1�I?�B�v���|��Lm u�D�MLZ�ʦ/^ni�o�&�e��Y��!cWUz��G�2�$c��w�����a��w��(�cL����u�Vh|��y(I��+�ۓ�R������]?��vb���0���l�=���'B@�j�[mgV�Jd�O�>w*T�J�����s]�0��oL����i�$�R�ZFH�'�&ũ�<��	�v�l����)շ�l�LdԮ
Wi����>��b��{�Jd�Ф��`���+���D�������&�΂igv�����zv�B��i�������&3yP�\��,}:��8�(���/5�:�8��;~���a�����(a7�Të�*�ʍ��C�8�uu9�5�#����Z��"r��vg�X��$ ��i^�H���8C	�݅�.� )�;y���~>���j�)Hl�)��Ԣ-8Jh����{��e�E��u�q+<�{�!�p�L|���ml'H��u�ym��� #�2kv��L�͕��4l��6��+�dV'�Z��g���Pt�f�l; ��9���O=XW�}y�:ɫAZ/	z~�u0R2��{0$�����֐5pjT���V٭�g;<�,��مv���c��.|����w_�k�����#�Ƃ�?�ag�<;o�*��<Ĉ��OOm:���a6��+}�G�c�s�u��D٤�>�Y��JKoލʳ�V����L_�k����+i.��t��K��q��g���������ϙq_;C,�9��m��+ۼ��FY���r40����s�V��Qt8p�D�3s�<�H��pĈs§�kh��'���R�㏘�8hU$īs����˾�|_͉F��.���yo�0�C�X���p����j�j�9��s��t���{+�7�-�7:�夁��x������pL�E�2#�F-U���Y�Azh;{���O��n��W��:<��7�!��N�=l� �j��s$���"��pc%�?jx��n䨨�rͼ[�<;;Ϻ���S��aR���1���ϋH��w�8���H�T`������� ����a!-��r[]I�	�X��l�f"��:q��%��+�,h 4��ۉ>F�j�&3D���&he��p��M�N��bE2���=�QQ�4C�w��uKdcjH�t��9���E�{qU�"r��S� I��f����"�j�4:w���)�F�����ܵ��˘+N� �AM�%��Z������v��^!-��Ǡ}}J�a Rf����#E�a�j9����SL�3��1��>�^�_5i�"��Џ�i��x�3+���=�s��{�#�/�}�,���v���V�
���q���5$�s��v��gO��6A[/`F���y�N�,IR����Ցb�Q��uQ(*���T�P�-��B��:�!Hc�R�O�j��D���DX��S&+�\%t��{�X�#̹|w}�d�=���0z�S'���]��	uۍ|ΐ���p���r���^>����]�ׯZ4���}����3L�3A�s��x�f�F�5�J��T�@~�'�3~xVAX��^�`������*,40ߤ
��>C!��N�5���|;�t�����cJ���C���V* |�i��߶G�1���l�����G�PԞ�gY).��r>�����3�MRA���KX�t�,�z[G��O=\�s�?Mٻ2��&*��8�Gr��.fr�&L��Ģ�gi�S���^ެ��xr����es��fFr�w뢮,��F������Z�q���XD����/q����K� 	u)XW!Z�{څ�M,҉�UKy`�(��0�]��bW�7mra�*q5�e�W�6��J��b,��?�o���~�p-Ж�f���ӤT3s���3�zt�3۹+��n�e8Y~"��o�^���)�9g�gz)4�
�m�kb/��3�|����K����ʭ��~�z�lJ�<. �,�KPl���
	�3����x��)��~�r'�y�A3d9�����E�Q"�����ǯ��]��D�v_|q�ڝ�>�\�m���Yɻ��r����M��\������l��6PhC��y`գ�j���*����|�OC��S``�������9����e�Dd��3�q`��Ѓ�=q]m���z��
�5��׼hGޮ>'N��@�D#��~�8�w>�q��+��(k\��p̹|Dców��m�E�8����F;�,F��d�V̓�<)$�.�]�t�g(�C��Eʛ�w�Z�Ԟc�0��{v���\!��Ɨ �]�WI�`_��4�ݠ�2
i�����~�	��UC��ܕ��V��<ʜ1[�-�LV-�Cř�	n�~��翆��s�-��ѓ`�co�74����o��M�o���l�*x�t�/��]W%����;�N�׈����m7=O%�XK���=�^׷+��Չ��t4>�H�
ي�5T�|)#�q��)�7�]�m��A0��-�VX���j� l!Vz�����)�>,a[��< �����R�c��t�ĠP��Q�'�C�?����� ƾp$~�L$;ݦ/?ڦ�֧5/i����O,�q���G�Bf���?���SS�E�o�x(AWȩ�B���{:���#��g�T���ڍ�5q��>���:ﹱlK�\�&��"
���
|������V�JG���$�]��~��?�^แ	^�SL���:k@���Ν�Y�%[���	�>����pr8buk>� ��D:nL�ْ�D�-�&��@,S��Y,R��C�T��eׅ�5��� ���z�-�4�I\�cI��OCåYu�/�<�ٗ���<EY207s� �\g��Ĩ�;"�'�Jڔ�|���Byh��cGF&-'�!�[H�����t�O�,{���L�!%�qz���z�����L�����ъWX��.�kCV���������7�j���Ӷ��q��K���
{ ��N�qǗ�k�/�ZUq�4�5_bK��B��v�&�G(�w4盻y��AR�q᰿~�P%�6�.��k;�6�� H/�6f_�[������1��k�v�>�>����_m<P����Nv����[l���3�?�K�Eг�,�ZOD�z���Ê����в�3���X��#��x�!3A'i �o0����;�`W���aF,�,��-�6�v��p2��]�,t�y�Z��{�/��xA���1?�Ջa������t�P�O��˻��������쫲�S�m-
��T��<�Mr@i��Ѥ`�4c�D�J��dB0�Z;�nBq�D�8��Wd�$�	0�F�|QܛO�a�?��,�?}�2���e�N��I>��p�F��� /��� '��1�u���Ô�C;��5�s�ۯ�&��SƬ���*�eflLZh��@p"ξb|�9����IC8ҁ~]��5���z`�����$긑=U��Z`}Ա� ǅicX��I-�V�T;�V؋��M����K6_��|�����1k<+V�Ҁ/<�j�.�fU#���u��?c�����)/�g5IO0��%ȩkaH��I�2�l�ʸv��Lk�B��C�g���(�&Γ'��]"0� ��^wx��R�y�,)=i�1�Xo��H+{6����9X��h����������^iLQR��Ϲ��ǝ�bv��?F~�����?z���k�,&�$7]�7r���K�v�۔�#���>�Rl[_Aa�T]?�	��S��fOO�9��a���³��4?館L��Ad���fwV�\��m_fF�K��7����x�?�j�Mh?
e� i�X"h2!r~��Բ��9�X(�BV�x�V�u�-��E�DVu{~�-E�3�N����h�Q�w��x��L������֔�ZB7&���7��k�c�ƴ+���
ͩ���͔��HMk�����ڻ���Y��-�p��!�5y!%�_��D�撌?���T嗾��>q�'���˽�fڄ�. "��W�J��K�P�O�Z�(D6�����1���zR�6��"d��`�e�
@��F��&��y|D1�9Z�*�KtoLJ|�4Vߤ���B���15&�t�e�yg�v� �9�iV�Ɗ[x��ɀD9�zDҍ4��-}\:y�U;o](���� Z��~q�_���"����<���^�Hn�M�h��Gtg�e��:�f����U	?�0�� ���������ǹ����Ɯ������}��N�[t���j7��gSSQr��z\\��J� ���R%N����^��W���9�1�{�Wo	0w�]E$i�/i�M	��Nj�Z�q˜d�f>�
��o�ӷ_��m�a8�FzG�ӌU���/K�X;��g$gN�غӸ
Y_VdF���;�b��Q&���Xx�Z���^��1�A�	c����8ǌ���<S5/�T���[:f��Qq@И����i��=���+%������CMiX�L�5֎+��D�#�_�5�%>!ż<�Df)��!�6\�d�]��%j���p��nS�2	���<j㳵`��f�:>;Bk��f����.������nV\I�x�����sj���z?�Qu*�֭�}c2���ؔ�+�p��K�x���S3�#k�Ώ�qL�-Ҳ�*�m�b.۸Bgf��]
��� �!���	`e�'�@�,mτ�O�q�[3V	�#�h��3��uI�sM�;��۴t8'ce���2��q��>��̼��J��B4fW�B:䯻Lč�������E1ac<3N�8�St���7�4#U$�����_����_��?��NH�!�{�<���E��\-��n���h���/q����s;�#���X�a�{��=2��1t��k��'zN ŊUEM�!W���=ysM����24y���?'
~K5�r!Q=,���N�YpH��ވHh!���|����Uǣ�DZ�V=Γu��X�i�3 /�u�S�ٜ3�͎�bv��cuP���d���-�:`"�����ձpl�����vA`�B�w�����o�i���DJ� ���T��AH'��Ùo������:)�T�mM=
w^�6E �Vա��5�\�������;�ۈƜK��
�xOĸ]H(p�<1 �Q4F9r{.կ��
f�����S�����$�Iĝ�R��0lʧ�����߮!�K��D�MD����<]���	���e9
TͲ"����"�8/��.,��n���!�����Wp8_ؾ+��<A���4���C;)|��p:��$?|)�N![ǟ��TAb�5�w_�hs�ͳ�B�̹9+"�b�7h���Aϡ�7���vܵ�>e�Ǔո^\��ȡ���r�E��\��ͫ~���[�*̇YbT�@p\&˝,��O?i��	�B>��'�cӽ7�g
�{ �~��m tlQ(,1������a���Y�a.�)ᵫT|q?��A)�7U��f$߮�z�*��ޣo�%�XIt�RԆ����rrZ$����q�'1�3I������%�7ug�2Z�h�x]�\�A2�W��|��(w�2֬L&�s趢!�VF��/�uR(R���n I-�ٓ�`!8���U���E]b�<~��|MR��j�>}0 �c��B��(�ɢ�&ƪS.ȐG�gt�"EG�t�(�K�|����\u��%
9^k�w���E�GQ:H����A4�{�r6p�}�D�Ά��98��߈����ӆແ�ĕ����S2��R�����ނ^ W��(�e������/]��\,��p���aA�Y�μtl�����R�|�p��5N��:-�#�c�N�q-�U��>�~p��i�ۅ����-\��8�ٲ�Lr��֠��
�mjJ%�Z�s��n�M�n��3����������B�]8>�0Ch+�R�W����G����!��H��K��Α�'�F/�^��~�-�ن~/)�~gFU?�G
eW�[R�
5s(]P>�)�a����BN�LF]@���CˉF�*��+��˦���R��NoV�y��0c)N�������P+���'=ќ���+�:�	;�#VN5�;�����꘏�� �����FG^�:%��J�ߨ��P�y.�#S�D~D_�~p��,1�c1�������?i���hM��5��jV��I�ꔸN������ ��rp��\�.�����&͑����U�6!{U���C�p��b������H�}�o'��� p:�ڶ\�%��O5��۞\�(����Yڸ�k��$��$�#v��
�����7!��s�9h)vS����@�/�Q)~yI��D�P���f��u��O(�Q��
_�R�;�\ے�9~έ��Xx4V�$C�X	�4}y	�T�,^��,�4}���q+�%X�k�kb�>t�YFnï�y�`���272�n���QΤ�N�U6�,G��K�)7�2�P�,��