`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50720)
`protect data_block
q1OBcnf6EsZNl4R9pwrxr+oGd3W5JnqVv0XBtDza983mj7HEPAJe24/vOCckTU0Uupba2xq94imV
zzSeDM2xnZpOzAcVnm1MraRBpMZ8oRXUiZS11N8VPtuC56Vih15jiuuuVy55FFRm2ZH22knSGp/p
1772UGMbcuVckyv2obRRWMZsuEaOt/QabjHW7SbV6ibyZ0jO7CVt88diLPQBJ+Q7Sp+IKjZVewKY
dj2z1HAElcVAPxgqLb46gzviWAM4pNkh8CSvgjfTV2q7UvVsPT4jqO0d5I9I45je4z+P7m8bVlqb
ZUhmhnx7zbqt1LCT/HZxU69YGBtSbKh2PdjlGM43R5sNQz3AqHUJ1qT/Os5M1jgQZxaTXjFGY7gD
fsKmiTLUtk8m6piJbFqqFkZUwBs3/mUL/QxBs53Ivv3v0h3qedtBIpWD4hCwhJNaCze3nD+JdepD
TAIAM2AVeCXrJ1sDzObPocF4nk/HXvX/hbDIW+AX+uZtIZEeIkNb7i1Og6qLvcPZFU0TZeR9tKAb
qaFp6cx923Wrgxh+PHXtui5aHWiwWXJ4mku99lx0AghVNlZQ2iRSzacTb9FHlunRkBDGIp7z2RXo
gUF6Ih+5xbNsXU8exEPe/l5Wow7BsBB17RO/m6FVLFWp/WHAUwxa95vnYPiBLY/V8esmXHH3lLeO
vG8oAw+uTT2UiPzEpcI8d0/0mEzmzbXNDmf3/P6Uq4hWHxpWZXxSMgRTAq3mBdeCUsI+mDWEplRi
1BIUO89oD+AMPsdtThJ9ppqr1GjAwy0/kJ+PyOWDKlMyQssM8cbMzMPOQwW/fSpthar7GnQRLKGe
jCpzKQ4j2ws/6wbD+4l/oa7JA+O3Z94kGLwjYnl/swb2X5hmS5BimHdcS9jXb0KTT4+BxTyEdSs+
sy+UEW+PtujKOTCg20DJ76+ft396p/f90SpDITQbFO9tcGAArBeqwRfSuI+/eu/OQQRDeK2j9+hY
2xDJQHWJwm4lMZt5QztLg/q8CIinUznY7yt7yprst7UKA66jBaNjV0jDJkWQw5A7i/5Yn9rux7yr
sX/+NmMQdF2d39n2Pil/DJ//FzQoSl854x+cXeOpWkASOKyiy4V1OtRKMj8SdkYJcZMwLaSW+8lH
1keOaPUcWJb/eI2qD6RyolROXXPaJL1VaAbFrnTgjqX45zcmT4mLz1aUns65EN8Qxu2UiUJOOVsy
R7rtVhHomXtN7nj3OBCDLLdgEGjewgGrr3Fo5g8BiH6NVL0z/hSWdbgnhBzrGSY9Pk0t5WHQSWyX
AI4C+GbxBzrcni8gZcwZsC9sSuRjjHZddDdcMR2MbUufGR776vM4NKV6/z0ZjGGxTzZsEF6GqU3I
qFKtrk96FV+wKL0NjfLm2N1Xl/2s/iwBWxK8G7OCXmGgWKlEXFcu5dn2nFm7RujPT3Ka2Xdfx9Nr
+imOJfc51T5iiyLX0WDBA/BrvXAkOTqZP0QA0GP6S5JQtYGE9WGAGmwd3n3YsDCYDjA/3eoKS3sF
wP60bRNRt4jRAepep6a364bjR7swh6P8ZRxE8DIXjfv89zAZN52FcBJt9Ift1mmYvVeh2vYijKqN
PVlXKHsn9Q0KRxQr2RoDF2QRQilWxbCSVVOnOUqr++RK/iu5UKmjmUPcGlP2w+RCCB+i9VyQhsxD
EnkXeWlnQzMo9i1hXg9+XYksoPs09qOk5gskNLpLVCBX6GHOhFXVzM0dBqfJ12COgX5M3z0goF1l
BAe1a6vrr/UMYB/K1jhcL2aRP9a83rAibtw2Y5zJGlPQX3vfHWDkJgcOSXo7bWojZDBMRPTc5vx7
QovtEMjyYyllViwWFjFQIffYHl4rat725xKeakVgjvhcw2TAn1hD6/8cVMNRIQD0SyZiE53Qggh8
V+1+vD62D24PPfELx90fIOlmagkbzDzR70vX6OiGZDHBSU7j18V12qsd8wBR2HYKs/6gh7wovJNO
DmpBNmRzBVYGa/fc33z5qW8vTFCmZUF+zh3/hfvZah8x5bl5HSqh37Lm6W2buh8/qc67/zyofO7v
2KgH4AfD2GYgh45eDxK2gJuCQQ9byZz4OQA4LV9gNfpnV4g9KdDZoJtD62/YeBmi9Zqa+wKM0Khu
rKbWQoB9NOzYlVeKT100V8Y3RrSqdpL/pivAzz/xOy3VGQgnCNJuI6sTgtAcrhCN3OQeo9vMILK9
i91zxA45jgPLRCLgYHkPxKNO5cuT6NwcW1JdI8YtQLRufnUOkOwC+RG0hX7RbAG07GRzYMkgvNoF
G91UBQsQwH2jsB0W5atUdB1VFpNgdTyU3pe4VxGfnWYcUzHclcJsG1laiwDrK7IoCphZKhG46CMD
Pu2qw8WcO3M9RYiq7B0shnNhAjnPWniCVthbKKGZMP5reI4EkP4rzOPexArvK2LJe+RIdGO8O0c0
EWOUpEsujXVJ9iS0ZLWUkWPVGh1+4o7oq3DG6fq5oCGqLiFACkoFLv146CncVVENP+2/FZfuHXLh
r6L9qDDeleTK1qoiGLma3jR5F5ancljiNZW/AsmgD3/4+dH8ygPqbTnYA946KYQGmJIpjFWyXlcw
7QuLDD38MIJ9ESvLMcuBixW8tWiFRwAZBXzccq5rR1ZYLZIzk3JXlw2nXjwkzSl0J3Pri4A0TzwJ
YSQqH/f8ZkHAd1hPJqzGdPifvNb6x3DC8sszNxIxAHYL4XwTE7OnGW06PEP2z8hzRc60Ol9jLGAW
SyiHEX/gyyB8U0IJ8pDQYFTdfJUeWCLCLRTnPESn3llBtxpDzisB1KGNvuNpeaMMxKh9YyPJ9GRh
NQmVSejobwmVKOaO9GS2mUSd7UGCkCnvNXBDFbqnmscu/J20unEx+AH6o8Mo6eScVNkIulOGMVM2
zuNzv58W2BI5a+8xYZ4A9ZQubqTgoqc5g78QN4HRMiV93U+C8tib38LQ6MbsZoXBtursE0ett8eB
8fjv2tsqMNEGwlOibhOazYOlsEOK5ajUkVhRntE9gyqyEz+EzlC8xExNHt5wKgZKrQe/z5laG3BS
466x6bI3z11/IFoRDh74mKbP6tRWP3+MWwG6juSY+V/C2PJIVEvF/IIZzCL320MPIxvB3HTBf2t9
gecHJgFmdfDOk0SK7xsG2YlOluphq8gktLvLxYzQLm7bb+YWViQXtXQI78RniMzUNk68h056yznZ
057CIE17k5gw4WvO+2wkakAQJ3M0EXz78eEmphlzY1hMXsIBPZiWqFIE/BVOhHkgrZh8FcXQrad+
XNJTN7mL0oYRN1W7oZmt0YjhzM1ukQG2TjKijCHAMXlDYMQQwATfP9LHPV3GZ54IffELwd0MdLmY
NmSCw2JcW87L+r4Y6qMHyuoYUOZNKC5lx2fahBjwWDmE9lH04sDTWrjYpKM7zwRyCMvcXoD6RuJo
rA8hrN0KWLwHRGyAAC40NDSSkBfcLL9Hk/bAxoffbxMl0CI2cxyqzMw1OX9kda4h0uXzuj0LMWU/
ff9UVNHq3A8h3z32RjH4qeUISiYqaCLSLcOKOU2aUCz1WyJpnqKPX3Rwt2q2OD3jX0ThXdMYOK+o
4XXyyse2UJMIa/lY4LDoPE7phr1kaEJCZ7wTHiK5D/4xBBPVRcpE0voifKbzRe+IpJr7MLubvtxV
msRTNEfQ9wIAvOaqUyl4R29wwgaZqg/z4xxnYyTea1nynxmD1k5RLpcaNdDp8iNIeWXg5k8U+PKh
1l3QBJlBk+FfYIkE7QP3vRy1LLsKI9fdL7lbxfqITFhuPuTYimy7ElK5qO+6FmjkujWxygF3W2pb
Wy/OZp+Rfw4UwzJyu1EThQHydG20CBBHLRXK26MKXtPRuhKKixRUvE7K8nhNvISRVJC+wvrv4ete
0utDijFQ9l4vBoFudCUDwALbjyUMVjOZZ3irlAHZjy3k4i5+988+wY7iOeSAJw8nmWQsCFySrS8w
hyInQtbtRfSurLClFMtz+FFcMCDu+zthkz6tZy2FRGzR7Y+iurwWBkewaitTDExDS054Akbp7jVY
qIZLHt+/AbyqPuNfMvSH9esiVKdU8suO/xWUovNePQ625Y1yUXasWl8bESaz8CeMmfU+KGviw9Bi
B1lntyJKg4ozhZr7w2sks9zvNxnfjslKZLOEBNVHpqnPh/KVyVE4Qph7bAtCa7zcXIGONdIoQXlT
v8Z6jCaq1n4m9zzsi0uvj+OW4++V1I6Pa6dK/NrF5FHVFkZHxerBhypjpCcvS76Ni/YFMiQUEIYf
ABeOR4z/WW8EbZeWkTFJe+QKmDD0gpQErmvtS6VyHvBWV0+O5i3vg6B1/L+B6qRn2pXXuiwnkxhF
/zluo3E1HZrN8grxd1EUF1IjyOYG9eW4DLAXbCDmtAGtFiEuOsz+uNifnv0Ec+8WPztMsxjORGPe
qqpSUE4TpOnnj27Df7DlFciwmKqIga6dbec7qpa6b/TnNqCICuD+N3hVuYRTU0Do6Tft4+oF9BUs
1Z++I6eEvxhBI8kj9EskZ1SgtzfC5pjTCwRopLixqaAvk9hvtB2E4V1UJbTcUt/lS2txXqJXXr5a
SmutxpwE20laM9fzDtB+wynERt68CseeCETunvy3OKbHg3+Y89qV0B9M1R61aadr9eJMeV69kuSV
P9RiZBjXe708BC/aHDRInuwaaaANmkgxj5+AaTX45lFect0K850UbDLRyruEiLgUFUzAUNsdyIm0
AQijzq0HSx90v1jLFudjyr1Ysz6XO7RVrIYOZ3xxfLQpILul6zNcWVO2oQx3D2aw14RkJdoIHnLj
C+LrL5ZkoTzWQegLptGtbtz3m73ltgfY/wTFy+ZzRuDURfJ6KAB2ZlqgtbIgi5ek8ZzxMKH/llgT
RxeNP1MRZnIN7vhIJgd8GURt/i8p9HJJlTKkQo/2W0+QQTRYEJLge5diNx7upqTCa1BdAYsi1HYn
iwV4ArVKi9hXw+dxaEhv7eGymAiNYQA1+W1R3JxxSERgpzxuWTlBUw/rm3fYOy1ia2xo3aZr7pU/
i9jnI7tLoqV4QSsOIJEQ5eywZ8xJaVADhstubPWNSo5vbVytVDAfveOZf8WQ2e1qCDOR193IcaVf
31GCvT2O420goCM1E9KGIV6L2YJ2Il1r0L8dX4oICc8CT1mbwzeEKty+VkUx4zMw7uJqWgixVA5/
HGBJPL0xMhYV7vT1NJ/qFtZGGDmPHxt5gxQIdHXZLXxsRgGfrJnqfF5XkOvuk8ecf7ujPM39LMft
bSI1J7v1lQwp8MPg9dvuw0yYGfRMYeQUxV4/eA4xdMZ7fhackXAvN9pvxHRRYMwFitR1Il5n2n3l
Qpm9IJk+eoYVxDhK2jc44PqHcA+5L2nStrb/SoHdGDoaHc8A/UjBkOBTtF5EVReNl4ykStCHb9dd
ftkhotn/v7UtYqWmDHCA+MiWo5DMgywzDvuA1R8w2IBu3/qr86d/vbxrHdNRZE2wBeybAwL5o8F0
Rr4BqX7ynUB9UP9cPgzaS/nGduAnfbPgSa7v6QrO85x4134PN0e5vHlk5BDPS51taoJjEmwlBeJP
K134LJJ1yxaSYKgM/w0lypaIXW4PODYEQLieV3no3oUqNXkReqDqueHVCio1XZwkO7EB8bwjnfEY
sU0itN1vQGJqli4TiHqXp0BqnrefiADayvIkcJ33Qr4bSMC7U867AH2tHhVvTV+OpmG31moyutl0
kLgrQWu3z3vNgTF4YjtfkQf4b2JyZuh0tsRLtJzh+l+tQSH14bVoe599XO9UzWYbZK0ZEVxgOb3X
xlC7iDjf4ZbDOCdXS9ZWj32haGkfszWL/TN3CfilCMizhiJdMxZGRrlrnYdLZ7TvyLJ4EkVEmq8J
ijJHoHWUTJ0Z3qBeS/DKvUtM6J0dxTp4vAH/ZfMzqjLL0fwI4EmDxKwvWdX7X34OiukKbgUZpAZw
2EeWPxTqddvXzfVn4+vTLVf5zhG88fLvpHtUTZJii3UMU/DPc13Zfh5M+evE8pD58yLqFSqkfvsF
y6bDJXiL663XhgZNvTAYYfAUk+4NS7LDtrczLqVMQkM9Ey70qUucKLV9E9vDvaE6LkbjhKC0AVCk
x/Dei0Ld4i2D+xUQ6ee7B6FY643l9+KNV6ixYbDxXChqS2O3/N6krStehMJ9V0nsQyqv2qjOIcTl
W3J3nAgCW32ym9oDHtAyCWX13kok+GVNlEjQyP0EkGkRK/p6ugejgrlB/iqSkzPu9vBaMTkKkfwn
26NCMGG0CP+F+Uo23wI5Z8x6DoZzZ0E2QVVw7QAZ8y/hDS8ixqUlzE4CxbciBHpWFkV8ZoMk8AtX
3jwcYbIzaj4RKU0RhOeTK95rERBvd8QOxQTvxJafwOnPAwTm7qLqmBC9ddy5CCZo/Qn/A/2yalIC
mf4sz+K7NQmW+6SSepp1x3ZDdqo7Djh5UoUEPdlCH5I4jhv/7WU8vOUk95XoxLnI+gqmRZXJITLn
hlcBJyZjVZ1hq+tDFGZBSuee+cAqGngxFCXLw8grKvW2doBYCFaDObOnuSNHiygfHJyjPhRvK0sa
Xl8c8AN8MUgSfeA9j8OWfWgrnRbCr34h1kduQX2w+wse1mMGFsHJ+o1khaXavwuQgKdhp3oXkLf8
jq7+GnLH/pOU8T9wHkTqwpWmtTBi/3mWfKl+8TQZHCHrhM55+7ozZzGBzBpVNfL3I6Fircm97A9I
kJlFsm2TbhgJUs8fLTD8yTF0IJJnIb9SPrnpeRcQ6ul9aa8D5GE+f3pE4LqEUcliSpEqwa2MDGe2
cje37olor+r1STZBxfrVW499ujSZbOC0XGkRtdRayFnJqQU8tWTO0lJFSsxeBUcjk1jr30GvN1rb
G7mVPniyMYd98GNVNEtr34UjEM9aeNjZ8BcSUzZqfmUMLFySAfjaVHHcy2ojFxzTDUkK95aJ396y
CM+ZSAAR953B9U8DQBuzCbgHuF41EntioRFZCHcjpM3CfEuxeN2V/J1B/zZjN6QH+shR/j0i02Iw
GLJEl6drPTATw5ojHZT0ygDpHrew/1VCOKTWNyDU/3UQyoKj4clGgDtMusCaHZzvXmOhKoaforZw
0J21Qvp62genSi1kLAI05YWMDIhxbng74rQrjHVdECsVg5dtBLpmNOg1e8do+OjwCk7FaswRxgm0
N8RPzGqfh3scaPDub5lkYenjdlI+HyOmybZV6UDcCw9QR5sh+M2HrGbAsHE63rtCkOKVTQty8Ov+
FL/Y7dsfbiA88YhgID+asOk8kdOmVmNSlDrq+i6S9GcycJEvUp9rUE6yhygn24my9Kx/sNAH994t
URqfJxYKsxklVgqO352424mCVsMUtn+G0L0fsFqrqFmFKr96a1VGMJ6toaNaPRPoi+4e9Ak4B4Nd
Qnr4IVSvxJBbgMVttJZPttJVVeBeC+8PHzseaSxKkkL1WFwppZl2dYAGAxgYC+A4qQsFWxsSFDjq
XawmpDBpeSKOAYHPZyOv6nAhzB6BsKxbNLJck91znvPxmhkliI9z+tDp89d+E3bIU8+QM8woZ5Gy
jcc5s0uR0EpciMOpGnElVLt9AT5CEtpvEa3CxgiOQCyRYje7PFH0c8EP4TzWlepDbZ5zYKcS5Nqh
cchf4hGoKAABk4RBMJFGifUEpiSwMrWtw8pIzi38SH6IRv0KCd73OVluI72TCaw05BdQ03e5DkVZ
VjKaYXFYg4qT+R0KaNQBvodA2Kxa3478/cAErU5qesy/04sSSdvTEUpUCxE2m9YsmsgfoPW9ESMY
V8/PTMraVoTul17Fp8alOcZCFgrWhEgMQ6bYLFYLc8a3B/luFrRctVUQtdb07JOHgg8uGw3L+u02
cNDDyrNFVX1089tJTS3tmaQkmrUkhV9ZBkn1A/LnMjtH6lzptNxPTgpAD4yhjX3Cdi+KZViRDy0H
AVziZLlEp8oA5lET9oCnxd/E4wMSUTpOEEQhtJDoCmIFperx7Ot8o+19V7XVr7swNbonExJ5wrfX
qH9HEky/hMKRgvJawIheFxGuK1ySpLnSpnvToYiwv12sM812fP4L4FaYWTGOTUCP3bbFdJqybem5
tKV/ZaDRND0jT5pcFGNslwj4vzvv3j0ygWycFUaZSjyWzSSVX2rGTcBngzrJzxwkELMpDOpZgDJk
pYf4DlLA98mf6L655HoyBLItc+l2/2EP+k+WIPu5ycZCt+Hecc33KKQM54jw+f9Vu2FecfnSuJF/
cIL7ssm7jtaCE+UCTorIWwb6x7NwLtP1ricXMT2CiffRK4Zve7pK2R9CN9xTyOXx8NezgZ10Qk4d
H9vEbDiG6vdeClhRNCQdcFy3isO49ALZmB9A5Rv7oaJVbuJ+tzswqYKEvGeEZddnfVSqizoQ9g6/
VoROlu3H3NTGpOUh9RJI60VIdMv1i8ZCTsJNhvPur9042tCBDB4sQSIjBQdoD8adk4EorMqYbXRI
H720cqqshzhgiRDtpA6ODIX+CQisD0rMIHiVWOnW9JG6ty/ovk6LgRpUz0Qw4ElvdrhJeprExefM
hu0cCs5urQdw65nbHUnelrzGjec0px2gEW8n9Waf654tIZGpQMJP7/VYnLxfWDvio8bmQhXJX5gj
VgKoex0QjZI1tGtJJSyRUhoSmmSFY4kYRckkoZIwRlc3zuICGYtz0tJXOVWlqv1R+IQdmkJ8m6EG
idmoQLrYMmxkD51HaitgIzZh5WUR61hoUDXW3k9HH0mQ6ChspLzBU5p1i+/Gqf2ntdqZ/Ayl9PQB
zIwLRrqLl0wyLPaIBrHQUjsSd/buzqkiqomJALSdEqbz2NdNkTg8qVfgMm08UvbsitvwtOFfrVWw
hbKUQ/6KgoHRUoN3twSJm+8CaswMnqfkonXXmQDjhqfvvXCUGipLP1817Fm85LMbys2qfIzkojYF
JzYaytH3bGZ19X6P+xyoSx3PEHrfgTjs/EyuF8HQ0POecngHuG9D0bnWRtSBbUvmY1IdlG5DgeHc
JjEh8CHK3rFtF8eCko9N5Ux71DrMPn2fN3cAUIkm9z4FJfDC1kIOeyHo6FMqwas+/PlkENnrVNlu
oAF3QpBBFmU8+70r87rnOMD9yEXlNxQYnZR0pBNIvuMwEaAEYGF1cLcsvjJXOk88f+w33ZzOQkZ+
kzORcZaszB9N2nB9SS+Am0xrwzr6bVX6lYK5Iy1I5/9X+0AOtx3k+25FBNgO9MrtSUtIfIRimvB8
HgHZmK8qfu0GVk8MaMFWcM2tVJ5cHPVF7TmVg/32w9tI3d6RhPHoZ2h7BEcS642Lh1jAFobUNEDV
oltDEtxF9L2hEdcYc5gr09Z5YKWclGXAL0GRItvCpLOnSWp5OEmPEA+m40ObhuwbILW9OgIXyg9j
Y4KBzjwcGUQIec6ffVUc0tHSTNxztlOjp/ie1pXaNWQVmiHX+RQKWDQfgaQqL1jVlzkHEonhCuVZ
xBsrSSw//UcN+7F54VZw5Q++9FsT4zNa+4kP9X8O5weY/87omvEbEMVzyrt6PqivbHGzMcDxSXU+
NQIlZAiIY4Uo1qDfPE12T7AQC2v03REBRLpSiyINPitn/L5wJbqo6fQ7SYh2ndK128zIjJero/0i
c22ZMJxxPAzVrI+F6eCsb7ANPQyH39slpquPnOd6+eX6Jhc6k0/OYsAvz4B5lVE9BrbTySRJRuqt
hCnqKPDKXj2t1g35yuMnfQA4o5P9CKjzDaNTd5+mfapw2nQriFnGtMmaq8MS2CLpEXx5c+/zvwIp
6DR/Q4wJPF0pJiGR9L3NqfYCfZyr3jeXFGPSpzL8WbqHPp0+wL0B4utpWVmAfs/rdaGZOPUZsu0a
Q8ELZCEFQbL49lw2j84VRo8fY7MM45Ay7HV2dcT6D0rrFJYdYXSHOXVlSk6d5IDh4DR6xF1uWp20
pPzoImnsVlzNothXT4SNZ9panmu1Wyk7SivFlB6cLhhtM5LJt4VoDO9uxXMObEn1Li3vYOF7pfMa
YWggamGQWevCdWVTp7eULdtbyryY4G2p99iNKXC24+zyX884ePRl50KFTAsaqkL0Yd4gCXaAHFiZ
onYJB355e5eh7Z+qECqlg3uNWqrGpyHANjFX8mQGZ68CXaW9CeMigOQyDahyTQbmrfqBJslioEd2
3jukfrkz9CT3jThg1WPUEEdyJXWOq3XEbLZK8mjXw0vrP7qgk/rL5YRhasEwZ70/xmMzEAiAjdQF
Oqk/ZMJQstSJxPxHUDtMw3sxq+W6SrXoAdY22p/+uyEDf5B+l+gbQgf8jwj1lF8KRgf9V4MfHk9y
BGVMIVJaWtEQtBRp1/BudpGbaBXSmXIl9cgSCX/xHuaqvSlTUKQgtDMkaGW9sHFmoj9SpwNIQXKZ
2C4kzms9ZHozcm9TfO/sxwpzxTyUWFFqsjk12lmKrMLF6cF4nHr9EsD8EKxo/ah796AAMcB36fz1
rmCQGuO/RFfCkCQ/DObn0R7hXRF9XP1Pn4HBTneQgRsVwpXES/mrqoeLW2kdco3G/y+oSWm5QT98
jTHerFKmF0XPwWUEv2eti8dbJPUWWisK86XbEQiRgSFcREIPKlCO0jDJB6XmrkK2Uk/+Z5NfLlto
Zsve0ArZiQZLL6Klxo/Pd0UM7pdZt+9IUr+NSlY2YSLNLKo3DOpDMjN5wc/F6jFgKp1Rn6r/5xzr
YVo6S4nmGUGqxviCM08p/305OTjMT2iDq/8yBFwgf+xAcJ2WsrJ00GJx0IDdbKT56vbwU8ji76qG
E8yAn1VYt0YSaK9uxGhWkfUfzoBkg0PRr6U9KPdkRAgGFpE1s72qyEHhATupwDU6zwT/Fs1Z54i6
cq7uB3n2IZwJtMBVhq6KpRqVRljoJR6lHb2y9TQE3GnvXX+39iTh788OpyQeKK81fyBPItiFBVrT
X8Hp77ZGmueMHgQF3qE0rtcZNUg5nmNSzJE8hD3cMf/sKQZRzUvApxcAGPH0FP7N/FWLuYFP/ZFr
6ijLF90vimooe4ig291k2tkJWaXEFUpf74MZLb0t+OF9jAGXY4yeAAsYosLKirdRvRn9D/c7XlfA
McYvXn/zXdPAq4peCUadxtnRhjKRcg5f7KPuNleFPumD2QmiwaX8FCww1AzMY4cUiqkHiiaCKluV
vG1K/w7R0f6VxClYmmK/cBbbKxs9sJ25NStkIsTKb8GOdsX0By/xoDvjNLLcCNWxpePZNhTKAd93
+REmiQHRtepGrMRBhSXOd9kUdVQyys8hVMO876+NhORSb/92Xy1Mg/aRaQb+oCDi79ca162lCOvK
mWb2StwwMiU0wDL6NPBGbsJBcPDFaAdrfyc+6c+6Ycg0aylL01dfpSr/6vmCGfnzWqik1WiDj58H
XYO9ZGjPYXO45nV5j+mHdJ48W9OjsTPRh3c5jTafHC1BG0qrkJLh8vuLoos7QLOMC7L4KIVPK40i
Sn306HAxh7trn1FEtl68cFGOBVV8rI0QLoEPYZVqrlGmo+P7Xcvf23VL2S89bVUPeY1QRfKOA/gf
AY8yWAuK3AhjOM/QeLFo95WKhrHUOWWkRDQPrst27XCD7yf2bGKeq5vaZOHszEe1hHhiVoKUx9Gv
4wPA4hQ2gmghSuegk5a/cn6REugWKzQxk+K4jdcUuzR1rJzHMcSvC2BZl6QKr9MWldxrhp6tLLF5
f4VZoWLsYDsgHoRPjc1Q0sDUpNSRUT01akqvKeoZ5TliNcXQ46UFvH4Boqm6V2/LwuJywQ/9wV8P
r89oWGKG2H6oyh2Dn6AAGomShAyUC1b0XMGGZ2bCdq3rg+EHmA8ejzZYoDGMIRpLai8c4YgkCADK
ZocnTikYM+d8wvZ3EpXymnivkNvfRULXDpRZ4e2Nq1OP3kQmkyXjwRAMKCxAYiTyabHDLWZActJu
JtKY8k0xtxbio39tDn05wgBi+6aVgQpaA3wje9usAH+tAsoC1y/vOYH+SEZFOP4O39rBN4klrzDo
GOE4Bj1rrdPrXY6wkhfdA25Ar1Wxf5JbNFrAsj3sLDKxUdArW79AOPe16B3UIPdQDM10hjLmcVKJ
90Jx6SWS7q0oboRjXjsLF9+LKisK4z8Fo3rdpG1N8VN5HxGRlveCkTOfqPW1E8Lo/iVkjWvGSYCF
q+NRJ0rFTYl0jJLIBnskd9vpZjdYUV5YFCKQQr+HvLHSgJMO2LI3D+cNuBz/wtEhzlNKlDEHv+hf
rajfAkYzWqE88YILmXPVyDdwAJV4kI8h6sYTK2OiUR/hANIfhL6YSk7uUAHTcr+W3J23OCFNENuK
bDTh2a5qgJ9Z8fxs9Kbtb7NCwhV03KwRBb0SEMNPFV7mnvJxFer25M4YDiAcWgPIsfi3RBT8D0fO
TkA428oVi1LmVHcrPHu4HIMQDbliriIwaZ2lHxFUiBb7t9jwvxrEA2gUfU74wmhx6TjTyszasEmx
iSScTX8Ae29McP1t5PuOosJPn7VCV7IRyyTaQsxQz+e9xq5M3bS5/Wf6+s0CaROIiWsDK74hZpkE
+3JDEEo+i/73wS5Qc6Dz5RHVxFw7rnFDZDfWKv1TfIM5iGc8D3v+GUbKe3u0hoGyFYRsZEFRf8DZ
IwaC6VmpR7jdsd0eriEOOX6rhJr8bS+LR9NNHxs3FItd+TjeKnJuZWwBs0Rx2jyMrHrhAyr+VWDu
N0No2P0wKeZDIykOUQnPTQcnn5nqJBlo+J5b35pzuUo+W3E3oSQj5uONn65s1XCnwr3XGv2XV8Mr
zv8w3wj3WLopT2a5twIkYZSKqJBkWw1vAN4zYSPLHAe3cumsvYLiEyX9b0Z8dLIfaJi/dgpc+8jk
Mo+MhaTjxFopMQMJ1Hwcqt6ZixVbMNnTiwkE/oq3vHK8qczDtxwHpx9HO8ik3JRKiVUWsWfrQ8gQ
75ro8lEVsTOr56QSzKOzxmpitqfSprsE89n4sxMgarIFAAOZY9JOm3i4lLuRCjqjEiSmXGduZj/V
6rtOReoh8L52G9wRUYRfUoPQra/wfcV/VL4MScW6eYf/XELyPF9LHkDCxX2T/4hlVn2f1xKlVofv
Y+42EI2jxcB/IblXvYCbcSOqWNln2W76BDdiTkZ5nTiU3yn2DtuLUjhjKbNW5NgmKpYgdK7F41ch
GFZfYzl5ZfE3/XaCy/n50CcRmfku/jmGEnK9JLxfKdVDNss/+jn/bNHaXhXze1zddi3rm1CjEG6z
Q3TUusqArFh7vCg35dCFEQCFkDij+end313+CjRFxsDOCYXhz2AbeNWFWmSm/xRs2TMt+WBLLlig
GZELqQJajn/kFxBpYtCTF79j8TFztYd8hTzB0TsZZNIPgQTJvqlOgQw3VLeM0WSnKN/jjeHqZjdq
LAgEGKC2I7C9v/MLeYlWHQVh+rlew9j66m/KbZCEnRobXNdeXfAczIbTAL1gp+euSkTu2MlHJKLp
PB/anzKsqmCEMI9Tikfx2Wh8UHLPBfslcaMpMURaT1oi5P2cAkHhgdEHAQ+YzPYcR7ht6gB7tAQn
T5rkrIjxGSmy1KM25LH5MxROR8yjavDh4XepAYPLWVypKOM2NsKq6paXHRh4eqbtmhJz9SNz7ojL
FMOubXYCqdyCnIjnelizaRet0GXCCjgM+0r31xXjwRLbw/D3t5gFg6ZhW+M+Jqe5a2ZXN//fliym
RhLF+hWTN6xQ2HWhJhj8A3gGbTvvN+7Z8Pb7sIwiUEbSTnfKqK7GFRKHLGAZ+AMmm5tsR1ZtN1Ps
fxAYinpf4Xgzsdjp4JGR9Zqil/zPJLVG83akfPsK3qyv0auKg8nh6GPweBcZyyT9wBYJ8ozadYMh
ncHvxMQseidMySKv5bmAjR/RNA3CfpTNd9/zbYYOn0CyGICZEyBL5o00/89/Enh7UU3IBpSRHZBL
a/hKJom5yXnIlw+ytUq6bLL//B3skK1ZrvvD57B30Y7pZhoMXBOTwqvX4/xOZp1nYN+ZMdzXnMBS
4COYMIbVIsh+Cv/yCHVBB7TMRAK17G6YQ2diwvncycYvkg8cX338mPMwef1kD3jHaRUsxwAbwIli
U9ThmR1vKOaRGjs5Xqzz968o/zwnyiVznmKbo+TT523wHw2kpmItsR6Nr6AnisFVfbQ/gJkbJYwI
EBhdfek+Kz/5SH0J3Ipv4LQSBLHGwdSxXMgsvukwXBB7CvrfqLD9JaekYvYqDEnnsAiGGqm8zW52
y2QdA8N946kygOCbbVpjfxkKiRf72FFSUaw8tGquPryoTNQL1+dKAcjL+lq1wk68vMxe49FXmNbe
zREz/W0txa1g/EK9tJRR5rd6WeM/Uct8BTCOXTwvlLAr/d4DRQTHdvYeFlx+mfiR4FC3ehJdK1Ah
VzkKK6mVjMtrg9P+d8d+/6/PmyJ7CuqWfE4QCcb5OCKYuRCPs6PMuzL+lGZGkAZLz6ftaWNAZ4J+
/uZR8T9xu/VQuKWnf8BYlv2ZQNsCgXDhqbKbgijo4lw0hgEPqTaeyrm3LYwLmeAOt3KoDF27pNhS
3T0LnGzfGkzCYWyhRZlTzBm61Rf4x30TIyQNmR5YCrwT9qvm3k3drft0RuP+KZbmntkkDNzPpVST
+oSjg1ggTp71JMx8u7k8l+YqT1khdZzr+yTb3IqfWDDPgHa5ktxezfYu75wTK77kR1r3IUZQyz7G
wcC7PYR+Ly+Nj1L8TCAiCNS+lJ8ZSzuLEtjMGBy0cRJ3nVTepjaobvFdoXyTNuHs6xErZNC4Kt4k
hiUZB8qLdStcvYML6rT7Ttpc5NoHFKNqlHeRNl9Tx7ouUc6bmUfQpLyJ2jsB/mocYQvC3iKPJZcf
oyOeJQKt/tjP4klmesUZVxzxwq8Rj/lbgWnr3HOBmUNQ7Oo1cshk8E8AUthwZk7Z10/gYt6bFYGK
GGcFfQpoSd6dmFBuyHJmw6MwTAWc3co3mDq7KiavnYPmvcjXoWsW/wDExMZb2YzHzGh/cysnBWjm
YOGakXVb8UQCNpGJoBdqe3EPsryDXkqbpL0hmbBRft8vKihu7DXiV8YI3p4HMYixCFlW5YPm1E5G
tRGI2tcTwYVWALEnx/5+xrqUZWIilWsQHzQ7Fd+45uQeKouwXQA/HQyKno0gwo3GFEbZgQo1xTvl
FPqgOi781Rg1Y106QU0XpCX2Cf55ufcMYlarMkKq6v55wIm5x+GeC8Aox8swWd0Qeqlgtksme4Qx
P3Tl/WkZx0rCeOoF7KL18bmGk7CJUywJWSCO850Zy/NTeDQATVf6Z0LgjXc4vnEp11Cv2mP5M6Wb
q6wR0psrI2uiOHRwIdJxM2vWoA2nvf417iY0s3rK0FOW1D9HIP4DkDF8aacH9zcOFGKRw02A4rrT
R2vupFdIoxiNti6JHMDSHU6XUgGFHwKUWKm8d6+uUldEnG50kd1fdVL1UDODmWh/ooLxebKwCY66
ZsBoY2xrQW85vwmK4KbO/6ESogHmzF/p4PhB+3IiYFkwoCt4mYsxzcelZfL5E/m38rPDjdNyLzfs
3HgFDrUtZDbY4KTohTo75TqRaDI1XauzAIb5HR6TJyw2qD7xy/mZIUNFiMenedGrn3bllmtqA/pb
cdE56cWAqz2sYvzfHlh86o8cxDJ2SeRZYiOvzwc6VM8XNiwznInmKYIiJ8aWA2u5fzg56JfXMWi0
SgFVKMkye4vIzYH8nVAZiEpGZiLcQrHAfOSQsZHr6vZHWRYIdS8oFKen6LbZg5mLNTYd6Nw0EBws
drTsp4Q9JwLG+hiNijVCnkfKmyU0dz78YzbmDxEM3Eu0zcQPENQoY9YY5XWerisi1eCvvHKlhSvf
tk8X/zxFjtAtOdbn0PWmsC3Q66QHBZVLpWWYEm0o2Da5ZagOIZdFtojCfABDWjWdR4Yn6ofdEfc5
Tf2pY2X/kItcnM3+c4XHDKpWqkzyYp7439sBMeqwd8sM7FTIDuu7cDXVaPTip4rzk+28KrManCSl
foQvg2cPyLHmZPbwzEYcHcvKIahvh5aKxp6dgkY2d121IXOnke3Hj8lHMDg1+/TzYI3mk7Am1Ah9
QwIfTQ7fb+P7x8zrdMIqkvmGfNVfLCWkvFRcEBQ4zuEf0eIImq5ojXDrQZ+2cutEvkzv0r69/MvO
j9RBAtucK+qDSmBnCk6O1BMx5gZWTcBZIN57XE3tUgUE1UhnB3EBdKpjN0x2D4/F85SxONlKw0vF
3fAnSpXaMll1Ro6bq9gF8sUMlUoA7ZFLOTO3ATTf93EWIoXsZVJ17TM1XuQP3QqlZ+PCfaSBrLgV
LdlQCx918x68ruIy1JBDL5tX+9A6Hm4GRZg9NMAWRWyAgoPABZkKV+L/o8KDYBSiLrngS/I0IiT8
asy1StqevpHz8IA/z//sGwiKT+uEwA9nIAx3MrJdB4/VeGDPeA6CGCBxBi61ZNwPZS0PAQ6uIn+k
a76EpMr8raRoMxnSkrWkPuOUQx+jr4d3nx1OaQrRKebkpbnur2SEfeD1iPpWiFHCnG6qLzehGaAf
h7AOsQdxLOBMyGWIllPk/1h8IfH3gvWQE5sWXot0Alv2enPX4XBFEmpgc3V3TYpVPvc1aAUbxzA9
gE1DJqAexEBaWzBjouKeczWTGb18FWKCYVTznAJkfpP3dJagkK+Bb/H1VHZ3X0mtvG48sq+pWF4v
8JApyVWDB0fEAJjdF6u2KHcsvDNgbBn1xoWaQbkYjUTEt5oVlxD+utJ8ouWAThf8442M2CZBzKK5
uRi7K98B+elSPbK9IGMVXwPkYhkpNmUlkjoGyZREpOpm/kqqrv/9ES/cKDp9nhPt/z3Vz7aCysD9
VCmyNyp4N17dl+RH8yFuSMFbFB1iqJ1r5Y1qHUT0y2Zc+yOUhCh1njtcsu0aXIgsjJCFsn5GQTE8
kY//aQCV871OKESS4f/iqLyn15Krc81t59Im4nbroahNRvmFl26sl22xHb9oy9EaYTzv8Jg6TqLD
5SqoIxeGfClvlrda/CsvEK5hiG9I7RthsYpYH6lKhguY3JYpbxj2lxGLy4iAdHzALTrcArRryCHp
gJ145tpP9Zt30UKZXNa/unlc5+217Pkj9doctBJ7sm7/zUl4NFk8DV6xo8Lr6eaOyth2jsAXzasI
Iz6sGMl5sxUf9QMYwqeJKvfzXxw6AHCHtizQJkh9osfegn0a3uDyCo2sPv2lg8IY8xB6e6oGyGsG
SdWoET9bT+1uHtRHr1F1wVSI2dc+o2dYM98z2ubwysWjhP2vbVw5wqolvAXxiPZN4lCaAki0QNhb
X3SxMcprg7qY/VlBdYSy8tx87O6kPrkYUadNkUfnDn5rkXCM3LYtsKHD6sgZI8EppKFg2XBKpx9b
dCPQoTY0AAFG23T2i17g9KTPtWYBXqyTG4rRILyuY+ZAyQlkImV0g9GK0Z8L+GCOsorb7F+AKSrb
6LDUeFhIMmTCBGIURkVzfgXtOVvnys4+A+GuoDM6yC3pf0eMjhFZiE8P84asdY9CVU52ZRkzKOKC
UT5xyENKS1f2N1xCeX5pHr53Y5QUVXvttbMwvTj9YsB/w58U8vqGdVvRv++/yBC9D2s8P5YFxhzQ
IMDj8Q9rvY0xXRmJuZk2EixSPJtZe5JDu8UIWUWwcf1ebjPH7efQhJbxGbX6sGJLFxCb4ekWgufJ
x4qNxGo6ITOnF5d0t2Q59JEZv6KDECRER2BZ3vAY7TSfpFeSNyBTB8cw1kiuNag9YRvyXmiJqPad
Giu5qLFoJanEpA+oo7ZklZ3sH4/m9vQJ8Pia0zEpPORJMde1g+p4vv2ijAoLtwEHwBVxu3G7vw4X
svGGo8+fcLu/Z/1+shWAnG0QQts0189OsM0lJ7iaixGlhcQxu50uRBUntJfsi6oIFCOxBQLj5QeY
KjuyRI1d98AyLwWBsMp/bBItd/JGnXdYNjJvZwUVAjMEzeD5dOuIBbxCbhxrCRvbpEpUusaFd9NJ
quKIvr6T6SVd1b5vEN9/8iHcPzC31Lvwv3DJ0qVJYl/v/xyK/vPhNvuUZPakfD/4eYxSzpR8DJTI
VbZsD7uk+Pb//ot9KjjnviMtdCoafNHSfVeRf35J5QYR8bgBqp+KNCJWZfJ0dKAqGkFwmqGWNR++
4NiPkXD26JNHKC8FBaYoTB86STGSggLQew9nz4eeFXPF2jUnjYHpDuk483RNRTQqFb4gPN6U/lgC
MqgBZ2l8HzxN7+i97VEdAqyhsk8KuG966YI7uTuFakSgAgXqXshW7xLhP0qNfGSe3LdXb6/XF8MP
zK8Zysu8EqOn4h5z3WzR9hHs3AWQu4tHE+7uIicCuwRSYCUXPorK8ykjSNB+SmkFIQD8qXOBfoi/
WwRy64NWunUq0whL3qzh5gwN1EuMY27/LFBl7S4fpC3VZQCK5O1cEQRks72KkbWRJvdnrBZHDWo7
jHN8TFBQ4slQvGoA6fDfcKNPj2YQEp1doyYMaKeROouADQwRC0b8OEiZFcbTpf6KVN+tC92HBNeO
W9CvOXNkfEVLJsAxms2HrCNB4YjN81rfxivDqmdtcR5b50pM+W2lu+WQ+ytvCXzFolDPacUn74TS
3rMgXqa7BN5ofhUxGbI8q+CGscTp1r5QWR24eRPxMXNPlPRLEX6LJFmMxqnRbiTJZC9zAA6/iMO0
oCx+Rkzt1SsPKrmu9UEoI330cNdr1aFe4E8MJZBWmIbgL+qlYjCy0FB6mN2m8sGux3BC1f677LEF
8Yq8o7I7BUz6RV1Li8l1sSW/m7LPJCpTJLFUBh5sV9nnxp5l/jt4rG9S8zqTs/JreNQRNg7PgrDB
ZdIaoti0ANNvesDAHYPaKsloid0tTiGjl+l4iq4u8O/alh8JJw74Uei/4Kr31kGEKD2GUyzoOIGP
mghfkQE3pDet6gFHsOEPDgSkYCLwr90UwsFsfXR6uekBt8ainnMHDUBl0DBOmPw4YneAwYZilZ57
BmD19ZFeOqWgCcUo6/uf2eKtxMe7w12oRpaX0+ImLml54Ds4hjXFJ+v1VtwtRCcAJN6aoQYaJRxZ
jYwN7zcpmgew0laOVgLJqwqq8mq9BxiCR+Tqv2WYcK/548ngiRg5rbRmrVeWN06pCQSmJpshL4Xo
uoRflSwjMk7ZbAnHoxrpX+e0qR0h5g0mEwRJ69gRHhQpEeQtU1WMPg0TzYf9LTP5CdwTUvWnZd8W
sE32CM72ifMZCbJ+vaBVVZu9/oKUZ0RjE9MwQoLYPaLtzQhE6uPrxSiCw9923uH0HjX5wyLhhouN
g7F/GNWTJAKm2guaHH9Aue8Wb6kJn3iAK8kSntQPQIvm5Jk4HpBsjjeT1qZGmjztFbLOcalaqhXQ
D2GswoX3mkmxE/JDp5H//3VZDSMSJ7o2Q8nTwOOohY5TicdDPhMkvkuEJwAeTI4lT6zsJ98G+fLq
C0E7tFoFjdLiPnVYz0Nc7z37aJ8l4ytLlnjL/HqkUIhmaPy/rwTMEVg1yx12qGdt8SDy76qJ/2C+
NHDuiSZPV0B32ze0FM1PMLRwoC09NdMsrGo0ZzuVbt0Fvd1otdgOFcYMFWtS6WGcay6asAypSHhC
XjD7eQp2MdPJ4X5XZU5DfBQMxQeDdaC6WF5DnLdBdXSnXrWUYk2og6YpoHVLWXHyqOcqT5uqN95K
6QZREDmv0ro5TZwi2z9ISvr5aWxHo2zb9LMyWcbeaAv6A8QlLDGpURxLdnMp+btWYkRr/yPyptL7
QiIlWCQ5eujIbCMP+MfKbWaSioM7LSbsDK6m3t+wBcfTAwho04u80mBuyQQM4O5ic1/T696C2xKk
if/7BaDOb0qFEhUulO6elDyWf+G5Nt3gKcxrdqGJgmy9y3MKftPBZLSmavxkNkDwCd5lSNCQZU37
jKxzaeCp7+yOH3+8Ic3QO1ymvWMDSIw1IbrLQYMZUHrcwGkawmBsZaJ8ljlIIWP5F+eVN+7dktep
D0B31pEjKde38PPSAu8FXtc1PErcqnnrIoF9h3qJugp3qiW4cnWxNrR90EROm4Y48EnaoGTuQfpv
35Yi2twdNVqzSxYcmM75N4SrNyOBY8vq2CcQaYufcFMOWXkC3xF+AbWrj6bnsY3PYtAiyokFE5QZ
BGx5OIRpjPC8MhFt/2tc21/OtKamxycPuzYzb0wHD3UvUUyk5lXxRZ1LyYTEM9f+EKoO20o5RSnz
vHgNWETZvBwGUUouzKw9S3xsMAkewADBkBR9jey8s737zghQWspOYyIfOXO6m9IihQDw+GpE2iMh
eN9mFa07WWIyQLY5kPIOm8OCMc8FvLUaVULNiDTAcytyWUA+EyUzuJg53BsvUxOQhWtf+mSWyOJC
rmC9Ewnp9QCwbIIOCxF62pgx0Btg7vkqwmDBAuVSPae8euGOaE2ZQkT+VWSLbH8je5qhurq7U8dz
mfo0w4+cp68MjqCJ4FtuYXu3fxWpL4i1g7c7qDFmabLO+Z5B85XVXA/dQtp7YR1PWZGG3DexUfK2
4s00ZvcR+b9Ul9oc2PtzOvM08YveMdkfIF450M3s58nnybxE3uLDLwdHjlFL/bl1wAV8T0HB7bn0
rhCK7E4hVcUg4OSs0zSuNsCZ0nMydp5mWEBprCxeDP3zmDdCKUgdmgLodfe5XnhvOHY95KPJcr3A
8ZIU9qANDgnUhyxl9Di00oZL20BYulRTk/LFV6GBSgis8janxtP75RNbN0mj29W6D/xtByaHVFwT
Wti+C9ZF15xK+v8tOtOVx9i2dWVrMwSBciLY0AiehDfb2B3Vo48VbEiJf9s6BHV4A80Ky0SRfda9
lItx0eX4ITTCbLHkdDcOOZJlNhNzePbgyrCJw9b8cuMXkFeCr66dI4tUSjeDNd4SSxDDMP/658ID
XzExufg/rsuErHXbWk1GUwcIpQXGNMH/C3I3ESTShA3Itp5qdvfdFPdgcf3z1bUWIt0xC0/m0uNY
S7saF0cBBULH9/xtVAmG3kXw/dIjOKfg3c0iL6ghvUR3Vud6ANuifyyU2vmIXMyu1c0R/h6HUxqS
PNIF4pNUJV5Bj73Gl9biV9liW1Jueub513jL2SdFNIyHDYQKbbMnwz2GZSiymB7RnwAs5SpPXNCA
0DbZRS/8+1oM4Xtojv4BzbdBXyYiv2nOnW/8CPw0xBrE7ziwCliEozH/QeM0umIGiT5gMvulZ05C
yzGwQoo2xZDmDn1kiqAm59xOHxMd/kgmr7EVBLkDYi4Elhzvet7tg9U9ZZKrxk3O63GqUNX7GkVA
haAEH+wvG0oB2ffWqFUF5GQV1AuU01Ku3/9LqoqyZ1NCXysPt0b3/eb3qCTFNHur1LVdl4NiLo+k
agD1kzZhOYj5LLdx/wZgERdSoSUQVeyDVBQa17c7CY+RjJLQkhe4WxJOCjjaDMfDXqBbKFufzSE+
QkUtqa4ILriVq4I0gCEMCmKXynellwtB9McbAtl2C3XkIQWFdzyVUpmKn0o1GR/66bUs5qeZ3EVS
EZr5fiy0VgTC5pnNQ+DW0vq7EzAXamczW8YprpT1Iy7zuwXwyyfymZNfhEFjgDU9Rs8PP5FSyPO4
pEg7n7kEJioUmX+ntTL5bE7ngXlR9UUpb3YXNdCCRiFGVawJJMYcG4SVy1/Rgy67KwdOfpapa2+F
OmYGuHz7bfyQufBk3ed7oOMSpCsyYy1j3hDWvQE9AdNMkrjybS5LTcfXX59pTtJsRI3GIcSXEwhV
k58muatzFTMSI9PBzBffKgKZLfLj3sO6t2bV2JutL/AC5KkA2tYTV6dz7eoyhBLw0VEB9RWh00Y7
kawWW7RbqdbXvBrOiOEL8G67Zj/bMii3YN6e6Lak/ptB1YNsOaYLjBO39CmATXs0MjvupeS7n5nr
i1mO0/8NCGrsnB72sazy2XexwTx2XUI5+VoY8H8V6t/loWgFQQnnUiHN3RBs0AoojclE0AZS1UQ3
YI9cYKHw795uVaFBwUmy1h7xZu/QLwjWmH/VSw38tPHQD+8GXlxta9hGgQgjLkl4WrtBZGazLqT2
1zhQ6PU55H4D6L8JfTnkPZKufKfFkueg99xaqJF8AzYS5MhulFkhsPABTHHkb2SiO8vhxSKMkDKR
+j2rfwCRj/dBjTwMRoYd5ilDZQvDmjYSQABs4zLJZ57Mjb/HtOZYAwH7HsQSZssX25wfJ7Ex1tU0
61DCrTqXJEKMA8aL7VJ244WazvTgRsLNaxhrt66Cr/Cqz7Qfeciu6pOhoJypBQy2vBRTtBMeu9Mo
WIAtXWS7tZ4mCA1W+LLFAzml/DG6rPiNkvkaYibHLedVRsIXIVOC00OdI0tNvYwedm5oFmXxkzDH
uIpRDXNGtHTynHyg85R3LnN4YMJmPbY5R8TIuB/2PJQsgZwI4mqkKFJyX1P3msauC3tvoHcSXRKb
5T0xLsjsW35ibYwIMK4ENof06YQb2tvy9hB4ecxiPjEASlHLMCoRhFOM8w5J0yYBXcuSFKwh2bpQ
YvUBQ/oLRgdCAjx706hHc/iBRJ9nPbumL9Ncpbo5gcUF/036jxyepCgNfdcq0q549RBUFyZq4zCS
pB4Um+wNtMGrCIli/Jaxc1QwydS/72JU1SDty6zwKvOACuCb3O0ImJ+HA2aBC+CdHX8nINOeODnc
9EqSK669O70yTDWYk9a3PUm2C0lulWU41Fp6T4NkK9bpAc7lwB8SdOq5qzR6VW5eqtVPYq1AGLmX
dJ0xfl2fUS/e4Geu0MhhLgRgZN5VFsY3G+LlPAh1C5nJGK2SkDVONL5QY54XChzr6EBwoE+svnWC
SC+0LXwqDVL7zIlqd2y2toXbLR5I6NnwrXmCsT74y/5zRM2u/KLP8m/gdG760E0h9Z7vKYbcgz5A
hupyqB25Cw5NUTd0VoRtbgAQyXEn98xuXzxt206JylejEEXxJPOsQzxfvZJEm7gm3d58gPaIC9SB
pT8nnjwfazJWfYulvTCbnKBL8JSj3x5Ow08nafg54Zr3C4xbKEho+IvHEYmTHD7A9AkRidzR7/4l
u1KTHmSbYGDRX6Lq6Oi+7WozO19jHd9NPUKcS5eJIMjw3AWZgZgIOoSnI3bzCuNffkfSmtzPJgEs
DyBhQjGZnGqAJMKX3ImhSJWmaUvHgalAEw2UX7jeNBWEfBtBh33GntiPfOZjGEFtmIpYXig0NOGT
Cono65K1iVSsGgv3Y+wPtj6/P/tk5YglW3tzu5QrACuU9ZLjjP9GttXGQzlJucRpLl3vIgisVApd
Ln+V+sVXYRgtRrbJP3+NkK+GGr3jFzNMH8Wy0Qw0OuWYp2HRfuT2cHsOqfu6U0LoL3P/zHkOeXYm
+1LkcGDYfq8+Do/oqANkubHM0tQpRcAFHI05r3jMDHAC2e+RuaCsIyxoGwInMOEDNHmvzZUa4pPP
Xz2+VzJGxnjMQ+TnL70CQrXFYECSQxlAZD56tR+4+BvsuSm6G58MwCRPJhwZhJPwRMLAYq+CnHFy
dZH3TVL1+e6odyXBNZcgKraE1qn3WDPkYPqfA/0OTSJnpDe/K7ALZDKsxAqRbh41Vb6xGvRJKYud
mU9Yijkg40wgHSby+dzni6ywo9RVb3vxq9uAb2OnTquk6T9//HTtlT3YZTP54Q5rEzF8ihHCHa3v
miK2kNbyTKjAR7J8PbXfMxOcZuhri2/R1crebLAhv5JEwYXOUL1sr6lSatqY4IVm2vJCse3IbBso
7KG6Gi3MWZgjMIBCptGFhxq3cchlPhZkk1e1RhrlFZxt8wwelC5HmJEcffYB3YlRHzLeQuG7SCA+
Y7egkEo20eZbKDHZGjZb5ojk8kLyYmDFSLvmaUyDi9KQYoMjWRfHZf4viThwJop5YrLtZ84TUtmA
MqXW5uyNguCeYZejftvvAN3u2Pxnk1itJAqER+zHjYtgkXMwWtXaT+4kUxARSDVplSF/OLYrKv61
LrBAb4AM/nu9yS+i0ufq3FD6qHuSZ7DmUSNyMqSbcBAXEiprQPFgK+QfPz9FLR4xU/HXPy3o5C1U
EpGslLq1IWEUkL9zYb5TLDBFGFe0Pj6rRWQLTuL9z5TYQnrsVT+103n5p8tFCVCO9hpoymrrz4+o
3Qa7H4BmChbgLKr5nC+m09FXKwSEdTxQAX2OUEHewestNtL0xypCi6fYLm2rneR27u/yKPzHSYBK
z3Du/KNDhmxnYaOqi2gAcNoZIWiFurf3u7FMdN7yZcrl3Com6Bk878k4GZu90idLHuDyKvJ/Xq/f
bnUUil+Hkuvb4SpBI7YOQG2B5T4cqj/YHwRWChZrPsZgkKwG3OVwtWuG+7t/EQdxD0f05Ez22/fe
6zsukW4F0QfgWBaD3+D9Q59RcABvgdZ9GcWmWIIQDewCtEHaXqXeXWX/khvJngz1j76LovGWzFgi
VHbHXnDuv9GDlJQHwoM9bhaegVBjEnFzLEjficeFLNnQk6i2pscAIGT/pA/OmAYJ2xAB/1/eLPxi
I1p2dPuXObkD9Tq4JGsQSCWnEYBiJO39T7FfLmFfBg9h8OyJaI4W4hT6mlDHoYsWhSGQ8Gwm3UQO
g1McsUC7Jw3/zxoLomRh409pCoRIbLxsSevc9qR0HO02CVVjOsXU9IMYRvvu5RT2fyv4lH4OfuV4
l3j/YpLtVhTRuKmpB5toRLCbc8sc8VmrOhm6rmyXGiAsfqVoS7WmQAA7Z6SNNQhsvkS8E6ZwE9RE
9ooTGmh7QcZZ/yt0m5mVfD5WvVR2CXsAQ/WpmQlYOpD0e4CwSkeGNVGO1SdbY9XeR92eGx/spmqE
ZH7JQnQF6RTWHlUex8xcaANjZnxcgm+7FUXrQ2houHx7Qjxm3H54DpEuWT8K+ALTZKBiTXF6IzOb
X6vHoITpn0RpJBM0VskHERc1XqjErwyxmn7r9Qtrb9GPMzN9Y/e/a6fQyz/+S8HfFiYLvdWDdXwS
fCjTpgw7dQwAVHM05TCQvQ5Qfo1sOc7SJ5+NRf+VUPSAY1VKoNqqLja8UehjBc2+GAxL9XDB4lcq
Nk6M+8NHim8skV1v/LVG1BpI4Pb4ozKLaqRh80Yf7OoJ98FBRjAAv8AOgguhCwDaH28Xc0GN5AzZ
90vV5G2KNkaYHQIu5qBnpD3YJnBukZMQw4zUd4V6vCxszgKJkmbNPKBpMM/02FZoFM7bZlOABvbY
feRRiAkhb6VSrDoFOmy+sNBxuHULipj0lI6wSYbTW12djObrgQHH+8Z45PqWK2Ef3LRdrYsRqznW
UqV6DCepR20kbnZ8zTwhVXyEI3QNJlM+6Dqnz4hF9dLlVtS0sgEPCQQpYrgfD5PH79DQ6UxqyIg3
GDcsQDOn278CjkKIRrQ3CfPQ8xVptY/RMad1o7aiUQAuzZpeGSfSBISanHJgdsvAf4O+NPSG5svR
nRUWsHQldKD/iHqifFCJBjGk8EtEoaLQU/PIUwiAwjgFWZXqpLhVJsWjZQ6STdZ52PUFWlZZNlQz
l0UmubOJZKI0NB1tWK5xd5yS72hDNtnNycAAA1rPQ/3tW3sN30RxL7xWSepFwLP+WQKCKFSX6rra
ENwo/yPA/9GGaC3MafW3I01AD0xwxTgHdCsyxfpd4XGEOJRzJBUdAuwZ6suoFFmRK4e3j+tSdAzu
Ko+Hrmjf4WO/T8QmY2isPHRoUYFJWaYOnFwR2ngAxHQLy5fawOtJcslcUhIXPR77qzVWpFeARk/j
ke+fFGnhS59/ei/bF4FzzgabW2ibdyikYOrM0WFk8u9NDEFbdZWMomHdtRdi2rqIGetne9/gbIlP
W5y9PlOy0pS5Ypxre/Bt3Ll0+oIRz1bKpGB77brIwXgsbj6Rm+rXYvEk0+Nucp7oszfJZyLVYZVM
OoxM0B73t1CvShnZZuyJxbKnfg95K05rBZCk2bLHCQv2QwOaSrDCKOHKU4ce+GAoaifInsfc0I/j
YLP/ckrxtvRA4I08hCzvb8/SrkiLp/VoaLtDexroZNQ/nrGypKMa0+IZ1Q+GDue/avn7lvWHkQol
+FUXXZ9mijk9bCpIKGZj442B/sX1dVURt1HIG8l4oAWy2vWrtZLwc1tAnXr9mAhaqyUmdyYa+uN5
t8RjOYyryg1JItYdZ8nyDqCr01OR/0CjUUogloply3df53CF3WLyVaNTsy82pcvWgScxFn945HDb
t5PlIisWia4vyVhCY6usaMpj4ujRQpB2hHPrdRoYG/2ndZBoZiLBlBM7w7g40Let2xVxTPIvILpg
ENLurRpUcoJCxwLyOZj9dGAV0IsaNoh7eob+VWOXa9AEhfsUGOJUEHbP0TRnzoWc8xaXaq7itrLQ
seEIy741CvQYI2Y+c6xFObHbAidbayFtQ9RTWUqFVbH/7TVnbAv/B1CWHPLIAOgyf1XFv7AJ99hT
1KfvaOY5ACZ45UyBrR4S61g8Jc4Pp+g57L5H8Br/6dOu2LEvDWaHlAXXiBfv2DHwDOe2YIJ86I1a
k1fZeP8efmUoJ1DEHCAAY6s0YyWNgoz7NhkC7oTHx+jwPadoe3qB+kgYzenIO8AGcApgNibdDpyC
K/Z8+TCAwMAO/EgzjCE14y1FX8Snj0ANjtq1JmMsGut5UXXqlb0pJe/8IMhrn711VMZwDVbWH0LI
dMSgNe4gBgateQJTCdV6dfMFiWBPqJ+2XZE3z/mEkGTs0TQ8Tr5+kVwaQxS6vQFq/iOYH8Gq+APL
yIb4eaMPjuN/JAHStkVzZYvnxnlflbC89Vft5/X5+Xgoe7JSo+eg2mngGGTdRiOV744ObKGz+Of0
3qJBAzPSqQdjeIiu1wLsI8KO+DsQmItat0OIXdc/H1otKKeITnqeycrZR845iA8FIB0FuexRT+rZ
lJlGarW5NEBx5vnuxLUtX94yptzr4BaEXJp0eEJuPSQ7+vmKXhYyU9mYRRs5yyx6M6Vg2L1Qptic
jTpmSTI+15xVKEWfZfB+HjMH0ruUNQkRlW5nc+nT74iKBw8n+EcPpRqdhDwYRx9O2lAlWqII4AbD
e8Q4mlSMm6MzoqhPXvrjLA/Rbn7hP4TyPcUtCuKOCpSsNqmFfT+xw+EZ9AxppEAkF0fdSvK0P+P4
7mN1aizFHC+cnlB6KbkFOyYcR/NdASGGBwTjw/HsAVDo2KhbU+as4YnuV7kuixV5CfmMULfwYdcZ
Qh5qUGp/Ft430hwctTX6gLAn4Abqo71NXw4S3mSHgdZFJH4a99RA5gYqu3loplvF3FuLMOCVRuH+
gNi27w+/vkMjO6zFB7Z0uplTCbOR3KuDThPq7agbBFwVviGBftuGPs48eO3apoux3wUsusJpUC/Y
YxcuOIXwfjB7lAeSiQ1VjeynkTf3GqMdJ1dWe7h4H90IR2qnBXxvIQdl5pBbc9rgeGF/e6i9fzph
ibZbH204Vsl8V59P1FnRO26284VKOrgfqS+Rl16uwJuvZXknFt+RJYeCRHt4HUApKsTUOB8NTowI
DxhRA3zuUrVggCvJHfWnCMA3fSBIJ2YXS0AL4seCD97TsXmSjoblP/SBHAipxgcyMCdMGUPVXBsi
CG7hx+waYcFQvsgY6mTFd2OGPtsBgq5BpuXnHLHTwbtjlo/PIa766crkM2amcq6N+1axPHcoJG/p
FRPRhfjoZOTAF6DGLTlLhmJwO+TAyl3Og+w0VykAUHbzAsMde8AvjdXw1PSBWk8njL7iTDzc2dMi
LGkyIAyKA4fXWHdfLoENpXlKB42G1EsuJOu6BLtEQeq29s7gR3ZJu4yDlgk1hW7tlLoCxK6M/4bH
2eXtg1SFsvOd8DsaAwhYOuK46Vn2jGocvFrNjIH56aMciTo/heGky97Mkuu1H7Y7V2VnFeyMmz9r
mTTWLDvphvqWKb20EVYRb8B96dahrlOv9DbCDipzJMC71aWp+EKnYJYqk5r9lMRpoWie6xGr9Pbk
8cxinaDgmXO/pJpf47qlymqWjS5tzcu1L3BHEEsXYB359CgQ9o+rVhgfb7yD8WUoExUGtmO52/FQ
nb/Mi7i0Vp7BH9feNG4YopzgSm74T58lNf1D/nO8B35U9UXsZiUaEarcWZiudnrt8Mjr8qLy7Mlm
gmNBpEN+ORa589iQwHA21kvLQtTNEtvHhvhn6dMdv07kK6kcYoPyFEBsEna0CcVD/ChbOzU18Bip
W2JWGlb4tan4ZIzkBsvuGYT5L0QM8V2SWyLYlRR7V88wyjESav4j0ttFd52X2UO0PuTBhMdxLdew
KJtzsfObazFscObyBDbHarcRLyJzlX5yMYyTDD9GXmoOFRvFIb8lUcEl+EAS5V4sN6zJBRJJxy0F
JFPUny9ZW22tag7NfIYfby8/4WPVFW3urab2VQx+yRiAJJ3j480jmDsij4/8LmpQTC8njyUpQj6C
G9uE9FTzry8TWYl8fqlvI6K37fkeJPhpsXGW/Y7A9tlml1SiiDkgK8sbLFt1uKLgpuoGQ5hvl/8+
TxX2S2DzNPeHqF+eRZxEwTiBoGuH6Di+iytHCK/sIEkN8R22jS6easjaQTAAoGz0A431TFY4JFK2
/4Ck7+AvISjEABjzGaPntjDcg35SqXX04YshGzJHZNR1qdRVM2wdKJma+iRDEJj7BVEwEMRqSQEm
SkUrQYM+1c3P+sGzCR+MOEMZ65jptYXlHZ/Ws/DmmQnvt9/06KppQjsrrQPT0v4vLMB2BQRxxfIx
k1jew1X/rkE5xMwlSL1hW9uCOJ1JUxDRmGBm0SNOBF1uZdLknx4BxTunFPg2orfKVxiXKwcMFETe
/VdXNU8LvrTArpttZ1wOUbl1Lybj2A47g4mC6ZTJmLlFuR9L62h/LULELR/dlnbbUFfu+ymcXLA6
AXvGf04+bUL4v9SIe4EYXxvtVnRy3UuWgkYPiYR/glhVAk3UY4+1tQCS3XJ4CM1q3SjidddduJNA
3PUPKOsE2QXfKLKjzI56zUOoMSCJmDIChCRyK5B3zJGj+MglvtqczwN229Nqh91G5zQ3tJ5q8yOh
IE6FV9aCXeHj1dL6qjnlPsDRwPWs2MaRecFMz50/w4OyCrQSKRcagl49XUJmK4TBDrxYPZm7zE8+
mHxr3dS949Watgu5RUcNf9tpq13tfq07yXSQANmgjy8HSPeYGTZUOY06eBKQiORChPy4SmTktzr4
/ys5Hxi5vJiQAyTKytcLY6qetJjZ/yoZ8/lZNagjr5IoN3Ht+WhrHqPIV4//grwHQotrQAiNvcnS
IZpD11ZH2Nt9q/WvfuMC8N8RexEdoyvx+QcvQAEWmEBQRCFXKmIDErJuxoAUq29uB2Bw11UR390s
QTwCKT65SZ9N79VnornYceCA5/sg7My+rZ9TUkzK2+SGgVxavImjpEhDTXrgmhI4wH2ubxEOTInb
yxXby2YVt4Ne82dgMhdar9tue00fc36f/Pc75yaSCwyBIV9yCic0Gy+LKVDKuajgpNLqI0ttlNG/
QLboQlxrRqn1H2lS4n1e5SH2AjZj/SySmTfh7W0N9qWkRk2cfCc+xgFEPC5ghixINsa3W8AdxWSm
uuFmWC+NrdrKRyMd/JwkYezIbe210O8inKFPLg7d+Qfs6t7B8a5ig2Ome5AA+O92GIEX4RWdd7q1
OL0NsGi9DBL6LQshTBOMRe6QIKfk6PvCf+aLGhCOXath7QtORK31wuRodeDxQM59VoQ97ex1wQT3
7b1zB8+xJf+rTs/gR6WkI88bZxehRuZbV7WDTeZ8bePgNOBTzRd5CTghMGW/eCcgdKMgEb3UV8oV
pqNZPJJ8DPk02jui6oPZhA2PnVpVJI7Td6ACaxWxBOlPbAOYh/Mo9aS84Gqo90xg8f0tWz0A/PTW
XOgQfSDlfuhpo0mWzYWDYLHeaVLaNKfDsCvUZvzO1xti0hKyqhWAyT0sZMi2TfpT4Rj5zhcjcc8r
tDCMs2ZtRNNsRUEXnHjrtlGkqJUB8I7W1onhL3hsJQLwlLZf+xo/VU4Gym1VewPzxhAULsSlBHrl
K3bgN8dp0nSAejl0v6tUjsULRqGcqG+ZbNJpnID51MkaBgS35JIMRGghjkjypf0SRkYZ+oWjzoyx
S2q32GIEjEPpJm2nzCg7D8STD1erDZcT323ckizmN1ms8F4qmCGRMzTBS7T3rRZUiCxE01aGF/ON
s9K32mtV13PrJR5wnl/+sd4nA9adeFctYpIKCXmsxLiRWJUpeZZDc83n97HovKuiEbs1sgaHzpRd
054J52dtTDU29DZ5TYatI676weX8ix3y+Xy7YgEU7ehwNv9oHgHtLzGBceLU+HUT0gZi2rsxPZEZ
SbrAppxxHFrMwuYXofKf6GswqejxnljFnfkklUA8HNP+0miloLILpWR621d44SUQEEWBCqcKe+3G
zf4S0sijgkE9xWkJj/LtQsZGL81IcgdcZVwSlxMAlTgKnWC1lZp6tzSObiktLmyGZLVOIrqSf5/X
w3KiefGpNfUFRuK8VKQIXqbKtbFsK3FQQqrThV+m6A6vWtxOcuPTIZojb769D4FVT5+youwzDpQV
FDQJur2UHS5/FPi4CPPa+FCbZOxZD8yq77/YysFQGyAEbgbI1tt22S1lF6ZBY1jLd7pEEBeV0MIW
Xc0BI1ZmT6No4Xa2Wy6IINNyS3RbCglpqDKye8E6uXS3q+y6FfL4EA5RQW6pleuCSRC8/z53Atid
LWbGWXwW2ASn2n7nX97fGdTURLEZZgfit7PIwAaHGuU9MFfWP3D+dx/0r0jGMgSs1Czns9lmbQJR
zx6gLbGBQH6/Fxz9FAmZaZ3z2jXBcJ3NB8ez4xeAIsaKGAu7jjfMJzJ/TZ2CLm50apDu64/bqXLp
+nRyDKAF+Ce+hkgXySeBOR5NdF5trxZ6jpLYabadS+PIWGHvnpOruiIxJolWSn54S5kmQZEL3S2c
XxujMDHnvpk8oxkBaoXVqP1vQlbYRcT4+IO899vSQLBRW9G2Fe5DGpQILW17zC3kryHWeo9IbRWh
lMogmvFch752NswMUQrcOs4C1eDEaGjpX6VjXz/WjfEreLG/DdZu/Ba2qyURngV9m5ZVx/cpiyia
6IXNbRHGP0TmT3BqBx/lymdaNA428QlDFfv1YSrcTxcjonlc0LN3f8CJsUkcj1qgJTlb9K79lV9v
ByGzfe2kYZfMu0UvV214On6ObsLUwEk0Y6qf/Q7wQTwafV/fCT4IRTQR2welNcXzuDTYK2Owr5vs
6zoF47Lqu6ETtXhCcko0Qp5xei+0cX+P/zYG6vIigF2XbqajBefbWyJm6kQBUBsNBG1HruHhvETT
9RCeb/sj2URM/v0Xar4meR/NK7sgblZwbnNBY+EcZ9BZZuzK1iDxG4goL6W2U8ZIuFbxX1XPjq8o
rLLdBBpvf2boAcBZ7JKo1W87b/pIekSH2QENwXwM0FN1i/360xDFx25/FVG8VN64vnOymttOAvzR
FoV9IOYPUgUiMGI8uxv5bYVPptSIttxCW9Oka/bZjCWzAQu/0v9Csb7bkbtln+4coSpQWm3Tzfez
FBKrUJsPWrexMLkrsqdyFcK4TXxIQXPSOM7Cq8iUP1sDS4qmwW5dk5RfbaqM5pmZcElnKoAP5fKi
lTSWkDqXflNxxig3AsNCQ1bt5P3EhLkS8fMzlhHTKbrFBK9EeCljfv6tY1KJ11i71aF50sU9OgzM
aAJLQHbq8FKXbmtSSj8kTu+AsezLpv54duaLOpUzorFeC3wsxm1WVvq+Xvd7KIE32NmCLIvV9RAJ
2183+gjl4LQZwjpIVQS05fp9jtItiGwUSSWGR6aLCouOGEz7Fs5f4xoNbjigX9R6GEuZLOK68Evf
DAm5+QbdhcudsV4Bm7/gBwpQXHydosbpFekgSfyWcYVvDcJhcsXadudlBRJqc5vjq4dwdHN/Xydb
K/I5ayIIdsMk7h03E4LHwaB5hOcX+mik0vHK392PivO7wzTunPum7q5E+RTWish+DZRIFL9lI83L
W8DQb8nUuRzLpso99AJFwFwxLNcXQ9l+jdB7WceYD/K/NPm78/KDRiLIl9k6xDadsy8+Ja9/BDNI
qh201J2UQrhVTdla0rX1g1PeQH0HhxH7spMChcJX+sXNFigPazfwAHeEkGj6/WN2fGbW9cajbYLi
C0wWPz2c0wo18gtcT6hgYBuQHLiZvmwJ+0yjX/jkyVds+UMt18U6mg5/dE2woVyp/1fy0wXiCPQA
pujId3wH07wHwGHVLndlhtVPAw1aIRJEQ/vq9jVqa1c1kHqVEzIQQi5stxj4HahF202pEOHq553M
OLaP/dGkgTIPO/XdeYhqGk3XkH4bxFd9nyhpMU6pcfbmQiq0OTFZYzVexICgSBY6CGZyAaegrRNF
Vui90IWO94tnpcv7EuGMMhEOcph3tgjagvxNDCVTckkupMsQ/f9lLQzbohar8kiziKUlOW9R5l5Y
/ftoGUcoi9eNa95Oh2OeIIkTtDF0fjYkcaEl+4ro92dPd8aL3d1aQ9HhEBcy5DasNFhxyhUCLFk8
7tPU+FnixIuXnOAZQpUN/I8pZgG+BGivQV4cAjiN0XEDyRcVplqFrMKtktuYww7PPz9mpGR7anMt
RKEBNWlYzRGw0soSHRQ9AAphKT+DJMMXqIQle+LGmADbSJ91xdYvxXMvHoZSJPIkLiYtN25LSTpr
zl6GBuBPl2FI/LjMJXEIw0cXxk1IkrX8t/0en/Sis3RRyzW+uM1p3BIaWaveL2KtsmCk8oqyVWsG
dx0Z80892ZUiJJUBAT+0Hy90XS7eaR30FD2XhaGWtmo2qAVJhzdDrmp88DnFpzRR+ElN8rBvEjGT
xHCgfmMYneCfYEnp7/6OdeDxxEwK65hitSZ+qhUd17tXFioT9bv3KqPP32GmT1cMwmzGqHq/umfz
9DknCdmh2X+m+qKyZw/U516FCNFfo5f7yRWbEd9Set9mcUzfKnu2sMHj/2jqEvx4ZJnJVRQWO1TN
N8H1f0jkojZ/Ywas2Geb68ijEF3CKGu0EsoUQJJpeoHEm9LnbXTq0J7X4MHp3KPLDK8nnJoyaSfs
Xf6IvNe1fIze6knFTutLebttImY8n+7K0hj8kGTJNdV760PEFqGWzgZEjuVB8lkZnYMf7UcNdPsK
bFjjZ+SMi7ciilK6JYq2d3poTc+6T1RHUccxVqWZpVxjeWXFBGr7y2TK0riGWoMgWaCYdJH/9Vky
zkzeTElYagtBhgRQm1fx4XRDxuSvZG0VCjFJ69QvHXYxZexhBTfSZEQ88bOcw/lZnoh0kyleK/zg
hIUA0TUH4oENkGafUiuh4GLEDdRcAWqIOddoJPkFUCqap+0KGDCYI3p3eccpYZoJ9130wqlJZPIe
0UvMoJw1qUtYVSMgyikIqe6RkXdXaQEL2TqYwrnM6E/Eu+VfBfMk+L+a7XjlQwdO9rQAN3Dvn7M4
00Ro4m0kwhR0/Hpy9SUKmRd6bH2dPO696/wpdUK0e/pdJdrfsWigf29fBsAnG83SUNCQtEl4Y4R5
ZbQgzaWOybJ1IXMR/211lFAkNJmgBuVAg8TWX0ihGuGhYAN9e4E5HudULiJKJGFBBoRuRM54t99u
9C+FfwPIZ2baAa5Bqoimctm8PIQKkIS7G/wzvrX5mtjUMswS7CWup49zWoIou8SQ+P+5Leh57PlL
Ipj0KvQXUedPZP3QvczLimm7msx7tJ0Vgq21Mcri/s+sWUXT5geoQ5ImcBdOgwAjF/ze6HidWaAl
i90zKTRYNdpOLqRBcr/bwyZMpgxXaERoFYCEulp2in70J08BYUnH2YM6LsY7n2D1BMGtjiMbJONA
cYTbAx3hqJiec86IQz3PrxvYLmGM+XlRXLgjaOLehusbqMIYQGzh7FoMUdQd+Rqntj2XS/RQ6+Za
HObde1FIFPfc+qVOcKmc2V4A2fwFqU8Cauve5vQKMSaskiuYqbzGkcf5gw+c9A9IhE2TwNBBoPaK
iJLDbRYpVgZjTSDfLHgw9WRvde6kVw2pthI+FeqSHrK3WOf7/uQrygqDOnXhET7GkiRL80s6s9jL
xWGCrPzBHPd1H3ZPLshZpzC6RIwdBtzNE9bPHTk/dGPoUjIsWva68FSYQxLrucucqdRsV2I+ZrmN
1iYp234kkUyBWJOtug8jptGBcEAWBnVNl6Nb34UjPCCb22bslWTNdNOmxY5QvhYYfSIxTUqvMrqp
qh1Q0aXyAnm8RSkfLM4bSWPjfsW9POio2aw1VddQpjrzVvujuUnz5aTurHuflTVPthYau6m9XODj
d2GFrnt21iCD1w5fV9Wk44U7dV7TsSP3Sdez8upUAMNu63DdqWVuVmGNt+cz1hw+0MsLjj0oCFLL
n/cJK6GqGBGFf/Esn6eDV+zKKvo+MT5asYi9CsAYAyq394FZxrgROkuPMLgRlUdRaEiE6yy+AL+O
C3SO3FqPMlJ6lNvCTpV9ZICZsDT3nFXKMOD4Hk2AkBVPh5lqBkGjhe/Jsyd2q1tlD74aAphkd4na
7+RscrN9CGnYf1iV7ss2GDjtzoGDiQwf9V+L3RcRnU3CgEicyWQjjTQAfuM3UbPVRKuLlpfY4DMh
4Bym/jJdQnYIruxgpakZm8kYHBZtaxEz6+vfmnqmBeKImy5BS6FJg/FvGPyCHlfUQNVcrz6SqXaQ
bkAqwI6GYWe86emCT426qtmchgjq1NzyX6YN0/USRtY8Jb8C8Gg7MBZbfkeBninL0a7wH3HISyKO
PUL2PqZClpt3Pl8cps8AiNpHjjSNpZJEmxsxK4j20zdki4Hyc4AK+pUNps/nyqouG9nCxZ40818Z
+ldj1fT5OxrtjT5iZN8oEu2BJr8DMEP3GjyuCqGjMip6Yntuq0uIToakpqZMIVIRg2a6skoeHL0i
nhfoxpd00MJsZN2ieTIkzwjTrxiZfKss7ifIy/QCNuiwCGMqKreAZuPA6l4bYw749CD+YDnzJUJ5
U2k7ZAq1Hcr/18QxYJnGZCusF8rz/V1OPFZzihsB/NENVZqcd+Wg29YhDw1nEhT46mNBrFU0GQWP
gaa0HdPsbd3uk37PXkn2QG/fpxHmoapFJw4jO1UPmQRwcx74WtL67hRSng3FFbnEBIZIpwTQ711j
Z5c8bCeFpmlrpmJMQuMPdxrb5ZNgTwrll6fKCL5VLRcRNIwYhlCVMtdLs6KiA6BWWvxVelGbtGAF
+kThsVxxKqq71oGChoXv1eoE0iQopxBOtzMzsKaUW5rQ4S8LZ0fyc9DALgvK/FjpHutVoItDSIFb
9Re92Ez3J8f7MBbO/OK15IuY5gRG9Q/NnVUnK8SY3We7B/tQ0falohYKdWcoSeztcXxIaLhajd0X
p2iY/rJcPN5VNsoSJgb2ny28MtNaQZLopwWe4I/1uZuGY3FaIa0VEEI9iA0qBHk8Ytn0C1Lr7ilC
VxFXCUgsFBdwIfZLiRzx5KL8K4yVJVDZlZ85xvfk+3V+7BmBHY6q1ZY8u2lps/LEk6VYSngQ+HnJ
/1uSbej/TD/+6ducKULv9NeKH1OAkafSaDw4iBdcHtyJWUAzT/GN9LfNBsiI2F1ZgcdQ4w1uhIgM
bB8DRW12qSl1FbxofoKPxN6qc0D2rgyNIWBS2yWqz/V+n7fU7nZPjWoIjqHbRwL2PPgq4ucG6WdD
bGK5k8g4196p9YRaJc+vftAYnFKIbE1LTOY1GSNF+P1TNucwFbyMiC01ScqRCsi1STfjijVplnvJ
PqIpFL6h8vKpcLhj9q4ANPuu2P0pmzJOk1ct2CMu/hMhub3IIZ/vUUFstuhupbv8Yd+hiPSoNe8/
xdJSGEOafIsbphTQ6/xYZ1CVM3nIy8WLazmkeTDz2ntCEp24cW0FuBOMAVPZqZDuFQgvSz7HrLLg
6hhDltAWne0g2a6xIGno8aXm8vNggCHsNMLlVRaX+B1GM+L55YUfLmBIvuBuEW1JIrqP827G241a
lIYH4ezHdkyfv21Cd3xAgAhJSlUUdnx//2B6fgOmjPmdM68vIafe44vZ/ngXHgfyuXPIcGrkbbOO
2j732/2hFH0SuMKaBsfvsYUMGKk48Nq0AJGdl1FRaWCmdh+vvzICFfZuDSryAd+U4sR5+Y4wHopF
u5hiPW/BbYUnjaMSoAXJ2LwxG3Vdv47dZyuj18JbhU9v3G4FeyXrnO0yASc24cNE4C2ZHlURR1Co
CUuGi4CNjtEQYtkPJNPOaUsdx1xCX/AfEnUMfuIaEPwBkyrfCVpV4Bt6tVN1WCjdSaGA6aKP5EHI
40PB/iw7WIFZF/46MbfWSCPoxNltDM9C6y0/CpxqU04f3BqUu5T/V03bndLqQ3pDdVExZcbP57uI
uHDIQj9oq8uaWXgs50BSFUXHmPOHhQ0TgQowphjAMAblFLnn1UJ17gQ0I+EO4TKtVukTuiiG8Cxt
LZ+KglAN8TeJ8Za0mWmKYbH0Nr9FL1ykRY1LcyCyGJOACL78hJ2FpqPnZ3iAf0/k8CDT34xCfQMw
F7wLuse6S/YyhmQFDHyf6GrgFzwJ7JJ31Jt2PALizrnWFW0CEo+4+/YzUO/j3kriErBGuNd5xorr
16wBvrzMhLtCsi08ELbSlwp+Id2+kv5S6MeviisorvqxTGylxLTZBhbYxszITTZ+P1WT2wVQT7gf
xIXwYWmPRj8nkUIrVgSP9TSqvTtKjFDg17m2uQJwuGNgfMF24/4T+V4vz/vyhMc6xBMA8Zvx94Ln
WlNa48MMdyu0oi2iNrSgivPkjNXbDoOZjl6ovNjuPd5Sv4wHS0UZNUVSYV5Edfv0pJEQND08hhLj
A5yhYIiPf6SZSz4y6NlNoUsEYG87L8uy186+BOVF9pXnzbJGLdayt8GMLz4AKKtpkuGzr8V8LJ/w
8l/aZ32/jeOfkdUsLG0d2KICRKT49MBINh9egq62gEo0FF5SQhGHs1vdqd97oDI9g0tFD2dC6UuX
8RwT0AMMey8tWA9LsHOtEH/hyeRUKZ6XB/VIWmEMO6NtWhj+lFyLE7aPEbJUOlqRAHU3S83yPJbU
q7T85jZbeoDbNT2R2xGbxAsZPQ2IB6mY+JmzIewbD/49sZbphJscPWPc9nuJU01mCBerycHit/Go
ogyyT4XHuVlI3ahaiq5OuKjofCTzJiAw7fLcQRCe17q5yobbNklbpRBBtFdxnDRxh7cizw0qYvKD
ug2iBHD6yBRxNTjRNp1Y3MwO8ddjuO+mGRMcN58qYtXUeYk7sd6TQaY9fSmhwauAmaxl4huxoB4C
4Lqo3xig/DhF/OlYQSJXUaS17vX2QlHaRpckeBsvlDGKFkA7Fegnm6D3+22QtAncJggRyCztQTe+
0NXJRHX3Dc/v8LV83lI6rXFRvtG7XulgMHCUIWn8KC+lSF9ngCotxz4/Ve90/ZrkEDVrBztp/qE6
bRn/51BlYFd4qPyNQ/zc7/ITlz1LQsbkNG/4cITgiAz9nQnRX5Ztfo4TCzsLPtxhp4nYFk2/KARo
TvAbinXbNDVgSLCZ9bgK9ACoEpTKd8/gddl3QCotSmlX2yp+wmbMrjQg2CvFRBbIpSl9l1+AyAJ/
cufdM0UDweEyoeoc4NN5WBH86yhMWf4wyq2PVvFmFhq1yKf0sQeAISEKtokFmMWJkGa8Wn6ApRUE
P/DIIpgZPlDjB4rsTpRVC6TTIWrfVsu7IZf0I+DcSnpUs4/H9V6VEPxf61Sjm14sU9Rptz6mT40C
6b3+IGR7ip+SrFm0oOaDSvyWCjyN68kEM62CW2ZClhemp7sr4pnySgV7bXlcepTSfVSmIgmfpFLE
+yA2rhRO4r2CGHQequIAyXbyZk3r6pESVwQC78gr4uLnZQs28AzV7M8X3Pu3H8nTJvb1q3QDVILZ
YygmFlDW2UmUznkMgqkxTlbh/4GBSFgjB3GdKjV9YIWEgyy4L9gzJIoyFj7BMDl5VNr5h/RQ61OS
a5dX4vh3B9jo1EpND41uk7y70QsFnQk2dX4FYHdfJySpD+1Lag9a0NBMt2gdeV7gd+rmijmKOjA7
dcxZ1gL53Jkd2xUd/sUEI43hY+OyGfAPe+RdHWZXHXiDIHSC+oeLFV1cWJOHI23QRHd2kzU2kEm4
MHeG11jC96liUF8rOaPTMbVjvgMplte5l7vyXXyIx3wU08nZh5NxhXTjS0omxyWpNSi8A1lclK5C
uAFW1W1WupmQJnMm9W0Dh1TQ2KOpenDLYDWEool4hf6El3X2RC+4P0AJfh3g820sAcNwEoUqKukz
mXQaQ9O730zYWPqm6Zi06yZU3R/SIee24DDK/RqOowwo69jwLfKb7wWRfpl00n86PnCW2qPISJKq
iaShQtsABEXMe/fQiV+6LvFDn6Ujdakd7/IlUlaV1XEL1zCTzDDqXyUqzBlYgAMCCJVH4AyvUhOz
DjJkOtd7X/U/J/7eazwr+rtdIm0QBQ9Q0SIRY4o92Ec3wHe8JHm/6NJz0EjNXfPpz4kRruWxDm4S
eiprwrAcTc+9/GE82BmRic1a/OoqcDwnagByB7V2Xk8YXTLbMD23xVH3OFTa0XdcP9+YhSugBXZZ
9DabGV3WdNV05Ia6Bclum3uQF3AQWIGIg6ExI/Ne4HCYD++XWUcfLxfcg39VOdafN1vhYCDIGE4e
4xNQCKTutH/tirDjwcGcrf071z24rUonscTX71mRjTGDHlZHzrHpE/tDZi0scUDLzCZaCBV5rsr3
36R6rhyOVsGwUdU3tyS8GvI919budIFJD1Yb8pvx9rNt0SHrKCszAuBrIGxJrp0sODCj1qMOPhvJ
HhoP9Igs9IMxIDOJt97UX0H2sp07iSjY/yAXOZhLS9b+5u0s7f/er+R5/KyYQKhscljUCBJXxv95
k9ktfD9b7F+n7g17s1ec9IingFB/FOV1Ck2zYWhq3s/5DaMQqA9qrZfCli3ySxx3M4UVoA+jm1ng
gNXuqr9eMDMq08YUf40gZ0BzHlkG5iLNIKZdFccIGN8FFtzth1P9xeZQ7tvqF4L73mxfeYn0zMar
i2pgzSPAhLXdc+qTYYCgNUDKxqN5BdrrZnlKs4kE/D2yKXDpdZIfgGG2h0n5or0CfaMyeTxjnKdx
4nCSTnY7zqX1cBGjQbNNlIEonErG1W7eO473gRzvwl4byLjcBeKQYN660skshb4zcnwO6C01L4M7
yH55ePCnA8czlA6Nk7uaLkkudTl2NaSq8vevlehgzUo9/VcAjFOOB/Et6ixnSIZ92NoKmG2MNbZ8
hDtEZR3+ogcltgBeTA/IXPta4RhGeRdp3flbYpsa+nd1tC24sVBz3ee850Z63OgadR4x4J/CJlnK
vDp8dQzd6OG7eYWud7zH07AwzhduALxNHaSosGntYwwOgDcEFsVS0OpHfwormyYDbZX4upedWkoC
FO2teAnmthBAGq0M67kKlZh1SowKxW8yizgcIbxnyTLxNj0QRqDidKEKoiEehlZqro+y9HMZDmdu
yTu2ubDdS6nfBn01njgt/xVLhNEsErX9CVjMv3PgftPb74cADggKUthjL6UUgFeR8hIjs9O8jrdT
5uDGVj4bToshbahyHPTYoG8vALYBHRFFtSbjubVodmXp2TmaunkL9P0j13OaOvLVvGNCKkit10dJ
I7L3YzHAH94vkrDiMMmULtZceamQRSbptnmM8PuY5PHkWMwKnenTNyxt3hFBPJD73jaaL0k0eBFW
3AqQpDggQZNLaLNvb4iXI0s22Vx6rgZV70dG4LnXEIbF/mALhmAlMq04mgUZQTgrMKqfT3vCWtEw
RwbqADzKAheVrBYzSqn34gT5H4MKvRFzTqxugCrEHR+++8RzkRYZQTqSNQ6xKfHRC3+2QumPMdMb
/fg2oAw03yZsak9agwUioCA58TrgtNwoPyvvrSqGeQGco8oEHISy4FzuhuAvTn0fhMELPqBQgGha
++sm+XuFW413a/UJQrm7f1LoTPdZD3dOlmhYqnGlGPuew1qkncF4Dcmk/szXQqdt6k/eJti8TfZe
sHVsoMX5fxqr5mwBHoYyGjCU0O2agxN/wHiEBjmgJpFXAH3wotm450i6UxCwIDQibaqfkqQ4V0yQ
HfUyiNalny59nRLIqMT+Pdkc/GNYXX9BTCdDSe5SfNH/6Xo3sED1ou+6uBQNmtYsRHo4DJmBqtnv
nzJFjRuL6aZdq4KpnhVOqhYjePrp8NRSxDb951UhQNw7EJJOSCMeq/0gjwcBkME+2gAcSBnYAJZJ
BYXidYJ8bLrL5bnm7csbt8osG3bGWWUrFpzxROoDPhHhejkdD9WRb6UcCRcDU7dVjkgPBq2quh/B
/QozVGClb7i5PS7JAU2NaNsruIxTVz8JuoRO9zP7fPZaNfKrgln2WomYuOhqcP2/SDB1f0F8+4JP
wIkJMEWR2qC/jN3GqYvQdhkAHDn4GEBTgFslhjz8/mJxegPTcZqgWu+j/bNRM56afeSnALeC/CwJ
IUbINTXb9mJQ15+5I4+IFYlKRYe8cNQnRV8u3cxzxy5gcoAt+Cu57g1bxWmfRv8tuF4iOv8PDlDi
p28qXbQ19tYxFmHYfRiJXkPPdlDsY5JiStCS0WZVgq8TMRYmBZ3y0fWzyN/nhJe/AaMEJnSlUXUG
o1kGT8+xOzjsYgzchfr2SGD3E/LT1hqFnAIzZLtYdWxEIeHfUTg+x8UEt8BEO83QB5Gs1nE9DMb7
eEQUyA2E35aK5GNXk6t+MIPQF16YKp++/n+NYmmILyiMw5rCyNcc+igk5KAfG27XhnlM9GbujE47
tQFrrpN/65spAsFE1UN3gHKpBo1vwQ/cOkVJZFieu4StA3EaaAH4zxxy4M54wldRy6CrBzbrC2Os
a8aS0S0y4vSYOPz00h5iUAHgbRm5IzpbcxAd/RjoiZYZngL/rxmpx/TbwhnvnoFfKcjCGZuueRUJ
Ie6c5XA/G5FvrMC5EskRKaeSnKRxKQTRT5lcXswN6XMCVqc3jENgHUJkaI3pfO3O3/LfxFxYL1mH
JKeYba1quKkV1/o4Y0Xhi+yHns1BmE1mOl54gtgrEwzJfxXuQDhI1HPHtZ34xQdisedHYBd+nGKM
h+gw9iYef3ofXRx1xb/m30f7o0sMvh7BTq+g88OmAtvgks1BzRAtZSzlMsQmbLrtHJCJC2TRwOpR
eCC0eUzCovE9YFCCsAnU7kj3XIqaKhKTal1P4v6LytOXSrByqRh5Ss+bDcDvuXaZPib42gBzXDpF
LiLvbttFYdncgvKg8mP20C0hibmesrDpEv7ZXbQfhGkh+531pzQId6tGcRpD4qNUaqdw4gpkY4sY
3fJ52qyIXjsk+SAOIxIfGxLsXFkgFdxowV+VypkBiIx1sLu3AGze1QatTU151yRFpyaNCTIetYxH
FrBKCGvMsZKXs5j9dupPcnW5yamskhU0J5RTIcAtbys+DquBzBAMyJ+I4wJ/V1diz9r5wR27y/eH
JuofjctwyNO+6z2s6Vvc78bUsjGWoz5AGAWsBWKOkF4TF52Gm20sb2thOvg3ZvYDRcURoyLDIH01
un3BD+RcbqASgAhytnxqJTfB/bk8IvrrlS0AIVC8gEKwWMtJXFsy/fN/P/mr5d/T3dyGE4IWRukO
X7va3krtjrhY8vRn/M7fM0nD0bEyPl949wHuLa2vsICanZ4c37Ok6PXtpBbsfjsYzcsJfrhwT3ou
jfma0mSsYN1ByftlWwNBeAk7CHs0X7WRdqOIauUF36y1Rv2gSzOx/aidO4UlQh4KZY5GGHcACV0z
qd+Uz7ZY7StDMOuOfEbTdpRMj6w5yz6FTUHRPy/r/kpnkiiYC6jtxFP703qwBFvISlZFvAE1uz0e
bouUgT831FJkBa7w1uD5qN44tmE8G03LerlZiVydahnplfXrHHGnAme6wLBg/gcAKAUIUXBIrJ1C
vC+XhwJiU+62CzsUpeayVBqGMH57KkTdi+xU3gd+SeaLjCK8NUYRmQdhWemAAybAt/2wE93bQmFr
lSs3CTqr8/t9MwjkuGvPtZYdA6hcVlB5vAFafRR3FP2sOB4/ZjvEA71mC8hDquCCIRNgdmX0XX3B
wRLCsU1oVmC3iiu34m8fd0SZyh07n7mAZ4GD9gAj70ftJfF0JR59IwRchxGRpnnMQ2pTF/cmT6MN
4VMxLAz/UmejZZFPM+30KAYtvbOBTzg+XIazWc4VLSRxhO6dnJxAVYx2IfG6pK2aLvj9UUL6kSYY
cf9mvkEJsbRVsZsM4FJ/fQJn4Usl4BnOOPG47DlXJsVQdAu6PWL2G28PqxltcIY2adqM83Wg0oTx
eVYscLE6FjlLFHYkmTBv+1ldAfer75a+mJS5rpciajOzHNWym2F4b8mLUl4IcipQplK71XPkfLVm
IYjKd2j4RmaKSBumYeMt9tv4c7APZDJE6tgFDLLUrP38fkVpBjgXnPhzFkb3PVyoLHd7TP81N/9A
VAooPGVw8ePcbuC0PWQUR8tI81/289kPuTRh4qqVapQ0ild38jhUfBFGKmM8AeCsxow/3+r+E1IU
hZI7FR1sadgoh1Ui7QtDP9Y2sI53peKACYn3UsaouE6GLBmYRSm+V1UPHyB2aADSbo2qfhejzd44
PJHQSGlgufqk7WqbA+OqHfgVu5EjgvZarebSS1bwQvW79bW1Hi/KjCX5enjH7cvUT/ghLp6XA2lf
CaayQJ1lkqMhMMUdW4uQfoV1PhNbMe0JNS6gVDFskrRELtO/JhGjPKXpa1/aRX7SDO7PvxfGpJ57
mSzcYWlWmwjhxM7/f179LbdXkA2pCt+/CyPOFCgdTjwNtaLbhZkVV9BdJ4Ab2GTeSc3d4NkzeibH
f2miAMYpRHm0i2Xx9upm1tbsPq6H/1OodAcEs1N1oelgBec6d5+XpjDGYO4wNj/DKwLOsu+dK3M9
/5bIRNLGNpKUoeKrOlRVHyuEy/JbcNdEXrI1vjVlQrC9St6jtSAxw3Kj3AIJPfYLuTsFk3t+82E6
zZLTLQWfJpf6nJqcHb1EDCmixYwuAykHDw6snErmVZ0s41tDYCE5zJXI9yt0x68iZxrmha37YbjH
OGooJWJfKBsmb9xhhfofpc0jdLNDrHf9YqS87Ph5fJxoKrn9coz+X2viDbtWnouETVo39+Cp+BL0
w/1Mxbwd2Zb6CZxHg9jbAZ5Y/vaY1sEeV+WXKXieMr2b1Butfnokvi0Jg60gIEIrl3kFMqgjfO7n
/dCFr6GdSuGa9l9Bsh89VodsuVM3Oj6HJ76hEmScXm21FHyXws/HmQxsGs7o+sEvbcT1WN+lhs7O
llYnVKDLaZBTtWfJf4UKRVMK/WSf2658jCVze1PxfXeGCRlgU5lW4tTD6zo6tYzTRlTGe3NF7+be
19624nT5jLnP7o/k2BpWkxsS2vYFLdMzBuOMCUyCshb0WkpwODDAnwVfV1pbhoDbB5fTxDq/oBmQ
/ico2IccB9wH616Xtcn4lRsMbX4GlbJcJxZi0Kzuom9m1bgqnmO6K1/qim2fm8ANmi57aFVxkcEr
zS49q4OyTbXxfjvrhh69NmQY09PTtehxtEwOwWfVhh2TU8qIxPwryZytnu7bU1PFwBeHHamudP2R
sAyIowIytO3qAXlDb2pVaPCwsgJfBpFIHsBJ0LzpFKS6MoxTk3RJ4Bme6MVFGGfaih71+dH5D0Ru
Tg/PWwMJGU7kB9HXXX3ledwfv9Ch8sT/kNKTEiBUD+qr5KoXB5SAwaL6c5SGWOkMXNMkdXWnFXtX
auZE7EES4PIgWmUV1CPIGlWNZLGiph52dcRMdCw81KnyRczpcZsmWylz3xRI7yk5SdY9DKnuIYU3
v8tihpmz/dMRRExBCgFq1NvDLOngyM5OtpKtHdQM2L6gMCV9tcY9+AOtkLIAgzkAC7okvg9buUB2
rgT7LFdEPRSTAZdv7XvNn2iNp4Oa3M9VaIartJACJF8YbjwBTNu4mA8DZk68wvMBPBzSL9oOX9YC
25yXFsoWA8o4r+/dXuiuU/tSr7M/THghxm/U0KHM4mnPqTpRcP9XfLFphy0Dj/2WF8rwMDxPtJBq
NZ3lZgVs4lz/dHI85VV78M+6nl1IGJEGgEgl05URY5m1m6M2IpIPzNbwMEeSAtUTje6eMWYJrGGR
Dn12m7vZwIWFf9eah9T3CzC5OF+pcmA4IY+U6cAUxieNpPJ4CF9BLE82kcgirZ/+hNnuJqRa6cen
Mr1sqLbDAYVCUwR68zeBW0/zFgCoFxjSRs9BdrLCS3iy1tGlDJRoOxCY3zOR3AGqgZ/7fNjKUt5D
BFRMO34NYPjMZXMjyWdKkgR5e62UweoCh8At4BFOd1LMeatIy3yZrrGKt6OfFS0wFIAlwcd2kSpr
8460SISXlP7KiM+tEmGNREp7BcNGImEk/Ru+psGS8wm4nucCPO6B81WGUBTKkaXppe9U/dlc86md
hrLOcn3fNfAeUrfl3Z+NktYyX20SmeCqS6FcwZBgXZm5CJvIjQkk3DTn6nl7VAyuuQffNObrNNfX
JUtBwnRQnzn5X3VVffxOskIYKyzIn+DuidraeTtetuDvQmyRLjA2RdHWzdeHxVzzMKCBfbtNDCxw
YF+7WejIazDigfwVBdPzdqeH8Zqa0kaZp8KlQoY0LYUDJAEROQ/JtwyrzjKf34MJwCdfUTdCyO0O
F2+TEqQnsV4+7TeJPlllQat6VwatfxLd5PmTqY49MLejIZlvF3hmh4khxe5/mPSmnMlSSkONuqVq
JlyK3p6UtlTsmT2eDSfncngMx+xNcB22uukyhBmkS1Lrgh5la3kIEvPndnNa2zw3V/AvLxiyc8Fr
Lmk4ZqWG3il8EDccKwAkt7BY/lQ0oORIHbElcCThyIG4hRBAha/ZBTqdAbyBo7+FnHphDpAtDS+r
MsnWo6Qi7hXXED9q/zAbsEfkwXunwwuFu4Pkv6pwoCp7cUafj5iZf4dy/UxcXaHVZ5GM/llETsgc
/G8tISVekJESj7e2MVjS4ZAA8WtGFMzPkeuoW2CGP9iXRMIjIxiXsg2FeNhNu3tQoOmPcaZk8u5l
8ZxtjFxH9sIxnGor0UUNDtgwINmfk98s4QKxbUJvEXMJhfLyThtikwXBYuWnUNoxsrHNvUwfHs5U
OmvmU1/pMjsjrwMsfnaCkrJliaRVl/AJGQ/z0Z0Pb6ii5V/lTBIpNX/kpltC7kZTjqzk0bP5ODkw
HdRZuYQKe66GFJpYsX5ep5OZAMXI0grdP9Jleh7IMJqeTat5R/jwmxYeeL3InYVEyKOt122tDxIj
zpBqXr9z7+FXcayj1Z9IGxgIYW7IvCpbKMls+wTeAl1ncaAZnTOoHyei05iZbt8wU1urmUXV2kqF
8fut0crLANF5WJqycrP1AZbccgLiiffrHFomAPiBzZqEd2DfZrFS5oyIrYTpDDEWjDaT4oJR7rme
f++SK/04qFXq87rJVU0z+DwxdVWSJW2oiMI/6XP9Jb67bxd9GMhq1P56TXI6O0w8vFoeQW56ZqnF
WvJcg4rU8GscCbA6M/p1syXwI2Q8cLsCl1/VlCv2XU3EEu3fsdye3qS2GMbfUCSXwbWrG0SJvbhq
m9aegAbQI14FMzUTe5ivdUg/8q30/AskCETr6vw3M/WnauEv+fIQSJt3f496G6okcgcOs5at6scB
p8B6omDauQtm7i5csvN3awPCoPU5qDt0pKb5KkKLBK/AFavPm7rURQAEYwz88D2BRal9SPZb9qM9
KfmfuKcOFd2tb0PEmukc2SFt/69b/KcB3tNDm1zL+quclGKymxX+Vzy1zg298KXFyXtZS/ljk0+p
3YwRC7LVan8oMJNpjvhmQ1/iRFfNQFS64T0GNOEtCkb+7advcWRfG/0WWisnXHmMLXcyMdpqFN6U
7CYYSFjs8XLWEwN3IywAh2jOjiQl392EFayh9rVnGJTg2jiMi977K3nDNHvHHkF7w10q/yeKOPD+
0+/IOnPah2AI1bSP4SoxjBY5XjP41jCDIxOSwR28tSTEqKBhpGPVsDh/NI+NDnEMS6ih6p7Z0ybJ
shQqVA382HVt7h8clx5qhMCeLUx3aQwnckY5tw/jJstUsnLbrbE9X2cgZLGl/i+um1m1wXm+tljd
ca4gVRlffaYhDwHG2tmduvgD+yNMWiWn8w7ZwlgtkXzJLPGZGybCxpWXS6/5+hOxwpumnoIHhxMh
Pv5K0EMghOVemllVJ2Y75abhksII2noqWs5A1vEH+ElASLuzNxlNhRU6fhHxYQLeSq330qecsnsI
q+mPlI4sMbHWPMONvXnNLFn1dQ0p74M5vsMYd+6WvFRAYXjYOqUZ/lxZPGnZoQykxwDuGiLuEJDD
PJX+fpnkJ2NIA1vj9K5FzxA8ohqyyfvt74S/snzSO3SjVob5u34amKbLO9uIqcQoSebKMq+rx/Yy
JSE/lNkVr0L9Dv2wKbYsAXBubHFkVll/L1GD7m4IhgDh2+cwv4f5Fv4TRucR/V/uIFRdGrsqZAlM
2mroS5wpK3cm1vYuc3xOzunc1HG/V+20QedgSdp9Rt/GwRQzriIItEDXv3NqiBfaiolq+MfJ3Ntx
ht29mK9LsTL2MurQOKvydaGkxD86KMfJuULn9659AdXyQi/EUYq5MP4ByBqVnzLWKqE46i8pY5T/
EvHN4oMVQ/pXi4eWYY15CI4kErHfdzZeghExQM8IjFhUQasZijZIeIySkbD5cmS1F5cYCuOxhpyS
8MddY0pUDO3eDakY8OAxAJTB2TJkFu2jCO2ag0j2MVFij/1Y3lX8+CqFTOf0gOqqLIDvTIjooDdt
VAdOlxvNxyFEjOp7H/2miU9WaqIzXWHnFsjEa4JSnu7B5hLB4snmwtF2UoPov7Gz879sTXmPm+Gv
tgnyI7RIqNbbjd34bJUavRZ+7Kz4UXSCUKk2cvry1ulHlTZerjWXc6kpDOrokuRjty+xCSJmTfNu
B2nzB3uje7PSL3cgLiDzWYM0APA0ebmnuxzIWCEAIT5AtRSx8kF+oI0S9v0YfJUM5Z2suOJTm/FG
ptscubewC1XC8pfiQSguVNRASjFoLveuiWOkOnj6kqfKBAjJ9c7WL5Dyn8HhKxf/hqkV7P7AEKkf
8k8MYzs63IRqyS8lXpBQqqnBP9wepl4KcEcNWnWUeQkYnjz57wVsUUrys1qTJbiI/R4Y5v2fJapl
AFPGNMpsj5Q+w4eLmoTxNGxiV8cTSjJVX4ehrPZjIx8+dDptSRIv7e1wSxHMuRUaHVGrNuRgaZDp
6p+mCBwxcfBs+x2fJ3dfH28Y9tBfNRpaqbKC0F2r/FJC+3KWC5TSv6YffrNtUlNMy4K39mZzrqCm
8yUIuVm9iWxJb2WO/qhyAaT2SVTf9X4SLrAJa/2TNklS5QIh/Jv423AxPHl+AUML/IM/6Tk2H3xT
xEdul5g3KZUgHISBDZars1CBnG6rRYdZ8oDABP/o3p0mlQ46BkQvlW3fnC9iq24QPByHWdbEmx5z
7iORy2B7Ng/hz4uhgsYh4guS16JVQV83PyVV1tmh/nLPY+1lQUJzZEFbEIxCc4F6/24+FqlBI6gp
IZ5ZAOmcWNkiEkqjyRH/2Vf5eiUm5UxUXGjdt4wUVEMy0W66726JBszKDeRrNztUyWd7JxKIFuxv
vY83GpXZxzkBJd608LEB9NTfzi3vtQYFPNwsFBlA8LvWbJWFpnUqAvsdt9Ch7sadmFCmtJecDCFV
crGO9CukzdmIbzdwSFEFNzj2dU1jPV5/Rw5GhAitmCbve1JhKQZJFDczODEfgUdhUu1LQx2X9ZEk
zOeaBpV+Y+fmTDg5UL+wSNBBin+sQaje2g/dhNXGBVexYYnyZQHndKjrJftg24PiRGEW03W8wH14
sWAvp+LjJqzFg9PiVRL9VfPdouGJPZmukysHF+cqZmabvGalPWyV7AWkbQuqcBWF8C4kyyvJ0bkN
vkesXh+o4Zz44sZR0/1UOTagJULuRY/rVRdMU+LdD5mUmJzRNIKwlO9zj/cJS9HiF6UiXuYaRpuY
vR5eWbRRDTMY84OPpSlHnOK2rNKK6SqspdRDXi6dv9LWkOeEahQMrE0MwOQtkr81fYV9ka3T7pOd
OqES01iJmqPgYnUVdUYM9LdS6aWjQJbMzmuJcd/VKb78ty6Yz9/v0GIVlCjO57clnAAdtLbVgo/M
uSaO1ZxImd36KsodR+tysrOkvQXoZi024Km1kOnqyHbjLrl/u1CQnZdwXOjslnaGZTpNKKSGpD8R
pIvzjyAiLhQlzFoBUhjyYLuMqTfr2xZC08dEOk3uGeQy9b3r8nFMds2huznShI48vn0yA6QW5fD4
uPULIbC0Y3R7/VDoOcBbWZdLpAxbnwuxiaT7d3oXXNjGmhGcsrogP0/2+unHJhajOEQEMUU8retJ
sLincfy39GXUGxGNq0bkeHbLKsQxj0GNB+RPQ42OCwsN6NS+nvTUkchE+FpC8LEY1aqPU550nF70
Ep3RJfKpCKgaCUXsOAaFwe0p6K+wkJr189PKa5JvJ7FmrrSzf+ur/KG0qV3GdIpEZnET+Fh2Jz+T
kJnfZdr5G4vbFuqWWTcSeCwSt/AafVwvr4nM/bkmYiR7Gq0ZIgNgvBR88IcMW4EtiIT79xB3CrwQ
TYWiSg3+bkEm/uqycFJrhnIyaIrs3G1+0ocZtWud3ys5P3H0/fu9J/i7L9skiE1OhcfNhOLAfnq9
VFB69mvqdZXMKQ9y3gc4+yv3EAAohrOx0iYC5KRSqXK/ptn6BuerTFCoeqqydN39a59Psx61iuIS
1OP35vEjZvU8MZvNQyxl31Ngpy/0tfj0kiI39Md2rHp6KbxPpZpu7ErD5jWoElieeDfA5Ya4CAoi
+n4MRlDY+YjIxZqMqM9oHAOKTzb90b1NJett/Wnj5nOkWIRTshWGcOBpZ0qPP1aX31E6cKFOSl1Z
J9Xcj1gNofJ3PbGpqRLzG+l6JIlq5iM9LGqaO5lZxNzJE/nTS8iUu7QE2MFWVxy2qb80OWZAvDPJ
bcAsNQee3oJZLVl0YJT3dZur2M1cdV2zWmD1b/rT4RMoRQ18r4wP4lgXrVM4+91Wxjm4p8lfvHyJ
S1Zu4sjqCDvj4b6nAUJPJrWjTbOwztmsw4gm7dTRsR6cDZN4S0IofMlI5Pjd8vKeyLYvi9FG5qo6
fatk2Fm4Qxdr5o9Fu6E2+2QEvNwXOVJwsM3sJVvv6uZGB+js42qWinTmGK0tZTDYoiecqq+Ed2/0
5xIFJBkpYv+GUw+7GcGacoo1QKfjIMDGkHMOTYlaP+KpiufsZTc+kuqQBbwJCpkLAAoinZjp0J1w
KVaJudlV89zFrlPo6tuKVC6/o3s7DWV6IwHgH5n6X3pEdYvxRytWEAE74LKfw25E4+2+LprS7zXj
kzaUm4lG0ouruKXiNBF4mbclGfKDAwzP64Wo32gD1N2hZgxnV+uiEbU75i/IZBKqp7u4ExvOZXxG
GYHZR3gXu3xuxldk22GvGZsbbow7by0Vsre9XAV3aX41z3KfUrXND0bdtT0hiTIqoFYvNdRye115
cs5cix+VVtLJ0UuY7IeC7VkW6ALn+3NoHfWM5rZ9xeKX+n8tHX1VOIDfFsQu5frrEKifYNot2zM0
rIsD4WR8VYaQ3FsNGDMnPWRrnEQInYAEyo28fe35RpHR5wdN4DIcPgIuri2REO7AwjJ/gevtInhL
pTSSapQXSP186FDlP7ffechGnDRPAmQcygZePRWvqpQVa2e/RE4gU1HL1P87ewQ92rpWecozAtgp
vdTZ+RmYjKtKu7x1mhc7CzAwlNxxuZvkphg7OAJCccKIDzEjZPd3GSjFd5/KaZXsh7ZVpr2m1TXw
HCDxWr91f+1OIxmYvb2ltyNTYnPEBP0EEj9r+zhzonE6e0VcIhqNqudW0AmwhiYlimr5vqGUf34W
GAnC7Kb6mXBQcWGyHbVfC4i8pi0h2IZEHiVCUMHi2fTy5I8CJIxCsHXBpHJyLkZZ9G0klntalHDx
DhbXxmWDhj2F4Ym7excNHjptntOBevdXCXwDfmOdVWne1P+KQwm/2ewW+uWyzkGCDyHa6ngMpJR2
Vy/fclxoXeaPeqZlFLAO9aDU++deEqpUz+eMee8f7ZiGwD8du/nzMtIMTk2rzmo1EeMlRZL+4ETG
At6PJvRm/PHoYQdJWVxjVKI5DYaV3YRQ3L/lcCcp5U8oFjz6c1zTiSeZdOenbiiSoP4FPZNAkfDU
yUqjgZpUbUEdX29kZEhxAzw/cZQZ1CHc8OvRJ0Cys4OuDNGsY0h81Z4+wryuEuOmMHichW570U2D
o0Vlt/4fYWrXJjsWnUTy5C6tNnLjs8VIykQ72xT3UMyS+yIbCfjjtQuhre7QHev/jH2dh8KVO7Sk
jVctDWvXA+lKaXVkV4uvBAyEgaSLDQQ1FHbS8qd6q3kJanDTmLK96hnT8LmcfSba9aZX11mdMSQe
fRiRlNLJ24P3GLb0exfcPtXM0qhYL9zg3hQ3/m0uULDI/1dojZ6ULTh2LtH1UaznlBdFA8BNCJj/
wqK3+VSK6Uwy7UslABfEagg8ylqxyQcQLjSQSUaok1IsRDwUwOGiDs5FeK1i/KslauXKnxn6BMSW
i7tDgnLZBqE6Y9xi85uPBANjnWhx+Wc2jtwnZLEs6zmxN8O3q+Tj3ZOX3KU7ArnLABV8GB3fql61
O6Z8tJ/gCazrqShxRV5vnmIFi4FsoLbPfKK7q4KT9blcXsJ84iuD+6eejf+sy1Ie8zLw2bHCbuPb
78im5Pew+t4tXumlYt4j1n1rJevXR5Xyj2hZNE4bsuFwXSTL7cUjg2Q9Qp2EdJvHbXMYjCNO+CCL
V2sIPxi8BsM9SDQilWkg+ieppxDRcJkzvgmaluaakRbHckS5OuTjIMNDceGfSG4LlQupNAIu0O4G
4qEK61IPlbz1lwN3k1vn1ypygX/VGstnEGNyNmAufYXdJvTxqOhBd8rhM1kA8TlfF7Qsxo67fsni
G98l2kpQKOVAe/QhyYoBVsMFtFR7/VtWSq6hXFE3kU9qrCD8dxWLHlkc/8KA+YobIdTwqgenGx+x
yrhLnFYeO5sZZUh3yw5GttbexYRmbDFLe9Z0hVKpr81iRIgX51aifcOFfKOYdTbVxULkX2V54+nZ
giQPpz2rQde3W+qfmh9XeoVMdFzU7eJSkJGGf+IpODaNbP60zOKhVJwxW/4nq4Kfu3A+gIa/VxvK
tepAgkaXM3VleVUfwe4vMflkrakCTDLNUsYgw1gC95rQMf53XFggdyh1Y5RJ4z6xkcNI1Oty1rah
ZFd8wTtCFE9/hCq5pIY0aG5n4WunG9v8Bi/VElTTxwa82fY+Wd1YUjyApA3EXfwmJ2/hf0qC2u46
HsNBtmJ2UC5BkWxPC+4vTwqwJ94fBoMY/gupCWaLN3D5e8cQqamv/tKIv1TkQceCdYNRGB8iEEIc
+Ri0hgEQuvXAOb9WPPwClpM62/boVZ1raEmP9dJ+RAsXbDvcVkB0T2g8HuN304oMKWnDL8ZnY2qS
QgoFQjLfYWKbEv9ppvLP+btBl9Q2WlIVSXb/Z+G+7U8BaMrSlBKgeQJhQtJUkgBscI5tlw6GTXJP
HvuqrsgL8SiLhjgh/xq3jo6oyeE3nYcP+xwOlUXp8MXRa7paGpn5m1J2xoVqYwUPTmvjUDa1ZYLq
Zj/1DjbSH2b5CM+4xOwidj42KMHKWNA+VZLCaM2XVU+oHKOVo7pPyF/Fg93fdxXNzLtbBHRG4Kvh
0E3G2Lljmg/7FL6V/4g3o/nHrpIyrkseo+ZGxG5O3JYLx8/UbQCNelK+NHeAUxCyEfhuYosdk5Io
VUPDG5QltV4gw5kW/chH+YOx1W7IZfVbxbwTROF6udbV5xG/LoGl8/zoZCDvuABIj3SgRR64BpPw
yZA/3oq4n1CPvGiW89LmcoLodncvTF1EIWkRAUh99eVUZKFDHZBIzBfqUNXjkvIUZHi4/2vp0C8d
wove3tHb76t0C6qu1/7n2s+78AL3B6fXRg3DhQeQFRpNmsL725+HOyPJ2NhWoaODuB8V3Qou3he+
ZvnJccorZNk2wgOClbZuV+1JvU8aQHnD7jp5x1h+oniEf4ic0gg1odr3sDXBp2mZnbRKHjczartv
Iywokicriqhiea0gNJR0uwtazsqtPF6X0P1aJV57QUUXLlB5x5BQQ7bFJIahq7wQ2/HPwtzLWyz5
RguAmt6M5P28CouVh4ujdz/gTpfBjl98nLwMGRnzghVbLl/TK/EIDKhIzdLypccJTVpSnDg3Tfk/
Glf2Z+HBFy2Kxn7VggwovyV/59ny0NxducR8eXFr31oLplhuSs+6lafhjw041XSFF0b56J549XLi
q5PE0ti38SfRNPKnOusRqal27QxfZGJpvHVueGhd4CJTodUJ1yQiavHm0xnupq3z9ibbj0dD4kGx
4aYNgSbYv1+ezL+G2qkR14rBQviOxxY9JaiJDQ2S/i7brDKjkJIZE6vJ4d6iCmYRcncRQ+xxBHov
Xfjkp4n6RVMdOFOKMeynFT/A2hfdWmjRd58aPZN8mRYiQyVN2Lkv+25OG9I/Uz8nHIytX4/6UHdv
jEIeHDGVVZMUrc0lV0Y2ln0MhepcajuBDxcaH/wg67h8vvTUpFIsRA+EQJqH5MJ0qEqjO8hd4Fa0
hWPkA4mnrNl87QTfbCSP0OsFvAsErbHBs9iYh0GmyTY1w0vdYWvm+6zLLuvdpwsJBCdAWq6UNUz1
uXVl792AmlnQg4wwgBml3ehRMG61DcBI3hIjKYqQljVRFDaVa9GTBjt60Uhtj6/SYRgtA4H1uCIy
46aUBOzYsOO7NUiL9iXDGaktFXZWXy27mYM0OJMaTHPy3NGN2X25jQkvgulAlRof1MJlpWXscVoz
Xe38O/8gaZC39/poXNLcJA9RvISa0JEUkK+EYxVZGp0sQlwthfexARTXgljEeZpEFP6Mhes0kFl8
1m0CyURBEVnDXOwib62qcti8LWK8CaK9WyfoVnlxWrXhB4eF+b/EAj/znAYC63dPIr9nyro4uRLv
KnBrYotO7BFZcRirduEir1NMWkuePjQX4heV2KDb03RX5Bm85tOsVZIiMI80xeH/x+zEwC3ntAQ+
Vl6w9VjPfOGy4qv0osjupZfKIh0+6wO/p9F8B2jNtzobjoBgTQoMUG6WtGJ7NyXDW7GX9dQJs/9n
R1kHUi+oHenqZPmI4Iwdex/diN7M5xiBqpMVqSy3siYMpQ4K1gehJu4KensOHoXHmLzyMRS0ZCf+
xvWoqpx/1mrH5eQxwxMyONBvxM+5IOHPXfv3CM3/POE/iP3wY0g4mteEfkilcRDskHzu+T+061ik
JeMSncgfhhOgl8Nitji/UlT1GPgspVED4DDjXmGYxEaN40EVNnVAWKSEdw3m7cT9xlHluqBKre3t
mr3znN/QzjtZauRYtZdQ0FLzBREoeAmNtd4j3UD8yUzYf7hbaDchTm/jKOu374ab2Ch22Jj8/CDL
Em86+0axeM1Fw1gmnJFCn0n3LdSpiDAC3QbSmZz9FJiv98kSGTc8AP0RTXxT1oDSlSkZBNc8uDLR
L5dQPmJf422gCS8xDNdIb5Sig00kmLwGrMznPve5B3i9TWvBeGqNfAAVc8d2GIsJ1qO9basCJPdG
+ojrgVjzfQPfx5DFoM01abHqXnq4Kck85boC8erIYVHiFgIlT7YDFICY3YqZKehB5vF1UzTClMmX
yAzU3Chl6yLvg28UeZFjvU9ETd/sf+cg4I3HI+PfTexbFdm/qjOZvhPhXCSn/EHb/yIXGoXGKnL5
hbd7gjScgLgajL/yDC0Pj2fqPtOeef6HHG0y0YCWWkCA5fnjkv/x+AmgqLDilaKUH2/phzg6kLfT
jqriEuCj5NBCTRc6DnFJNxXXu1M+bCSKBKgR2q95uZ/atDjBLHWeZPg1mRx51GJfVOPY74LW+Fx4
FEKW97gOLuyIyJPpxxMehkoOAHt90DP4Ep67ylG3gIRZ/CCCVE10L6otc3bHqZgE1+ellugGzc1L
umzXoLZv4bOKIt36opwV0LRtlKPNA5vJqqNb6USGFWcWLJ1IpPyOXn+rPueawwZXJIwo3ayGR47w
Ov5UVV7jOq4SMKPX0BrslarMelMrpYFdozqUWIIi4grkkYAeRTg44OYOgAdO/6LPXGaXqPE0rGIF
mUV5nMXNanWchvLpdwJzpJ4E5/Dm1y/5BQrQwOn+IQKPV3CLSRXtDrD1hd12rw5r+vOYXp2ige/3
hnMgOcS2baecvQHXkp8TVBAVZhtIpspH7wcS4GYxTUwvGlRvYJyq5mynTdhu10WF8SrhxaxidyLG
xzO5mUJ4A9wfeHMHaBC2HTo0azkB/zW9o+Epsedh5ghchpwpwsTrb/47RZaptcowUHinKCvFjhtv
/VdZgIv+UvUYX+Ed3B5b3yQqnHdCzi9cNJMDxVXHS/VrZ/fnp4GofekXplRRZKRmX7r94Z5hkRPM
9RBNQrV4CCfnBg0vd0TMFMOmRPuhzzYwPmvFSd3QAudmpKIKB/PAeuWNZvh7O/V8APEPYhEdAUyn
tITVEvVW69hoIiV2PS8LVtQK3vh0aJZEMpOItIibfhCmBKwGuS0fobChbhzJe6xsfisjj3z4ybH9
KW/jOkCRbXG9Gu0ujeMXuI2tiqJAA8rQ70X3DQv76XZFATx2c975TwNaRFZ7XT5hbHvBmlT1O+HI
Q1gYnxq+6efELd0nsIFJ+iRTQwrBjFW6MYgzamMoCKeKyddTw/D+AYfNy1xIR8Jk5446qCGiyzLf
QqTWUpH1W1bavHFIO5BsxZCPnFUbTO14rF74AhutgAjuAbnSLn3IGNpItVez5Tn3s7foXPoBJXXp
EFuyT9bdgYPp6NrTniTxG4PQI1j/LYtbluiNnN+4R7dgyvf2WGqzQuxEmvzdQtLiIuPLdzhnacoA
+yKgekDSScQzmYwRxIX1jPnK95Ia9YmtsKhR846Q70IP16/2qjHtkWdB3aXxaINNqeMbYK+/ENsr
QlQk43UI4KPmVdEOMHvyqlT3C9vsalfQtAqoGoGhnAoJQafWuReE2feJ/HM49pInJypbW08bRS5e
lsu5tCnGKyBEYGK1KQ/xqD0OG3q6a1sUGtXLFNddHGilmzHrw9I6d7fdBZss2cN1wI5h/86oZkx6
XQGMC6xfhSUWFlV3BRvK0n6LSk6meuixVOmyk3ohl1CND59cfcvSwqwSYr4ZnsDk/SE8uIaWf4qv
08+yEOFhHONX06TZDr+lN6gQcVCFDQp0OE3O7VYDTRNdRHeqlsuLcbSzO6ItkUB7DoGcDrzR3Bs8
sD/KOxxleIUXLe/p+ZNlKyLS5hbWuTo3bu4+p/37H6+3uG001J4BbJuRn/7QewDycuXQIXU1z59G
/n9xKYALxDLMerayR667IlmURMewCKWuG1dH5+A3QJ2lXtXe0VryBB4sjWnTcARuzFN8iRqnzmEe
SLdtcRtoRnxy5c9GfEKFMRgHynqCjUSpzUXMNXjiz3qnWMX+fgZVawSuhfN7N9Ix1R2RNSGS9iNZ
dJ1YENNyNriMbJ2R38JgGaiSuTdId7V+EFR1mwNIX7w4VBE2NoEoZBkk9CuIlpCLRWPlbU2/WnJg
g7/Ekx0AJR9C0LMjpjIPqyeVjuA9qNRR50LL0UogO0HiPPaL8oPcBpM5miK3tuy4OTQr5vzh0Nu3
G+236eg9o/ZcnqZKxzRnX7PVnpCr1xvM79MnXTmCNKRA4Fxwd07Dwpd1EV5VfnMsefV5718KxqKK
s7lr+Q+YW4YhH7STR/jEOdoWiTumKdPjZhWwvul4ep3uVwpygWFSdR5C3k6/xgZN/cdvkO9y8S4D
VNqQP2yZ/gQufMRyBe2CWh61CIxAgvmUhAhk3gj7onl+yVZHGKyXHmOYCax6m9an4FnGGiX7ljIu
HG5y9Gem7kUt6tPQYng4AQy0oDFSt7kHVQk3WM2Xk3Q0FJMwAOJkGp9eWmB2rWg7NNCQBPvjLkCg
XKIFWxfOnEPVkMyWSihwplJhVPU9U88XgFKHTZjPUhpqOaiFeLgauPGtvQmYQHeNZ0LlSr71KRyJ
OXWYM8fxzq2m6XBp7Kn/EQ1TW7DdJRTlo9t7FzLuGuoYSyXQEjy24XB4FQvTboGgw7E5JYdv+100
MNufRlfyAPXvEmls//RkQ4H+Dfm2Bjp1hCxZPhLj/ZKk5C/iLzpOl0eu56MVbe1/22GR8jyppRj7
7COM+GOLNGLOVf1uNcEtASwb2hyZAqay2HAZZ0NfA3NjVZu6wztfRLZEjS8NTaNTh6yn2HZiB7Hi
X+eBJSaNDorSclBtURysfFxMb8Tl9ZGKKV7KWUBhxjK8UoSfReS2j5BK8YQTy5cwrZ4KUII1fSNO
s4OreNoW9KoffmYv7dSBidfD26UX621dGyIOjMyMxGbnkMbmZVOmtgHQCg0fD6b7BN+1RbdtSvSu
4E98k451mUONykNAjvY1WZPsoAChVlTQjsImQoJUFlOrf1BhlxiL9qaXoxiLVLVVY9B+ezhMvFKo
bQdcHwu2mkymrvA/UTVlU9WfNM+jNbeZEc90en79MNQeKUKUFMCh+tos7Klu9OSqSFB13dF7je+Y
X9WQ60d2pU8CL7rMu4YiOD/zpQUcWeF4pL1izXJSkic1JCInXfntjzkqejzHe20tcJcZCquNl+UG
jFGptXPh+eunmmiUwbIc/cA7aaSIo3vbyrm9aiB7qme9BohM3uuwvkhvB+bubI62ObF1dgytoy+h
c4FfGZMjt4zbJzGyUqozNgaH7LLxwG/a+lETzl9SDatQpRpuI8UiTnkFZMEoFOvtJbFqhX0+yiwZ
l2QiKL6uPCFgl05ZBVgTelJWl+VK9aPOUvWH+edg/XwN3dRkQSBU7RmsdCGg/ImtA3DSHvaxHiks
gnORbKwzLoy1QmVipocehlYyuC08wBj+dAvursw0Jkv2YJ4qND5LthTPtdZ6N4nIEUe2OSXkZyMM
WkxX76XmgZ9OPVRFd1XlTh5cO7so9OYdFmUrEbK4VEsI0N855bvSdRiTEApniz4Vf2hfW6KeWTre
2x8WveycRD7gHLa6QgxL+nojjSGd4C95294BwvEhYG3c5MTdZOX1CIj5AhdncyPBPgT893F6ERMP
4nXN+ptTdOnfrQYCO/RApOwv513JMnXGM6OStuJWA4r/wwo0CwWAyhxsM8xulY8R7O4QOcoZ8IXN
ERbdk05+G+3GN1XFvMf3c5sctOwOTeD0eG20LulRwVXPV/D8PmRjoXT7Y2SSZlgQ5u8kC+2mixzZ
JitEelj7V+nIcqG0Swkkf8v+kwX6+NAWG/wmVMh85+2SQIzSriXH9aS2LwTiqiiCD5WP2P6gZYmz
7jYhR9PRyIsCe2gaGt4pBm3L4o3+S4v0JNIa3+VsIyKn4Cl1l/zl/ZikEDYfrikRFuxQV7rPhyJ3
Ma3zpQXeugBChJWRMgGwHkndkESSFuEc3B3b1GSR+6Hol6qCdd9U2yytPQBq7pGF7olcuG/Hutzb
CkHC7mVaJOwjOwbZOqEB93dFsYHABwujRH48eLMhWDrgG6c7xaCpQCyhmttNgdmAr7s4Dpi8Q+LC
X7LntYIczT7q4XL5gExTQccYJ6quuozUBgzsgtvy8v/PCJwvWg5XEGB1CEbHMADZbBwEKn6gZYvM
5q/q4LWgOJEeVzA696/kYSaUa+ASiwmNVt8dfAIg6N6xBBDUszQPkWD/g37Nbv+bnnl0NXCiMB3P
rXFllx1zl5vG38T9u33Qt1HTTgD1dv2MUmFHRri6IQGlIK1k+QBc0eKme9K8LM+21b3LnPq28iPL
VIZL5p4l2ocHPpvLm4Q9liEDMEzJdQf20cQ/4w5rvOb//XdD3WGybt4FhZqJoCS+monV/GMi5pVG
Z40Kr5eY2zbZx8YeZQ+6BDZwKI2ZOBnISEBSs7mzshhuDp8QlVucE8F43lC8ofHR3ht/7IK1oVro
CJhssUu0i2mVo3hJ/BVaw1ioVo/JIuc6bsnApqr1LX6PRkqZslJpqwuBppA14H8R7DOE9gY7CxJG
J8Drg0cFhP9z6hTb32AV2IXo8giWlPIz1FDCvJXY898p6CLjtXSWSLPLYqNskNgosGqzf8w4pV2R
64vqjx/nHPWODHw7bJsK1pB/MGNj6L9kBDOUK9+KNDLNUX9Yd+pQRzDxsY6rJw2N0MF6TpQR9r2q
ygRuRUhV36jHBufrIlqrbtD8SmBsvuQzIRlinKtnciyY9LkPsR1DlOKSTH6Xog7koTa7kb+nToyD
fGbwQtc83wkkJtA9Bso3zkKN5SHQ2rRcJBC5sSdIqm8Y7y8RXYeB8SFORSn273f/JG+3+7xBmw8j
/bDvPCACcZ9uElrCD2LRSmq1RofUqQ37Y+zADIDmmsIEArDLBr/buYsUyyyidGxDKnyMPlMaWCnh
fC68MswzvGH49mwXBu+5B+IwoD3Qkc/LSxLnkmUvz6qlDti5282A/x5bcX84mXRcak7FdYwWpzGj
VGAL1j3MWlFKWyMqycZmKGNZ5+vP5R/R0C5wM21tP3VeiQfJbaZL8IFdgThkP1tqlMNBGuaPqjBo
bUzq7KIdl7X16rdLPTLBl1buoxrMNAljK9KHlXVQI+d1rf9e/GdZtVGNpmBz8qk2TmdG3ELf9Yn5
TcAWjEHPj8oJDtw3m/gfsjfwY4P5M2cTqcpYAG4CPvvUlfD25JKfc5Gyj+mwYJotJaWGApMyumgl
xV6zhLiUjNrovfiERfHOXFmCrr5ilbI55nQClUqFJy602sB34RT1VpAH60/STKUZV71ZULFEj8qV
IvGFmeSa4/DXGEeEf5zg1vxbzZ54xXA36YleTgSWYlbz0RfikvNmLRL62YeU1H4n1DL2ezlO8YdA
KeHMnCnpyYHvCkfSvzygf/6ho6pvkuNapkfQNjxdkrAY5GBX/DXe45Ml1VO0seP/FmoISm3zPcXh
7eTPjBRMJl15NIQiv15XjoOFTvzezRR75YdEwIaxGlqXSXuUbQX5h96HnUapSHZE3/T05B1qSBjQ
NPDbweTfSNYdS3DoT2kaVIjigfQIgqts0NQ5fXKSbM6azk2LJVvbgbf6AtvURT055hMPgG840rMo
WtU1DzTOtfGrZfuEGIuuuAfjrH6uffXta/aUJ465/km0TeNahZLXdsSRW8pIKk5rQpk+jmnrkTRR
xx0jfnFVNNmQZorhmWP3sURye68da1xPebRynefChibA81tkzraqjltqgNf3lYzfk/y2nzxgRzIX
8lrjwmLGrrSRVBCYnS96Vp6SagdHDNyzwPalh44IdeSATuL9r2SfCndvbt/rFcNnCcz623ItchAG
FCAsB+JsUMznIuBtRW2zg2HT12h9KWFHTepG4EjFqWJdlINm3ZprFwCDlmW32Ymc6pO3LKDG3fL1
k7Wues4gwdKnihgJpt55Hme/4wbVHeQ27pMzFxmDdmcAGEDhxh27U2Xicj3YR1usvYC83wu1Pa5K
PCi+ps7dWybFrl7qjhem0Bt9h4ea2dr9SfABgdKCYmz6s+MrTcfJzkRe2h+F9U/qoRPyp9AnwqB3
4hkMmPOA+1peppBd7yJqywEiesCUU6du0aTifwhqDiCj60swYyJNqPj7xNqsHsobyaS7rnIl8zhx
XtlpKL5ldVS4Qp9lhOF10gbmptMh4GtPcfl2PcKMr12XDWeB8m4b8Bg7cZTQwp8OaIJo1oHUgOwy
JeaastN2qS08GRDSS6Ifw2DvQtDaUeNLvcrgDod2ZCQX/uRifhdHaNl9yXDq4X8Mj3+7uMMkbOpW
KDTDIvHzLlifnsJ0avFQ2i6R5Ajxx4uoJB47Mrcd6Vl70GVboB/CegFNrSwqW2v/L9iKYCgdFFnO
VBeK7RqEu5fE7EkXTX7xuqB9uC8zOpM8AJjEsF6g96JdI1O+ejJYnuJL04xzyDJ4bMEqJbYj7QDf
gM1Cu+FBE/kC7YidHzCbEG4uRuwm9meKiS4nqrh7wohkcwLFY5z4T299lMqgxWn8tPXOdMpADBgi
uPe5HuYwYi9WfVgAkbSwCOBfUt8B/NuEdVgVNZxgjXKftBz3UpbFiTNr/sB3mrUcEepDDftFlKmx
8YgNX6tWIau6vjSRbRW8D1xo1EVZRP6LbdPBwNTtyTaiY6JnKh/e7HtzroLzIs5ow3rRpc+J4Biw
L0LHJIWAAgjHBe+C469R79g54sL8EGw5obOqCvHx0eexBTIBh/QsF2Q/dbTPvEBLJNn1IjQWGjdQ
xacQmjk8IMfJAu5BkgsMYIZaet/zWHdH5nPvwo6XKdX6CwIDwe/anr6MkPGqmpow9ufPxsQzaW4q
h8aglmJijNkCPlHcUcAR8EUabKIjmbbYtwHjc3SVmpYLPSVzg7YI5IAnTTlVLJBIkyOVO8pKNeVT
NSAwNpLuPLDKYlImHimtHwly8K1EAluX7N9T8mJ2Q7uSgvBqD2yUEuEySNMtDzrJ3pCOHirrfDND
ANEZEgK7LPCMHvZR8q0Bh9Q2FOBvM8s5gnL5hl2hQ5M1ZhDdlLLZne0OM9U5HwQU77omwNF28Pvk
oZCJPBBAh1zJG27J2rwdQN3GZu6AJiBYhE2qm5DchxJ79u2DzTaUWc628lXog26n2iCf5NIwIM3p
GePgINcWfuE3HuAQ5OJ3rxxhB15gR05hdhewzsNSwdflbv675KsNXHDzEhwdsKzH21EPGrEge3cc
ZlzT6C32DPWHJOzhf5LBEfai1XCZkPvD89D+ApsMjDXbZz99BkglrK5xkOGbuUU96QHECnH2rnfi
B0VJumIjiG6Z8Ss/jQ/dVOKYAQFvspE5V0yL0L5DUAJM4Gw+BhueAIRZ7fkTjpq/5WGMidSEm/p+
qtriIj0rLZAFMj719xKd/wN0yYKfob9HvmmE3m/ZSpJlhymvQZcWmM66NgqrRZaa8x7QXhV32gUN
xF2LBBDyrE8kCuS8CG8urWgHB4gSTf6nzqaRjLEy1i0Lbt5VHXppU82ONApR3lOuQR5fE7MU/1hr
o/Ka+5r0aL7g7v8Ls/d3Ww9CRhCrBPqs8+gaTx48Ex5EiSUHedJK3C2ECrNmBYXOUlayJAYVkPZJ
bC7Jpu8j3OW/svVTzVzTQV7q6hUGMTgFxLZkOdICjb8n5wmxLuwKkY5pgXem220nS4ihZkzZZPwo
uga/D99cIKhSwzdx6xDcl4SXVFMWesqnv6iMdAYs2d9uoT65GXzeffmR0Q++WHPoKHjXxn1Q9U5H
HMOCQ3s+oFWUUszFq5qfsRq6HxGjBkMcgs0N6hSRnh6v7+yaJNiLRwV+4wzFjw/3Pw1jRNMP6ggK
VUBjIp4G0CqbG9WQrfuSF0TUoZqe0UTamPTW0y/4XR4oDs+XoXwSqH/EaquXU9geK0DefwJ4/G+L
QyBFQwhsZ5Zn6Rm0PGXeBJi7wuaoQ4VryC7LjT/psxNtd/+zpX8ZP8AFzYjf81PfmsdqSsCTDvVz
XGLvzxkBjanR4J5BuSVrOaZS9RjXHpNwEY44/sHEEQN6bgaq4he1Pg57oZuIBwHZG+P2bjoPhrb0
QxDoKr6+Y32I7T14ZQuhOuRZ+vd1LeeOYmykiRJfR7WmYWFcL8QF8VGzkEmkPeq7148GRkx5Gjeq
UppIXJBRRckbCoBIjEXeZeQ4k6WrpOkKcmqUC3NlP3umudPfSqGU0c6lQzFn4Hl1+Vv7cr2QfaXD
hMjccqocYlUYOYK2GwR35xQkabtMMA57HxcpaXCNjP3uIIbEn6BeFxI5HhXS1P5Ay2+/JImCKF+L
MJrdKToLmNNp9w29Ma4UpM+apsf4FQc1Rpmh6LO+tb/Rk3bAgnCA2YssYAeJvDM0VQt6ve36Ewj6
f0wGifaMRCmMbaiQv6AWmq/B9nLxxo9vqnK4X0mFPUhP/Ht93P9Qg9lswEwTZ4+u17qnOpiwAPmc
23+5eBTv1VMdWc/4Lm0RpRoTpce95/MwW0R2FHRgOJ5p8/Rhtar7fks36Rqfn6fWC5zZc8b+Fh4e
4FGOT9sPVXTRmT1p/u4B4otyEPND4FwLsJB2w4xsS6sF4ySyw9kZhH52Fw/1hzbJnMbDCUiJwFhu
Js1csf79dNS8t4L1H9vVpYGiO7TG5djn+HGU7/faXYe8PEYrbGFuyixDSfPPEV5TuGMHQygqWpWV
gbOaJEetBa3JdFD+BMrnzUivHjSxoe3Fy8oVlWiBivYe9Sk+aqHd08boTBeJvx5R0htyNc1KsTZV
fFaghVudRjM30Nxuqz8IapqlWuP4EcPMaGtTGTuaFk+uLGtULto2kiE+eFBufqKgSA5BVGntxMwo
AQcHCXCwcZ1hHDQrnwWRIQ7QxMP4BOLudg4but6AaulyjZOBVUqtNL5h3jo4HvAmXPQGKkn/YpB6
gzEG5zENxGhN0DNcV7D92x9ashXEnT4VF7bx6t1jLV2axJ0AWY4R8XI/WNW7+JmqyookBr/0R0PK
hR7KDT1qrsRz8QU8BSiCYLsiJWC9sKcZgPuRsI/x3BO0Ks82SG07hS+2bHMIM41fTLnngdyw+eUr
2TCD9O1zZO+dwHzNSrHtR2cNuFNiKZrJYjGtoy7agLmF2PBDmqbTOlNfscFUEoiTDpzwDRv9u+P7
8pYeXVzwtmM1RVlvBInJpBLQJv3DLNj1VKGT3hDJfSin6ac63CgJNOq6GsPC4A7EWI87RPI4oUrz
kRExloxfbP3FBTNjSR5HqwpIvnm9hVcDvXmSept/DUSbTJcgyFeanws/+J8NYft/r4O0pnMJfLMq
vBAUZIZwHIBYXIr8euUBXMETe0pQLyjTXrkFckLgVdgvH8a1P70ocPJ9RLSXq30QiSOaAnWVlpmG
hMD6WUiT7QDgilzzVhzFgKychUcbl1uFZ3A2U3d4rUshKCb6y/w+IujBBdbXjnZf894cN8P9g4Nz
dzWFtWC0Q0UlpKtM7lbbR+8+mXHDmsp6KsdTjJ5JA7+REUo2IKJEV3+dyx9T+bqcaSrF8HnX4hLk
7PU58IjwQd/C4UMPpOGxMDMQ91YWtoTMf+1agh5Ck0OMo1uOSTizTxX00xzHubyvw0CQo3j0qYaE
k+f717gIw8SGGdtXQ9gftHVD55XpNinCQQTV2LO/vPqtc0Vj3idxwYuVCxaFd9Z9K+SE4k57OgIZ
F6qeltVbfgr0IGCJ+40Olfe6OdA8lnQy9/pra12VxRHX0fk0j6Eqc1BPy0d0ZJsAVCGR5ZwHUhJG
3zqYBouSPqZQdy4G77sltwRefPxhp2JOoClmVAGxbA8NE4WlAlJUjp6blSe3uaDEW1BczkEGrJr0
0ZcKdeT4M4bKfvABGo2Eb+gwtOqmWwrF5Z6bOwg+YUXBpxbO91EhJdhvbD1Gm3w+rHluwBdFvVax
/+krsiObBVGcxAsIw6GLktRbq1LDrZ8WQbgYVvuMTqP0CC0C9/JWxLmFy5a5S3/58i7LTJFLdXH8
qtRRJtjIzVDCQq1hbIrAyDQ234pEUz1GezPCLhF3l5jJNSEwHgFfnlmaVuaB9w5H4Mrw2jUgFlG2
hKgPXhaMSmHWOuLrfiq+F+IyUHhG36OmbxrvsJkJIkkzJ+BNUxp1Er9dN90s6osxSwmPhZivtnpd
nijqN+DTpZoXv+P60WaAuf7pA7pXCDYb/Qq9nWwfxefWnZ67wf3BL04zqt1pEQs7rjEjEUcAxsL5
GtjUMFmhHiWCbVpLU7OwZX1pybV/lNnCe59n9POY1L5N4T4ExICTvKVI9eQNXmzsnzq+rCZ8kgw/
aF+MClKS+r4kXUGAr801uC5ZArkx7u/RQQQTtz2jyhK6JepUD8im1lE9rui2PmSR40tUDYfSg/pN
h5pWps+FdPR7CdkGp9njNvlakownha4xNs7z9hrsqjNjeMNYAMJlOFiaIxsFQ6MLPVSu/Mad7uBF
joX+1P958akIP3noVjCrGx/OcYq7wkoPA7m6yNrOjr1YRoxf8CHn69CojCs/fN/kb7UXQLcktuzE
IzM9Qs4016Wgs7mCIjk+7D1wtLl2fgWHa+wERGkKqwl04N5rJz8d3tGgrPSr+PzuENgD93aAFPtv
qJgVUOFTz/oW7nymLmxkbQHNwKUnhmuoZtrl7bdsZFMqT8jD4ObveLzEF7Dk/XaKD1DoH7TvYdkT
tDYf6LmNASajDfw1xOwX63WFP8JFGVGKy1xDpO56jxNQKVkHvdPdQ3uH4e2DkjDU0MoBAo49sATQ
6dW80LjvLRDLLTNjs5eWkdxKSjPM3iB0tXiNe/zI/fIPiWBvjy/xp+uXRfTT71Pe1VjGGa0MgBm3
L/raYUzsImOQdixbYsZjTsgLZQQBtU/AA9jpsrX8Brc/tWykwzeReuJNGUr67VMmUWGAsDQUD203
aCXgfq6+f2mryAEE25sfq2YIpbpEUJjCQMOUPjwpXeHpY1lWJJPbXrVhrrnJcM3oFZaUlooVsDik
E2pLV4RWQdrSxLx3gfN2LPWxl+c/vASN/USDWUFljRT5yqdG7uD/jAB3/76MwgGRje7a2rNsE/Vz
7zyPpFBIm996PV8azW+GGu3AvcYYT5dJBxOnPh01fNzmAvorFmD3UUu+Po88z4+9t5pHcEnnyLeK
9FKAsSOfGsQqu7fnhEjSZEnma3mM0KWjDhBqO5jvtRarAqlZefJKqXFakMXBqYgF5oPSkdgh45NQ
D6VYqtw5xtGinEISnhdn7Tyb80JOASrZBeKmVeKoXRa7WDu16TW4gMrPhuv/uIwo5edctJE2ssyH
Zs1k6+BRiBb199blJ2pWhbhGX+wXA/6BTiJEbEQS8QqYdRAU9KPOWGdYyzAzD3Yqvp3fdlPTpQDH
yLHrlex0bkDEgK04uFK8at9pMn3BvKpvW50sgiWcc6KaxHN+EGfC8v4UBNz5J3QYYMSbXz+sacMY
yCor04KpmVsXKgL/lAix+fhFc1WKGZSwwl9EnDfYZpKDSw5ygOXk6I48qabzzeMM7l9tcYEEi+xY
xWYrRCc08CSUWie0iB5oRUZSGKg+jKIQOGhkZBA9iHBr+kiFeEBFLpSH8+q5hmdAPT3W2y1qxbLi
cHWBJVk8BHZoBgm+5RII0mDJHPOEja7/dhvX2qEGOQj1kjnK1Knu3FnJ1rwUl4g+SxV6YOgHoXTG
C2RUKnBiKOyHmB8aWxWS5Ob+QkTBS+DqKD/EyZ4v7aBTsOGj0diGf349BayQGaPQJ2uGMUMkZJ5c
HV0mRqMSaAwHdb+04jdp47sHruZ3jLtvjX+tulVb1ggzbK8gB2me9GPcPagRGBQka3TaMsAU2Hbt
Ad3W9zyJUwilUzzg9TxFvZ0xCd2ADqTxHF/9iBSEp9iNcoQjURPQ1+PtkC/q2TZEj/GaMv6G+hU6
7rEx1RxS7IDBrzAiHk2DxDd7Svr0A/uGNt2yea/xAr06xpJXBmUP7GMlRz2pcHnncbG7DM4UMLW+
e4mMCLbC4ZQK/mpXIJawH1i+l0iiLMiRMgCAlftvJ47aGts8Cpe6ryHE3uj9gSLaG1G/6JB3OMLb
aywm8mTxSzHM979TfuWXXLE2eJPs7V0na/M7VAlprZ1HDt0ef5OVmiWRDnb+TH/ogfeZSPBIN5Iz
r67Ewuhfm4h5Rt4N4doxaooMOJX+Umr4Xk24qbf42SgGvAM7BVh5kk2vceoP4ucBvR6+wH0qmW/R
yEk41EtK4sbD7CfnOyApCmAJOIxMovGGYXLIsKMJEYwVngU4hWNbPj36kl03EP8BPmTfFEfRZ+eg
VDc2AOOqJfkrawOsBR+PEO5sMsipoEWu/NONzZWY3WgCjpjOQSpkmprjPzIve6HNM7SJ7uLNkVhW
5zglCUlqlCug4cB0PJacTY+KkA2CB+cB0Jsr5eqA6j7pIcmjciThuDK70bisvYsb+6DzgaAjO4zp
k1k/lehE1aUMpfl1NPkJin6hcGtnzFIAvPTs7XST6DuvRd4hGA9gRVSNE78dxg8Yujurf4oRckRd
nqKRHtnqJH1aLb9XQdX/pD+grXXE0ACF3HcgWMDe8WU2YoFhNpLnBDTKdUFxkO+g+mBbq1LinmUC
RKDiocBhJn0RqUKeum65uMR75PFnd8bDuYfRCvkDtTClIwscMY5OAUlq8aEMGRE6t7kGUfhkA5yb
ml0OIwX+sA8SVW8jF/NX8TKB4N1cNgwO3oWuYAZKEFjOoMuoEPikqp8NAE1tZkBmXYjUXPwiLjTp
Vd1UmP9cFna2qE3LGN8+PhJDpJNNsic9zhPHwBctevqzgGhEmqiNL08XtAZ/OWvGYOvF2I6jJH5d
gIslOjNE5+OxguY6DObakazr9A6sbr0cAw5MaWDtxlih4oi0VHc/DSD9doxHWM5v6Xu99yLUALWY
ntQvWeYlNCWcFz84sj4b4i+2r2BFMMjbS7m3Yf9cLaAPWFFCCcyL+guVZOIqagvnE69wxtCRMfGS
EpWwkS/QyjIZM8Stg17t9/MYrLmPQSuwU06xhSyiN9G7WvtXUoTq+G79aWoxiNaAZkupNmGkhva0
wBZyHjV7zIH0F2ov9feP5iT1TpEpQ47f2JyLJCzfEpaXlpHcOBGoRQ+wbhi04GtSr0E3ZjfOCw64
aaJMrw40RrZ6g0DB+pXJQQvhdW32jcqHsTzBazMn0OE3BZNwwXHXsFlbuP7YSgEPNooqgeIJlnKm
UfyGPoKht2ssTN7pZoRs0MhrMrkV4hYgiN20RlFRSxxloK8RkOJZ3AGYR/YqRvlmc3EQuwUdKCeL
YMK3rwSEvDwn1mP0NC8YhBHQiyTABSJLuiWPiLkBOTlombhE9vzTXJZoqbjDA+3tQFe5f0by+JI0
aD9wTYfhu8nYO4Wqreit4ZfIvEhqcqbGtlQLArx/DUcN8AyipMKicG6XkBe/2L1XNMiqqfPzfV2A
KG1qVLPzHj2rA/lNKv1kidwZJJiqEnY6QfqC+dmRhaet0zvAVoTcycDEwq/TWcRHTAPoaO9KnUdy
eRB/7FSKeT/Wj49nVf57fNWq1++Qjf/zE9wWVNH/e2M6j9MfvhCJ/dfwdXeWN8ClKadQLf0Rp9RH
7vUPJSPuRn/6y21Pm0D8dhyxb7F5eDPiYlbVfn7NiVz7WxWZeFgQaaNgGVEOvSwwcelGhAwv1ms0
h90CsTkZ79gIp1j4rel17hLTcxAht5NQmEdFtmzV2idM/flF8qkpTJLgONrKQODCYB5OTbWQ5cU1
YbplCv4NF8Bm6vHpad7jOtV0h6GHUb1m9H0MUePawY2Pu0TjQ6m6FlYntEa5yyKFi0DtkI0hhumI
YCw234k8a+uSbk7TnuYWYn8CeT8JKIJPXsLfFKnR91P4uQKIgLWQEKMzF0NQ0yM8Az07dDx7GPMG
/7U5ZNMQcKNL9L3l4UJVRuD0NpgGTwIQtaGXNf6NmzRaM0ezcP5DwV4B73ck6XOG86+6nxd7DFut
nfTqYyWam1vh1a3iNeP5OceqFFttt7rHjLAeDG/IDciI4GyOA+cw/3rKOc0ImQ/F8coFL48NmDWL
nM2lmGjHFB7l9J+trE4V9larEZA1XKwh+6Xy9j3I7Wl0Cr24et8XT+/KlkjkpJWLLjkGcz6VzY1K
3U2qPmeLMYVMpB6zJt7C2UotU8EeHtBzDS2hLeEGoNTPELPDgJpIvr+eyp/SV6aHlwgJ+1DwARyq
FzMNGq4CHB/4hzTSia1cJNHT485YTYZwpouoMi+aYbhxOYp7u6MrbIYXIjqJKlVuT+QiFxuEqdeF
gPggEQcR9iy0kH/54B51zsQoDQN+i+c/toIgyKSU/rd6x+hM2K0GkO7hsszWKOucF9Sxi7sStMHE
21sOnEeYJzcZqwJIO2o4D4Vxiz+u3T3OXURT/YLVblBLDNT/rrJjPrWmqE6f5+RuDHxpRWvR8wUP
5TSp5i15VoQ6nTJtw2CY0GfJINq88mhPwOd/sGxW4ievBBHf9dVAPpnKMaR3jdk=
`protect end_protected
