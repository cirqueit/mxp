`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7104)
`protect data_block
N10a6KKWT8TGJsK7twucU5XABlMELuyN1CYTMFxQ2FcgMQdQjn6zQGxmgbzblCw8kDYGsEOa+bW4
9xZF9tN8wxuJIY+MByfds/AaC2oXUr4kyw0/W9w0VuKqGYb79qaJvs+XXtwKwFRtilKgyKZqU5EY
YTqqTjTlB9iOkAzjELCogSSOp3+/cd0a0JkE0RBOHhGdMPiThGPSiZxvCavsKrqhca/bKx/GmZrc
ebQiS5AhGUoozSFEAG6DGbi8m2Cy0w/9KjrQq54NW7p1/IdiTYOZz8Em82jsvbLFBATM+cD9m0mV
NhMu/PIs+mIz4AY8V5JkvadC5gkN4ZSyX0EWv3eAmEzUYbFojjqqcl64IFEG+XMMfVzU6UaPzPGX
J5oe8IXtpKIacb0SovL2O7le7B3gVqpgBYVoVDra5JRNpfeZOIjnGMtMHxo8YIaiRs2EOuqKDw/4
qCdzO4k0g2Z+Lk+eapevnK5cRyFSlFGff7CNtFtIoRR1zGgZujk+r77VEqRMzjzmodqg1M9sWBaU
2PLZlhccUnvnT06ZWLeWmcfp7bOcyiMEu24QMjUqnwbm4qyZWT312okHy9CeJ4KzCrQsOzVFuCT0
4Er4HmfBivKBWVAfkIyg/stRfBq19NhqDrJ0W6eceC7GBjD+JloYUyFu4xYz9+pooAsk/hViXv0J
Zrt60pUAlTDwwJrsZolw4Adku6NlfRtokGwOP9n1NzimTRwsKH+sL4rxzN3VHUCqENEw3s/ogBOv
sd9Vgtc+qrmF1hXKpkFogTiqnW75AYx2pGFmOpS6ULCqynvDXnXtIiGBe+CpOGAObdnShrb1jQ25
FZ0Ozhlrd2iNv7Hr8NNo+Tl/ipFc03vXwnhhzSfFH4Y2Zkn0A4anJ8UTcW+khTAiiLbAJxiMLwEy
jS194bAkFNsh+Giy8VzVD3/c8LcaCZJmKnwuSo59r7HF1nOn26L++sz9q77lIeUJBZE+Ruay30NX
8vavU7pbzp7xpO24MonAKp7/Weq5ofJSxMn9hab6HsUXyYUhFNE3TJov/CHtnmIbV0nudATKtuND
6Ebjm+fKjQyiBzE29ePvJw2NjrRWe/3+K3wfS/T0tfA5wqbDQuOY1rTVYvjbQv0GhGauhWa/CSmD
LwO7qyisiVL0Z4sd1pwcLSXfzqsE5tqOcWAMUcL6Bwfpz8cwoqetabVOoRgTtcNFbAaiPMD1ZukI
tQ2QK+65LIS0sPLIgNfHEebMmttqZrJr7sGny6u1N6C/e5pxlDJ+sW9ItbexIXpAi07kTUzcSCFa
Y9AXqI0FteIRC70daT5KkcRLJIWNWJb4jhuUZI64wmj+EV+6Rkm6mh0saXAolU5ZjuTXEaDEhrvb
a6umDV1GTdjKKvrr+GamW1zmArU7GnVPtGWrclSgmCubiInxIjmVQkhdq+U7G0PZqVyVOEm0rTgQ
fpiS3LHLQoZgAbMylgHOj8EAXnQ545fRhKh4X6ioZQoMgjBchuCRTHnAXruf577xTC5z/AMSPzRv
YZOE6oekTIQCS8aUZxaS36BMcGbZ19GVgLOPPaz9CzkU5WXedHRYlOPjgu7893R736eAZxt5BQrA
y7bTPOP63AxGwYy/b3pxWKtUAp9IxANjIfjm+cgKDa3sbXYjktWRWIjUL7PcEx62g0gnH5VZVimj
1zuqOYbeWJ74riZNxtAuYiCxw81WB81tC3HVz5I3k+0n/fa89FRH7SSzJXGShBN20j0XIshIZMcp
pwxVGb4AdaypkQ3P5SmUBBz5MrNluadeQctYjZ21P39vkVchGiUfR+cz23m6jMeDY9DxgnzqLyUw
mgHh4vKs5ozqq9PQh2zf1gLXM6QXzBUuOsxgkLAg54x1fHznoEX9dS+8864pDp4KvJrpIs3+HS1e
l6/iRVLva6kgIZLd0/6zjjN9aVZ6pSPMBDV+eIuQ4xsfNSRdYMsAB4Vyi/7cnMrOHAJXo9M1uUOL
GCj1gYkw7mX8jQCLcgahSxJXFsxFYaAl1zMmdueqRfytfIRNWflKtI58WUxoMiD/zSTjYcJxif5Q
Lslb1z1nbuEqhsWarp20AbzkYuWF8343QnO3f5IIJhXoo3GNWMHPqjnXm5MlW2i8HR9JN6kC182W
T1SQyi35GIPj+BdkV/tn8vZDdH1JK7rfLEHyUY0wgbPxa2oG9BNs3qk9r9ebDd7lv6i1bkcak4F0
6mwJqsby2JIUdm3cK+fGE8m1tKpu3MXQO+zNJgaaAHuQuH6eJa3QD9Ew857oWY617Mh6thgRd0Hu
5Z80qyj0d9W5xwf/EYVY4VjRsk6Ryp5zTVNDehSmd5DvGVlez5riIV1+QCxVk87uiv8kvyG91ODg
AoYEwttQjm/5mlPYab8sBaAVkg215WKN9Ra0SBHAPkbBHwxwTaDqIOJYGRnIsBGV8uX/lkms/34Z
3jSlkttSS0D0mX7H9td015bzhli+JKgWRdUg133bUVfFCPXz7/rKqGzVMSpQPyItWvqlYbKMikjO
aN6/zgKIJ/7sBPOboXmaMeshhxIuznZG5sBp+E0nZ3LqlS4EHKr1gU7wkJsnveT6nrLXorHoEE9A
ClQ30K+A65iI36UAFhoB0wIJqfHS7jiLUwKoCqkvxdPQrUpdbCq/vkF0yh71L904ZdEleV1ULRey
TVa4vNdRuf1rUD1g6hYLx5Wa4kFbzUpYUCUaihq38zbnZ9L/0RtaU/BuGJ1f5UnfAjZCtRrk+6jm
SL667f3Ii5TDwTSogKPdhTe5z8dDENO2vqhE7GU/E3VvbGXaOHjUnc+GtsFY+ysl8Ro/pzIYQnAq
gAS9HyjTmmS7jHGFU+U2BfBK+/KGRDMTP5O3AD5OQU0cU0kgMN4vG+cautcaIC2KE0d0maRycjWs
Wzz07TqPH/Pkg/zfMlh8EHWcpoB51qmx+xHHGdMY0Mygi92iNJr+2Dtjx1bX+pakTZfsRy4Dtquk
B2DCocPN1RoLdmScczQFVSQAw7hoapojS8ss/sTScvSGD45/YZbMY1QnIlE63CUkHyfQcvzaaH9Z
XaQ1ZGLbwxeOKyUvWoItatztMkdW7l9Eh0cOhBTsZRjJruFSZLuVm8pwrzsDdGH3eu6aitnVQG8r
V+9MjIPgnqnR0iU37H5VgiQHjvA1kcF67ExIYTBIk4M2gsAo/eMmcSWP/pnH2mFmnbTvyw8Vqdjt
xomlkZ2FiZPgY7h6x+rhH5hELP0RKIgwrYdgz89BGELLKRXjM4I2Ymjgb/3lpD/dEy2WYecVzlQC
4JtlHY8E27aZlQgi/VVlc4fAvsrMillUeSfN7WvCc0t13Y5GZFOk09nMtOi4VjEQP1VDCHrqQSrg
u92MiqtNefD33IZG1NxJZr1JfUm/Y3F/vvgiW9d2S9Mkmkf0e07TmN9z6ZVnI092m2axluJM0ITw
Zd/y+CredMHrkcCA3pRPHJk5rjiB9eVD2j28UFcghVrw56xGCr3+G5SrhjIAbdTXDyG3LgxHfry1
lidtT9rxOMdnydLaFQeK9n/SXaqZBgURrO+qajHoBUoRIOnzRquUiFeiR5zzVGdaDu0fpef2LZKw
SeCsBTaNE7m4SvizDTVMRTcXagRIuIVpgDMRyIK7s58gaNnETnG6kzLbjcTeXUEXHI437PBQffEH
DT4yMuaVGGAQEgsCPiS35ybRVFfHjD/Cwvr3g1TMD9o08JRDZqU43mpJRnm62NtdC64O5lDHO+gI
KddNZ4FpQWEKLStik+3TiW1GUql6TagJfZxnLfOxzXqHFMrZmby/+EnAA+V3D/VByMWL6Gi+A9m6
7Zu+SvLLzkXQEpTtBjV9kHz+PRHPsohr5lon0QZQq5CZg8io+tNejGli5xlR6kmFynXHsbqogjfJ
UFqtrZwJbq/FxfMbrn28qxXHGt33m7pImHnV9TXX8BW8tbahu9Y+LN5VHB4rx3FqT4Kh7uBE9vA7
JTiqjwYnXdWwMKxTZsknh+spPjv6rqF0kTSmK48cxEGZUaaip3GDfrissng4/vDXzKNd/EglVWxO
AbLEAbMNdKtsxAR991pK9P0eGj05U2nWH/3CsJQVdXOCOt3gZrGv/aVkXYu3eDjWo0vE3zoJMlf1
xlRy9y0yIazPHXj5MiItFnruwY/xcO7bPKXAQFauAQFa6RToUkt5U0l3lbt/ThXaHgl4NFKB65ZS
3nbbiBpgFWldJLH12+Gi1coYPnAnMFhci92OivSX/bzviWquYTio2r9fjUeIukbaub8sLuvq3EGe
M6WS8qklj9IlJtpkVKyfTuL7ikiEJw427c7vvwKZnIWKBofgPrksOh9lfxKW6RGKtj2MdIc7UZ1M
MJa++VLszDLEIwqxP6k/TI9MMtGMjlk9ZabAS+tToASNnk0/GpJ1RDErmKA6hM8u/Y3m+0HGuURo
o5hXuL3geZS/NDRDRtLQQmjs1BT9vRJQ5vXznxmBrUSVj/iv3B23XN4cJEdn+snhUaCIxF00nqVS
B6RmFLDF0IeLDu/7wDNQQ4IijuzakgNrpkZHpi6X+dTOEsNHUwaNhccVr+fkhieSQ/7Q6hEEJc4o
G0y9k2VgW1CJ4iRcfehqgDFYeWowyR97yQScDYjW6y8sWsVctOQcB4DfkC3WKd82mWnoPoOL9TUV
Ers1T8zQdii4chkEGsMoLErjb3ZdguEjSPAFKUc7S1GBbMYIUE1BjSP7OXrfD/FegXm05G87YYfB
kz8qBuOZyEB4KixdMgmQIGp+r2gczeHqiV67dJ+vNMvZ7H/NwsA2VSs2IMZ6Wv36qnFi9o/LBn8d
inZ6fe1mXG/VIKYMqXkib+xXV/bC1zABL5809Xxzy6sS94M0bNFIPnaEpSP3TPj+FPxgDvRGsiD2
XHs24hiFGMQFLg4Yrh+QjMJI3kF6uTI8fhxIXcqnroAJNff4sS3Ml8xtq4WZH3DySvS2sWc3KB+J
mbhzN0ttV8NXezNO4xZrShcHWDwzGstu85fe9Xb26ATOgl9VJYgChqJaiIpHQMjBmgh6jteDgHpz
TeZV50ue8KOR6nWWUwOOLEKqfTmDEbK+t2OR5zKM7xsTOhfLoMHZVazO8w9JRAi4etqj3Hw+hxuD
DyBdshBfaiiNnHl/p0ST73Qe0ZzV4Ub/QC52bAvf7BfIKQqnfbyxRxBz2ZvmX6aiAyZB6dZ7GKpq
l07dGoAWF00aa7/2ZqhVfZKPuqrmP5ELrRJ3gIaXkprjrztXPyOkjvbr6k37onyYQijbT+jYZ/ag
j2JjfOmjU6S/VSLmNIHGNfKMBnwHX/Pec9i30NEg/GVt+kUR0X6+b1ThDB5WYhVe3jAqxkwFyTzw
tXrGy6B6Ld/6MJyXRUoBe4oRabliVO7CpJONPzRtKi/PqnDrdbtvyhuLFRQDpw5bqEdn0Pp9i86n
psB5cOoItG5GZVLMjrtBOfHuh4rTP4W6mvxGu1V/i8jNcaUOEy8dVOpUO6yfsldvut6Y3PbHojXn
juoieAVC1IY04lGi7QekPpOlDV/CVGXRJalH0etDP+Jit3U6KMy5fPgCfk8alHTHunXR8Kal2b5q
P+ifVpi/ZwKUkYPMywXYa72JwlmjSIz3qlZzkGMZ/BB/qu28E7mroxK9+bA//QU/tghv4OLbYPgs
Dp3fC3y6ASL1puZ/92KMkFI+w2W5ButZWUR46V5s9ioT4vKBmwZvQNhDDyw3dobCTzUNF9PNbQNE
6+vb1GjeuKGgy0neYfpd8vnubjdpqK2ZP2+Hbly0P2xSb8qOxeXcCzO/OlbL5bL2g3AXUMndORUn
nZM4AxwovkTBKI4JCCJc9/r1Qy9x48nokR1R/3VZR8Bs7Or3kcvxYRLppHEj9d2Mxy6wt6OaaI+T
CaMZTD/W2paDq3ffL/soqBA4CaHSiUoq7PyNUPSb1cRSZJewjMjC1xI06Z/js6giN0MBTewz1Bhd
RfXuZlKr3VjFEK41VvH/xtCSF1F3mZWT83YdEwnvC4l7px8GQ9Qtvc3otHwuHSsZjIKm70SSWeL0
yH9cZbMKMv1NVqCTUfMv59H3SjaNBJOwHdw3tycpLOxMv/I9UTNZ47EQ9nGcP7PvRZ6Wklr8UiQc
ENWK75GJ7YE9bEk7crsCOYHIFUzRWsv9Sd36MWEplq1ukWJXGNOhCEYUuRJjsEH+5sl56tf9c6PD
L6dr8pumoIkdd6s1jYfJR8H14c9+q4hMqOTGgdqvlTwiTfbCKOyVOpCE5albH6iXy0FWBUTCCMW/
sa2deWGwK6yBM4yddl7Aa3L8Q1AbVuauPbDvbFiU7hrXMlGzDTitOaU99SBe5MbNWGI9ESolCpM1
L16k1S8gsy1DGO1q97hNVCST1+F/Eewr42m0tfCnvtmECqFkzpzE8Hn5StnCVUdphY5YqWxRFVul
3Bf1lnDUhSBWJqIk3G1dWK0a5IbFJP1kIBlupJCfIG96CFrq/M13Z9mW961yitHHzsF8QrLvRRDu
WGLoS9AkMdpS1hedz749u52cxrezI64BPz7QYCe1DkUYq5JXMHdOSUp6hJW7rvcUqMmzzUHgzUW5
FOUnd6pL2jA0ZMiLyiSprwlrQ5c+etWaBiqXtFAuyr2F0570d++gpS9Jb3nBXz/cAKzksMQ8wQoI
bweMvQWqju2/LpUuFL/S3DX31VsSTvNVPhlasMmbmbF1WomS5Cw5BqWAhwaMlB2L4JfqplcRz8JJ
oIIUQI3wL5NNhi38zKTKVSIaIfKlU2A4mDV4BvcnDqU9luidIhhEoC+Ji9pKbQBtwII0KHdJq0jg
YiBNxUWDUBjZ/+7punM6XIF8h6VTun2VD3CgBINLqLsjKdJ14b8Cs8HgmvRybWzzQILZLkVco0Gh
ToYxWH7XnlTRANLMU4HTlYLiYj2lzky+zHlUASdZQk2NY7K1PkvRqC4BJLzhEnqF3hQEmyNVFx9/
bxZW1F5E55Q1KdpVytdxw7sE1P8I46J5L0upmgvctR37RwlWkPErPpKYsHXAXUjye2Hx4A2IAoZe
0a3RrecH0L7FSuDMyNIbD1Y+dTdGoCqWDtWs73c0qIF7jSD44YW5efTbnAEaxAS5PFTjIE2UKFOw
IpzVDgyVkkT7TySmVnSiPJVD1LnXaFzDoKdpgv9ameodz1ZTt+UjXj72Pxk29t5OGDbbYcBxWNo6
oOha6jjIfd944AZznSSoOk3+cCLjxXeZWLhzm6m92vsdiyET67l8ch05EkBdO1epX8ztdP4rQNyp
SoGI8GeaM5aoSKECuT23dkD7vWMBZn+c29B8dzWe+xrhw+jcZtMlCb7kEw2N0CxVWizkRYQTsVIE
XVUOh8yyLV9ph5aNuByFs7HeZfMWZw7LvqiFOx5kfxfdFKI6Hp3fCJ7+lSwvGSwqjySWA4P27+8y
4rhYINp+9btx4sW8IEURjZjs8c+AWXjy5d0M/TBVhWOn8EgwJBdeROUSHhwv59Koe7B5b4wk4pEz
gXI34ld7y7FUiBOznkJqyzE3C4wWRK9Pk0JV8ydoomrzcYVYaIZ3EYM/Oy7hhdx2o5Kgv6anhI6b
zKd9CKe2XBNjt8q5oOcRkxKlHVmgfO/hRVepX+BXkQRUT7/lNZ9wNxwcMyrTQN42HKuFi9S9OenN
DDq8UchhEU43o3MM944uMDQ2Y62I6i6h8WkTfq9mx0OWxsCa/u3q0ZJlnL8hH8ijEpz8m1XmItcL
kt06N3vbbisoBMKcoO3Ho8D69kcSg19OLXBoyrPD1Yo5bReJLOICbUd8718uywRQVq1mjNaIKB5z
aE2oarKKUxMqthp1YWLiQ/hE3yDUmjzx0kQclmECK6BPoE68ZugdsDIso9k3JJtZCzmxhZP47Qnz
joOnNSXIB9N6LUW1HBtB2XJWuYiUva828I8PJ9X7Vn0SBJ1CF6tJMrvxkQPswM9oQfJDLyAo4De9
kYi9D09H7xZ71QQSf6KWlB3/OuWKLwHmjfCcmAFYTSDf4SZNHbHXcptADDx971lRnm4QyU8iwuJ5
BHgRJGl+j0l4E35oH0VzJMX4D5bZvIJV7Mq9QfRINbW41pDz+HGo9/aeYmUhZGIhKY6J2XmA43X8
naS8xuEJdTZtMCn8kX734TNAeg2ZsG6ZXpI9xYC8FSvo+OpBYKbfat/Yheb9OAmlA+Xctfme+ZNZ
r4p+T/PwXOUYA/rN5RXMdrYKtZo5Ypq+qpdD3TvrntsO53dwCLxppT9D+eCev/fij1TztucCe226
amqqM7qT4ZZIVObn6q4drqZkqd0XmQ4+PrFUyO2ti5QASiXGebh6jRmJonViPdoxUO1xWmBJN1RZ
4cz58Wwf0+adxVTAZ5XOscewGbSFUfgkOCHuZguNCZgEd3si70LFW0RTLE+s8a2/mwoI2vAHTuWP
QPd82Avk4su/P16VWDD2pvsroY1B4DM5KdxdfkQ98am40b0GLurUxEBp86cl62QYyIJZEm+v/CqB
WJc9RIAqrV3PoL4H/I6f+/sfenbrtWPPdn4LPwjvEnR1hFpOBwg6M5NCqG+uQcv9RfcXCmtd/vJe
U81HwmYv8gKlmUB5Hfi6w8wKkELKcSGaefYCqllo5qnYanJUJVYDq73Jp0rHWvmKYyeTP+khsKti
jjYDCetMvKzQDrg+jl/aB9ZpN6o5bXNAh/fWroDtd68lkU/G8pkLRCXrq2NfY9nne5UfGWR+CI7R
9J3QlgDBcfAJ0bZKBTkoEzHcJomr181rJZTtehWoapdWUcqM4qwyRjiKRmTF99oROu93vUE55+WA
9ZRScLAJrAkQmnu49UYeZKIlqInuH30hAviHUVXx85/PcWVmghI8jUEpItrUNEmd3sMshZbk+JC5
S7+2CDDG+UGMosXX9MlIb8LobPDXx6RiIeSJMeWv+JfdDfppxR10nUbppbl1v3iRNZYydL4DCMpt
9nvDLYJzcNCqafj5omJFl27TtS4awacjTkm7r2I/kOnegCfNpx91CJQ68ci+9kGmFD5SE8Zg5JYQ
+Oovs/j/E38fkG8LofuJeTmWX0XyjrrUmCPlp1eTs7Nnx5duAjPO0oe0or5IMV8tQ8b7uuSsd2ln
M1ogPO2gTH3Xb1hWye8wlmXKpim1IUeOQ2VV1p2n7cUMR5lk8Bokz3e3P49wN4AIYZpGSD3+2g27
4XNdJk37fSGhq8WcV9RSudkSzx+xF/8/5NNYYHUjTF8RfPS67JcBa1UEE3E36UZoWef8mn6s92A9
UcM6776ZPWI/scUbBlBbecl1cWy88Cj8rNuANiwAFaa1NHzEmu3Dcw8vKbnG4UU+d6xb+dU2F+vY
ZzyWOgBi7K2HCZZcXBZd09D70CBSFVGYnW5YpfCG5zp6LMdhMhqEbiJFWKc3GFuDJ9l5rZHeKUGT
3t25iM0/LzDO8zbAnqJVlQGUj4MR4OBFzAzHYfFaZshprjLpTE/e4OSlrkt8UVx3FTIav3PCP0dt
igqiRJyLw6IEm3C9DrVfYN5z+We+moYETNPb+grLgrWHnsi+
`protect end_protected
