`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25696)
`protect data_block
rVMdHTffvqkodplsvFgr/P5Y3ywV8tV+PcPATdPLL/vd4oJGe3GbGGgwOaxEusynJpcJTmrWfJJG
c+C96SJmlo4lAqr2dHnpxcp6bqpTdr+PhJbeRM7i90nvpA8AxyX42L776k3yvHKNy6YFDbUB8TYV
/X3zRcBFaG++MWfE23ZxaD8nheWpzyu8qHDtDZ7nO6rxpjWYre4jwZnnMIfhkou57ka2ho58kDv3
SjouxqOIPq+yH6I63Jgn79gkgm91cXDNZcy7q8DwvTmGN1UkBeqwhTli8JVB6IIZwSYOvSLD1Q6+
YYrl4dyNsLFMRM0FJRWa78w42ICRAXfjRuU1I+a+TdQg3GjSj3IKT1kpEforySqPHj9xE8oKLd5D
j/xViHA6GlsavzfieEaX2Ak8+XEi0oVPTNCsowQHpZRuPM78ua+w8SO768WBA1ln4tcEuLx0tVc8
qy6jhD4EdMpIWK0Kzq0TgZ7nFPXbqP94xHaV1pEVeW5VdwXA6tKlLBHxK2bVLw7SpwKdZAASU0wM
3eA5RxWOiCassmsrTCj5vL0E0DYqGM9KrFvzRlw5vdMVkoqgMPNbB7uccPVsO/o70rawocGXslxv
tVL1jgNYL4u/xofK3zjBEs18Ww0ouxqfil4hY4hzZnAW+q8PL7ByOMhTkX13FPZ7BIjyKEi7/8U5
qUzxkejya5lBoZiMxWD017jNvd+22urKPZGU/oRdf57h2f4WZcuyZZgo76zhRhgOAg+j4Ot79vKU
W8kYeOQjtuk5/olDf5x/g2mfN3Cb/ZiDiKcljCMIWLryYEQ6ygmvCXa6kr9WXbQX9i+VlEZ80uZu
0QkAnT/+zqET5g6JZro0rIiOkHnLSDui6+pOP8d84xXAZB4Xt2FYbI7NoYsDCHMJjKR/rARh2M4h
WWPOzH51qj1PXpTQ6qorVy0NxhAXPLzDRA3FCpAvzvTt6MYRO2iYcw0U+2PM6/iFJ5jX4CkmV5qV
pLUadq8ti4CHbembj97R0PMz6wHkaYXKlF60zX1n+vpXysV7X0u5RN3UC+ABBKUy5CGNasgOUppL
b2O6m6d0jKHF+6UYtRqx0hUo2mJR+TS9k+FCCR6Xhia9qXqQqEJ14fbFwrMz/EH7GSEwC8gofRD3
Lphuy4KuTK6mO5XlWw8wfTjMg/DOWE3hpHRaX+Deml5LyjLf4WZCubYZh4ODnDTbV8qWngtDnbDu
silgYldsOYqH/pJcrVJlzlF9/WSGGCl82sQHLlLTDlP2iVzprkQ1lvb0Hc4hdPDK15GuHYFDjGer
55gEF4FUWMfP6y29qY+N8pgVUo0ULRGbXdn1fR/V9sYqgQg+fwBmJkgpYw8R3RKsZUmemwMbUmNk
wOSq9vfAzJdIavaGm0nXVcpzG4eVaY8l+kr3tukHgF94LoCBX0ig/5Cvxi1HaJn0xz0uaH1OFnJ9
r/3P62w1YzbmetJU0tEwEgg01vhGBPUhgMnk+6Q48I3zw1YKh4IpLEsESDNP/m2S/PRJ2hFJIeVE
xtnpidyRImUiZw8TAUvvi/c9F0pEKCrqXnKwfuo8IgydXjpJk9TPo3YqBgHS6XcEwTEdmCZI/QTy
9qckTrhd9TS9ABoVqv7oNPz1Y5+ICCWGx9nOFiFjxpK111lTuTK19p/CTrRdq4/Sr8Gm9M7bFc54
pMXub2uLTYNMYnPivAKvG1hKpB+mKDIyzi1gm/yyhOJJA4suOxjBSANzk66ytq5uZGqo/9Ho/Y4S
Vu7lj9OVa1H5VRRvp9ma8eKV8XTjd2L5NxgSPA0BdVDNJs8vxcZog0Cxzy38gWuBIwbdlVn0ija4
qb46b5o6HJJZc1XwTTryNdk7M3yDH089DEkW1YP7YrDCVa9hiXe6RN01bu6xpYRGEPanWdRau3b0
lXgzfxZtiQD1am9l/WV1fAYLHv7mJhO+RS4H5mn0+u/cD5r987oC3yInjpI2OAlS3de8q9CrXOnI
JMR/Eo1OUVQJA9e89K6RBcKDVuhqis7WV/jBah4XdW8DygdG0rHBP/aC6Rwn7jigo3+9nDiGr4Sh
5TVR4olJswpKZ/iuqx1Z7En6/s4NVmjbQ+dk0GwDpC/2AQgRew2bRpgVGMk9HYj1HCQvjr+oMc//
3FZF0hxTCKfUvA0E/Zi5qBVraaQ3PmtKqhW1CGV7c819Ai0ySDN/+9qQGrs9rhqbYhI36zgInJs+
3AeOMihpJY2ZjDcsQT5U4xOnTYapA3asG+wcLwyMPZ/GB//fhV7GoMpZPMoceXE633FwgTzRZCW4
vn+qC/6MzTZ4WpFNMJvmCJZg9tfqt5PUuTk/qVw8NhuWT+aV1ZLE1D8rX2U+XfT0jxOAj4lcYlYF
aBC3k0gmzXN+/HojiQ7SDojDeDJVWukVrS/I/HyF9q7hbl0DnZL+VexH3RRpwvR6FDR/+ka33kqK
po6ySpjYssWODOdzoc+L5M2sKYHluKgTgP/oyGO9MOhLuthWmDFR2SsYvZbROal1vYH+mKIdAifn
7WOMHP0qTMwH46q+Uy7DFaVaG8KtWqMuJrRGckdTrPET076LYQ2L32PlFifhV04pkJc2I7w0afuL
RSYMSnVIT84IENtjr1OoheGW8h/F+KcBFrueiow2Oio8LX7NGn1wzJbeexYKtZhXPZuGZE6UhzMS
keX+dgXRqKOwLV2tTVZ0gYIPlWUCoUsgsFhLQ8EZyc9zS8sI8UppSnUHMBrk0rbXMuzW9jIUhBdM
YXd6XEZgfl8jT1MExYvMdtSdZd3DngfTipkkt0xRQl6ksjxZXNZhDfHgvcW/w+1cVIz2VsWeVorv
unz/n7uou4aS6aVQh0w/0JTlrBOjtB+xjj8rrozZBaVNCTbyHAGw7JyH/PoR0I3SJJboCNpw2mM8
zi1WjBxWi+NHwVbgXdjaJVhfFn1hCm0Cx8jGMGjxroLR8Hzy+4P2QrnUR/0fncACISkt9mvLiknQ
HGP+ji86Kqc+ioQbS9ESRfV1yLAXSexONIW6w5zZNSoljRsL0D6bNNq69uRiqQeyA6p4LXqEOgSd
+lfK80hSPaMWf5+1umgpL+QV06lJQumdWggbJ0YhM1Tnho05mdH9si9dgfGHHfq8UBL3lxBaX0wR
PuewoCuD2qTPdSGpxtoglzqhoDUxvtNqAbeQX75UqYcGqPOLbzB9+ijKQudIkw2FeqtTvfCkedjw
I0HXLFl8eDWAYvDKnTcblGmpQB4GQbUFJgY/N2ACk6Nks7LJEIQa+fp+d9fbhSj60zDVNCRxyPif
81NOaxj7qJcAxpa3LAb9P5FgfZ1BY1y8zhmYz6vKE8XeeiuAM9fRLi+5q6B1H1l0yMihN2NMylvW
guwmRGIO5koCNT4OpFIfy8BFRGRr5WU6H4aAsQTr+NYOSbKBMPx5+e1P2MQJUFyaOEN6Hg1wqBRo
XarOZ2lZE6LOi6n8p+nfzSFYSKCvkOCwBuwzlfkhB9UTRtPYkC7ohl1ncKKMqxi5SO7Z+153ZS9n
qk79Vxe9Ajg/3ISPgpxGA0mZclpLl12H1c7WqMvyddkKrCiRZkhaMtQ77VeFbaUZInyF/fr6rUUv
jDA2yIwS4c4mMipJU5hliFZ1HST466s/sG38zQfTB/mMeybr/edAc94yg7aRT9u3l74p4kJsmRM5
hL/ok9r/tKm5JOEczbsdhspz9RV9K7FghNC17eWnqk3GKgygzogwPpj8ud9yJSsRV4KvLkIc/UN5
r6htymjWWHDct6dMcFYop37CjgMRZtclNf8BNZir+i2+T9hiqVFNJrxhwi3kXzrU5DiqTbfFwyku
ZPvVKheIBu1rt64GKdPzrH3aZblO8IXW4pmq/dVZU604v8rf9DabzlkE7JYIv2zD+oU9IiNlAgMd
Ic6CEowMYIxVRaOht1EMgOW1wsyoGgDGXRxl/JngnjzCz5c7CiQ+KQetLvfpOMAbSO+P91zJpSid
Xp9HFPyYJyuNO+t/GJnbQntNtxfXAycd9JlKeMgFwy1iPd782CC71DP2pd7NwMsG7EzDYqnjPgPk
0w5c3w4d7yxjv4CVStUOEaOdNizw8vpHsz/h6Igb9lkFeASnBUr7buRe5X7XgoAOtgU7FGJECs1v
qfzqtMZ5rC2mf0beR8mc3YOtM7FdT8UN26YWePNJhKl+PIzQdH4T/1UIZw+aEF9jjsJj23KZqvlG
NWrS6Np0Tsh99LQb3sb+Cwt8GGe3YWF9xqpS+uapyZ4gj9SEp31SJHzB/vPk/ErLERrIbI+2otwj
o1zZgb3vu9zLi6NyOEw+C3xlbUn5nz9ZwZCMF9KOc4TvRlhWOeW2NbwxMDVdq7VLl6yLvNvZdAuY
H9AHiYk4+juU5+zGiyRfiLbNAretY1JmaCAtK0IqApH0WsicBj0Ld4JRHrOrMCBqOh6G9QvSKiEl
UbUScTcZfvcZ1srjGyLbU77PKxGTlGoGSMrbNxLqAYe2tfn7aoMxQ4YqEzGObWDrGp/9dNgTupYZ
6f9RaLTiiGICV4KYCVK8WgPGpLWQEIStzcPltk5Vc/QWq6yd8RTQi2L9DEf19CcsfbJJMole3zwB
o7UbOtCyh/Cgb4Vbq1otBWYPr/I5PSnI/ND8c52fz1h/g1+XHeepf+6WyCbGhlIQlxXWvDwo03RO
EFaSl314U2EiPqu53aDc5QgKe8Pz777Ah1i4SDAdfEt5+5/QGsZDI1tsiUHZS4QfV5uMyrOheIpt
37/UJG9gK6oiqOyBvciqho4LhowNgDNrlBNYZEr8ucW2iEmIczgObHDaU0Rbf4fRDsLyPYo3Iv6K
sw3vX5n7/4kYI4BOetD/386WUL/Y/Iu1Cl8gPRmGf1zwps4A+ZslvZEDd1NcvGP/vvaf8L1hZJsY
Y2fGDhekcuhpcYBam16qwqA1Glp1+n6AKKUm+Lv6KMqFmkHElpjOaMATx9cyqH+AIRyBov39ArYY
7rLxDLoV1TUQxOm73nUII+YVnRZso8wV+DXv8QCi7/T+k/1pGbP9STN0p+dG/6xKkelUqC2AtYW2
VXa3UBeMvJEgdynHGRYkIxJFSsDEem6NmMDZy4k5sENRsAVyBvprVsSHVbQzZcUJYQxETjnPZAwz
h/48x/QzZQnTOaODbI1FZsAtPuHp1K4ZmbifU+QhF+dmODpLJvA7/kyI0gYPFWjk645U17leiyZI
Zyjdje2PLdQcIlz0Ylzh8dUX0JNslD1xpX+WCEjJID4mZiZZGQmCJ9tDcC4BRdjbKNkhzM7zMKNy
G5xVGSv99gEMqa/O5Sgpaa766lATXWb9sP5FrGz7zTpSjS/yzyzaFjcgzIevJbJHG1/fZRuCIc4S
Xd85pKFn2vg5uGOsYRYoJitQNz3F99f84VD/hlzcWFGfNMjBEfJtic9nt6mkvbGKR2UI245hFyI2
Ns8WK7JBtPdmLNraGzKy7G4DjHC3sDy+aJ+redd7/9sWj1k7o8DhbPHM1u5XAIrlZDDzEtSp3NwV
HUkVJ5PpxsFe2IY1rOb5lEiB9FLSwgbSe8je4k/+pe8FTxhPEArG5wXw/tkP9mSDPgPiYZHvT0rp
j7jGyZy4Frs/4MSG+nTXHosms3hrcdmhNjDbmTwJYOyUGZ6pRCord14iDSxYQw8zu2XLSKI+A1Qo
nKHtaDeXGVQaeoKfyUN+3Bq5evNcJL48LdOoruPvhroCkVAUPKuSXn7ywlaYd5kNIYqNoI6Ujs1M
H5P/wzd0nF1BQ6ny2MRo7Al5MeTCMuAo9rn7YhSesIKk4ziWhURmXwqPbb6XWULTq61i2gSQz+md
MGVIjhQ6RKZjv9LVBMO6SISoBGlNZf30R3wsjmOAxUd2n6APVk7Grr5YiICUh0El+znpoKzA93eR
XlKdySnacjATEWQ6hMBMCd2E7Jwcg8zAP0/ZlVGXukdDC8tHcW2MYcTi+txSwI3GVlJHHv/Cg1dL
RdF20oEnV9P+5mrYP7bcXgsrKpZJwsIjttOPhgzOnDVls3RxCdpoCYQbQOyn4de5nVjI8EI98KjG
cb3Y6VD2NjTerOFl164fH0DvOjWqh5a79mUn7KekjfxOvqg5S02TXOJZ91lXhxxLPpKlGC7q34hH
Dnt7RO6oyGxVshZXX4fj4e+GAHtzZ9Dzc+bLczF9Gk/vGNhC2WdP9miVNlVO4MCYY1+hk3XsQQIK
XQO3wbpkrWK7FjGOAqc6MbaHTH9B/OCILYmEpuxYKDjxOgm4YwrMLakCKqLDsGElQw8YSNqSCQrF
gOeq+3S7vlB8C1+7ZF7EaDgQJWBBrkYCJv6XH01AwbPnlzMKK37LFWXr1F2vtf/KNodDipcrZ6jb
9Nn6u7m8XWoapbm4vcUfqvoWIHn8P6sTMuluyy9G8etWxmu138PGoekSAoBhOOg9XaXJYrp+lJAt
LS81077IdRiXZhztgLM5gaDP+DQoP54VrlLm6yP1qCd18kMHmuuHqY6uzjLQxMGPGaZd5VJxxtnN
w+NYhgVWYBsBXhGUzljInnWYgV8WctZmT08YbdyjCRfnOXM/hvPRl+4/utC5D/eD7VyRlfYb5UOp
XXtXFJ/YVDUZWmuCWKJCrdhlpXxPWt2vibZiDBV1FtQN9OG8wz4G+QRPrrH4kSndG1QisnZTiB3w
AhsRCX6/74i0hCgVD0V0gXjElqvnt0qLYIJWsEacPTzdBoJ+RuBZBb47xRXZ0MfrqpshZJPFMkxh
6LU/V6d0QCJbl/QuyzO27xk9PnwngtE+x5KdibiFr+jScoCJYzdkLoQkHkH9U63Re35NNitkbWwx
pTNxrQ2WB16APUdlCBVF3DxMzF9MRa0mkuVBJlVFMk+Ay7fkH40bvdNILWWBw5cGYyFDba9fyRX6
d5UDhTG1YgC+20ZxZwTglNsDzY5t2WjRHuU0uQt/vc/Hu1yLl81q3w5LVoPS+uozr2FDSeMECb0X
j8AxTSZt2SYmCWjJ8gbi0rqDc8BZqRRehXRuTC68rRULA0+1rKEtYlcTG5OZzkXPcncLUAFejbEB
iCTbFhVSATcMNCQwhEZs21sVX7uuzY8e87qELBhDCYIug+v0w3EFMk7qalYVbvu+xrkM3pubSpGk
7MeLuLCc0nYx40c2BpWxlkySQaenj9It2M9StPH4m9MtH6cOhAXfFB/3IwbcfNk6Tf4+PzEDcdxP
Gg0HziLOBIYFMnV7XGQw2b9bCbPDUzBIejD3OwVdfuyQOaUh4nOf6p76kodwKLFaHk8moQwvhxh1
hCYuQuKHKEnagf+iSn9IYWFwFSaiD1jp4pKGH288N8fM6xYKqSZOKHOrmsitHvn/3Wkpfd9jt+fR
CfBaas4hWVlxbxCPkUMKSacd+jX6M3EOsDCT5wAbpKw9BhcoMCuRD12O65NURn+JiGf6zEVN3915
9HQnDYbV8sCMzYP463h9yMNzD7EXpSeOXnQOp5Nt7Ur9ydixeLUB48wfRjn0XLiQLpmQS5tmgjvx
hN+l2oyJoa/a0v57CnlTkP9TEuAH7r4OlT0Z8KoPIdCTvmU1SKKyD5cLDpwlqDZU25Sxhi33nSXr
T3pu6mzx70c9rMm4HlZNMUEMC6GRqypVDRcXTebehgD4zPwPSi/O1C0PTEwuVCqjfisDyKSdr+zB
WuGal01yllVL0t/xiXSY4Qf20HGwV48JnG4IJhzjHnkWitMIs6E8QIZE6wGpRTvyIizJLYlNA6Df
wRZCr7qpBwMOK5eLSQm6fkUXzQwT5Ro3yt+yBGZNduo2L/2jvqxwgjQl1isf/c/69OmDILxabrJf
LjOrRxsT186adobypbD98leiZf/TCJg6B/gvDKHyWwRpTWiuqOyo4nghSYAb+clbaI27Zh7ApDwm
UDkL+Y/mRvINC3EuYqikZSqQThemsC8KxvPQTmp9d7EmeZK1961jvuUeP9IfNG/UQiwrbJzl0wdn
HTbZ7Y48hGznybbzvLn0QqGuiCZRogHF0/bYf6L/kQtF6T/xP5OPMKN/7i4xs5c8eMM9vbRaL7nu
MGxzTsDBeJ2sMVWUp1XqY78xHcdkUoJGojijkDvq8qV/s0qncaVnYLJJ2XcTOSbUfjfhhTAsxndt
KtIBBhpsi65+5SWubIWab9qWS5Lbz+RwflFsdJ5eYIuEbUsNNBBz52yVj7Gnfl2PD9v9kD2WproA
4CQahC95oyZ5yACVJXkl4W0+zqEk/iH2MAME7EubNSFBhsqRPFVk/wbw9v7v2ZrnP7dfrIEXLO1/
Ftjk1gvpY9C59NpAtgj8/I1BfsRFbkEUjzmO4gAqgf9X9UewOeDsJ21WOBH9PlExv/2SK1YaRMu2
zBnpY4nSaxCHWiu5aBVSNqAJP+tY0vuY3X+I6HwVe3S/ierL9sD3fa1L7apiDzhDubN9W2KuJKLf
LIJ3ewjEqtFeKpNmqPFFEPfgx93/pRqstrav1OMS+P7k29wDk4W5c9DGCOt7ZVe6hEcRdUiW1kph
uqwa8KYotcHfKubG24i62Lxa4CbEI3GF7jL7Ae2Vozk0wvaKi+D2yLyqH6VrLvdz2J5glBtMZyXg
fPiKQAryRplDp6ZGraF6OTsaMFkDqr86Ohh6Gz4E9/KGr4GRcWo2fAXJqWw4XVBst8noCCbzNclW
QxJeSs5BB6jo4yB/f7CFLqvXfnd94CLJWt1wDqHbjO24kiKfAUcjvAAuCgm5xf7SpP4IMzZsfG/1
lUHfACt4TZB4qfgkEY01aGZW9/NHByMGZXaC/G1s0IeHi8p6U64Ji771S0YQVAQk8y1toJcWwOv/
GZix4xIKYvb6mjoRfLNTN097nCf9+BMoOw5534mV4ZvRZtDznlzrpKfoZkkUCZgr1JebdubQzIXT
hUmK73QDhdLw0SkcdPytkcOcJ8Zqq6JJ6uDIcW+R51Zqw1glvdMm3hsnCk+GDDer16bx5bmRQ39X
04E2/pGGD0KCJiInPc3/dGAJooMtaAeLUkRREIqvVB6b4EoacJJs+dRttGy+Oj5V8obfdoeROT7Q
DMvzd0LK/pXt5mW9bfj00wNrj+sZQZjgwG6/FbifldTs7jNEDvzDO6aiMa/ZPGVgWCgz/9/ZyAEY
VRvpFcYOnFPHc8t+EN31zrq3gZ2G9Tl+wFoVg1rFqA6Ot7EomSE5IXBZ4BKk5c9IyIdqYQ4dB9KJ
Gss5310IL8TO1huHpEFp5dnTu01fZ+0F2EEcDq5jEW+g8AbVat/hyNyn4wvQbrwKgeu5PiElJFxt
8HqyQgAEKWDfu4YUaqPi/2bQynIQ9d0mr6OLUzgmLReF5hSOzg7YvNoPEcU36ELVa5QfiUwzTxsu
EptnMLRSLDDmc9ClXuavSYuG5VZdsudRbV+vZQIyatl/CkAmqrvckR4eZb/cIWikg/CtOvqMD5ZE
tF5DROGxSAkc/z21yFIFkHtp1p6+Z9uDT2ENu/LubRMaHtWxuxmJhKR7Q5KEn84ipoftYA+ogIyL
SyIjXelJypJHjHCHdgMlE6+seRgUuNH2/sM6Q/D9jFheRa1MY70FBrs8l+NkG9SS4+0gZFK9hfZc
1BfCclD6dne/Pc6tFZ+HJAOLizPC4NGIZJtfnlBVxMCYTeS9BJgG8DiTHY4QM9+hgTft+MwH+rfX
fm8LWKgXQCe0RwWBC5gheQ8mhasgEcOPNaVKtpGENNfTEjwRqVpjpZQPTqiC2ZyJtz+OqHiQ0SMn
D7YwIAZFmwogfYQN8mFq8PXrgGwUGd//ZMntTpS7+R+X8Ztwagx+SbYJxklaAYHDKraZd7WovHs0
BRftDfdXrVL6viwLGXmwFDJNd9vYQLZvwT7UTBWZk0mPVF7K53Njork4Br+irDQaKsS2yf8DKsBf
sr6KfXy6SJCOHhexXoYmQELRg4jIarK11pTRCiHkG4iXgNYLaskzPWPNRKp4StK49RQP2h95o1EU
N4JlZ4atRYb6TtpSE+IQUem2dmcpN+ZE3Tn8wCqCWrACkVDA64nQsy6Im/x3fl0QkWv+RNQSrzDj
ZUux0qexueZZuHwTO9DkUWEpf4l71OGs/V83PyvjowyaWjMtL4hZ6U5rXepo1yM2Rk1W8csIuTTV
8g1wTbYbqqJq+UWoqHneG8TzDnP4EBF6ilFz0NlGfTRg2ra7mneC/dFsVHRGZyZMJa7i5vrfcHH7
wdgn6MbHa56G8dXmfuVVAuNdxPSSYUh2NaMI+W9FTRZwYMr8TwmBKRMLz1BoJ34Yv+ZR3ZgOliZM
QezJ+SEDYpCR03fKIkjUjHq+jz5qAmfbD8Ze8MBVIDs9vMGPyBjssA71uG2k2S/Ok6Z/xUXCz1qu
73QVOgdBNcMklcyNpyUbmq8GBfPwW26mWEIKWfWnVolaGuEzwbXWB2hQkLS6nR/MTYKZrySxos+1
x2zswIqbZPPuJNEoSJNxO1uMHZ8WE2dcEYKxReppnMSorZ9Zm4cB/fFaPIvKERdoWrGMveIa+K3v
eRFbnf1bkFo+vHRlr8v+oC5uMkNi0CGDpVUDXIc9ryy2ThlbdsT/Rf5ZDqd/DRp6cP2zIECSdwvR
NTWDECUtGYGxwAjJuJRxs0A08aWJX/erHd9u1maWEV/of4WwlrN8rWUw8r0DndiwjChHCMcPNVyB
/v1d6My5uX/x+arO3hXWwSx0+dD2CU5D7h7P3VA9KpY6BBkQns8UGYFCHhyTKbLAKx1UsLPNYJM5
hCJReMLPABwRPkPgQw+6/RnofwlHsc5Rr+ccxoFhjH74rcsXvGs6MFW6fhkg3g2KtahozhS3+YhB
8QSrix/hHonZ0F0JU7eFAuJ9hkZAn/wKAcjwozxiT3cZuK4C8tHqnJx0M9EC1xhl6sVXXt3LENaR
iikWaCsPuUurUXWyd6Hr0AzKty0kne/qwpmwiBjiE/fPQe7Vb5RMeh8KrPcx+7svUoJIkoAR70Dw
qAWcn8FH6dc8XKEMiiDstYAJcJUUeR3tMSjf6/timsKIeKNFnjj88KsE6W8KnvuQw3QTdFt8p61Y
aA3pGG1ZXsWKopCpJqH3m+ROjbORI32MPIjgMdub7VzIEx1VH6hoOJuxEyi0lDa/NS6cpXRykh54
2lo3682XsZoCmvk4QqnRu5tX44yt4gRCMW2zs1gPIAbWEmRmjyuT3hviiaVlxxLk/GJUyl8lhWpP
9nfYTWXwRkEZ5bCKSMuroafRddVv2NlrhA4QrgsegVwXzYBD3JP5Ug+I6+KcxLuQ61/VuyeWb2pn
lkXDfXVc/8Tfm1aNFkDlVatVTzcNTBSLgOGfIWcFZoqyFKH/7qFWM45kD0MeyipkSDfoAv7UfXwu
6a+FJR5ijZHq34E+k04nyCRNaHNnc3OL+CnA8mNZ2En31b0EusELqsRqJ//g/eeLpEb9zgxE52Br
3nsKnIV83BVkLNtlxDRzHp2xEZMszetlLMsO67yErOglPW+HlJhvN1jHprRlJ0MPewXDTKbanEwh
PLXcJrZ6KfCISmLvGQu8qi/lkK+KW0YXRNbBgjPAbZNqMSqhRxAJ7FPJ1CI4E9pAdvC37v+GF1md
gaupQkKedvtZskRibxBM7Dhn9jJ/xAZvVfB2VB5UtUX4TqDDhiCKDsmHQ1ZrKW0nPQOYH9x5xC1a
NlHKKXxIrRvjS/cGkph+hqMZ713y2UzL+4Fj+d1dkFjrm81rOC1K+jIyQqLRQTHHs/mjgX+lXI75
ddmHkSBREZ0PeAJJjCLT/+kn1v5tJfDcSxvU37ZLO4gRB03A7iXVL1BDeRRSO8deyUnjyMuYN/xP
dMpbduskBI0424N0pUtLud2+G+tGFzSrxIgdNAF+DcygaZ6DqjE4McB5rUoQHbhRfda8AlhtJGg4
j+jd67JzYvvboa0WVrRNcQ37n3r5TvU/L1jNtgqJAygi8VjhAkBLP9CmNKM+VDsjvLM6LrCcJqrL
Dhd8J8WLZsPUC0V/qW8wHr/2VRnfyOsJRaWvQq+kQD6hGplwvGciaZl5YGL/hOlCjDl8RRK2Fj11
UYm1hCDn7KZcEkcmuQz4FpS1wg79wzlMUIokQwVmTKKnz8227uMWvyesHxEqp74bJp1CkMRUixv/
s3zgK6WnsAz3PUZvSpWW0caVT5/MzDln5ASqoLxHx6YxgNjR3jlX6GOREh0cXhlF/0JEyldAnxD3
HcpxKzaraUdiCzczsB9fPhY9kMTMLBzgl/1dHJoro7wL/U3QfefQoDDG4rAZIm65K+9GK4nJ28bQ
ywlsauat5pWdKqFvrgGP/QVLdfuHVGmc1ukvRtMXuNTgRQ9LF54Xvxcno0W40AJbAbcWov2Y7+Dh
y/myN02nwJIbgByOYa5GKrLD55tRhDBghvbVhCMuscKHziAeolr2AYueHHeHCdrHNZVmtmzJ9MzN
+lln0P6SUUGlAxEA7P8xdeE0JRvYj6RRQIondhiWvVmUhriEVYn5nA4OzcL9384LDgq+21WP0AEp
zjje99O9YdoLO4hqvwGCEEFDQ0HXkMNHyQFYV67Vwn0fJM4LfqBadSwJ+QB6x7+c24xBsEmicDp4
IXuOqtiniDrhOM0ZmBBYjDfNzyBzycptQ09/1ePCl+vNs/EGrTaYTKXkana0ud1yNGnOfNk/df7e
/DUKT5Qo3+9S3pEvxy9aL5845iSI6u3nDi9X7QJyy98jiBZKgDn9LAvTXf48qzdnNtugSkBmWZyw
RPYKfNjxCdne5REPR62jftfFJKLDfOakaXu4whdn9dNWk2Xh7mQCy8GguVpwLAuGtvVYQVQnGCeS
hI4gWVDMB6B/F001HuFhaQPIXJfkXFtoglCTlyHEn784BSr8bixt6VA1lAu7/uwnGMvVU3NHTrkx
lIHx9cgZIbhYmsoL+l1fiDUreLbPvfDiN5vguxJ5xNFpxvo6IY7ijN/tmjGEZL0uDxNz2C/RfwCP
jH/9HEyVjtgxQ0t3Y8DHUDhiS/uvoNCCkzyOYpcyIzvm2uBBc1oFfO7VLBlWOwUeDvpFKL4vIFcn
W8Tm3MLOtYx690rfpCCAUnM1bri1UzGdptkYo1oRY6zGI1L2QjY/zM4ySdwDaz0zN7DFdnfAZnVK
zecmt5Nfzaf6TrirwHqQVMo2fDcBIqarTA/yUxq6VaPjgx/foG6+D8rqDMrc5NM+2gxhOwfpOVRE
bjX5HRoo0ca6q0dApgpV8v55XoxHanGCIYi+O3HS1HpFm/ifxT7rGFniVSfFHsOcKsWyow442kqY
wmwtNwpHj387iZEgL4t4cv5DL0mhkeMsHLvH3ypEz0ZUxxvQQaFzwY7fcVIuGv16zrjbCrkBGykE
zET3K/1+SIXYWda2qXl/oeNycks2B9nlOMoGtGOHKi91g6xljdbPFi7mGlPYGRHD2wrXcTDrpSeE
nbuYneUKYi8kT+4c4MnjPeBzd4hdsapeQUZdWPxI0T/ZUXH9T5VLWwspfBLJOOjIK6oidwmCtBkI
eBeDtXXZMcUrTtGY3aR3cpMATEIa/9wMSGz50HfDOYHAnhLCVL0AJfsqR3lMCT02aRR+NyGvXbts
Zk8psovbZSBoD4BUA3OExyXxn7G2SX4fhPLENMvZug7mbO/3tXPxPyaVAhM/t4ETa7sIt2QRBSPz
YjayeKEbdqpVytLmz4F7rBFbQkcw/yy3Vg6EJUbDGzvIJBfxtRNA4+HDAUujEbTqs0ajnCLnnPOQ
EO275Ckk0iOmT43jnzS321xiJSVCM2sJ7QtSlOotyHPFx0q3FCy2DCzQjjxTWt5LzaJzdrq20hV5
jJjuLcpdEPHxwBFsigdAjwoweRq+626FjZzlYDq+MSzHgq+LltNPBD59PUivBM7IIgEXYD9nWCJH
M7DwqTIo2OtdRMGtHncoFQYO+Lq10MyPHiHhjej1x+kTXI0NgUuVvz+BM7/MQZSVc5JZWKEE+Eu5
r7XlSMJ5SKHn9NYmUR4Gp+wwNcEred6G+a2iwfdIrQAoCfZ/Z2X1vwZ/0DZM6epe8iU4C5Z59Cj+
B0a02RbV88v47cLaKAtv1WwiZoRDA894aksnSRAslGFHKa57Wy5NA1NncdwdhfWtap9ljHhMM6pP
4IsR0j1Z+xtoAmPpRNCruk5Tt4Teg8wFnOLxYiLgLFWQAdf+8onTk1zviA29uTUpE6Ef14OlOG8p
x39rvltQtCiUG3bT2kYP3eNyLd/S0C6sONsnXtL6ksXYZmyUM1Zg+BnUD07lFXH+2tE70MF6VC2H
0mVzqsWYd7txOTeJJfuy0MAkfsy/ouA/FdGrWvKnxilJUQD2NhiFmku/soJ89gqy53sTIn070ZIx
2HOXZUcTcAP1DVxaInf29kUG7SStz7LHaGmusCgRyE6CqmqzBYtg9kpgQn8rCq8f5aMyLkYX9KIB
vRb0p68BDGr7+vFu+OuhybLHwPRwSYBGc3FTNTzLtimWGERg4mN71whEjnacLR/xbIjcS8a8LAlD
gPnlKo7IC7DHq7cmhTkJdq1NRSO2nR6SKxiIi/K6724Lf8dCw4MrC7PB7BPMsIGE5dE3lpwmSXsy
tEON1KJZXmOlIuFaKbibyMbeWJ/OLowTXPVhdpXRGo0gzjbWfct+S4SRGt81dPf9IyJUnn8C6eDl
rCQwQVRhMfEkc83OEj3ibDJQgy0zNAB52MSbFdPC5ovEcQpxMuQVgww9rzszvVbV/L6c1NNjHG2o
weQkMPOhHn3ZYkEM3Ze+/cZP8y4EgO5zpFDxqC3o02nxJySzEoFXltBxevTw4eb0wWTZtUFcOUM9
FNCB0pbiDOlUiRwScf6zL6LvQ+HLBeWi9ErLZHwo/FQJ5PscPVgiq1BZB5XbPZrTGGug7ROSgJfv
Lj8NVz+ZgGLpfu5CQ+OI5X3ZdOnOv1ywQU8/bxezSxiVZufK8fALTNyMOTojmU/KjB+Fo17D90LM
jkpfa6+bT+HWGjiai+Xszie5Ru8KqL64jPHvw7wwDVEnTA2LXM2/aRHlQwlD09bS3SRY4Lr03Aot
VE6+hHa4YbQSbB9jmTWwVxDgLkvpxtHv7ELXOO6trgmErLzNtTRGQ84aLEg6akNqG4cOoENYc2zF
BXOtp6alXUxkvxDphFYetX16wXPiLl+0nrxl1broWQRm4I0nWOBRCsiREccLfLO1alPoVGHJMZR1
rI8+pG/YEhJ1Ll3e1reLj65nWViPV81PkDYZWjrB37Lb2kuSwcLKPn6OzMByWz5i1rNTMPnpTj61
+oMBnFS4r4OO+hR24qn+9nGu2a+Yp7edmPByU0UBHuXabuwR4GRMkBj9ZPTqi/YnxqBrpSY0Fr4W
avHYD2xHo8kAtfvh+d88Uk6wqjVIpfK3GOaIQS1xGQWP640I6vJxuzO5yvUSX4dHYLQFO2w3ltgt
B6n0AvNGcfzl+XUAOlpixXqOcSHX30Yftw9ABcuw/tujcCUF/JnCX5zWEZJMBalVLNMBFoXuZAnP
5NPXICtsyA5fgErNgA4/QRHNymO2DlMnjN8q0S8b2ULgdVEacl0t3V0z8K2VuSY1xMBzVE6RmKQq
HG3NOSWbvCyyiMbHNwd1IFEcO/+BrnfBGKCHgq45ddnupItmauPwd0/7IL3vpzYEQSBaMHUxJOig
fh+v3sJCJVHVLTRfvmfOungnra/TAJS4+piBFRU41bzQVAXmeVkbT4yEogNK34GN31PEAxAIjcHa
diP8bN8JHgSg0rX5Uvuds0zQcWkxEZ4/a0Af4RiFNrdijWC6Li2Ot+VkkbUFFhHJXk+Q2DajWdyk
CexJTP5MK+LTNyncs0DxGuaE1o0kcf7D8I3cIFxzI7//RTJobpORhtrNDXjGp8H+ECID1DT+ZRjP
00xGbpB3ATxUe3F+TN/USS9pylRAdQPXFdN0AIR1rTUy8G8MaQgL+/lUYfU/v/w1zFi4fLjd4SiJ
SQZU8rqsbXmLgBkD7xBaIjbOdazA0eV5SeVwpIXAMPF7Xl1hteEcGQ/uhjM0sLYbzX2rekKrrkv7
QDuRlzkIw46BcOsRm+xRSY2CXQ0fTBQvwtbaf22mVxa+OChzp4JQrNeS4Ao8J6KmpFSTMx0Y/KxF
M1AfMpfa/rO4Pjk7hqZcwwEJzohW1JihVW2jspTdxdqcnJ2vfFGyhEJ+k5//UyeOVzCj/dmw1exu
ZMs0OeTU+P+XUZ2BN5Jz3eHctBsDUoEuZCRRM4ocQutG9ypPfaFx5lCDpOkKcwAgEU580b3epaDX
Bgv0jWIf/GXF0sBcPlkqrdnIykk03Qd8hbUZYNsbAipxOOaUccIjRf3gZTTH7QKRavGlfK3puDEQ
ms7nzjgKsqN90/p5qYOX21yxFiwwq0eupZIi1aQngnbhkT07ALwTP5hApWrtK+5oqV3IlF5iCpxk
6gJhyG7jy0t+gv0DiS/bZlveUk+Q6rINlP9SwV2EU5WD5tF2g1VSgy/KrEuFwcHhaArqvxhWEj7i
yeIlVLjUPVWiewY/52aiy//VJbOwpDULMkIgXr/Fnu0Oa5UVx/OlDB9PEWw0n9dMs0VeJmaPKyTz
d+FWRBP+IoQ7NyeQ8+fowUK9c2LsOA5P6Gi+rBkJN4qBwKnzZY+YiXVnQLLjWKCd/icBzWp68sla
3wlRDskofuQ7XMOBlliTUWRVzBL8PPkyurj4ilem3jgN+Oqmy6eQwvNx2FVZopElFyJQpCOxnMRq
Nn6fR9OQKIAUGBbkcyoK/kQNWPiURhIWxsjTkRouzU5MPU77m4D96Z0hzUbCAwHLmNigpOWDQgME
aVfksOwCYJAqpSUr3p75D2gOYI+ZsylUM6vODaYMertthufOSsCdWG37wzuf/liSNzJwndySc4px
2PycbeuWtZQd+yiWrzS5fWRTv+ld2U+q51t0RCQUI9sTLaRdBXUMECFFYOinzCseJPvGuzbhj63y
UJvd0ZLcb7BwdZUssKWYWOyFsLB026k5zsPMWqvQkcnodDKl+H4ChnEtRGcBJvUwX/D/JY7G2gvu
jIKJUrg+KLW/eWVbOrAzABoId4QA7wgKi3EgRcsq1bVDvtH4iTRJYZkdan5eZCDCabaeZDRz+pKq
YVRCh7ADEsD1RSX0KGMF6nZNJYGYzbysJj60nEabE7/gZsACg2NyXZpQCVWQIKggXMxxqEc5Y8K6
cCOnumQn3bqRBKMMvFj8EmoXuHaTYNhvxwWJ38NHlsfG8G7S2X6lye2IH0xC7KsbtcNZ458Ue6Ad
mCJbs4L5QPfkZS42u48j1iW6Jzdvnzac8ZnBcSPTuWYlOEblCVCMpnqhJ0qPfSPBdfmPhfCV/20D
AK45gih7CcG3RtAgerPrkK5dbXRohxcIIlZBDiIfqyYRj6YEg8m6b76UOdUMBuFZf4vg/WG2beEb
fundhy9Bdq00CszcXpRaynj2g3Zffzsnc5NYPekOO8whjnOf+GCyK9uDrL78bUr9bMT8i+S30x7F
9U1kb82kY57maLlKEChQQHdJKwZqlyZGiCqq/1FmpomcTjHEWmCIyxl147ZMoY+i3Uew9h0We+di
sxozkcHDTlSA9IyZ5vt30sidrsoC+v0lgiKB9L/Puc2FUVQzyxozHE8Ts0W27TO/tJm6EJ5AqC3q
larrnk1d1IREmkSaLG+0unusvIZgZcbI0lW1MuCwNStj2g9UlDTHWQF5u3SF+lj3rSyrQdRfyMEa
S9Ivm8LXehLEs3Kg8KncMGJ0Zlgt1d0Yrtt/WgRoRfiGCydW+GNO8S0iN4XjPsElf5wDff6O4XY/
afAMaqd9tnNUdTedvyh9xzjLWMTF56MQ6sM50oTAXAylY6ux8GNMIVgcwiznqXyTPMKhr0Aj+xVx
NlbSOdv+BXKv1F6qzdD5uG5SAzwNjQcvGpKbVuquK+7q6GtaMS2CQ4kNFRNeKRtjkc6E90bTd2G2
IFjIbYRSnxkwiALGPKSx7jDlx2H4AxihxHUua/3IF9rNQhCl4jiaGeOhLtzIruKy81eE2lK+XktS
7/dX1QJPHvvIZFcDjK4sYywdqLzF8pKlQLFEQ5Ff0mMSFenV8m89yCLS+QMrjEyF/ztsxZYtqFBK
XxygyDCGZZ+OnoqrCAq6UM8zmqsznz5cbQhI0qyRUGvPYTNxQLTaDVjysmQjtaF+c2koXpAteJP1
RD+2Z7XBMd5aqxnX8gZbJcls3OOW4oaW0YciSVksLkHru4yYcagFSBF/khYTJJ49T3oxCSUDGq3c
u8yboHpTvtlGtjnDxB3VX0+yfiJsibCuH1wewXVW/gOept1wcBsx+1qV+V3799yXAMLobwg3yBzx
oErQfSyr9+ee/ZEEdCKt+DzkFi8MZBi9Sixgli6Boj+HRNNA1aM13rjPW17gJyOHkq+UxM4T0lPZ
iMWaqr1SiJWqal90ZcD2fdXus25NkscsEtO/DOrAobRHdLlKzQph8WK+vWbIytG6RoheGjo3oV3H
c4p7kMOAz5P58QJu+uVg1NwiG+j883C+3klKsQnrXVdMYp+NA/F2dON4ZQcRRjVazHAb6Kzbx78s
0tASVTcUXXdcchYdZe9AUh0KZc12QGcDq6CF64xqYezs3krD7VsA5up1FOoHDhqIJ31ufqUb+RuY
BuHdRuwDHLJVrIj09FWR9peM7+C5oRsqOOHbqHLEtb2vFlopMakrOWEoZ+wqRd4LNDfJEhAVy0Sp
YKUwFrAO4cY/pLClEHXbgxY7ZhPjSaYO+3J2sLC/v46rA2eVfVZHH9sFqrmB11F8miE6wPxMuMbx
ch0mIvkqH6WTny+Qmi2w/t0kPAv5RlOZa3AOHBZyp08AHEHi5UvWu+DRCDXidmdMl6hJxOFohxcA
dKi/YAmBpil9NuyPL9ldW+HDw8WEDK4/4tZLDeHfk5c8V4KU396k7DlShDKvp5SBHWvA5WT6ecM/
CBI+07N/iK+TzCZvTamBBPXizq667pRweqbSWASXe4ma0x6L2ZQr22o3voBFNpuh5hhhicfTYKSS
4BfObM7I+GKNGdwh9Ci9Pp+dpF2xjmDbuABk3/n0kIu42gP37+Mjstlib2DzE9EtmQCXAPua/Bs/
sPtg0HCWrMXCAGF3gdKTFw+uXeCetO4ciFjM65OPkHPYf0btN6IcfghnBefmU43GsCM5bxJKA1AZ
Tdf+3yg8X1OAyCrkv7fsUNsc0r9jjrusyR+mvHwA/QDo64ib3rJhUCTheoZ0+RdnVmotz3G026wL
XkGD7kqDEXFTSK2lVJgDo793Mn5LQlB6QZDA0CxklQZhxh9eBGE3H67JgDnpdlhqfzGfUpkMR53a
NKC3fwPHCoGEaH5krNcU+D3YDl+TDr0HaXawo/EQOX51y7CnV08Y5wKCDn6DAMAz0+2fjZeNGKd8
bFrc6Z0t/nIfERVg/cIWgkwiB+tKnl4OVW5nehUJOCYX6Fk7QJ+NLk2B9DekqDHgNTQ95BOfikR0
wNYSK1U6qPQdd5nffZLOb806LyJxdo5NArnAOjJzQOYaQnWqOD5L99hFtRIo+q/2HeZDCQfxNoo/
AUvEmduMO9Q1ULxP6dr7lx6+0cWorQwAlSoWbFVBN3/tnY3vawKl1A615t76csZbygCYH4CYHArE
73mOFNdU98ZM98XAn2jk88PNs9cYaVmXHUwAtMuzWMidEcqaeT7A1vnmqO4GKn07DUUSgXuNaf/Z
rRbk5igL69wdGwRd+ilwn/hT3ujkzTaUX6FhAgAmrMzVQ8sEkgy7az8YDZUMr5Y9yw6hFw9mwMpW
WQ/Ci9pTTGPHeEnlpTgKTO2y4O1DwPhlHyLcSjfNwNeyU+VBaU28KWlcotiwUmbA2K/i8T4Ld1lE
LpieWvJEibbFSXFGlBKH1hlXWY29B+d99IquT9+eTS/k+V0tqgEuWUoKGg6u3nLc0YAavfwhJv6g
rhnFQ0SCDTkLsZygaMJsMHoHONg8JfS/T0Zeg2S0jOj9YeMu0Gk19j/cE+Xv8Jqa6BTaIJ2Pd3KY
EvSuiyinWCs0ph88wUW2TquK2r+3cY9QWBg7ZzlOGBx9rbnec8uik0KfuftpE7Ex+6+OtouZdU7x
JGJrFStaQZwGw8zLEl6eku/AwCF1Qe/Gle7g2w/oFztd4M0gHYF5aCBtVxItTai3hpV/B0gZQoGc
/DVEb1ve+dA7zY0XUYsLHxk+Okka1QJWKD2Ei70FYygmoDtheMcAkY7aoFFNLn9qQIp12dUDrL5H
Isz8GmQgkHV+X26rueEv5PMMv0+BxiFzaL/pvWLTu8OXSbqUN2cxsqO/Z0xJj5xzZoA9iHTFF9WX
unpb+AJeePh7TYW5T0cDLokAFANxMnVDgQhJNDnCd49yoZCdZ3cubYI6hH6HuDfttWkOmPUGeC5v
4XHu7U+mQDstood0ImEfzhnRxFlv9ll5PzNQquslM6IcY5SCfOgQFBOWyse9sot7nmo3r/JaJrAV
ThZgP2IBXdcFNQOjUy7kuNTO0ICWTOpfjuCg1pvNZF1fX4ElOFbWgfoNbSiJDZyYsLg7cF1AVbwz
lwSC87S9i10ZLEknj7WVSPJDV02hLM4jh43HMz2C1iDMw1UEsYH1bPHIjD/M8cOQdIotCJA8MDOB
Fgw/doTL4+Ta7rox9rmBxuLkBKN66T9QaLUhytmR0iu65onFzPlmbA/UZzxIdW4vcdcmubn72BEK
J40iEv+JXeK8pDrXg6xhYEqX0G4qEJT54ZZbSVbHJwaHerdKk1K08roMf9oXOr4qpqFFMlZHORoT
F2WgHpNHmjFYZ+LCckQp8yBZeByy3OYJhcDqdclHIAbMifvg0FACcPIlOp/zqdx8gQ+7OkAj1pXB
+MDF3TruLfxGfWIfLHOVdeoDqlcn8lMssxN0M3RYUyrCc/fIJHHLpvp5Vuw8K5CSfsqAqsH1NT0i
DmbfIT0UaEEtsqiwonCH8ssZ5Zxh9TbrQyO7TooZ7cOs8ezhkdOTlXomLLd0o2cM7YnApDTHK8BO
3OWOi+cXVD87uppvx6sgLqhfAL99lgPbepy93zeTMNRcewuiKA9X+gnkza4imCIvtWW/CMJe09Pw
ZS6IrnvOsHa8SPRXBk9Vo61JArSMifRp7F0VSqkrRVDMLWuVXapgyVl3cAreZmlRCj7fxECoobH/
HueDT1Ez/cT9k5NbJE99akgtn5yX9L/s2/obZ7d23EjHq1DC1Wh8I7PJs/5KhtvdCvD7h9GingPF
G0Jy090+sgHR5qRWpKWi1nhGew+d16LBDYseN4Zz9uX3WH828Xrd86NguQSF9FB153TE0xRYCOl4
gFatu8l0CwFxPL6EOJI3YjcaTZNVLK8mUTUVBewb9xlrxu12QAFcp/ARjnv/s6VRt1eVTuaiUZMf
uWZXYm77te2DzXwUrWzrkAkagIwfxKslKnxFgry99CaPC3DtSNDoIumcN+VsqSF0StIemqFq4dAZ
V+ZR+D8GJ9v/eme7Qz3pWu6z4eSt4KkLjG5VAW1A5Ni3Gh138RvJics60tKEivX2HCCb4I9IxuHO
qB+KeTysV+8xwTkB1KWpZKWOzHq630GDPKKcDKN/qx4iH/5tW2o31/bcrQTHPcHCegJVYheungFp
PVetqef0ZHuy0QXeCdCCaZASGsXFu1b0RiYArT7ZaYI99lRpIFdw+Ub0cc0r5YtOK9B+s/p2fWNt
0AiFKEPdMs5yFIB/xNtl5oVB1N2sP0hxv458nvWTamhoSXlVJK+gWvek7sCJbqeKSV2Q+m+7iz/j
01eh2bkeq0q/TWSsvL1oxnQmNcQ4gYgnHj30A93omfgTNUCdeCq/0Cz51oEbkjp1rUi4lAx83XoY
zbfrXSg1cVSb1ZS4w0QjxkaE4aSO7YvysZfaTPDQCUtySrONrppFG/8/P0XIwDhDeEnjd7Tlu9my
906MuKx/DohSJDwBsWUEyNooc2DEQRnwj0BI9OlbLWHFmsYr7YoHz85hW4pH1ddD8EFR1Jm2Owtw
oHC512JFQpD3Ya3/ugVPS1Qoa0SNe4pyX6NHJDlEUmX11BZK+N+NHKLeJgZ7XHoyYaBTF9O54+OH
VH4nYKvj0LHZwXmFJPh4mzo7lcRGuVUZiTOOiTR17zaNEM6G5xGuBFiaA64OHl5+5Dsh4ceyefrb
84fa0QWokTJ+zk4KZ9HCl1K4qbmVkvhne0bTFGOsx5xtqhw6DZgFTssujCF6Fjjn5irKXnO4b9fi
EQXaAdKothEtwtq4DmB9MOvwqfCqm8PHrGSoqEWQO0+Ku9ef8MfO8gpZ2pEev90OOl7h/HEngmEx
PfENntHBF1XGAoJ5wNvjA3Z7xGf1GwuORxqhZ0Gx35scHMQEKpqsOfP8JVev+Rm1loCRIc/1HEaS
q7Azd6ANNgAxgJ0Whh2C8GP6gD0Np5c8PTGaJJAsh6SwMeCMoRMRGelZKCbAdhRx0TJnwIiSeXb9
O0MZk/00iwH42sQj7ShIb0fvhOy7hJ3dvnQW/qNEDgnmEbNpmKrSdfEeNFEKWZtg3rrqudS5XC9V
aYK0RaQtLg9F1p7A2iXWyTNviBtP2zEYNhJJ9N6oXfYQrMP6TIfu7SDsybDMvi73cqOLqMy6VrX6
rEWVdJbEjdYS3X9Uq3nanOUGsdXKXgq/ISrNPBj6wYCgJiEk3b52RnyDDRPiwL0uXISj+EN6w1UB
Pe7K+vGCvIqoVXcTQcIrIqWAtSxf5i9LBKESlNPStlSJWzXl9dDTnnNuMQAb+WFrxao4zOcNuFE4
riFSC9+K2rS88vk+nGJ9/CF3kqF7UUyUvflpGHvRZ/KwADgdLebjlE5XVSQyGb6pwwWwSRsd+uXk
XQvIRyUFf46lETuVyzfj0QHyYQTZbEkfpQhk1Aorj3mS8M3HueIjH98yGRZMEEw2jz63gq2rIkbg
8OHBAJNx/G/Jr8v2/MdfEnE9+mMfv21nDYDlKf8y/fSLihpOt+IM3ufUAcBvPB++jU7d7EIrGrAE
0zZIeDfpkSeyZ+aQd1IhGZ8+GQjS8wyQNaFGSiUYrM0eUZFSOtL2VEKK09OERl/GiTD27m7wWkqA
W5DjkhjQl5CJzo04M3Gj4caY1Mlvm9ONupzgnIGz/kN/eGf4d7x79LuWpth+nZCbTDBi+FzNMsDr
feZgpbyB22UrhlZhmJyuiLOC/mGMmr4cF9GVngjEckLN1AaY7gVQb8VTInp1LPMtTE3gTdDwrqFy
4WlPko8jdDf3/U07Iq2b/YF5xzzTjxPNCRQtJN8xJ7mdb0GaoqrphNj9ShkpCVQgs2LUVd5zf8TF
CBX1Mq7LcnumvNQMMmn3xhwwjQLcwZ7HF1wh8hg1EKKjXk69qq+1Gb9PNXQ5icQAp/deUU6d6sKo
0Lw+7ZmmnkAGD9LAD7Pl8n+iwoDQoNd+L+evs3pkQ80MoLfoDJfhrQpgNgnUQAbj0JRixZCgjjz/
XESnsIu7SkEc0erDxdomx/c8axCL36HkshpdxakUuEGJfqt9HE7SqONMubhBLeTCd3XJ4TLzQhNK
28d9MOUZmz47171iNiBITtXjRnKnnp4Nx0jhj3U8YLj1V8uDwJ7lyWLr0lsnSJYO44JqlTYiOQNd
44sEYY33Wp6o6XIHZEWSIgIHto4RjlueA+02M7GOd+Qu0lHqWxdaIeMH3jktr9zkJtnHQujpHwWU
Npugs5h7i+215cXulPx54PyUYhVUnbXAYe+7xYu3V1jai90DfNycuQ57jOuhqS/K4J/bqRkUwV4l
HC7yVoqwJLhOPVX2qQkNwPg2thmhC6OoXTazOs2pTDI4pzPMUoIiKkXfbpfBziudzz52R89wKw11
XvgCw+0q05ZsuwcXLzTUasJwDhWRUF841Oms6h04lAHH68nx3kv14LWapJN1oq5PP/cMgystV4oH
eIY0zTFh1BVmp7UDivNZ0DbPmVY/EoNL3im1zCcuKQYousbNYmpPw56/HvtfShsggmmAymnnLZNg
jeJLXK/663/7rE5XhwZ665YsmBAUWX9EEeA9VffXwEVdRzPP5z9QDpuKS6K/LvMgTddw/aU13UuU
HlBh23TIksV0E5edyOu45iNmdugxBbTB+35k9wFMectP/LCyy4TDRDSkre+Z27W07anxmCvxKeZz
tkD220Xk9G3pcab5NzwBiTUdwFU7OPsGwLo5esAU8ksBryUFmGrYQIZUNjwAQF271AcjxTrvstCN
9+xEwd5IdfWUuYG+MVksSqBiUyByqW+5XBRyu+lDic/9e5ulSnBlyeK13BwfJuZU+ecnrjxh5vr2
xW+BweAOzuoK4k6DuEnmNaZa8iKcxftdLn80OXj4OLSpx8gapsCY5YSHnWVbAmvbq3BjPWKvyEqE
LxvmpQraTYsvUy4Gl7vnqH9ZAfFZwYbunXHj80CUuTm12zxAAvN5yzqqNfsz/zam9aOYDq9HXzTs
1y/boREZW3FSyKInAe0nU4PynO3vBy7lub9irHQMjluKc9snY8zpF1wmc/T6KG0YGOehEp64pryX
knRvpFkMQ0wYK94p2Mp/zfLeiILQVLh11/n1WL0VL4T+Q3D6XvDxnMQpKYzDPnbZ3GQU+gV9yaAm
vI/SC+RpST2EyzvbWKS2rvz8UuBJi3mk8PunYyn29YlK3Lqnl8YpombRmEHOMWVzDBE9LInT0Afj
rpByY9PdaM9WRknPQ7KFqWD+uJYOIa+huPjt5Bb3UQQDVoar5ZeuxT7mqgkBW+NKbud9yE72985D
M1Dq91M13pRHyU2qL1BM70IMiV15gxPXGBeZyUYpt9+vDZ7wpIKl++c9ZwRmblkkdpSuSBQmC3AE
0MOvNginyAjhJIW7vsV7CCTpERigJ+USmCh80Z145xXXovkFJPRVbQz59PQXWdNs1Fjf39zZq3I2
TJrDuIq3CVLlXwnlJPsV9JDkbOoXr8AmyrkqLlX3l1z4hB3rfcBO2oQw9sblUKUx3p78545JDD90
T/0glajhVD0Gw6bTEzTmQ5mBoxEIubBPelKHaoVAPlo51yfkUi4bC4iyJMTL9wvRbUCx79aIbLD+
sv97iyLdIkbbxfIs6Asz5tLm7B2AlZOtP3qdRalfe4bBYxQAxEZBbSid+Wet2VZDi6s0C9SDUEe1
r+VjCSxgDbRiD1hYauR8HkvqspJjz4+K3k3F0QUulvD39pgN4Z9UV7Jjs+4sK6GzkuYoFrRQONtV
VjjRBAI+7RhilQvTCPIxRi44OT6Yl55HjPGoZTvbP6tnA9i1pH/l2N+8oYqhg58gHvyuCpszwOYm
WFSqxi4u7chppKC+OaRToPcnyjt1Ipn2/UizxN0PivLSz/8oqbhKIrlDsPMFHcUtVFPY/dQ3gUdp
3SyS1OeE6SNselOQ4hzFZ8ZMr/YXGuxazdhxDj+W6t4ue6I7hlD25aZ8QitwRyuAtb5lilTHjLC6
lHYtMZL9ThhUrFN+QMbxtnzdGa2JCFupvNVUpVYTk9DZKHKSIOXkAnXQ3mt8NrcoQuGtYz+1pi3v
elyyV3bbk5eGd4mBDjuq0c3HX5BPjbfLt9kbWcoaOKn4Dq2rmuGdZfhPOqEW6MAvo4nAPHxFtyF1
abLA5kUwx+Wf/dE/COxap4mZG1FNWh64DoonbcroMbbLnVo6wyjAO2BwnfNUDLA3bwB0hcVc4+/k
uIRvmcX5GALgThnLgfdsm8ZruY2foBrcHVVqiZiTQE6z2psU1B/33egHgflSNohhiT7FgXjljyLP
bYe8NDdX7tbIsO/nR1un4yNd5VPacEF83rqxlsffnip61Tay40OT9K+YwjdEyD4upGogvOlbBIue
tlXrfJM85ygpJizkmj92Cut08LIZJzZphWqoUfwBeiKpMeanCvFjNlCELE207cABGuLxdX7LuDKB
boK/zfyT6dz2R8BqRxXzHooFLlVrS8t82JGH92SuL84EhD6fvYEcCBRRLhqE9JBvtky2ez0tsx+U
Q+fg5DYGpdywsPix8Aedd6MFp7c2togkqYN3oV0R/0JlPMLOdBYeJREhgjnkWuPYnISBs1viS1qy
V3mPqaUBxQ0stY1jWOsdSC6HffWdTHpo3JD+FRhz2E7ksZjElxCl2bca5F8lrB0aVvazUAWceGCn
YHvrtpKykh2yRAnT6PPTGzjQ/I9iNk+9Fy0/p3AUTmk/+LYpFCNXWdnQBHae3BaIgVyfa07/7D5k
o2JXF/bGPeQ8Ska5w4syaYK8nh6dnZzzGS+em+B09eXzsziawQT25jDg33/DTzL87XLdJ+c9FtEd
Yqmf2wa6TzMDxdXO94Ec0aZY33Wa+eTkJxqYwyic8BM+bZ3Q0RjOrtq3rQiqszfnoU8FvLnd7PNu
NezCyLBo7aA6Qzt5SaKpLG+o/LPjo7PbriazGlJOM2tKv44B0MlFTm9WnGKdKbCck7ilg/4jiS1N
pD0FbpGE/sb+jP0J9OjMOhpbJpqRQulbYZx5s0BJXslUHKE5LkNkfwbFYHmx/TsFz6bx0qx3oo2b
MeLcqaAtc7p470MIO8kVaC54v9bPFg4OsKeCdbR/VzN0ROPjhjkBsuVgvtiz4j7KrGvjwVU437FF
Uk5PeAWor2mfLQImOxHJuW/KqwtvQv9KpeU9lKQp53JiD6/3HFE78PAstpEgfmd18k8N0RMNisQ2
KUFFHMKcBN2AeXXjgqIKyB1Nr9dVP+/rZpPMLyTlIumuuXUw4hBpZTiV4R8hlZFONZrTf4r10sMZ
/IqH20eO6f0EG6ABD2+tY5SB2oYz4rXP+Expc7vPTPlTcR2SlLQzTCS5TV/dtX8CPsvghlI0DSSo
LudzNeBFbIZ6C70ZFMmrEsHL7CVkO5DDTqJi69RZ0+cyPKig4wq6OHM/Vbid8ELog6rUt8ZqsCl1
e4WSJlO5Vtw0qd6wUb5wxsZNL2fFdUDeI6z1bDxIo+iu3BE4tDgjlTfx96lFI+vx41NSXgr/xXeG
L3BpDoT3xo1KTKi3wacUbKWDoUo4gVNlbN2OLc9TlDV3VgF1j3xy/ju1vUHfjpirkGqp7cCcUgkh
gxH1mVYrBSbWmi3rvF/ItH6PYRS5Y5Rn6umH5YsHUzdM0foRh6ehefnM96TCXBzkwvThx7Abfeso
fsR2jMa23PrLnH2Lpo1DUY2VuuT3jEfNVIZSIfaHLJOO46Is0ioPpk4IkKcQsV6bws6BE0vpRAwU
LAEgwhcRY7EqQ/Uv1hZQXrKJNn8bDTtXE16tSzkt8I95i54rjdX5LxwFKVSvwDE2tlzpVtaEUeD+
B7rREC4WduSgFCC7ee7BDQ8SekcaCTOYtL9z1wrLBJYXfwVPWtKBLNIHnWvLJ+jakdDWMYDTUAMI
zvBbM37fm5ApOKJagH/KfLX5JkYgLxS/9xTH3fsKGdmM3chqSVvL6WJZo2FhQQJ8uZ+1fojGeOOA
/x7JLWNQyhxAQrYjX8Ysh8YRoXF3OtMUo9h8M9qEodspvL92NduhW99LMoQkpb9RnS1+jlPBB1Id
m4SPwfJEsr4I8NnZjlpoqsa1yhXBUWIZtHYK42GYP1VUJOSli28BxxuWOJ6F0EWColBMOlB+8W1Z
s94LF9bfGYwn2GmfSbC/bNy7q+AZ602iRHZ+I6k1n1vrBREVssi8Kr02vWFwwrSqsEuU2mVeu9vu
fO7Y/SqbttQOvySXGiDaxS1Xyv+2lLRsFOh5asUEt99GKB6MV39Dlnyt0lvbybOwrtzNtUQ/O8c8
eGyX4HmJrY+D9bq5kAQJ/ipWn7oDS93yC/X4G1SDeG0K4Lecy5ZptXWJ7NPXkpMJYIBh4evQDPD5
FBSxHE8gcdxfRKlckWgHxquANyBd7tscEk5ZzBBF0tRPbQotUB0/ybB6jCbPEm3IBkMDLQjnbuah
qmN4cB4gRy/f+gKPT+kOqaWGvI1R7V1LMViH3Q0IVEiPpWNGClb74UJH6LI+RQg3gcsSP/Q5tClk
JNddk3mzN++1A/hhoOlhhjVWEaSxT81soYaJx/YAfEyT/mMjM6p99jGMPT6kNjin6S5dXPi2gjdI
7z93dI/ZO+mSqNgn6kbsFzaxYUxCC9qIb9sQi0zbgjR+AtlnpUwZPReFPC5HVddYwvHujUnhpL2c
x+iF1yx4MXsoSi2D5mvonEisYcpwL36Jd5SvGicvzQarTb6JPpwmF32K7KFl6nOUXvgyRoffuMLr
WWuFP6uFbbkvvuCDsyMCCYEU2qfROd94W06JXKQS+cXiX2+cnQ406nW8V+rmQ39ul5vICzAVDO8+
UIFAv0IDiK3M8oWt9x4tnXv15F72QbNm652ybYSON5oWR5ULuzQ1U1IbvPZ98Jd0JSDgM6hM+JdZ
TS3gUBv0S783p0znJaPcdpA6Cpbe1zXWSa4aYqxTlGd3HXbNdXJKrrJv3UfKURn5qZCN948IUB58
oiAPvzV5+3KNNjofzuSNnpxFiWGZNe7qdG5AtfRvqQE3QYvJvVQdUGfHLwFO6KFVrzoIIuMApPHJ
TqICqjkJ11OnrAC3a4tJZyxIv2S7jad7YRh2x+yfEvu/bU9v22ceiYMcpFgvqn0DSHbqv3PZCZ5p
HM6VLVAzK0DGTIsx7ET4duy3Zf8iTAfJDe/XhH7aA1kxoId3erhwOzXs2WgyEXiGKErm17bhcwFs
M4+owTWaqTV/Z0NBkmAxD6PZYegC+SKqLWqLOzrFYrVHvQGHLpqBJMMgvsRPvfHRV9hGbY929hXG
PvWv72j8zJaO0I4HaUGRjqQaaDCPFF0TKwy1dpAsXA00A47wNPqJndl5b/y3fpYV0Bl4df4q5QSw
Qh+gY1CZuAJzn9Fyh3h38G/KJ5rVdfVXIR89Poacs2p6Z7BAHeMZ/kmyAsGlxoedeUlVUyxvbfKk
Iwb55irBTdgy+eEHlGWkuQWfWENIrx8wim0PN7pXYipO0ikWfsKTLsKUQxrfIUdSCt5WUW44zT/M
6kmZsTiaFJcTqY3ebRRqYUKPmcWL87wxaM+69I991k4SRQvcbiwPxAGXJj5lBKbtk9Xw/YsabqTm
cCMnlmXT1p/cJSi00fsusiFduXXf7W6M11/e2rypN8OZMJp39sWUDkz7GSMJ1XyQFMJGS8Lij4W+
+xmFPDGGCZVoPCIrckOtCAFYH595TzXqSy4q51khCt773nTTV/uYpVzblRGrH78hdejeyYWHpIcx
Wlb9QYuAzT92HULZY27mvJdP62JPXh854d6YmOiKY4WCxYJ5C37RpuMOmNWjyHjxppxcjt8VmRnw
vj9vQ+3bXzj9G3U9zk/zx2Lg1fTvtPkUQVzU58l1sh5qGJXiJg09BaZ+D+NrcbrTxh13VYFOAqCC
5fX1OlUBiSiwqLV0FEKJ+PhpUtttujD6xoOmtAqHK+AqP4bKeI3AoVHvS09GWn+Q7mNm8iX2IKWq
t782VjeFN2SO8CrBpL6CjFFGXoHrhD+Or+ijtgE6hoK1FQSArYF4B/pfi7CteEPl22HRgl32oRsf
wrFVL7XqFHRYFMo+gOp9JdhQt4Yw6B0+H53AEhR93ExkGTEW2o45BBidXLeXldmnF9WsjrUC/rJK
GY+PypqQoqOjpxr5Z7H2cr+a32L71+6YRJNP+MsUVdoBoSJsCG5CwanF5dUS9y3QcT1B+c0v+3Pk
Rh+nYDa2hCXmqphWYJWKWfqVkstobPkKyTeluYbzZ6wFw3oqf4D652vaijj9f/tg6oCmESTuuXQj
VgZQNjeZG4x3izoe4tsZH8WAmUIEOIReuYdsMN0e73rCmVAjNGtQxi78iSgZC0EIFIHwJCLYXa2T
5EaA0GYbbak+o75RIQO9CXCs6e5ehgB2vqSse/4RqR67INg4BM72ztENQvZ2z8ZUYz41q4mBymoI
sjJteO0bisoL8OKY0FRurqqn0d1cq4nHGejgi4mKKvmMaD9w2qAaRlKwPApLHhaa9r3faL/9DdNe
9/U2cz57+sU0FSlGi9rExVaE5NsE2F6+AuArPtTDEbCFDNp6vJ624LGKN6/10kmtzbdyCalsRwXH
mxod4BKQ8ZqYV5+QRphymm/1oW0bQy3N0+tcJIEdZVmFA2hz/uqi3IhLjSnf8eiNfu1aVNL4wK/b
O+SyRAW8vTsqse/FYLAsLK0Va12J+a5Up/7HPdEvrCLQvNlMLIc+lQf2hYTBYXMATa5LdSDmKSrd
IRtLZ6vAkz9OZN5znPVIjBzPCpVV04MUnZee1ZrIS73CLdwSD49sEUE3/mi5nZSHvacJX0YFUj9o
+as8rcVn8pDXnJcThZEZRcKhoY6RVTnJAJPsZ7506OYUCz4Ojycte5TZp0rWa2y8ZvyJygnnG3gS
/5GGHzjMPmYfvEVpBV8p75o45Cwxblaxsv9YwIHmAPeUG17kmb9IMIpnN8bvt5jRyci+/KhJenaz
ooXGZ+vi3Ki4cW9WnhXsVu15H4y55SqNGm/HBG1wP7csUGKX2U8hDLJ3Iwf2JUqzdKS3ZmXsasEJ
TZE19CZHnsRs/ENzi7aP426gazUmCNzmq+XX9FKEUX7HVNxWHfmeyEmwJQFd1ciC60yDtysu6THr
ALPK/olmS5W4T5uA9yVFjpEEMYbLTnke7PYErMtqw7L4/ZFrbz42fYzkdIvjY00vQcatAXg8NkWe
VgmY3zBzE1YmeyuMYUfEO+zRN/DnVeWdk4qXc1FRdpslbFJC7hx41JehBJFqTJaaiMAxqhKSq/BH
pppMXjOtz4YoKNoj1axP0gP1bfCuek7SUckXt+ru7LrqRvbKrgiA3eeiGbQZ0qOe2WOxLGYwGJne
cXeU0eih2PwiBwC27gsApEiWwVrJ3yuRsXqHTiKvo551usiBjiiw6+dLsdN1H9Gmy9U9FX+lBESR
tR77FAOybs0hPB4W6Qs2u72dj8kkPJm4FOHv1ut6IMaAkw1i+cYV90f2div94QijCa+n8kvs9CBE
A4ipu3dw7NZm8i0YcesE3wwO3+SEJ9YnAOVJH2KNwpzEksFDbsVGcQaqNhSkX33gaGc6D1sHv6yk
gjgfshD1yZJc9TyumQOxX/2Zegnw2VcFgGfqo466UrIQkc1ApjFV0nkWboRlTisfR1o+FoYhqXDW
DH9ZAR8kGJ5pyIYmDjM5u52Hc90lRJ4b/FgFhWng2xT+EWZYd8LlsWZnjhZQWOVMRh3C8BqQRmaa
pGyqg17Qlti8Qb4JL5pByy0idyotsZ6fhmBhX7D7yENGGp9wYcOIovixgdo9gGYz+ItbXmZvU2y6
zl1Y6D36Sfrsyv5l4rYMeifVQLgyo9CpVHujuewLJ3Rx33yUFvfiBOiO0HdHr/J5TvYrT77xfFl0
ZTjw7O3u7m9y3vX0J7aFpsPlydx8/iOrDJVgtXnMthsu80Ct8rfrQBXuM8n6KIcFXGxiyw0wWxTS
OGRLIhNcV4bZLJar86miiitD/GyjWYlvLT+caPyDKujcVZ8ywJcZC4DCCfMUiH7qUA0j5N8VTbg6
3Zwf0BzSIq4AmTYbWgUML5kraOds01mTFAP3lNpyrxuVgvZwQIZEWieOlVFmeiBNA61ZJFD2R4dL
K94Gsp3Kes5ga+SSLYd/aGw51JkDcKMl/UwpQeQXK1y4YFKHTvCfpJAXf7IFp8RuGYyu1kekp7HO
kyKo7EwvknVdlmk6PR/3Mo5rS9jCaAiqHXeFZ/0An+52vBL+0C+LR5e0yCiPEV/IRbCuzKblztu7
qh34KC5FwmsJbEkTl4PVPql2EnUfBCPFPrUkYUh1S45qoQbm0KNJHBgiHPgi7sfbd+2u0gHNb+3d
xgyqKswfXJP764Zu/xYBveN6itoPQ+RFWdvlppVQq0G2Mz7XCFduHcrIIwmtGu9+rObQQf8bNE5L
GMr2mwFPiAmruc4N2GL43/Xyi+/dIttlajtkLaKktBL+JQXPJd6lBBVQSIOfTqwxgOsRyjSsZRAU
DheAB9hgX4bkPezOc1zhh5H8sGJnUGSgiAcvXa5fWNjyFrJP+/RI7ElLgun0F9hEwaoK8sY8t61n
CsEYWIHSupO4OP9fMe87NQh7LmJvpR9GFSrSmyWtzGaX3t4BZfxjNpDuA1/4787sSqESwKL4fnkr
nvAO1Yn9CaE3PKpP/HbJgb2xagSRtXoHhtKwcMQ8yUo7pYmN5Q5WWsxMaHmMZH1xwKv1z3ytJxoU
sDy850rR8ChJC3naIuhPCwVRzIiwHLxmL1oVecI6wXa+0gegv4LxG/nknNoNMSeCKg8M0OqDKD5+
zOMs8cPdfrFHko8Ol6svuGSotmnG5YBTL9tkMf2DBeMNz9QmopND1EyMaKRYuQG60aetBie2+oOm
qJtPKfUSttvr6lo4xJ8GmA+8gACAQE9L/OwF/ZGmPAsjZL/yBduj/Ved9SU8wt1lG+V/bOilr4Js
EuvmE1SoUsO/EAM7m2eNjzamC0uMWe5ynIdX6YGNFeYM8w/5swoLJ1xJNCKRaLckGJPWiQef9o/1
3YRCa3bwItWG8xl70bGKli8YqX4AVQ6uqvPm0bPILtzyzlPow3LoUxdMeECBzhg15NPRYfuWXNyf
eICQJYTeHZa+GGPl2LT0Ts/DKSJH8ha9GRgfHtYKx330eKE3MnMNFgk2Cj7bsuyIFwgWkAmvVUkN
zmcfoLGNe9uEiTIXLuuaY1OdUQ5Ix4A+neHBqv/1KhhA41cppjj6L7dz46fxfMPpPLmFsX3gRwPG
quv7BzNLUHNP9s7QIRRGXnpawnn9PBUVPCp1algWhqnb2/nKBagknpvlWMlJA/KhSS/7R3idnB4N
XJdbHVgLwknhodPjPb4IWVWwBh47zJEF/arbHENW7QMHa+SlU+qxvZMUdJcixkpKoLiw8bRuU1sz
YkaHqGQoCrdCDwKKualeaiMSP5AUuEyH5i4UYFHohDwrndWrAjIhMV6MIlNhh8ZzmzHVg7n8T+t8
TX5+vBs2W6CY2qr/yHG7a4j93zgwja0Xjx7rvagMyC5Mdjhu3TE6Tj3ae3mKus+f/k1TA8zCaws8
pvrNC85nq94pGeq/ajBbeVJRhh3EEgg4IJe56uFw2MbMzty1+Yz5jqRy+rMb0ARHBCpcH5lkEMLo
F8rbPcH1kelOUhP46+epgtWMimM+dpGdme3ajZ+MhTWW0egEoAZxpAKlHuq1bp9VWNVpsjrbNG8E
BEvOeJDEG8H90u2sAgLUn2iU0v40Dyry7Gpa8kHp5gFDSSo3ZqC+YdfMXey/vDo/sggsTmF/bUtg
Hp+30UAj18MW65z8eh9XZTwwdZL2KFgUc5JPQXcq1ijCfup+RqXr/r5jUXDYi5qonb9iy0DhxtQw
5HnrNcASJXVxTExvNxMvvhPgrWkj2CvHyBkvG/juBb2yO1QuikfQSYNVvv1uW53BFz3gDJS1zdyh
NVa55NRPsy7tKNlLgI6dPVRxvN92ct9v+LFOZX3TJWkjdiNWS89nCrGi+R1P93qlY68MV8E4z95D
WlST39Ak88zs59eNb5WR5wUP7wTjiEqgR2TfT11y8P4u88/s5DJtWdd7XbJc3jIYp+V0wB9a3w44
cZq5+KoXtnH6SN+Peb2M+7IBr5NY0knupWtK+dsyvtbr3yIOHCJXB9rLLdX07P9T60lQ5d7+b+1E
k/CczKLxX2eCzVJvo6XZfEur63cAcwhc1Fa6vTzNUcc42qr7wyAdLd8dMnsa9GgLcUsZaU7uk37b
I/Q2FV5nImDN+VXegMve0jckYnpSoS6YpO6VTAr7zKu9mdtioL7gJoQvc66Sq7oDMkahTNR/RNgW
c2JRc1kKJ8xhnP3musvB+ZNmq6Baz6cLMkO/ZbvUm7QKSS/578g0Q46k8bPKKtA5MR13e89HQ6Px
8HlEpXus3MdCKqv77UASj/JJvo+ZRIiZC148qBYljg0glkjeLzH+8/OISU6HXkSEiWYNe1XeO97D
dLQ6MG2n4aGulo5f9jVUItWOLMOLPpx7menu7FNWtpuQzx2devUfd27ux2xRVFWaenag+3g+CdJF
0nnEeVafHikRjXk3h/s61Lpf9M1r9njL0As2RYrlwKifhmTGCDjPBwObQ04+uqJsJtunaPgOp7xh
3U/u5gEI8xjsY1gIPDIaJxs0XjZ6sJrGDNXqBeU0xaS7CtOmZ/jAQ1hRh3RBTa0EbNJOZl+SlF/k
QoHlodtmTC6BNc3d1rf8if5tpPF1gT0NLiajb+oFp8dnTExk3DrGfCl213HGv4SpPMgVHKo98IS7
zmXcbrISWKzicQVKl1w0oXbM5izlhmo2pMfziBnSm8LWZVWcbNy51H7p3x3yP8bLbwTwNWY45HFA
3juhUuP2KDGiqWa1YYnqo7Z1pPW/rli75zg4oLwOVD0YsDUS1BuqZ9tmmYlbn/IqrrZYhazu9/rl
+YubdNTGaiW00tAoPY5oI/qoDPLfmZDFUQDE0ZwSM3jv35FzY90WwQThEeL2PFgtPTI03XmaRRCo
vjascUZ2+xxb1huDoAxawstAfXb6iPV8AbCF775TTCnb2PBu+btOXZ1ifylPfA==
`protect end_protected
