XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� ĳh�qA�fp~���$�����}b-s�m����;WT�xK���q��7#n�4�����sI��H8��OQ{����-S6���d�@I�s��A7���zCo�^���՟E��&��G+�J���K�>��L��B�C�&+������Eb�k9EH�;-`,�1�S��h��<��ߨ�Ŵ@�Oֵ�^@�Y1x��k�eMv@�(�㗾��8������\0�#�
���7DH�E��x�g�Ye�,��P�/�����}	��L�g�����7iB� zkL�#w8�j'�#����}�h)�Ԁ�s�bӜ�P�
��s Q�kNwδ8�J�F�SEHk��{v��Լ�
n��I�i�� ��p����-b�b�͝[��h�B�����ps-�/�^�_� ���LR� ��/��&\����*���p�n�W��DL_:�!T��a����"y�?�k:�τ�@\Ps��,�&��$i�	tM;�n�K/���&��y^F�G��K7���4d߅cjǴ��0���Њ���>D�����\�g��[����-9PD�_�����V�S�(+�B�@O�����L)���'�g����%�=������W��.���M(
<���gr�P��������ɝ@�^��\��m����W�;Eх�m��<��F!�s��gx��^#����D�\��/���l��*�3{� `J�),Wex��9��%$��pИj�V�
�XlxVHYEB     400     1e0t���g��(DӚ���b��Q��8�w͡���#� ���|�#U��h}�Ei���^
�m���k��^�"s�tJeb�i>D�1<���GR�Q��>�k
 T�z�<Ƙ�ͽw�(Jc�%��Hľ��f-�ĀH�bp��k�f���l̕��{���������=��:�]��`��fr�B;Y���x��K�	莖�]��!��&���[�����/Wj���Ԝ7@NY �B��O��D%�٦����#��l��]T6Xz���(¾=<Ȓ�Zy�[��\��!�	\LT�eZ�������o�WRa�#װ8�\@��]�9���,�<H��-���	4�'R#3���m#�w���8��#&IJgD�"�=�+�q����B�==Ӵf=Tƪ����ۼ��[�82K��y�	uB<���<��]؏&�GR�c����+o� �{���w��J�XlxVHYEB     400     140�w���I�Υ6f%��rFF���r�Y6%��&�����e �u�K�_�K>�d��u��l�-8P.���<���N��θh*�[g�%W11�D� �����!D5Q@���se���.S��^
!Xqa°����^��F�Zk�:?��5�Ak��:S��H<�d~J9�������UY�P�.�7")�h���^΢��~��Ld˿>��o&�-E
�u���5�[j��r��\@l%	6[��B��q���D�$�&`�|y�N�`3�@���:�[��=�BA �����88L�a�q��T �bu㌝<J�D��;�(��P��XlxVHYEB     400     140�L���p�����n��p��d/t/�s����KZ�����A5vg�F��	�^4�}�I�S����9|L��=�Ua��)�rP���P`�hbI'M��Jk[)�KPQQq��`�<^>l�A�~5"z�O������u,�S�l<j
%&d�,�;9i�<��B�B;�c������T8E�_�FU�J�T'p{܇�QC1JDNN'�&�uqA)K,+�����m�"$C��E��~�K>Y[x�2E�QOk��|������Ob(�i�s��1��	A^	�3�?�T���ќ?/��}C�8Tt.�W���On��ݩ�XlxVHYEB     400     1a0X	fN�f�"ˤǮ�EL���m2�{��R�x�nX�z��M���X8�*�5�M�7���|��*=�jdov9M���ވ`�ٝ��<�����;�y�19�ZZ;��� 'Պڭ�}��ȶ̅l5o�r�5�A6��m�f�9=����*��F%�{����FKߗ��(�U�Z-�lP����5���Gހ�N���t/c5�I�f�`! �F�!�_S�{���)�^8U�ݰk���lV$���D�0^4���u�)O��C���jM����,���L�*�%��Q*�ģ�y�9��d͚�(E]A���VzSӫU�jM\z��L�JH%��[V�z��x�g7��V�Gk�J��=:�ބO�B.���^�m":� }�r]�I`��h��꦳L�l��6Y��-�R�� ����pXlxVHYEB     400     130�18s9P=-v')P"'³1�����{"�2Vr+4!!_�����^��봺���g�	���������onfڠ�r��.'bw�n{�e�E���e���~.W�2����E�F4�#O7`���:�Z��U��^�}���K�E��U�׍&����/X�K�eT��̠�׊�>;*%S�O��
�|ב��Q��/�\p������
UN���5�u���.ɖ��)��S��%|f6I�r�c�?!WnͿ���2��A�F.l#���%�%	B�H7E{�)���lKx���!�~�@'�҇���`J+j�vzXlxVHYEB     400     190�9�'Z���J�cb?�UH�K�o�Is3�#��ݑ�L=���5S1��G.���po��=a��g5�D�?����Xn�'���%@A�����_$�λ��,ڢ��m澄�o
F���~[��Yff��x7��c�=~W�LW��UQ��f;/g�:ךʪ��Q�.tU������-�'S۫d��UJ%�u1.I0[ƚ{�i>D(+��,�T;��yf��;-�z��ܐ֔S�_�bW(}6� �Ͻ�����S�� m��S�!�S��}�}:�r��`�x���yLaZ��x�-��2�h+`G�"�,��/�*;�0ou��o:���8�R����9Z�&�5�m;��O<�n)�Y MU���YʦVܓi6�9@X��bu[�9���㫣S��U�XlxVHYEB     400     160N��@eN"<L�C�v�ƞ�Ql�nYhtc�6;]14% <34�(�=���ؽ�K��	�^�������שj%��,��5dP�5ÔĠ���9GA�r!�5&��k,��Qֵ�J�s0����r��A���b�VA7v�JR,����.���(Z�����G��Q^�=B.	,��&1A����(��*5[m5��e=��:+�����.�G�}��S�	q��ƶ$�`�����{#4�s�iDw����f;t��v�|����}��ݚd�2�g
^*����O,]F���돭	Gp�M^�UD)��A/X7���X��K�W��B%ݤd3��}�Z��9|XlxVHYEB     400     150(!��Y����X�Yly�k[o�3��x���?t"��8x�J��Hi���G��BH����)�j�o���Lf��QM�0R��=�4#�����L!J�ۏ�����������T�Ł??�]
�JM�3�gsJGx+�4��h����[v������w�-L�R��n��'�|G��E(�7wOP^Fյ���OHO�T�f�S�A��$��8���J���Q;�6@��r-���;���A��[�]0��*��,�v2ɿ���Y���`�H��eꅸ
�\"?F�U��+_W��m��x� �f��CY�G�MuADM>Ǜb���B����3�k�y�&(}�XlxVHYEB     400     1b0:�Q����a� ����Ni���������c�9Z9#g*]n��HI=g��v��;E*�ir�+́J�yv�^qE�E��~�~��6
�z���6�ӱ��﹍�����kK����$�v��]ƜȔuH�qĠ������U���6����Ȅw*�	E{�/N�)�(�{��]7B��>����'�&�&"�!���P��c�{=3����;��\fϙ9�ݭ�	l�ꍝ�Ns��zd����Z��/�:�����mQ���_1���3qX"�e�P쬷K]U�x����P*�r�'�J�`L�ߝ����kօ�~<E��n�x�U�
�,|��D��@QΖ��ԫ�6}�� �V]�UPQbj �r�C��]ӱ2����1L&T�ǇK�ݲhK�OO��D���:`�١0�B��@����z�~��XlxVHYEB     400     1d0aǆ��(aO��=I��뜊���k���Ut��r��J�t�wP,G�ws:0#{e�b}��~��$;� �M{�d�v��M��`%��E�}k���O=�!#w���w��.��SBl\��� 31��'��_���]��
�zI�!��K� �:�iI�����[��1��0>}���19��O(��狄��F@�'t�Ŧ�:m�F,m�tOjX瑽�p�˔�;XX���	�G:���B��=]8�r��S>�i,(��"��x}���W	:�@����lRR��8�eCU�hl��O�=>>�A�xv��9ԺR�m-��ٹ4NTE���}�T�j�W%n�0�K
�L�9[D7�Y�_��}c�ti�0��%��R5�kc*��a%�r�T�27ܙ�����ã�r;�ͨ�s���0�> (f %���b8d��a]�$ƥ�_��o��M�i�g4B*��	XlxVHYEB     400     160�� �ˣҏv>����>����V����Fd�(l�r����Hw
^�c�i�,�G�;/�r��'�5�����FC.FY��.zaߕ�s���? ���`k4������az�T��ӿ+G��d�5E�0����+A���..�˓�v�F٣�
"�(�G�����E��3����2��ҧ������[��q�&%J������F��xdy��57����{}.�I��������G�ڈ�屟m�#|'*_i�������pk���?9:��P1��ˎ;�+�Y+��vI��VZ D�1�Ɏؚ$+���tj�J+,O��ڜÒU�?�����q�r) ��0�J�d�L���XlxVHYEB     400     130ӫ.$��� ���-y��w�+p�����^�X>�����K'�\<�4�,��O��[6à���͏�D�q��! d�6Nu�=v�תG`k�}E3����Eܯ}���Q�>^�(�.8��ΈLH�"�~ѕ����r�?3t�Z�gbq�J�a����+e�\�[0�$�*W�� b1�Q�D��:lR˖q�\������xL-U��G{�U�=V
[��(n�M`-����,TA��Û�e�Ø�������y���o,�1��m_7�E&q�	?�G#HK�%@*�g��,��G��>V M|��6���}\�XlxVHYEB     400     180ץ'����I2 �`$Y���w&]9�x!���2A�#(� Q�?"�qۃAY�A���( �x���C��t��=��oB�4g��e�g��w��" ����A�3�E�r�ѐ\z�(6���i���q|v+��W���X%
�C����v `i2��@n���{�:x����ο�,S�����U�A��x�-�M��{#F�if�nӐ�����˺m7U"�o)lle��QXm��+��6B��͢�B�JNu.��ƕ��[�r��W~k�3-f��f��l������#��b������?�άN�<�&,%�)[���5����O�� �;F�!.�r>`y7ڐf����Xu`�sBVz�/`G�d�L��Z�%�~�f��wX���XlxVHYEB     400     150�G��Qb�<���qx�&Ʃ.�L6�>A�� �l�5jb�r��y*��r� EP��	�:XH��f�MMs��|�J�[2О��9��$IW*���hS�[%�ڑ�7~���J��$�����R���v:lk�bR1�lD��O�!7���5��e8A�6S1p�^�{�����N\��f���Ҋ��Q�3����,���m�"�qd,�m�WI�8b hnv�E��sUWD��3ۓ/�=eO��5��Y��p�������H�}0�)Rωv����<N=�I���>��-�	��I�e�-�|`�׵b�m[�J�)�؜ �g�P�XlxVHYEB     400     120�av��G�;��o�7���(�-�k�!3Z5?�KSz�'q��GZ�V5�<�z'�Z�^Ԏ
�3��>;��ktt�%�f�p#$�q�0_�����h�╿HI�8���h# �����B5J���{��V�V��rv#��
.�؄��K*� �?�(�_�=��0:�Ulޱ��~�B���@0�ct�Ve�K�LhZ���� w�.�p���hA���p�Wt�<�~�jB�Tc^!�gS�P#3���B݂i��2T֏����ҭs=Z���\ X�n�XlxVHYEB     400     100i7�o��p\�R&@�GCy&��H:���S~AM�|�j�H����A���/̔|�AϢ�w�*Z̯!B�&\霩)�N�Z�#�2���#�5�@��b몆=�R��٦��OFC���sڍ�����0���o{X
d*oz����d�d{����/\�����vgYI���F3:��sJ��Z�'�iR��CO��4��v�С�3��M��=�>�F�ڼ����o��[�cP�R�W�ѥ�\rXI�����.?�&�%XlxVHYEB     400     1a0�)�yQX�ֱ�5�4����$YE�y������M��ѥ�o�BՔ��SW�� Ŧ��e	�g�0=��<��nH��"��Jع!��W�Ŗtl�o{ߗGKj��q����
>��i[��:v$74H��[Ub�<]��ŚP���}�r�7�"�|ygn�����DJ$Ka����~h�I����ڔ+�۱�n�51��qnQ05��Y?�)���1V���8=�^ ��4��h��(��[Vv������ןu��M�>���n|H}��~���v�Zu�{�Dd��H�
�5N�̓������O�����w�aG�AkUQ�i�N�(�S�f2Nl�΀}K ����ͽz��,��
N��+�O�q��G����-'F�~�
I�J�51��Ԓ�t��`R|Zh�#cw��7T���ʊzXlxVHYEB      27      30ʡcZ����!M3��j�}�`�������`I/BE��Bck���4�