��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��� k�X7���A��y�Q&�<L�`��P93,Nb@a�̊H36�q��OW�ZC�����>�o_�}Fp�Wvi��cH0�d�_�8��r���sE�������d�)�]\�\�(�6þ��u,v�����F�`W����#��7b���r���(E��1	��������mKEۅ�:�#��[D���;I�)yIS��0b!
�/�b�:�n�k�2�$�+μ�w�/D�w�1_�4�r[�OdlBڷ��q�
�����#:�AH-�y9���H���*��E��mR�8�����s�ѫ&��N�uvv��n��G�� ���_I����L�{�ZQZT	����gv��Ù��8��b3A����f�����X>D�cH�� j\ݵ�n�,𢌢7:�![h�(XOq���:4HUZ/=�2�RE��z�^v�0h7p	����������@����~�]����A�Mo��-��# ���J4O��¾SDZ�e"ćS�Y����~�G^-��/�I��8%i(|�t�o��[OG"��e�1l����c}�(�P�^uu���D�c��5$���MsJ����2M��e ��`��L�>٦�M���D$���.��W��-���#/�Tg|l]J^_��C�e�cntk*[�$^0����iD6a�#1�	��;FB��o�Lb�Rd�m�+�� L��%釶�FW�ũޢ��.I��ᝐK��UX��^�mo�6�Z�9����C��S�1�e�V�Qu<S�O��p����w�������)��F��a;+A����)�������V��&�lbC�Be�Ҭ�Yݙ��3 _��5n���Y��R�u���P��ڧ�-�����(�*?�d׀n'v�D�Ѫ���Ei|X���mZ���R0�n�.?���_��03Hg���g��h���1i"wE�ei��&�c.?f.�Jb�� � �%�ԃ�=!=�Vs���{�1x�0�4o�v7e�yT������U��7/�!��z�H9X�%0���]�N �h����ڻ���ì�����Z�9/�f6�0vq�\����&[�Ӑ���J����S��{x��P-M�z�Wr�f�2Z"ְ4���$*-��&�l4qf2H�3�m��D�>��5B��AЍ���(��6[�i���yz/�|�-E�>�	�5@���/�E`�34�==�k���__���+�S� �,ݡ�����!y+����gH�r)֒��F������3�}���O'�b�����Y�j �	�̪P�j���\ȉ:sd$`F�Né�vU�v�۪�D�&������K�|�7@�������5�bb���̘B�c �zB^wt�2p�)�/�)�^���rFN�ͫ:�Խ����2YV�mS`]@E������,8���E��*Yxd�u��hgDy	�h�I���v1+��m)�V�O���w�C:o��n��!�s�ek�8���>y�:]3�(ʭ�Ѩ�wH�<\W׷� ���4Zl#΂d;x[�N�,��&�