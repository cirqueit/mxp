XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����C�UA�x?�կ��_[ij���N7bzW_)�G�q3��Gt��������.V!	����
�u1�(�⸅��蕒䨔W��c���$1�ݶw	BH�Pp��O�E@���)��}13w��L ��GE���ٞy�z�>V��&¹]���oW�:���^+<͞q�©��M�k�ȴ=}IdN�	r)�	�=�V�Q��R�8�)`�����ܘ�"h�p��<EZx� ���L�_�����I�	3ю^Yۄ�zlt~�;҆�,H	�[�;G&'J���-'��X�քBژ3�(�������u)��Z�������P� �D��Y� ����l�=#6}�^��q6���TN��������r��=��vk/����ƀ�XѨ!_������:�XOW�g#�uaߓfQ��������4��Au�����5}�;{V��)`�-��ECZ�U�Q�EB	t��MyfA�;X��쎛��g
�PA������
Ҙ|�d�R)�ϼ���9�C�$]�\�a���*AU����!���e}ϕk_4�WFi�Zժ���.r�?y����?G�/�7�Y2OT�4���)|Z%`��L9�afƙ��Ym<��:ا�v����[7��{y�U-ּ���
�.��D�WB�7	z��O���o�UB��<�VV0u�؃�Ixrb��u1b�b�h_�ǌ�������� ެ%9����<I�P�G=�mAa���ɔ����_�o�0>|ܳ8w��"��T/<�~$�XlxVHYEB     400     1d0{"��ى��.�jfY��mM)z�8F�l0�R��|%]���r�+km��G�ԭ>gC�=R��XI��ޚ&��03�<��(,Z�Ч�~�4�J����Qai-�2.`�.��N{r�`4�f�)%���m���ZO�%�S#jҴj�Z�\ێx��<Q�`�����8㰛�����֝G�����6����~�Ư֮��"�6Q�4�#�:5�}���^���w��I������������A����?�ʖ3%�W�aV� 	�W��0��������DӶ���C��S&k�al������z�d�G�y��TxU㳰Io����[�	���ʂ�󩒣�+7�$J�+";eS}C�~	y[p�����\���M)�i�B���}��ҽ��Y
�`���k�R~�5�K��1��7㵺u3�v�Z-aX,:��u	^��<V��y�Q�rdh�r�m :�rXε�+��zXlxVHYEB     400     160{���i<�]>����İ�6����/xc�$�u��>|�xg���7L9�ps��Bjў�f�,����We�W�4m����w����c����q���G�=��T�Ic�<��,\���bӻ � �.�$��(��w��ˌ8������Zb8�{վ�1Yx�Q���2yӇ�"��JG�����
U�y�>�t*�$*� �mu����h?�L�ǧ\	q�%�����)\ǝ��{1��g����R��̲/�R��0<:�=*���P�8g  xe��2��*C�C�l����O/4�8 9�6|<��jE�P�<ڽ{��yP;J�@,��B!����*�M�@XlxVHYEB     400     110+��v=/6PK�o�vn�2�P!e���K�fP��F6��״��o��U[�2р��8:b8W@O���未�B%�Y��T�c��$-�c	:/���pш�ԙ�C��<�c�}�w�FK�-_�C��¯5����*%�R�%8��t=�����ʮ�o}��f��w��G�.[�����/�p����"�?�G�$uVc"�����vS�{�8m��T����Pب�y�}/�i��9a��sG�?�Zd���b8C��
�L��LXg��IlKaיXlxVHYEB     400     1100��+��i]9�4�.��-���^�HZ<�'����:�P�Z�d<R|��3�δ�d��~ַ�F���{F�<�
��:1���N�	�s�:�c�0�=�Q~�:Щ,d�Uυ���2z���o�	e�65GM0*�BR�� ��H� ��BH�&2�6�w�'G�Q���Ú��h�C5`X�N��yAB3H+��I0AzT��`���خE Y�B[���A������g�&;n�6%�����d-G�#"�
�(Q�F�vư��
�c�}Ro��XlxVHYEB     400     150�$���� !��:�D�����ɯ۰������
:?��{� �㞣�ܬvA�w�H��F�$+��R��m̤r������wo�3���������}�r��?ю���pO��ҾM�ApLqS�+$u~E�w�{�M�ns���U�/���I��u���K�S���IѰ����5�8g���Qޏ�VTr4���r�b*���m�����N�s��.�T��Qs�h�&�O�P�N/���V#ӈ��v�ءa��_�suXU�8��t�.�H�16�g�o`��J�5�cV��hx�a�m�c�۰dqIߢ�+Z}f�XlxVHYEB     400     190��O� �G ��u�`qllT��{NCP�FE%�0 JS1�H�����/e�}ж����+
�O�|��:�V�,�r�?�q�����<�?�9>�>��� Y��B=;3	8 �4ղ�7п�D�}0�����sF8��[�sL�R��-�}�U{���M���RN��$2W#��7�tv���K����Ĉ\�4�J�Q�F�F#��Jo-|�߼/j��۾΂��X�H�eŏ�	�M�0)�8U�s�[�&2�mXe��^L��&�r�d�&�!�%�>ƚ׻��l����� w��2�����[��T�|+�-��pW�㘌"�v�$�s�v�	�~�5�����a�X(ɚ���o�l��Z���}��� JJ��� �WR��"��K�� �8j:P�}���XlxVHYEB     400     150O�v&N�����'ǝ��)�c0���s�\�[�F��.��Ǫ���B��f_�b�
Mwm�d��4]�P�M�sgF�q)��t�zl��Y@�K�I´��+~V�Uz`�9��-�"X$T�x"��D��
�w�R��{��T�=�_����%ٜ�{��e���4����ҏ��t�V=�-�[k���z��@���й)D�V!�(Χ%pp�U����x�
�n��+�n�&L���J�G;6F+�{$�����<��1�����7'ą�5����U�ق��E������_�&��iD�݀��T�9E��KK�J�5�]+��uC.�DSXlxVHYEB     400     160K����Z�?4�xh���f���gyQ[<.������(�ҺF�].���8%R��;����L��u5���6��B�%w1Z;Y:��� �����abX\�O�o�Hld�L�ZSD�7R:h����|>g�N�Eb�u�a�7�JLdo��G�ukW.���3ɗ�u�4���UI2�	ʙ"�E�z�a�v<�j�o׿/I��(%�A��&x{�t�\AvC����1hWW ^ls�r�m�j5O���z?�:��`�u9������W����(��<pӞ�5�퀐@�H�$��'ғ�4��~���e�`|���_���w5�#�#�\U�4B�S���w����� �z��&�XlxVHYEB     400     120;�+>Z�b^�6F7��3:�Pe���\�"pn9*
 ��07Ǎ�W?�����i�AE�i05T%<B���h����"g�B>Z�8�C���0�n�y-�э����2�a�\fAv]}"���j���&��t2�Q�:{�g��MNҡm��l�!�p&)�|q���G)�[���ް��&�	O�� ~�5̸�{IC8-�MRU<|r��{~yN=��p���:�A?n�Ĵ��Q�®aڧ8��ۢ��c��TVrk��$�k��Ղ�e�zۯ̌3h��E�#=�H�=XlxVHYEB     400     1b0S�3�֬�@��М�r|~������JV�tAZ��Z�� ��Rl%��Ȟi�G��O4�Ǯ�W��8��uQ8}�Զ��>ȽJ�F��A�M�CtC��ӑ��q2����Y�g*�A�|^�>.�B�[;��6���O}�j���9�0� ]7�V�H�S�󵿚�d���ʇ�,o��W7-Z@�Dg�a+��;��b����8;�M`�Ii�^:�q&��vc(@�冖B���3����Ot~�b�Rrl>qu���|f��ޢ��<D=��v~N&����R���
��59��y�t̛79�-�HH��H��t���Lr3�D�ث�0�sEj��ĳQ����Ǝ�X�~N�n1�1��s,�rk|�i] D��m �d:>�G�U�.���deD��#�@��Q�(z������܂ڃ�sj�Y'a3�6�XlxVHYEB     400     1b0�7�K�9�T����I9��\?��4�����6`��}$��p=�nd��ٲb9Q@�D_	�x��"�S�)�3��GC��k�!^�Kz����������Ԕ�d�G�o��)Gv���M�j^K�EK���a��#�(E*����m~Q�*o�����-�G6��|��J���^1����WI	!6�.�%OuNWZC����j|�pc��g>��$��v$��V���$�#�62���#IC!����O`0�{�=t�L�9���θ�/��D��KQ	R�9�ϩ�q�]�����J��K���3�q�|��h�.÷CSm�S��q�Hg=�n1�4X�9�tT����;ICD���������؅�MWQk$��H� ��\׉.��㺸\�}"ß��mu-m�&s����
n>���;u�x�^��fXlxVHYEB     400     180���?Er��х��^ �����1�1.�L+�+w�j��6���ZK
'h�*��@�!��������y�qp:�������G��v�+-��
nK�~��dC�,��q�4o�LN�z3ބY}?|����#�׍q��{+������tDx�u1x<NZ��iF�5�߲Ֆ_%��n
����,R��Zg�ȳ#�����<�$ ��f�SR�,�ӔST�����y�������Ϩ>:A�>�� �[j���Ю�ը��o!!�/� n�������3#2@�)2 1u�-�]��p�>���R���R����c�t����sy��)"Q��6��LQ-�65�V�Z �
����8b	z@bm/��h�v�XlxVHYEB     400     170Gl_c���ad��蜍%��ϗ�Fx�N�n�tlW����K����N靻`�2��3G���:I�Pv-�UcY{|,�����dZ�����X��\$b�>���T]oI�؁��i�Y���3�8��-w��K�[|5�Ly����W��=�ˊ����l.Ŏ2J(��o��~��烾�x=�ߎ`Z�R�+�6�6΢�q"�(E������C�D��^I�oT�t�#7d���#?4�b�-��UE�Hy�~���/�7Qt	)�ߟV]wOu�J$ՑuV�uK��ͬf(��0��l�X2wA*ԿRWA��4��[rb�ϑ�z�2Kf��c ʓ�l{f���D�n!�󿓁M�<A�C�z�����"�J�����{HXlxVHYEB     243     100��}Q����ck��pC�dNA�/�����[�?��l��/ �D�C[�2�+��d\�g�ĺ�z�X}u�~B�'9�p-4��+�?^kV�-|Sm�9�]��@�*�u ��z��謵R�үȍ$(>w~T,�{7&�tO{e�Ek�a$0����p֠��ꌃ�Cn��11@J}lЂ�NPٟ����ӈ'<�.���L9'36r����Q%�r��:�V[����}���0�����K{��k