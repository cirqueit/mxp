`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3088)
`protect data_block
M1mmj97bjIk9Y/mx7/oi3o7EIpB9AV/OsedkTXdT1GmmnIMFOrYvrNvNUufJOzU9ux8CdBPvp6PR
Etl1JIfrHKrqgzPDq9k6XNmi81awJZZUfwZX8+bw/aV9JxA9KzZtMnp0pfmu8cYxPHrWyhzL5LOS
YmNt5VAHnj/lSbWMjIaR1R0jI6hUIaaqdcCDFibkvcaGHHL+qFnMfAkRnzKnaktStQLZ25rYHOAo
8+/tKh82OQys9kEM1QCyfEXsbCepyE/iM6dH1PVWGaXBR89UeMhkSAtuhiI3T6F1QneyqN8HcOVw
nAuQmjP6sH/TXjPGrNFjKl62CRlrdIdy6bFKaoDh+TSiKSM+jVY6wD2pvYZPt0KUowBAtOMskSxL
9zHSv0xl3QebSAPuElAxYwCYpLbSQbrIxsvab6WUZrqBJhBoZWls4f6vlDTXClu4aVh8ET20mVJ6
WOin3LfsGYITBkBJ/JEJkW+PZ+ZbMw77G3Z8pQpis+YUKZOc70Pra+xV7eoaq0dcgK0S77omHJw/
kuwJ/8cJeFYlA4kU6rJDsfiFhkCbnWxYxrW6okV/LQEfXkOwvcZ9Eh8JRd+qe3cIFS7+v2otL67f
S3RuLXi02Hex8IHLTqs990//MPgOLcvTuSr49QKzAK4AbgakST6p9gqwQbriJ1PbIqoYKWLu9Z/V
q0rfd7GtGlj5NfqHeHtOWg9UFwrXtmnJCPXQ18e9J7fPmd+KTWf4rkaOmB4XZ90IdM5wDUC9hRJf
YDqiJyXwP42krPRW8CyH6x1lMKG/Pf6VrqNCOP8JZ++VjHvfDyG8Zg0pCg1I0sjMIoP/7+YR98BJ
WjxHz7qctrMWynRr94R/CUeZmm755oD2kF7oOQW/LWs8JYZbUjkolo7LNgJKXPWpKu2M/Rd6lO5R
4V/d1XysB+i18wwCzuAhSpHeoh1AwP+fVukv2DfW62Zllofi6ciu62Il7uvrU9gXqaefd71WIFOC
D29tEtv3EVnjtmlyoaPJIAEv6T7lFy+OMZP21AdciK4N0CCg0rNC4ZI/DYsY+2H1YeYtsm18AsT9
yRC+JtZA3dxI+w5jAHZ4+fF3kUHVHFWNx+dKcitwfrihOpODgK7PZGrMCu7ElWGfA2je/sf8n7rI
kGt7saMwOnI16X8BkSJPNKh4keZtRlgVptZi/NkcSS4pps8RnUaVz4F4fEpm5kifvgO7iwZWXvxe
/7RGDNIa7I4K00Hq+GfMvcmdazy2IpWDEAFcU3jX3xqFbyL++qfHU+WLuxdgMbpg8INF6G9cOL3E
yS50LqgjFyA1fCCNpp760kjYrL0zekgn9ssUSEOcg7yGvlKiyMi9zDVnjxcMhZCDteC2PewkA4uS
RNkju9fP/DdWD7xcRx7ePzBI+ukI4RkgfCTMijcfUfb5dioklCwr5rDY8RmvtuV0cpSCZgHY4rhz
G0+uydwy7tHqEkI3lciJMw2mCMmB98VWDDhYe1Q9KqV/LzL2td8agUtRQz/CjaQNuAZSQOEa5DTI
znMd0iRnvcSDIn23ufRajycVvIZ+RS5hJrbG8AEzFrr8nk/dmFF3QgHdgpfQEzg/llFAFSa57vG+
87CqiHtUS5stMAUqrEaNaCBoKZ6XwPjADcIGL15l7uVTbAtooaDd0gpx2VMXQhAB939EWd9kpy/S
J3fT9AaJl/1b3U7Ee9HZGp8jJROdTRNighfBeAtTXYIgdx7fTfc7TzmAluFAOyA7oFSto5Ald4IO
aSTyiRK9o0p/ix5DtXtCUUu2c5odPofr/je6AEk+vEi3MapLhAggll11/gNl2c1dJmzmSEXQ6AIr
+APJQHYAxYVuEKENH6kTVYgjuxS5ZPukFGjFCHIrsRsb2ulKc+8YSpjarKqjnKo9nRejahTT3WgF
HiuzkTZXQ/5kwbtZmxnWq09tx0B9fN6dtxzATb1CEBkdnJ51WzbdyzSOP5yGMpx8DKLSKviJTVwI
c7Nnlu17irtrisedT8QeaG0mOEU7oNPR9EAIL/1cSzWA25C5GBhi45ZB1mMjM952X2CzqQ/pR6sR
mmHeMgdQafxodTpY9RPMTqlHeEHvXYqnUPCWmMvYQXs5+R2Je5fetbaSFOnescGoGO2P5bZsKyAd
eV5PHSnd0bbteL8UQymy/yzUAIjUggKEowhooaBkTCLhMlCb0j1ID+BLTgiNM6RouZ/hmsOcr8Cc
SysBXgAM5xBdvJAHoKwIAw6lo76KGlhIRqzMNhXvZkXzNmP25gMH2oWqS0RVQYuUHHblDL/DquIH
Jo2viOweQKkq1RK4I6eWt4AkRNIHRxgBHpYVihUW+s05DzLyOAIzx50j890J+iNUtTRdjTAoR77J
1Cd77fj9PPza2fRoATGJ/UaZj1pUrzhiO1MUVmCsriT7SUMFTgLzHQSPHxxFyzwseC71i0YHkRyS
NyZIeAlF9Na0Sw7CTJOCxW9PW1h7c9dTEwMrXf+zyI7gDACSS2vjqTjOurxzk/KZGv0s7ZQJkxwI
7JzARwbguWAxJ4NW4r9m0GMVKaJolQR8CF6yqDL8H+/iI5SeVzAP3Ee7mRZTNwzeeAkM0fIb47hD
Hezi6LaspYm9DZg7h0b/9it/KDHPRNb+jU70cnPsUSbXPjT2LuhcJM4cxrcCQZiAf/6RypmvF4bh
VI/BIqoA9ATrnrTOMkMks0OMw3A690cKGpF82A8Kv2TPV6qxXGMma97gQuv/fp6hQSmeqmaVcQh9
Mnf4ZbTmYR/0TWEPQHLqAhO6J8Eq9+ZEYaxtsl+GO9gFcdqw5Sx6qOoxWt05G4Qmo5rXg0oxa603
w/KwYhIq75aXE1M6oVwR0ozWXKEutd1Lxaf9wbMjFEClHsIzSdsFBIOEoEmICJeKL6QryH9rrRoy
edSgTiQUSqh5FQeI03URyvVu2mGkY9q713f/9UUYSGKn7GEjs2DSKrgUqx2obHs+XRPbGUU9SiLa
t4oaEKvASAczAzBMaD/93jVBSmnVoRZkNxfIbVQeUmeoZiB36wYDEmcFhR5LR5D8KbsyDRjqoWx9
8FrIr+rcvGpD8QKr+Nd/n7qJMyjUAymmGpciLMOHFlSW0b8K/53BCUpwyTUMAQqNN3cAkPY8gd9H
eVcSprtNsjQo6pANjzc1EQ4sj0cEJvSCNVwc48X95fbNuVae9H3X5A/UCr6rzZUQo048TkYjh19X
IFYQ/IPUbCDWs+Vz2wCTQQvwTvj6d3z5PX+ujO77gSmd/CKh+LYeSjf/o7eVJz75sqc1+o+mXlzt
INFwye6p6G7ZmM0IDP0Dk77b5Dn4s5p0LFFJvLpD2+aOfYUv7Gk0ctqvQHGLPVsI/dvFLid16Kh7
JpoE6VcO8zanuV3V/hRsuzx972Ag6HcTZgC7o2habvdr5J/smkBWISyuwVEvlda+7SFKj6d9bRuk
H5wYvDJU8kK70hJb0GdgdrG851zqR+iIjKFTHfTH6yOViT72mX/4ZQa5kxeifmsjs8m6Mc1KPHQq
osTy+0CCwjDTrv+wJ961+i1CT8X8QI08kEVYmI2fskMlvL1o1hhHb9jxbIEPehgcuXYtlXnwuHaj
49I+aghZW3gFZtllcBLOIq6FTiqMfrZL/SYJ0s1x5uxJ4cneQmohai2LbGK6jCl4PVLj8lQPMvUO
3Zj69RF80T+2YwQl8vXCqsob7xR6sbIrMqXb/RoC/1DXV/pUzrnity8vw6ghPqmybzJRUVLrlcRQ
BJyGMWm0Lpq69ZxhyvXVQJWv/FZZd41QetxR2Wq66xPeCEHVoFIaEIHGfCvCunWLlc7Mi7hL40jX
IL9BEQYCmFtO9e+oYbG98wvIIblDAwZ2sYFLtqyLVwvMnPWTqDNzQYVgxnIusC2pTcWEhojECIsM
2d/naplX5vFG6as/tW8etDJOZGQQVkkRxqhXL4yKIKG9j+fQmkzb5OawkQXgIPjn7QCDtT5fLTZj
H/zceetRo1d+vw1LAa7FH4hO0d3QW+ikJLVN1wL+HHo0zVxi2nzz0+AVF5XqELdWO9ekJxz9ArWb
TnlkZgpzwLGZRGvfTVg/Fyny6MyNp+31cYlb1WtQ9OpzyDPSjvJN2pp7sqZaYteJCz7qyFytwgnF
0PxkDDJ5+eCqvQ==
`protect end_protected
