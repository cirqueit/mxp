`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7472)
`protect data_block
El579DRdD4PBMUVxUmtLh5nLMGmkED3ZJYY7Hg4ggKaXslLR0Os9AMpw+PvG4fO6GD2VrWUwtmyU
DN+X0GrGTpxA+TIg6h+1IwBswgLWTMHN55XPMvA6ExuJEUrcHXPIkwCfZ8gN+ijRHtpzVvIJZpcK
gRbGc6haAu3ivuu1f3bhlHPhckdZGzcJAgkmyaBrPy0VoawKc6ynxe6Pq2SN/5lv3ccpiy645jmh
NOhbdsZlPcPZI7rFTmv+Srj/YY1Sm5HIam1kho5AXJyoLR0TAhMQl89eI1r2LUs9KRWbJ4Q97V9w
+oUHDR99qwmBcePILMHA5/TcbKwU8iK1xrXK9rQwbmrX+GUYaw03M23qsQJNvwnnD5TJhPaIE6t1
dDCqi8yP/O7OQyUNrJHfrQQGIo8zELdEDtr5aKRHz1mISA0GpDdcus+rCSrtCDTWxNKGUER4Wezb
C1KKCDzX98cOSZEk13gorMq5lyRansmRuTvrNK9tjfJjVUV2yljl1PW6GstJeu4lkS2Xq9WTXE4N
nfeoSBqmVO+PDnnyV+PRNSZDmjOqGQ3T/oPffWWUq8iJOKT2mGFKm4sm1WM11HzQg2fopm6reorx
8eig74L1yDqCJHo3dWQ0/fXDDZ7Qw/h4A1iIym6bpPqWfHq+moI8QyBxmR/O5yxu7G3p7QuHgm7K
PR8Vd8QvbUbX+Uw5Nic9P4l1eALO5CjDLCFl8J5otCtm46lQsxinZAqZeG2W8xyH2koxR9X9ZZVL
blrKFUadFyuacUAs2iYNlgHa60tdSq8cADTxXJWGW0LWxbVMZOtVuKJrrCghxyskAF8b0+/NPywe
ryDWkCmyrT3rWNAGIlV9yAfxer0mEv5zAwk7UohiS1MuUBuGEAXdDmNYcKQJ0NF2y5e3rn2X1qq5
7+1AipcCfirwYayY2pUO6UO/Slmtpwjl/WbrNq2k40KyhVDuvOiQt2TX9Maj9ci4nLphK7GcA6+h
/ugu8zn9qj2vh0F3Xvf/9/j/4RhnikDHrRpO3GP/IZTYg/wd2Mn4vcCWnESwouID0f6iWDFbOAbP
D3P8+S8VSm7MHX68eWOVevuFUOxyIRLW7k2rN2rWr+Ll0dacH1ryElcd8igxyPNL4iyUJAAf2HAQ
6YrlV4FsmsK44V9MqM7xSbmU/K4+GdLam58aOgsBdG674aTGMOhi26D718id9Pfy6JENmTujwasy
kXrNfjKyqmw86mPFSCXZlzTKR+dDBuvE6+f2y28Y8L436R/ChR7+b1pjQfGZC2xegBxJVmQ+1I7h
eZoj/c5tmMR0r8v5HtuzbZPNs0elik4223gQghpxcz/4k0xfK6NXEE/cV27CGC2ke6RlPbCMZZ0K
U76qtBKqMHFcTqC0rIpmpY+ObtdSIeBKPpl3kuI59S3eeYv1vM+jZJM4STsUt2eSibj7Z1Nlqpbn
uhDfzIO6H/r9r6XDzwNjtCkqQdR+NQT8FMoKhV62cjV3IEtPef2qt8ChWUCjMQaiiBZFvRi9u8ti
BIPPDBfvXb8jxhCt58hk3XWGFkDKo8K36aeHSYflR0ulcB7nQ2McqV+jwIDUcyqrcztCeAq93GVF
vjrNGFO516djorwovTwCagOP/PNNpZ5tavDjLX1Dqj3Zi8ljPfUX1cWruDc5gbRjlFighsf/dNpP
R36S+pf3smCg7UK4rJZ1bHQ1byz7zHXDq4Mz1IeGa7adfgWFvvED1cB4tGZcY/GSGhMOhifqv+vt
s4i0ZmVzRnfaOWhKxZWdlmt5X6DkIc66MHjCiW5r5BAFg/AbLo7xG3/g+Fi+ePmr1HAC+6950rnR
89uhsBviWBoNdCRKSanpxTeJee6lHUpJDtPXVsK/eDwoKbg6z7hVe+Cl1TBb62IKBjuOrWkfxD1M
A1iBP32u1+6DOeVx2968HaQRdCl60oeKskV3Rs9lqG1xJjtrnUAG+eXQcKX6qwCaQnMi+TkngjtL
XNvkbk8WLkOQbVSfSZyJY8gbs7ed20uvy+aTgg3u6oibpn7hIrF3bDaFp8xpKJ9ugP0A5vh+WeBy
jH2jmEqFEpvt4qD54RbkePk7Xtu0PmG/3ElgQhgSn9lJ/koFTrfaiY5JsM0PklS9yahsjvkPCQrL
YYliFUqrT/HVO48YHdqqGJywDBRyfIJdObldIdY8VcidUyAqZVdme6AI+R/WEgoSIChf4qH9HOcq
S1SJpiHwd6jctNM2OXL0bqSJog/5rOSkHmxsD5SZyiiQQveafiK+I63luqUEhSVoMNgenJaeSH6R
zmCXz/WDyc0SpGO08nugtKeX+Z8hQohJ9tjH9XcXqTeXJ8JBuLNUrkiMUU6pQf4zVdLf9bZdnZcH
dA+mxL2IX3eC4GQNNdaOJZdCwI2DewMyqkEKhAl9gSWmdHb7VjHiFG8egtADFkDpI3BumWqiBUL1
gsvfLKYtPsERZj+iAUwWvAUZAlywWyT3YBFRy9/0NGZ4hJuITANda+m/Gihc6z0O/xTmiS97Wlbr
AWqZMOmR+5QIxYReM9NDliYMCtOu2aXyeBdV9a0bPRlWXqeKNLUOdy2Ky4ctzJoUOIy2akNzo0pc
0n2pusvrBZ+cph3q08IB2Uzgc+KkTKQM7Jp3aroGDLALwwPztJ/8/Ntk0QecPoNvzA/NXotWX6yq
zsdN+z6JDlA+FEscfB88+bPxdJycAUT2E108E7stttB+rZkOEH2cIe2XdP2oz5tO12HA9jE3BUYX
NSDYsInWQhRN4NhzVvoK828FZ+Y8HcyIdllec6R5GBRhXC4lypjPmhR8rJwGSShRYjV/HznvU2cs
rS+DIJnuJvaODH6CTyQCGr7uYc1YQL5F/LKvALkj+Q+DL5+vc/uPTGfabw2jGBs0I8oE8727P4MT
7n1qNqv/I1CzqE6UCMEZN2jMqBZS2+a3GEl/+pVfOOFWowdZ/AHMLANy1eH4rzrO568l8XbBrAPH
4JsTPC5qFRH3O2Sz0JL6iqBTYotxHb+AOTliJtbKURzjvTnaIkFSOO/2eead57ReLBk9Xf2/yG+v
ZiwLUhJYQQTa0lz8wHRKBtYrPC4tr65J3sWHi55gfp5y2IAs8SaQI1TO+CueUqjOQ+XlV5nGEmPo
+BpdJYwHyX4BotInbYLcx9WkJLwgFOyaFfnOvgF6zq2sOdYfDwBoc99USeED7jRlWL+hjJwa+h8g
Ygo5RkTumrMTX1jlBGtzsxoq5r1ah4eSttpKGijt7UaXiZX0wPkc/vgB9IEXUviDt1AumHWZ9d3v
LGSf7S510bADphhKIv/0Pu/+Hb+9Q/RVjbj0w2919fKaRm69q/FmDqvmNwwu6H72+lEhM1P1YAR3
gsILqCSp6eVER268gphL7gtuBBCUWJtzV0iXPSl0CLtblFPig5WneR0KPONAGrPNrkdcqgYh0z+/
7B0bwOaPq+lWPa/5Xu113QspL2SuvYJVChh8z7ONN+ealzDPpr9+OBVsmFnQA9pO6jbKXrUty8j+
mo4qajQPwFjaCQqYD+IdIMcEgrkGy2MHHf4YhjJhyf9quDS4p3V2lCgF2yV6HZlCm+PyvICmdk7v
1HNDOsspNQcqbyzJqa90Vmc7CjfCLQEanlWDs3gXC3Z5Ni7Xdl2PXRzBmA0ptImyjBrPfNF0JVsO
0VhCyyR+CLCczVXW0kuGjX2LzlYX5CBEoFqbcay4al15q9pCW28a6lnsHh71PjU1z+ird0hgIBKA
4PruNjcGVX5InGfPIELWOTSbkHRMGrZeWSkUsxct2s7SK5HX0EiXzqaBbjILvLrUMS9z8fs+N9RC
3w47SsvcntpX4BSV/+0qKnoQzDbU37zgCFctenv2k8KmH/Ykp1Ej2hRx6CjOB9aYx7tnJvWwlCjr
T0Mpy5Cmsx5O8qHnRlIS2xfMclgmkfcgHQ1B7VrzCIx97GdVqv4wztRxtIuvI9yyRCO+5A19Jvg2
JnPbhzezg4A4xi3pj//Hf7kxVK/DoWgOyQWTvQdQ5dVeNh36VDhR6fOcO9iUJwfVmNkQcHfqh/kH
fW1rhDdELJYnl0l6rCh7hiq0MRKHJkV3wvJ1YhFayL+70F7GeofvKN1nAlQczM5IkeXFuYhfzj/3
i8Iyoh7Nz6gYPjfWBc1mC++shM6JWrqrim450vFRC5wUk54N07YEtEGQSl1tGuMw6EE0HqA1IDFq
dx29c9bw2uAChXkrScJU/0IPV7zV3pQ91NPGknN7nvXKOeRfxfXpBdN0YCILGh65G02PV0B3HsXP
/SV4+J5fdPnm2pXIp8u+5D/awxn4QUpOvbhvGd+KLHWYyTmXipEGuKZH7afmw0pZd6EUg8yTLU1r
nF0rOMUasKV47aheORylVNR75Z/iF/It5jhTC6xMeeIM6FRJSBS4aZVuWHAJ6fErJkNHL66WNokw
11HA8WHBiMsAF2Tnx6pG25rkbC97G7+Z+OztAZs6/1JS0VULSxXgScH5FQaB5eh2F0mEcyigZcX+
VpfbO7V4Vc/k62blOZaj6YyDeCeXA3TcK5bUfo/qKx5otuzrIuCVBoWFGDIHWTp/6AfkslfLYene
THrvdSqvghNLQDzApkitwJ+pehZzxbWdKLE34gRGpS/UE4Ovj0RanAjcg7558b2HQYDfvqM9MQUM
ODu2W3gGJdwLtZSii/Qjgbsslx3O6LSR4ccnIgu5odMP98an/f7sgTKR4Wcsk9UAKNP3jrfQphMJ
VDAKhFcyo7ia+Ofx+PLBHAnwqCUT/r9Iz8zwubEP/Ig6hfcmSwzEJoV1NnWHJeS9NISN34TbFHMH
w8VwUorh0HSr8VSJLAD6aBBs06UPEFPLcXLpcOP0WXBRYYV8NxYRwP5sbVkPHHsefDeMGQuWLvl7
zRAUH0o+F5x9yr1b/wKplHUPWe58B/ICDQ86JCldwlQi58BdpLiTfLYhkMm6x4uje1IQ2qOaFiNm
zxz22fxVanFFj/nx6GbzBQXVZv6dX0mG932KB8qcE39qz3pw06cIsZK9ve390Nyh5rOfw3S7gvFG
P6gqd01P5BpAA4WmVGywrn1leLAdQBABKGdTLirhwMgLwqturA72O5TF3GKVS2LXETkDo1Lg2vdm
ocm4r/RgWPDEToY7Nii30tkp7ckLgM4GWvneZFpvcfmJt71MXHPfSy3KhH91hC0VbWw9Mo6klYs9
XEiNp8eXI1bHfrCwce9eppKUs1piCr73QSy8xdZ41f0n/03GVhvQ1v3Wag55HAaegNYQjnpzg1XQ
gBNsqn/Q+zD0gxH5FZW7guVr3AUkCs8HWW+5FaYkuwUqZXKyeLRw4C7npCjdmdq4p3kVSmGeAV0L
A1d3jLoDQUUViBn/ZTqPDIhCx78YpUuPVckiw0MmkD5h+M6kBDhTJ2gtp0V8bXSvs0VT1ydrlFfH
OzOboYOME/Ex3hVyK624o7lmPLik32LfdgzNBP1koW3tzXfZOCconK9V3Zvv/BuUltShShfMht8d
hhTLyGNAcTiyyY4eQmy3Uzov4ObJbMytqjZ9S+RmN8RGdrjKO6mYrPHoPsEPLW0m2yZ4bkSBdhgW
MCM3sEj6u2hHR73MvtX74fQcz3Vcwt8B6PEbPzyNPcGVquUowr6AXpoQfAWBq9vVgqyJgQS4qczr
Ap/d/y0nYx62fkrYMWLc9JDh9ErSW402q0MHEUduLM/BlQV3wCzHxNDB07+W14QvTItjWkrJ/LZu
p9+edSDJPgIoMpEpLybJRMgPlIhAIS6akE8Vb5+iYIRG6E5ko/n9kTr2/L6Zml8z/uPMBINhb91B
hBxMDs4R9yeLj4TxufMpnR+brdsr7twhkSEhY735FIPVv6IAsCaK6RwfQ4CTOUEqCSvEvtnq30sk
ImgLIofcOqtD7B9e332K3Apk9o5b7feZYMpOQ8tQ17tIxhgqMJfcyywrV8gWVyc4EmCH/pxS0fXK
dtpy6zrnoRrpfsjGn6jccqqMBm3ixuevSqAbssVxFQ4A11LkmJknHkZsASGJdR3Xr8qEnrmuSSm/
RAluj95gdcuywv16Loc+2vn6ATAtIB5/CR04lN1pZjPlobLygqK76usUwtxaKLqJtqI6Yq74ZYCz
3ZceN2hcVMLtP1lDDRVvSuW8RNvPMITYmTKhmc6c/uCtD2vXAXUDPh+ALdiylxVrjPBI2P6gzazr
e0ckME9XMZu++87PqjwniMeTSqfihwltb+xxNPH1Om+DgncFSPRK7TR5de8qKsD1lbanqOtdeyFN
ATqeUIrLVWLx0dyNpVSWb4WmpoIBk58R+r7pp7pRZdLL0lzfoAggWb3PCOhyujwiBZ4iXIQpIFiO
Lq80vlXxqWmWWjNHk7UY1SWuEIiNnhA+DPL4wwPOFI5E4/TP3AOevRaDIF0cr7VUxomAl3R4CK0G
fQ3hMAEznkFbmDLvirAdHTomLeaSPKI1GsOvZH6qcfttD/U4F8SnTcML03wFPVtsfg7zOjt6WzdV
54EW2sUxiiE8yiqwafz7uK7h7bH6uQ4WBBPVOrHrCXY3DQBPt7m9MBd4vQDr8fYyphVB02+gK8x3
vWHoDC0tSFkl1zFCT/If3SK3CAWnQYIf3aGPe6oH7Ar8wmYB4OSLgz7UQpe8KNn0wvHug7HsxZ4W
QAYUOQS6K1Bdcb2u/e91j3N5rkVQtIx2thA2ULNaJr8V4v7wbHP2w7T3mU5ZahLcBmHk85ioYpTN
fDiyAuXD5znFQ9C4Zyo2oQ0Kqh2jf6HlCzrHOtZsksrnoqp467ZVEIkj99QEJ5+edZlVfhX0fEjs
Ykqmlii53uQPUPBspqwL4jqg5MoqS4LUk8q2sxZl7IoAHPNBiv4oq/+Uo921adU8MeAIn30v34Ku
H8+nxzmFfYtNK9AAm4RKrBu97tLAKf3S/xz+KQMM8sts+KVW8CtS6WrfIp/Cqm7FxklYe1mgpIEf
R61S13EoXHQL1yRG9fZtgBIXl9j+I9zRZm2GTcDyligZnZLW9Ju2Ji4/iQjtziz1XVPDPIQ5ScOk
sUheQopeaIxkJv8raCgGAQSoL9E5E8YMJZQTtOuCR3g7uht1tVn6k3CuAITC98BOiZFJhWkOGUvX
HD+6R9w/6lxSH1wCRKvMEm5gvFLZzb+yGNqO5yPU4AJsPZMmnb+sEbgfLL88XpxmAlyq5YzYeVW4
j3IEt9NFzAEmDz4AVWN5jUwwL3BOrLQDRm1AeQZU5K9Onkxj4Ofk7aPbJRd/NfV8MT17xGo7Q+Ix
7I52sS+ZkAokZ8x/emWI8Ls2lA1A3LqFC0EAXx5H86dpS+HjUMkn7WYxtPt/esKsKLm4bVbmb1kO
Rovd5AmngrMTt8tbt+U0I7JvCCX5c19ge0NB9r6hxWoVdS/jh1tqIUIlrBAkSfpkEsmzbZFANyly
aXdfj5LSYO+9ie50G6QbsDS4EYSh8pXj38oEv0upDinU2oMxG9ZdNCl5nTzILFLnYsa/XhqoZPah
K0OrLtS/WclSWOl5tmxXAJEh4bgUFc1B0SV+XDQ2uagp45dyaTIAiMavgphjNj2vQAG1Xe/9zQg8
slT2SELrC1jqsmddb0UgyqfmBXX8DFhP9DMAF5RM0YiTHuoivJFwUPf0SHiFjqseKzGWz1qwc5rB
I/95x5UTI6OQeu+A5IKPdiZL4gbrF8IqjSw/ffQJOYqgWVdm5WKgMelbKmCGRXGoN8QZ4Xt6GuU0
ad0XY+ZI7jNlc9tcOEtrkvALK1nm4K/PTbBg9X9cY9uwnMpiFMaM3f2M+JOCSFQPLHIwESB+LVdP
JTIxRCuKyUtRa9yf6ER9Qzvyey1JHTEXfyP/CgS14CFZMH8d+gGp5qGfd3oMVYQzYevXUyRk0ZFL
oS6dIJ7c+Nc7dubsZNMmBcD9vE08IDrW6Y7qDdPde3IaC9t9FplnhoBf0aXtj2lCHq0fzAqsQjHt
17Wa64oatG5yYKw70vHGdycNcH1Uj6r6GsSrPnd53ZVKdDHCogbIfzYc1Rd+o13/cknuL7F6cK1f
EisD9z5A+luJlxAYT/vyoQx4DSMuNqS00r6bXJypwSyj7VVDQW5X8pxbSmdAlDbgKCntqXgQVuef
cAT6cU0XYAk8p6gTYb37W7JKQNVUTFmEhcEZ+XIoi5w3/FOhqM8aM3Q9SvDrBPorbMjGeqc27uBY
8P4f/6qdGDn7fCSGWhDEYeREJ1MKHy+Ksp8OLndeSGdR2MSZDBST8iD9ohMqPShzMEdpiac/K7Bt
KApoJ4wmyGDebXILoU9yCf/KabE0j61hbhOOISvjhPOqVkzr9xJBInlsjVMJyOJIC01/T0z7qZ5g
XptNetKs3LQsAytYBSD0Y1lMuIbFYOc/V5qgoo2tcL775hm+Yj81euZcxTUVEv/hDoRr723EV2ha
S3EZY4Z182pcZGsuVKG5AN+DNYahZ4NKF9kJbF3TLCBl3zhah+iMaMVS1PqLtO2RxNNJ3RmTjU5a
mMBx3908a+/CEQ4qEnCiiu1sVGXozS0idZ5WDeBPXKBDz0wM0b3y0R91XE6qh7E5iZKIKXls9bwZ
B3vYYXea9wnPFL11maxpXiqe3ZxF9+10NykVDXQLssMHPKwK3JchMp3DYipEXBVb3a9x4CY9beDH
e4awy+rNqxajvs8WhJXpr/jCVs9DCndgN0lztw/6z/DKs20IjgH9cYKFm3dWjQndSUs8GLtDiJ5K
0FfftW08EyV54QqJCqCnBfY5QT8H+9CntWxRqr8s5fzv3j0viDPj3oBG2R6PlSU6E0NrjK5SO1WA
ZMkf/D1HqHp6sD15YURwH/d7Ji+hmf+KsQZpdZiu+iogeFXKX9Qj54kYYfoFmAGoc7xa5BQTODpn
to22vrsOfPxMReOnkIgiYwL0vxm1eyw9Ey+lajCVT6etfwzAgujpBwdSzzbpegMjRhUyPgcI42rj
lpQLpKPMw+BClyQEzmTpoiawv+qwTF+z5QVliADMNNFEDjaVX0gy1uPekKy9dmkGvf6hZHOn6ISC
ogzkFRF52zjAUzyL0RzlTiDH6d57/ELSW0nV04G2hG68lrzA2dOSqNnno8m/uW7legVWClfRAqat
hOv9+5C1qHN6xbxwoQmyfTQlQ195xrT8GNKecmLL1zBIu6q514k68inHpBPlbAw7aQfStcNprnn3
du2JqX3g/9K6UebagG+avBRzGO1eOpwCsNxWv1RzpF8M2F6z13Oe1zqoO52my9MikHS7fR6E52rl
tou8xEKtfJhMoPSoOKhb9APejp4L4MxMYIkrJflGKExHErsDmiqInxPvRrDYYUwyGOOuYbrvbCTo
HgRHiogC/KWZcdcnEs6NsuyLpF2u+W39ISlkwVnkrVIlgLfcK+CADYrgbuHyDbvOgTOg1DoAMWpv
Mci+690HjJGnD5ln1o9Hc9D1TTNuDNewMtNubdFkG/N5DVKZx0O/T3yaDfZbVfPOOGuVQBNBFLjO
Q2gEfyFxNLgzw6cDTzHb+LA1N/6QzcvSIiah9QaZ4541RwwPybyDj+HdVUw78/cp1rPAI6w/JoDa
7eYj9apHSjRk2mgL1FkEz8nkVDnIqCkUkDFIk0IpuLFtRencMzGny4Sc5qpSRc7tAiXtrFWY6BJo
h2qKJALvOkhzOZ6Uj5wJe3vj6tuvP/OLWOxRZAPSX80KK7W0koh6YPDLRnvvWid6N+mKlgqxHbE8
JIXjj5c37RU2c6LXx0lEckyJTtLM5xaDgUy/6PfKMcYk7p/K6D5eybffiSzNTJ9Oi1cyamOYy0Em
343qvoPxO3gl0MEc/AJ1JW1V1xnI7fEBp2baq2ZFuFRwe5pRs8J1aHCFIXKr60VC+28nqch8uJLi
UsXLtaXOO6Lh72Lu0CKI7CNoc4s+ux9NEcSERwkFhD0wc7B7UpyK/VwdJ3UbPgMQTivuOE1j3a6U
sboIHRAVfv7LwJWkuJtK4ZKuW2wir/AGVg/RjAKkpzlZFSrZQ8DXAWBxkypfckU1gYzzIleNvDuX
eAYtDlM=
`protect end_protected
