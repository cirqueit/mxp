XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������l�+��X�����@����6Z~����&L�t���/s�.�C�..�6�k�qi���R�e4�M�����@��;Y�U���2n֌��̯�I�q Ƴu�1}���{���ؐ��ۉ�*�n\�zWNw���4����ߞ������h�*�������<4���N"ƈ�)��c�	��[;��^��
-���aV[\˟�����bN�̾��|Z ��@E�z�W6F�pL����H�PPU��Q���Z�F�ѺTf�m"4��b�?����o�Ya3�[�ȸ�-7�����x�&4Q�L��I<Ӏ�҈J�H�ur*��a&�o7؞�3�u1�Z�FE�C_�3y�iմ��)���J�r�"�b����Է4p��a��~�.;;����)~6����1�h���\z$���1��ePtџ����W�2�Z㥸Zf�2���A�S݅�ȋjM�Vٔx�>#�	*��+1����+�P	+\� [���i��	�'b�_z����)�>�΢x�3ԲPY�������OO##� �	P����	#׭T/(�3kӗ|�A�dL��=�
����"��rk���ŧ�{��`F��,�5�Uv��YJ���<��bZ�,0rXBf�q劜�r@.3��
zM���x���1�K�#J�f6��_`����Q%����@�%GI#����6�|L�ށ�5c~�w)�V;=�q*؍��+�|���$�JK��ȅ��4܇O|R����ee�(�P���#8� XlxVHYEB     400     190OEm"3נ'��DN����Q�y��[���A�У�>�	1!��f0�XX����м�X��f�m�
r���|���������S}3� �����a��6�3-�T�����l��~��mm��J������ɍ��8���Ϛ9��h�6�>��2�!o����5ong�����6��9_�8��E�r�h��Zބ%��U���L��Y���;6�ae��`Y,Q�=����K�EQ�$��6���?�»�̆�P�*5�:5�pjiHIt���d��	�D��8���K��qE�Ғ�=�*p�B�w&�G�CW�>��%����s+s�PuNJ<e̋��HtY��2�S�Μ���* �07���2٤$�:�J���0�<2�Oj�N�ˢP�Ƨ$B��R�㤲Ml�FXlxVHYEB     400     170�ptؠ��eZ]���+;,���c��o��}���jU�����rK/����͵c_��1!(H\�Q�c��tS�g��i�I$�v�,b������C
s�5ɘm ��M�1C�B��p��;��݋�
wr
@�v�n�,\A����/�$�N<��F?؊�29�t�Tz�^&�L��^�3��Ȫ�+.�p��55���z!�8���p
xXS�Ml�Wq�[�C��v�ߓ��L޸��z���{-p��F������%��n�ǜ��*�u�/���ϛ�+_�ڂD�%9>1�>����a\��0F)4}�EI�U9T�5�k��U�.2J`���l�, �9�5��+��hXlxVHYEB     400     180�a�'��uJ���⪱��#f��iv�)��>����Hq`I�9uw=H���Ɠ�W%E�D��F8m�e��2��
[ۈ��y!��j
 ��� 9�Z���su1�S���A=(b aȵCU�����g�I߾�V�b�X�,�T���ŋ[�E3W�c���˔#�*~�,M�2��;�ҁ���^�'�'�L�K K� lw0���ܸ4t�����-(����9�AҼ/�����#.�}���=S���|�
�/0��w�[2�oygSCQ��a|��J���.�u�G�tͫ�`��	���;4�j�u?���rD�G�I~NUO�=��F�Z<�	�3���΅�#I�Y������@��!��k�N�����6�K���}�gXlxVHYEB     400     150�	ůw�M�i��w]9Q�&c]�Č9�2�<�R�2�o�IPq���wQ\Չ��:m��S�\Y�^��vI���ւ����g��2~���nq��U� ���G�z���|�<���E���Sh�R@�;9��p�nU ��?f���{�|��FT$_���I���u2��䱍�
��ύ)m��%{��~�e(��L�Q	�\2@��(�ٺ⦵eiߪJ�ޚ�b�+2���� ��eھ��e$��2�/���O�?�Dǎ+}DԒ�w~��lvn�SC��s�aH��s-m�i'4�>���&�@�������7����bpXlxVHYEB     400     170ͬ�o^V3���["%�bmA-��ck�d��|�f1�t{���G8�lh)������5(h�pYYL��bP�fCh|gދ��D%���	��/���&rR������Hx�D��6�[�>$r���~�8[6���W��]�������j���,��W�N�[g;�\PQXG|"�%P׸Z2Ƽ[~�OvF���za����u�h�.i˃������$�4���4�̼p�G�l�@
��bL��r��`�[�@:�xH[���l(����EH��#'�}�О{0<���ֆR_iХ��ө�ݖ��Ѐ�����M��y5���Fem(������a�>D�di aถd�ޤ�>G�m}n�<ؔXlxVHYEB     400     1b0k�ҭ���[���):���o\��+H����(��������\F�qⳀw�bHR�h� ��c���d|�^��A�:�_9C�����D�T�u��
;W����u�[��E�*X-}?��2�&={����`B�D �٥�)� �Gb���إe�H M5N�8�����bRiWhuάGc���&�5��˖�ּ�-�2m���u�%3�觓�p�lt�~�L�~������V���<�/3ө���P1�E��;�"�5~�ח�P���Ξe�V�K	��u�$�ɹ�O�H8�N�X�!��|�DY�U�� 豳�@Iv\����ޝJ�(ξW�����)L�ҿICR�*�����#� �n�|E\9�]���# ���EV�o��"S�`���B�*���?)y�J�̆����@Q�i�XlxVHYEB      e0      a0��+������P��A��\[�r#Slr���v�]�	B�Ȋ���օ́9�̆_�z��v�DҾzj|3��A�}�ϭew��A�y9SA�
K��$�����Q�&N[]����N�w�k�Q��hT����%��\���K���;�	����