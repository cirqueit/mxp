��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���g�"u��L�k��	R�&N�Gc�݈�
f��U���i�<����Q�j�eb�ttt���y�lo�?V�-U�W��(h+����z���=h�*i�g�CS�bXpc�M�Y�x�Q-��{|�u�� &����5��wHmaU!�%SP>��YA��tZ�wQ���>-�Z^*?���*�;��^/ÅA�`��98��ܪ�Y�K#���/�y��y-o>��A�~��j�d��ΦT-�"(=�U�?{���)'���kP�5rI�6�,�y6�H���`�='ٜN�&j�B���a}jQ!K��|8>�Z�]���0p/�ąiB*���^5&RHG��mj\�o3|��k�'��,��4�[d�2z��+j�M���=-
�m���D�	���������J.��'P�i�-���=�z﷊�i��!4�A1��k�-�AU �I��`1�y}�+H`0.3 A!dH���b	R�����GI���?W$n�3ͥF���� ^��=^Y�_��m��a�ɤ�73h�[>8�������h/��wFJ#���W؅ݯ6rbRR	��CߐK*�-1=T#����v��3g�yC��������B��<G��9G&A��\;��mE�ʖ>~�y�PFZ�i�f�~
�iL�52���+�,>~�^iX�j���G�%s�b,�˟���Lk��=z�g�/�Tv�,z�l���ߎ������v�;,>?GtF�v� �9o�S�����d��n0nv�G;�{O~XH�6�&oh��1�i 0��|#f���#��	�E��_�l_�'4�]��a�C����E��T[�x\�h��f�֠Z:1�] e�8�.�zV�!�&3[�����H��i ������vp&�L�󷞫�Z��I{���1v�K�+�x���wTos�K�{��D������$p���[�O�������������ut�<Vs�N��9�6�D0�e n����*L�d;�����6��kBaT�o�3�L����Χ�Xx<>��{6`j�y9s=�`�v�|Ck�[���t�����O�|�4��:����O/]��I� 'ʁ��s�4���s�Ŕ�!!�9j=�ѥ0=�j+ ��P����:�OHb�}�l��ִ���4�A��l�	�+|�P��;5��6�.��P�K��V����CD��"DqW��rF��MN%Q��W�t�N��k�LC������f׎����5�{����^d��6��v`�"�wt��g�e�Ƹ<]}BCr����>��ɿo[�o��D�0q��/��7��b����Z����xm�ivmv"E��<V7�?��ۓ�D����'�>Q�`|˳9� � l�Cw��u� ��.	T���/T�,I��Q��(a�<ȩ�.�@P=p�Y���:(u�����BlA�T�_f#�^�0مRV�ԛ��6Kw9*VTle�c�7�*�h��7�����?���"�Ϩ�ˏJ�����P��a㈳���E���9��ά_r�`7�����o�cxHBqmr�����g��E���n8�!5�;�T��[WS���^c��m�3�>���Z ����oN��n���T];�����4s�(�BEQ!��aN0R	^c�Ŕ�d3e�d��yӔ�+8���ŒH�,9D�Į��?��E�}����|�B�.F͌zr����[��$������<���s����a���(��gg���_tW���v�8S8ޅh����D�o��	uJ���C����kf=_�������)WU;tp*J��t2�?�� �-�A�~ِ�R�q��ΖΉfq[�Es�z0Fu�F9�/a�h-�����Z��߳�h�?�`�i�l�������v6���"���Gw��D��Q��س��d�;%I#6B���E���2d�7��V�N�J�Z�	[4�B�m��L��-��a@mo�H������vn��2��#5lT��1��_g�?�'*��S<2xs�l�[󻒽���G:�B���7��g�Bx<���j��AܰMy��L,Г"�/�b6P��y����+�?����t�sZ��|��G<��\ֿ����g֣���E=zE-d�*�_�'�k-�ߐ,�EX���d*���B!��.������5����8��x=����i�o#�(ţ���Q>�ꊣ�R�Q;/�*�X�,����ς/�_����*�ts�0F9����a�a�� �K20�ɠ82�.����i��yw0a8�&��(�K��AC�P^RK@I�̔���V8N�}!J�	�	�YҢ�c�"�ĲQ/K�H�0]�i���|D���	�;o�'���@�i��û�`Mq��3
����"@���j��ZP�.���绮0@3?ؤ��)�P�vˎB�lL��l�<Z�� f�Pط�l�������ʏх�Cx[��2��£8�k��)��PDX�-�C�"�*G<,�9v���N��ߡNy��3bu�� ���cVd���y*��IFtϒx�}�:o���_�EH�OC��tl��uA�
A�L�D���6p3r�I�Y� �<�^�����a;yz�Rw	����A���1���(��+���n/!*����*�T+m,���)I��3�߈2��
xm^��rU�j�]#:��Gx4�"�O���ZEo�r�9�,��qI���t���x��||#ƃ� KF�+��J����p�0�Al���|°t $�:�0y#���xe�����*��5�>�+Ŕ`��z�R?ʋ0����o�=8�G�*S��zټ?�eh�H�c��"2:fU��sp��l�A�k�ݩ�5prEP�EVg�6���
���;'�7���qg��Z�.��P�EZ]��������qG���饳�#�fU���v��K�%���@$��ڬ2{-A��{1�A��X_�X1)��2vAl	�I�+�R['��{��9�_�W����쁘�v�1�,x=�o��`PxHI���_�ѱ�M��^����x\�&f;=�|<U��:b�b9���'�t�m��ظ�w�R��Tӏ#ĄN�RB���$�v1S��R���~z3��Q��wj��Lnj�����W�.c��*M����ca]sG"`����	��ea��U�Uf�	K�}I�g�����G��S=�z��ӓ(`��s#��lr�R����}#���Y���E��ѥ�>���+�;�r��U v�~�Mщ��@���	±��_�[����	�[5��� �L�˝/����)K�]�l)K �"�#��U�C7����:_�(dN̝���W|�EUD]���2v(!L�4n�G#�d�\3dj�xRq(}�x�� ��rz�������EX��J��3&��>��\5� �XQf}*���m4�w2ڧ�i���W�oڊ��VO��?��T�ë	<?��YZ{<9����		4��R�73ն{�R�$|�KC�An$&Q�Y0K+RzLz�ܠ�Ww����@S�D6��=���_3	��j��x4x�孢
�y��O�K;���j�D��"�����n�_nvRr N�R
ȇj'��1�pa�Їi8���ݑIvv��<�q�򵉸�� ��l��Db�a��)]�l�_䎽�M/����z�Y��k��.8��$��W�i��V\C	j5�(b���̝��ն �u�v̀��pG���1m78��!���ʵy�u�tB��7oK��2"?-?n+����`�T�r3=�OoB+��:l�MO�w�b?DSۿo�fc�p3�Qn9�-ڂNK�t�mO@M+ߦȒ���\�F�ű��4K8QC����^Z��8�Ul�*���gE��y͌���B�vAm[����2C̚���(ݛFZ�o=�GS�C.�M�і�����1��Be�����<���]$��~o�I��;x�6̑�z��Z�/����mKe�$x��-jn)��Q�J\$����rz\׹�hw;�yUG�)��Ƚp�:�m���j�w(Y����bi�J��r�z�ʈ�Z�j����	Ҝ���	;��y��+Ӡ���=T*M<���|64ړ����GW �2^ ~'/%
�w��P��������B��gWczu����Ԝ�n13ۮ��A#?��E�4���PV�<��c���(�6�zq�\�]�y�C[����K�ro�@��p�Yo�ϲN<���&���̈�>	Z��q]=OH�&��Tm_���P�'tW�?Z-K��>�{&��*�\��B.�.h�^8'�&%w�c�ǨrI	C<1�[^ oLDN	6�wl� ~�۳�j����*��<��hyY����C�/:	4E:�)a��(:[��:����Y�����jO��&�֨��2� �ږL�X�4k+)#v�B\䍊�A&k���7����A�Df.�Տ�� �Eo(8�=R��P&ڹ޿�"wi�k�"41�H�S�轱j���9�_%D����� �ʪ9{&X�����ĺ�*,:��FiU�-D�l2�c���q7��W�[�>���!�{��߲�4�F3��=dh.�v��� ��rL�k��o�I����i�[@����e���S�R�!+٦�
$O���u�ϑ�=T��~'����{S�jsFQ�3pvp�\��7���W��@�p�ɇ�E3�%�"�k��LFU�N����RR¾{Ȓ��|��:���-Ơ|���jT��hPJqh�Ȍ6��������?����v�r��
�j��%~h�����nɚQ7���#���V�A����rfL�����-�>��O"�ٗ��쁢�v/�sK��Y���٩�Q�> 3�w:"����8����J������T#3�-w8�Y<80�흺�pBA�K"g���t�k ٫�M!�B�Eg���uܱ��1�_M����9(�9بH����Ϧz�o�\�K t
yn�Y؈#��a����ɢ�*Maz�7�\�%K�u.Q�2 	ay�Ψq�`�U�	���[�L�,*� �t��O>��	�*�`��n��+�N�l���]���.\K����;��ľ��@��/��k�~`R��$C��f��V���6�0C�Yg�,
p��A���11���S{x��"��n]i���OCX+�d�����l���&����\���N���+G
ؽo�Ls�Ԇ���ʈ|��4r��1�ۇ�x�ԓg�٧{�����i��k��k�����b0��A4�b��N5��x�25 ��f���g&�%�|��O��f�+U��h�Y�*^��q�v-�.av�'g:{>x�[�^�����0
F��M7�tb��_��0B�ZH���qgCџ�\%`�_�;����{F>���I �	����J��
x�(��`M������я�ޞz��1�|Â?5��ߩ��>1u�Z�iq��zW[IH�w4Qq��/�~����Wr�i�1k�CT���O�ma�]I�M���~,�=��a���gO��Xq�r�r�S�6c6N�:�>�-�,=z�0i�)D�Xs�vʆR�kk"��E���ҁ�v�*o��"U�����վ�A��a��Z�P��5!�w�Z��Ej�M���ZEW_��H�e*�lKl*\�\$�ggeKJ��_��%�dl�'SP*��Y�|X9����w�J*�8�J湧��8zJ~;*�WZ^�YǱ�!B��?�PU��ӹI+�U��,5�0v�ӌ����b�0���\��ѻ���A�Wżf;!�2.:/|���z[�p��&b�?Բ`
� ]��P����~9�	��Ѯ-��ir|�rS��avcg0z�l#9���xx�zаA��J�1�_����enH�� �U\�a'�JkL鼷���+�nT�S[�R
�����t^,����?���^M��}+l�6r�M�8��.�Ӂ��$�#\���a���ɗRn�zM�v�������$�m�Ot����*/Ӂ�z�#�,@=˖O0[E�o�:k��ط�4���zZ�Y�>pZ!����0�
X�E��1�,^�<P�D�<(���r�vr/��G�pz�1*S���Z���[vR7���i�PmN+!��G2dcAk�Ӌy�TC�M����!8`�q'��אk���ȿa��z,!d��E�5U��/������k��H:e�Ґ��8����_�<��i<�oZ�o+�����[�8�'kx�o��>,N�UJr)��B����̐n�gg�������s�SG�@_�.@S�h�-���⹰f��x�bv�p���k4��n�IJ����/�,�i{淖���u�ѩk�b3�����<��$�,%s�ݙ�Ma�͉�8t!��\�'5	t�q�=Ś�	ΓFN�ܵ��M[K��""����:����ɗ��vI9�̛�+ٜ0@�KӪ�H�`�S=H�'J�"J�8�[�V�&9Uj�r�9XX!6{�Lc���҅^���<Z��'ݤ�����d���ƞ��nd���/���l�ӑ�u������	����\p�?�8�����%�V�F���v�-�v$ʻ�����@����I;4a�"�v�&��+b6�c��M�)���,��#�.��7c�/�D55������v�l���S_x���e�P��y�~19��_���%U�U�g;��$��=)�F��EDzɍ�����(��JwT���}ӑ)4��ə��z=�p�`fZ�h̿�j@{^ڄ�b�[(�mOU�=#0�`�1$'�>4h1yRK��9�� B�Cᢳ|��F�81��pL�rAhc�tN�'�qcGC�T���=�(���br�2��*~?/������CÔ
c��qd�pˌi�X��:��� {��7/�B�\�oEEe�J(��D��Q��S��	�%�W�4x��ι��9mRթ�&:�X]�OW�G!�{��'�G��6�߼�{n�%�G$�X.W���ߍ�_��_�8��X���!��e"��ђX�U�5��ṳ���v^j�$��ma.n![]�n�;���]y�s���X/貌��-Ɏ%�)����`s<�:�;D;��)ݎq��K&�p�D���P�i/�Dz�]�/��!~���{�=�/�3T��f�x1z���h9���Y��r>l�Gc?����=;h��V[��=��r�Y����Wh?/.�$�a`nP���_?:�(|dF��{'�q�ո!�2���;�*��TǑǩ9�W���F.�q����x�?%J@�/m��xT8�q�ϣ�3�r�m��82v1E�h!��G�s轫�L=�^E�e��{����2�J@�����ذб|����@�,0Z���^� ؼ��<�Rz�rԋ�]Ȓ(�6Ԁ[\>Y�I�aoX7�	��]x���1԰����l���"��H�r�cz%#�s"���]rv:K�?F;><Y��.���D(_���}9�c79��`�!���,��}Rn`��·l��]�B�ʬlױ�Jq{�$e*��5�r�Ck���`K�9۩�!���5��'�ԧ �l]�j��a)�i��	�Y������`��)4���x�������U9�nf�� n��icjMX�f\�����#�,t����Z��[.'��o:5G�Cm���պk\!p��^g�%�o�܆|����qP��v��׋o�ı�2_�\d4�cI
 cw�`'C�p�C��]�>s=I���������Y3���a����� �~�����Zt+�r2��u,÷A�Z䱘v�A��p���H}�[��4o����M�?q��گ�]YF/����إ��\Y�L�D����;�_�1А��YqPs������6A�᛺�̉S�T͹Sm@�<�e����+R�\(����G�f�rB���m����m$�Wk~�B,��	o�.�`�d����F��2"J����Oha����N�#��y�ֳ��/����U�}�9��D����#��g�D�|E��O��}j�����0��$��\\�m����	WY<�1�s��x��y��*�r���ϭ�oK+��t�''��Ȏnl�b�0���%@XC�ɴ�)�4x�A��h"��?�3«a���c�T�i/U�$��T��o��Ai,�n��l��d�"W�?&~����)�`���&�*���c)�#�.��Fqh��9���D#�~����tʢ��KK�s���|��7	�F��sk��kc�7+��نT��i��Qg�;��7bS͏9�6��Ӛ�\�G��+T�i↜q<Xw�r��r�B��4q5��w=��ܻ7\?7�FD��Q����qS����G7wμ�btg˞Lo3��������kh2f�^�vuOФ����d�M��Y� �G�4ͥ�.a�O�}X�R�iB�C���:u���atá����r�?k3���a�6h^h��(k��M��s��mO���=��ƐK"o��#4ܶ��/���ȵd�.)-ŋ]�i�}e�5�Z����i/�l����o+����ݦ��s��PP��jsD����n8E��#bK,�m�]Q����=���Yr�諃�j�p�ȥF��NKkG�#���,oǃa6j�;�'��;۲���Q9��$ۥ�P[��D�S�{d�.�!�F�����vjS�fp�r>D�%LC#�I����`T�9:��^s��|����	��@,�#X<�s\�ӯI�1��P;���?�hW��X�e)׉����fO�Dy�
���v��8G;QXg?.xs�J$�rdY�
3`�'$˖gT&q`�9�7
�:4�ÓKnN)�o+���|� -N&�r�Mx�����>���6x5U�Tfັ�:	Z�Y��e�-�r����x�kY�S�����	�7.�E~�[_�1$D���/C�l2�˽ʃ��8���'j8W� ��@G��r�o���z;�\��PE~$��)�f��[X]���|�Z�+ ��J���Y�n��_2�T<�f?(�hF�O ^ >h��aҎ1'�*�������[o�u���I��4[��L M����቗�TL-8�+�w1�����M4B]�R�yI���W��i�y��%�� 9$��/�sMG��{4�o�x��s �v���r�ń��o������n��4/P��6v�*�r�Ӫ�u�4��1��\����i���ד�#���A�'��]?�Nl���5����=���9�բ�QZ����D^����p-������fgm*�c`�íV��]|�8�1�C����ң�"WH�,��i�B֗;�2�~�1�:���E8�fj�b�����*:�ޗ��T��|�� �o7�-� \��:w��J�^M�u��o��]��:��W,.ݎX'f3m��<.��Ch���$�)��a<�2����AW:\�L���c��/�[�O�XlGD�K,�/=��
�����$Nb�^�l�pM:�����V)0u��
 'rnq���yRUqj�M�~(olr��692�E��[Q M�#�V7�u�_����&M��Nז��yռlW���RZ^�4�����+F�]J�n��W�?o��������yK��M�)��s��lUM�=��*�0�k�.@h�H#�=��g���l��d��z\�g,ҳ  ��@�>�J�$i)U��_c�ހ"EH�|��e��t;r_֙��cV�˸�Nݺ�g/��]���ʉ=��˵�=/4��.�v[����s$�X�Դ��Ð+�mw�x?\n��+����;�"����w+���A��1-���;��g�X��Q��A�]�//ņ4��~6��:�"xZC�I=��	�e<��w G���9cY�\�z��+�k2�r�ڭi�ѳ�/V����ZݠϤ���J�h��?)��-�:�C0�ufOJ'�٤�1�+M�gw M8�"�h0�.I��_�@�Jl+\�쨠=`ْ���`U���C�.oΫ�������q>Q4eX�zJ���q�(�"��a-*����:�8Q�������A}�k�x���I�^daȯJtҳ���YjLL�=�;�P������Ӽ¥��3nKѶ"���?�`"���k��aE���%~�8�gS�ִ�v�ѠH�܌�@%�� 0��"s��,�_��U����-L�<빞��J6옩�e1��&�A���۫*��Y�wM���y���jXx�	y�,a����tra2�[|�׏�GT��w�61$
�Z_J�,�WO�7:��'�,��b0��`�^�}�J1j���'h9��s���lP�q���^�jS��K�@�]��?<��Y���?�y�o�����c0>z�r�!�ݷj��s���!� !Ռ���ρƫP�o�Q;��VmC��V0�f!4uq�no���p�#�㒻* v D�j�3�C��4L{�[�o�G��|��߸\*
�2k���K{�������N�Db�ח����h3�ű��b�@_0����C��>�P ���;��#�f��hk�@��s�lD�[Y]!u"����]c,�0��8/�jC��U�*R��H������~:����l�2��٦�'����0Vqx�b���D�۱���6�K]ă��b���3�Ov6�4��p-%{�%���kbZ�d Ǭ-Ѹt!�B�17'���6�M')��e�<F�E�9�4�f���n�Ɓ��ll�[:^�u_f�S���Q m8����	�3����u�5�sR�e��x��QR�:L�\>�s���v��2t�n�8^�R��]���z�UnW����%��8�_]�����F%���">�+�0�R�(�it<h��d�Gt��e�ZNT�� ����+��TQTX){ōk����~���):����e�M>h��\˲� |́@דk
j�a��G�@ٸQ�85�;�M���yYw=+��Ҩ�?2Q-&*�ĸS=.��E/^���,A��o0��Q��	��;_x�#�0�}�̊���i�f7|)�#<7��ȼ-iU������|����ȹn��-M���̹B�*���}tN:(�����䨓�?tS�2T˶edǅ����U��ﲏ��M]��#��%da��xb�Hh�me����\�6�?�iy��\�ԫEE �����4�̰o7�ڎˉ��f5���Ģ58n:nW��5�� KqA�n�kXG�k��� �X1M�1��,�����k�.��.^��'����O��tnmv&�Z�Gash����	j���괇�����k8u�����
K�u�7���Sbs��H0���0�M?<U �oed���f�rxr �m�<���q?q��p�cgH-��(5�'�J�D��j����&E��m��j�*4I
Ts[����H�C��,=����ݠ
�c���O*��CՉ&����8+H2��b%I�
N��O �~A1��x��!��έ�m��;�$����"��3�ӟ0R���\Pj6��0��f$AB[��*���;��㍜i�Wt��W���<!�f�:���M�.E�p�J��Sߛ]�G ����� ��r�o�ȡ�U,,f����*���s	pcK�-epfȾ��!"5�n|-y������5�i�k!ƥb�I�,�9��� <���aί��+���\�i%��Ξ*6�Ź4���0��'��Jy+��Tč����i�Ѥ^>ˏ���
Y�E���-��j���Q���s���` ���'�Hq'�F{t�^]-���c�I�Ȅ8�����ɯ��5ȀZ�K�Q��1�q���:����E�����ܐ9�{�c�F�F���C]���ˤ�:8�y6����X@C�_056�jE�/*�.�1���
�iv����,�kOY`ީ�ug�VM���"�)KZ� �ib:���|��ߓ�ڃ��=hV�[F��y���u|b(u���R�D�h���`ᗂh�G���>S	W��C)F���ˇ�H#D~
���#��� ���(�$3"��;03Hy�Tl&u�h��Ou�2���\���}O��y��Q��ZW��s�T�얫klh��Wk��UNe�'��*z�kR��H(�*�P0/�%��tJߥQk��,ѱ�)�w�.��w�d �D��Ub�е����`E_\%$!��~ހ�OZ&��q>���v�?i5����V;$zv�-�V
�u[ћ/���	O[�cw��R�ā�V�t3�<�ef2�x�\������!�V�;�[�����@J\�)+�D���G�̶\����Ok�`i�U5Vz>�W�t>��$,m(��*��2������J���X/�Ճ;��C�   �U$�n�ںS[\i��ڣ�!`As+W������qK3*�'��e�G����v����Y�����i�B ��PF<�ly���I	TG�G��k#�XS�c����p�jo�6�~�#�v�1n�;�paX����ʒ�UQ��>���pb/A���9���T�e#fO��&�(��è�@�aMF� �B���:����s��C�L7�"E�K�|w0~��~_+=OgQ��V�U����b�E1�m��s�&J�'�;$�W�������ƻC���v�}q+��.@#t�����T>�x/��S��ڗh�c^M����8I��Uuo- PP5���)��\�w��6�R��]ʳ�k����x���r�="�,��I1�@گtո9�����"&M[s�_�/�@�kT�'/�[�<1��އZ�/��Y:t��>�&F��tL ����E��W��{�j�<X�)C��wyH��l�2<�u��s�;;<���e1ga��O�%��n�c�=��i��:d�z�K:��!�u�����&u�j��4F/$���c����Kϓ�O��!y�mPڧ�$���6�Z3���:V�a��nʲq��-�BBΝk��bAt�C,�
Ν��i�{��,���1q�f�4,D�P�*�f��R�+���M�G�u�V\
�I:�5�qa{���3q�e8*��or��.A�F�4�4Ԝ�7��8 �����7Ҝer)��)�� MI�E���~)�;P9��p?��td�|��6�����D��G�n`�>O�]��Z����i����)cyB�d��{�ն� �}���v���Z�Й�R��Ohԡ�o̮y0v��1k���z	QqFA�d=�����wn��Xl���1��zїiP5�k��A)x���dOf��3�)i�p�09<���&��N���J����E�hdײ�t۞���E��q����`Rt]�W=�3���^i���i��Z<&*$�U��аA��}u�'�X|��W�Ԫ{�g��k5�8�]w���v���F�=�*����
*�կzqeit�"߽� t]����͖���ȳ�(��Zz�Zgڕ��(�B�����yS�ɲ��*O$P~��l�-����$�nھ^�0�љ�;gR���C`�(�d�C-6���&�j-�˧�t8�i�� �iv�픋`.K<b�y���|ξ�H��8-�.jIe���0ϐx��r�ox?�ꈛ�'gNaL�+�;�����.��r��~9����E�oۡ^��3hea�ߵ���mel��s�P4[��̂�5�����*��e�~"�֖-�Wﺺ|��<q/��3�,,/��S��[�t�lz����Z�ʾd�7 �y�B"=���L��H�'���	��_�����o%3��P�ďms.+�;�}Sv{^��R)f��Á�M����{������b{��ۅ���7���\��:ɝɑj�ց��<�;+&�ĳ^�̬y9,���t���E�F��A^	i���*K��u��F��'��L��++�z	�A�?��p~��M$�p,X&�r�ٟ��IL/-|Y�c���ZG����1L�P��ӼM۪�$�A*a���@t>� ��nd�� �cv 9~Z��G�^�����m�e�e$� �eZ���O)܋����H�����OW��u�sO���̸G�ێ@W|q1��՝�|(�2�i�C�=P��:�Їq�:8j���G�[���+�	7ı$���FM�P��Ҳ��"�	���,�:��]��N��2��h�)�O���=�L����x��M�up��i���2=��O�:�Ѵ���H��n�=�_̏6ĀT�.��������"�MIf�q�4����j�Tnp��>�T��Rsh��q�
p0%�D��	�Y,0D��\'������:D��B�7@3	����)՞�����=v�:���i܃�T�z�T��r1b�g*5��ŗ��رz�X�\��Z�<"�r����K��x�W�,$5�I����	8ǐYQ)����88�(�-ġ���w4�A�ͳg7���eiN��gN����:(r\#�B�g!L�k_=���`��W]/��^B�z���j=�JU� "@7��r���7c�*TR�l)�[
�|��.�t'����bd�d����I!�Rc{�L�Q���j��X���?&��,�ǋrT	� ,�
(��H��Z�n���2�"��]
򻟮u+�њl��(C<�����U+���X1�X}�~�� �����f������xO��C�rQ(H�{�4�ǎ�D�]��{��]���o��@���Y��z�e-�Q����F�3 �=��b%�O�$�e��ǵ�C~�a��h�tT�CO��ڷ�@�-(�jf5���R��q;�c�PM�ԅ���e���`�ï:�:�������ƌ'AΫֱ���귱��S\oW�l�`��֐d�h!��m�*��4i�ض�3W|�Q��Gf�s2|�>�)n0�T��c�k��M��6�@^V����a�2��4��M|Z
��E"x]�j�$�o�|M�Լ��2�KQ��"N�)��^u*�)��Ÿ�?m1�[K߆��1�&�	����Q������'XV��t���L���w+e��$g6���g�s��+�D��2�bV�;[֡��pq�4O�����0L���-3���U��1v�{��H��we�n��XԔFP([Mf%D���b�,��D���jz����XiuR��	X��Vi{�v����9M�(.��Ge����ٝ��lM��"�x�o��TW[A��zCT�g����B{�p����X��0��L���TH�n�Ņ�.�k����-+k#H�^B&V��h>�����Bu�/-lbF�}nS����rq���S�\6?I�!&Kk��Lzد�JQ����|oɗO�]SM���8�L�Н�Xˇ�\#�O�И���<@2�~S�㕀��Z�L��UQ@8�p��9�"����
HD�G�C�2GU�]͠�� 5�J}�{�Q1�^2k���ԈP�� �a6�#���|�΁����Vc(
,ŐD���P�ǜ=�,�L�&�u�	�Y'���|�-F��ɕ�QnEt05�z'�ed�޽���qq~�D�o����+("٠�p�`��|\<G�������g���yq� �p"h%�� ����G�ѸLH	[����z^ƀ���~I/��יP�8�H{v�Ι�^$���r'�U���\�� Ex��5)� /7�nj����l��:���׹�B5�#�qA���У��}簌#��X[R�����w���e8ͤ��Ҵ5��R{DB�A.�i�35Q������R�eߠBs�p�x�2!��3o�i@+�&�7���s9�Ҩ��P��ۏX1��V�Eg���lqR�M��
ȁ�`�72���C�{�\j�+���vf���m�r.�T��������Ĳ��}�<.���
L_{�-���|	�W�6�z1����w.���Dw�Ys^��+:޿ҹ}�؇�����ǣp������L �)c�e������ް��s���r�C�d��)���.I���3�GrBKJ|��"ԾYx��V~�P	f��N߇�1po%Ne�����H^"u����H� 2������U�ei~�7�x�ڍ�Sz,*u�5��.S7�G^������#P�Mw��0wwr�LЎ�RPf��LZ�����j�ۛ*�1�Nk8�fP�� 
$����~̤?�`t���"-Ϯ�4N����J�=�݀  �"Z�a���Y�T�mؙ/k+ �U~�������t�i�g���zz3�5���r�A�*�6��Oo�K��e�q��sQU��K���[\	.rT��x���=dփr�*o�s
��%*X�$&�m���!��h��2��+�3���!���:7����:�Tb���!4�͢CƠ��\q`�P��:fF����+_g��� i��a.�<�O� g@���!�60Kz ��px}D��@w����\�J�T����Z�t%C$��7�wߡ`��0��~�"e1憗��,@�M����cm;�[��f򿉧b=co�}�mDJ��(���I���>�$W�-MΒ��*潼?�#Գ2ה���I�D�T���9� h�u��`\tt�e�H���0�}	Y/��?�l�ƹI5�������,n=v�3Zw@�o�4�aLVڲ��'oNߠb��Z���Z[ffұ�X^=xi�cd� 3���	 �����Z��zr
�oh�.�H��!s15�5�Z��'(�V��A���H��ۏ���_`�?���iZ=|ïi.�� #3G(	/��!���ň�-�ڹW�'� ��J�*�0�>��G����F>�t܁�,)���tJ��$�B >����vfop[WE�
e�Ҡ�^����ž��`	�B��
��	+�r?�`��nbK@�z�c3u�_,��s�)ɷ�2�	]��]帖���Q�%�����C�w��x:�_�x��Eh�p�o���dO,�Ŵ�b��g�+�9j���ST6��{��vt
A���~!�c*�O]N�,�73M�BZ{��-�����2�`�։[:f�Gu����Vh�72X�z-A��C�{80[��D/dz���
�eY��6�o//�{��,ZÕ��H��|�u��iR�5�Q|�I���:I��d5q���zL,�h՛��\k�EP�s���;k��Z�1���[���`[]Ǿ����֘#XYp��D#q��6<,Z�Y-���iA��g�.)��i����SU�1R;���N�1٘�z~׆O7C���A� =GI��S)����qkF��N����$X�����+��5��(^��U���i���K�E���3��e���Žq@�mwf�_���)��m�2ǐf!���Z��"�M3b	��1�¶%�'����y�����+�� ��Jc��(:����X�yDѧ�x\A���ѹ�Yh:ۊ�>YL��5�Q�K���!U�&f���E}v�i���p_��D�!T(p�8��T��:�)�̩��|c{:Z��uw`e(�t-s��upe;����"�DV�ͪO48 �������%�|����7B��qpX|�A�i���'4�`RХ��k� c��n�m��\�L�Y��;�{P�bT��6P#��
�T~��Zx$�JI�øpL��`����O������2�t��[��v���̉�1w 	l��\�IJ�џu��[�"��x��U@��(Wk�j%�Z��̕O;�t�R��^8s��[�֏�1��*�)ʐ��۟<}A�>44�����+���=��q�)3�k)�JS%�Al�&��!��1�I�D��A�7vܞ_.j�'�{=bҲ]+T�Ա�X���i��}X�t�c�L��ɜ��Fj����2`T+�cRk���M)�U5FB5Ӫ�N�Z3��w��T��#�kdG���KBNP�A�?K�_������}�&sF.a�����Ir���O~��W�qS���x���o�^���3���V�j�$<�EQ�h�C��<��S�ZJt�ܪ���U�.��I�x�2s�娞F0%~p|N����]��%�d,��è��<ݼ]Ŧ���[>k�v��Rj�� *_��?H�T��S�<��mc"�>Pϻ.��S��^�W4X�(;� ��1���l o�b��.��͜B��=���3tV�?�*�����x]��~�ҕA�\��jX�q|�Hs��` ���}�~d�����	q��dQC�b����4 �7v�j���$�ZWc
=�W=����t���B�W�u�G�����A�qPa�����B{����0���/A�'u�	~�P
�ǆ�{�"��s0�E^�)����岞?M6j��4G���3�>���r�+�,�;�7s�pԃ��-h�Dk������XW�� R	��$ԱnŚZD��`0���Ɖ�"���jݸ��I�q6���l�f�n����b������5���e>v�3
]�
R]Ko�p�6UJò�N�^k�E7^�t^��B1�inn�[��?�����ZܵUY���w�n(�S[�{*)2Zv>����������o�:Ah5�I �.�r�^C"*9�`�����I�6p	Hx�81�4��,%���)��ϣ�
���k[�Nc����|��O8�~�̣�z�����O��7��_(���U�rxB��?����x�l;�>��Ksfߕ2z��'^r�t�"��S�dm���s?���lEN3�5�=vJ&� U`��9��r�Ч-�Z	SVe�%29��!����T�ȓ�3����QVw�e�u������O��C�t�4��k���ᄼF�f~�r�/'2����[j��eǧ��� �mr�8�2%���O�����A���k��TU��w(�s70o�0��b�n��#f��O�a��~q����q}g� D��sl"�����:$�K�_����7[�C��� �|�(�^1J���{ܥ���|Ȱ�l"48�M�7�)���:bp�
�oK.0��7���\2^>���T�T�w�^"�|�gդ˗�
�s�Y04$N��;A�>W�h9?��ٻ��y�g����2ۨ���G�L�����i�H��ݕb��n�W�"����7��K���ʀ�N�n�ZST��$��#T�J�o7�4D�?ӗCfW6�1��cK}?�J�i�xǥ���`�C��.@{ͨ�R���y �eQY8P��(�̡V��X� �ry���5�ЏKs��Y���"�oȦ�J7���y,D�c�hD�6I>b����@���z�|�c�L��t�b����x5�� �[�c���P�Ԓ�X���fq�L���������w�+;י�`� D�7w�O��y�5T,���c��7P�j�g�82f˺D,Sv�ƍb!�&wbXo�8��ٟ_I������X=��_>��/�E������'���<%	6GD���etz;�9��:��>�Ȭ
����u�G;٥�� )��=�����o%�
�e� d#�A���O�(��H^N�ڐ3*�s�	[�b�^�w�x�o4zK�c�k�#��!T�`,�9��C��X�u�vd^�,5�˧u�g����g�L?C�"����B%�FG�>JT��3���E|�WX���&<�a��~s0)�S�/� �^%�>K�O��<M�[7�L2m�v���%y�Ur��H�YG��^']H�sy���3�Y�koU��x�4wtn�~%�)��$�Y��m*<�1>Y��i�a����F�$.`e����0�"��������{�o}��o8�5b�*'%stb� "/�h͘+e�����]77�v�z"*A�Ȫ[��:��#}R� ]9i���mY%���_!n϶�_>�=�/~4�î51�%
8tR
ȌcYC�/D �Њ�?^���)'&����v��e�~�(G�7�m�I]��^�4re�?O˘)~�V^��o�Bh����AiQ��h���h?��h�[�X�hE�6BO�@��^�g����ǦezDulp_c����)�b��]�
'f�๧�x�l���6��Ho�C�l�c��3&NH��	T5Ye�U	����}��n(�� �����^1n��2��M�͚���^���' 7���bM��˃��W��X+�'<q�q��q��>�����{t��V/��*W3nz���o5�u�M����U�>�#?$��>��r*g�_r�y�������t�	�y4���Ro�vmi8�w�T�@��'�Tv'�o�3A��i:�Oh�\Xt��O9FJH.ƅ8ZZ�L7�{/��ù����bp^/�z�I��$���?�(� ���-ta�R�s�������aţ�����Q�|���?ы��tXj�[��"�d�5A��GQ�!9�O~�����Pc�����,13�6��9��ݤ��-���\�Q�m��Oo���J�*	˖IR���|�ƴ�2x<q�s��֍[jC_����F���?��������k2� �,��K�?mju��"�X\Ut�+���2�[�+Iz���dБ3��K��rj�8�r�Y	�?_Gp[���Ղ��N�G����yI&15n�V󯂍Rq��v�KV�D�PpB���f4��^��D@���m;ٗY�m�*uT���e@���xBi��{iT�.*5��{?�튦/����+��*�.:61!�HC�em.�\��k�S:��2�CruR���+b:U��j־���{����b|��������yf�O�	N���qLt����"�чl\�A�K��{�)~+8r=HUģ�
"vS�ϕ�"}u�m�`ӿ��T�GL<���meM���T��(ӭ]��X�>f����R���)��&�a)���}&|����\b÷�<$n"Ik<0鱰�Z��- 2�s���(׳8�>�c�?1wdT}�t�T8��E;<�a��E�ik=-�!r:�;��narb������n�!�3���`�M5�g9��N��O�9L���Q�sv�|�ІD.��2|��������WV�u���r큆�I�<w}�]�j%�[J��"Yb���N:�~�79��Y9��f�PEr�"��睌�SAb>b���B|�Rr%v��0�7S �dO�)a:���!1\�]x�m�b�7W�$���&����l�;|4[GM����D�i��oF�+�v���??�^�ګ�骉��y�!ޑ�@��f�*\�yFq�~!!Ɨ��^�������W�.YȎJ���y��t��`�*��-A�M6F$v�����_Z�1���å;nw���I�z�W�<���(����g��ev}�C�t:r�o���K��Q2������<Hdrkk,��!��q�+�Ɏ?�Ձf{��辠M�A,͝�� Kg�� ~�S+�v�µ� ���$���6B3d��������;�<9��T�����/4����!2�f.�?�6��?�HN/�WFv>T��_�iw��f=�Ӿ�9k ظ�օ[��+7x��xG����Xԣ->\��j���D��VX�I���dk��pz���Wϳ9#: I��I�@/�+<(���e;Kk�U�$�G�o�ܛ�������V��Uփ/�q��#��t@��ny�`���}
e�C��wH.��\B2�_�5�ڻ�>P]0����l��Q�����T"U�{o�����3+i�9C���dn����;�6c��)��#�S0������С��u1	��h��[�����@�<��@��,M��(��Ï0U+�Zu�u�x>ISI��H���t���n0�g1c��ϓ�mL�I��*LN�$�8ez�7��&tEs�zeh�l���PC�p�����J$���詟[ l�Z)��@��}�	6Mif[y=��m4i?���X�=to��
�٘�K�msz�o����Q�}�1�L��Lb��=ck�8�R+������/C.�K@ծ����]R�U ��+�m�T7�+ů�ͤ}����x2����b�q�Ѳ@��#�ϝ�9]�q"�A�YS���nݕ(�*;VF���0t�N�D�U�����o%Z��U�a����AkZF���n�p�ԉr5�yN-<�.�8�2��^�hlf<_��N�Ǡ7�?�����=G53��ȃ`�H���a!Q��NI�q4�v�	�yw"��"
���Z�%n��yob�=�w��հ��<z�wU�;�l�y�.@0vm�\���#�+������F����շ��-o�,�E&�@yKZ3�V�%0����/�(�rB���q6o�2^=nW�]O��&��"�0���	L*�s��Q.z�*�T?�r�e�f�믒�0�u8FaJZ'��$tkX�Փ��)z����e�)Z�@�J�-�� ��'���~���[��Tm�D�� � s��?�<��A#6a@�h��E6�L��w��X�h�A����OlcKv�n���PmO�vR����V���X;�kI]��o�P�������OK�m=��a����~JU��Ik�0����f�)\�om`�\r}OT$H
#WI�㉝�;)�,a�*�f$K9l4a��_����	M˼O��W�ݷ����<H�B��7�&]��~��冣K�_�߬z��#�Ch� x��a��*єYj���5d�����8O�%�ֳ�
�ں�h��#H}��� e1�����j 's�[��c���Mg�ۏL ��$jȕݙ��[<Ty*��lP�$���I���|
!7o{w���SL�#��}F��l�²�ųv����[0�nܪna ����k��9�=b�Ru�]T��E;m�NmA��5�r����w�����Q���/�����/;�:y� C�g��/N��Ѳ���[`~�^[B�!#�=<�T5���l,c��:�92 �*�E�|(-��eH��2HP[tC��KQ��Yn5yP�$'7�q���ا`�؛q�[�s�Q�S-����
~��R7�|�CI�6�P�8l���+ ݝ���B�h��o��2XY��qOS��.G�t]sW|�� 	���_YW-��m�9L���z�#��67�ەG���Y���-�U�����X5(�/kkd?[;=YF��¡#%�!�@ݱ̇�@�M:��#��i��Y�������`�}/@���Y����E@��K��`���)�r�{�&�t�����H#��z��5��8�cQ�l��;�����~B�b��y<7X��G���Glx�5�{Xy�i���??l(�IEJ�����kI�F�âFR�Xk=E�<����\�ނ`��eR�Γ��E�6o1�X(��~`,`s�Ɖġ�F�OS�Fb���.My�=ʿhk��#y��뽧a�#�!j�;):�����8����� �)xq渧r�u�Jo�<K�&�pU�o�ݗ[O�sG�3�1վw��!�Q�4� �G�3���%W��D��_��(�2��C� D��
�㈱Kc�_�TY�{�I
�W��ћ���Y$[nm;"l\i�uI �1gҙ���p���o�{R�y����}{���f�퀙)N�ңLؒ����шmz�Y�D�\����}��sL��,��CC��P)'-Lb��:m?���ɷ7E���?���`����R;\��x�;������k�G����4ϩ��q�HPt!� �I]�`{�)�3�X8���:�5����t8A`�|w�䁭��3��7xa�	�ev�d}Tu�ϣ$2c4Z�
�S	/d���d��o��lb�v�~T@ �����I���'@9�����k�n�f���HZ�G@fo���׫#�+�����>*Je�A��q��R#kN�� v�cW������([Ǩ�����L�Z!��X���5d��Rð��/0�7��W�F2A��J�,��X
F*C����\1��H ᆣ�ߝsf�
�=����u�o�m�:2�J�r��,%���& �2g�-��T��ZY��-�*���-t�M�LKgM��G$���ɹ�߁��ܨ[:�Пl��T�� 	�?OK�M���U�u����Ӳ6���0�H}^� ��R�+"~_S�~uB�w�)W�j�+t��e1y57Gp��&�F��\`����[KHPV�-��rq�^�����-,�"���yE��+�a7$�pv�q��!�FQ�2��.yk�VD�}#��t���"�Y�$�{��� ��Y�%�쓏�8�T�MU1),ÿ�xXǟ{�����
�1��kF� ����ݿ2�:8V
<�ƻZ�ϯW� ����l�t�X�uĲ#�����W�'j���������1C��E�����|��FT���G�Pҫ�n�25q�P1��b� #�չEJ��V��JN�ܛ�qD�c�Om�L'E�V��t�t�Q�h"�W���Nߣ�W�8��"`��.�ˀXe��r�_�(��Xjƕ�U\��j2�D���
z\:���Q�D̵2i���p��^�>��1�X��F/H)�ZP�ֳ���I -���hZ���,�y�ܖb���ځ���$c��ua$��������h�Ao61̣YG��H���79���$!�ͳ�猫�u����N����v�3�ID��L<�!i|P� <=���0�݅	r��R�g��+22����>X��[sk/���村diM�]�΢��'h��ҽ� �Ϻ8�m���:b�"{��<��<�gE%1� �#���Vm��¬�<ۃ�%cot�,&���- �_�a���U�D��s��ad,�߫�sjKN`SHI;�猢Xd~�Q�1�$ވ�\e����xߋ����PP>�%F�$ָ�C��T@�P7�qd����aJXU�<wY�ؠ�rUe�?.�����7��O#��ǛIp',OJ2�ݢpT2̒ ]� ��gw�ˤ��j���s��Ց�P��~�H9�C��^|�P��������-B���rL_E1����'A^#�T������!�2��lZ�6�m���H�i���q�@�������\�:�;|FwU'΃��,ىny1���7���~�$vj��,�����_ɷ�L��$��K�S�v���v�0k�o��ɮ����
��N�e���10�4��="(A�������w���݀a�� �L���;X:*���AS�h�)ny�����}Z���K�ۏ��3&v��#��XРQz�a -i�HmqfóT\�-��U9����eq�`�|����ws1 �������ﷆ,X�ݕR��GV��D9����k�<��zvzt��P�x�q�3�!�o���Ag!oA~���`�������+L�Aa3����=e1����Ik;�Q,3����)- Ǚ�MW��ԉ*涹k�o(VI���ks/,��M>%��x+oj��=8%f�opSB!T����[0��v���U��!pz'
k��L?���;?�+���ђGG��5Xx�'�˱�ԋ���H��m��\lۂ>+��� uM_���d�+�b��)�Ŋ��D4��8?ys�;�/�H����I��<|菈��X����W-#-3�h�9�"A#���%�L�N�K�cL\r]��F����O������L��o��8Ĝ}r��C�]q�?�8�����6r�uKZsx��zC�$ݖ�\ �����h��u �5D-/�Y���~˱w�p#ܳ4h�����h3��H�Ea#��T�YQX���!b��/�L���T��]A��a��]+��nG�t��W�S��"x,F#��K�ߡ�Gd"S��'�'���Q������h�q�T���@�yC~*�\B��<��q9.�'3:a�f�30�k�W�u>�o�z"���o4���/�Mz6��LB��}����w�8�0J=1�!��Jp�ƆLMȒ���0����)ʒ�����v�蔲� ��.լu%�Q��G.4��M]<z2����5�ۨA��+W"�O{I�������b�̝[>݌O���z0T��W`+�xf�`-x������3�]mTj3&��;a�D�G���E�tO��׾��Q��A��5���-��.	�/J\<.h�"N r�D`R����l3�W���9�Yʆ��}n�m9���OY�v6@�Cֽ�yHfݒ���u4z��)��<;�٣�7irl�d��T���`�Wɀ�J�:q�p������Aw��F���u��`�;�o�����X݋S�j�ì;YM�q+4^)�fK�?��Ddn�͝�i��>��ul`q}��=�7����[RH���*�V'$l^wʎ
���u�;��fν��oۡ��*� ��D���e�c�V>�+���n�z�]�2�0���K6�{�7�⌠���M������m :��t�x�t }cNE���=$�/tJ�q(���{3e5ʛ�S����X�.LH�lD�ݴ��?/��c�}�!���blE& oJpm�O�L�G��T��U�Y�gN�\�������B��p�R�S~�L�z����i��]^: ÷?�T��XF�h�:���h�qr�>Rur���\�9�VpLT�4�B4�,�_�JqX�;*.g���q_M�Sf#��8r��R)P4��F+��3ކސ�o9h��	��Y��T�����ݻ�x�A��#�0^P�������k���s��Y��?LThT`Z4�X��g��O�ܜ١h��V�a�⹀4�p��i���e����z�}ӽ׀s�X�Y�G�li��~�P9iF�g���*vF-�J�js0�;W�2[�E�5]���"�v4�v�<Pw�i��.ֽ~�ٌ2��z����J3#�1n����am:`*pn[أ�D�e�i���^+�6�������<�9�`�/;�X1��{:����=e;di�m�H�כ���S��M)A��-�����DKw�7ă�EZ��W�O'��)E4�'q���]�5�՜�*+����y\:��@N��i I�YW�J]D6G�#SmY��Y}�M��[a��=���L�;��7L��{�?\�F�N��,�Nï)�
�c�N���Mr
.�� 8s���el�X���_�4�URL���7~��Y;�j�����-�Nf���Ex��[nJ���2��U�Zq9=d��L�Iؼ�b�}o(��x�E�KC����~�� �ď�K�O�j,Ig��C���s:�h*��n�`��R&O?�ڈY���߄�ė�r�١���ֆ������rz�i7�
�p����*��`����f6Y�̃�~����B����PM���a��W׶')�K�t����Υu�iVY�2���'�C����u7�ûz�T�����0Li[LR�z-&mm�r���-p$�Bzee链 ʬ��N�ݰH[ci�N��)^�,3K�P��"����D�oU�Wί�a��\����N���:e)��e�Б��}ṵD��F�).����\��С>K��ǅ��H�3�P�&�頀�xד4�<�������l���bHc0G�=���nV15�mKX���^^���2�������ax�R����s�����������hda+�;� �6p7γk���|��0{})��V����ڶB��i�7��g�x��������/�H����^����x�_�Z��� ���h#j�ҽ�m ���0�>���%~�ZJ,��'�D�o���t����&������b����*o��6�]%�͸�T��,l 9����\,��?nƅ[hR��,�{上ah��T�$�)��m�7�C\4�j��n;Z�\��JW����!6�G��N ���ry��&�	N5A����}�����l��46�^r��P�=ǽdK���>��ǪC��3���>�i���J�p�3�&����Xg����ĺ�Z}�1��gI�DE����kzH���;�[�=��f�E�t�'e;]��4L����QUEu������{*���9�%���S�ePA�vQeOwP&�@H`�u�� �ϩy7,��-�ʚ��b.�I����i%pQ_����c{y��x�`8�Ӗ�\h��+����1�U��t��퐀O7��Q|kC����4⣽A�� i~5Q�V�!_�����?�D$�ij�m(0,`�U���!����q�K��ƞ#���yB�P���eO��K���B�56@��0�p0��B����ۨ�Z�O	#9
-skSJ4g&�A@%���=��ko[��h����:3v������f���$W� ރ���7nxLj��N��5��:�K��w�?�ْ��G+���:3���2**���]��ʎ�n� 8�����n ڄ�ze"��%��H 3Q�3��׼�TacY���<"H����k�Lr��J�3�FT���\�i@��$�	ӿZVx\��;IaF�(?Z\G���Nq�\2p�3����XS8��lȦ��x9?��7��$r�uUڨ�6�ܠ��$C������:g.�#�Y��p"$����t����ÑZc�dc��L��#^s��&���n�@�0�*�6��W�L:�]9���]=�S^���W���wtb���_�jg 8L���.��m�%)��X��C۷>w���cx���O��A��g%(��)[Nw�ߣ��Gb9����?^�:�dX������G2?��<D�@�uC�j�Y�J�LU�h>{�cV��U�GX�y��/䴳T(p7I�9}��4�V�7�QpO���τ����[��V^��ÿG<Ч��D�3_n7*�[1횒�:���>M�G=j^D�(����A���-��ς��[�r��\+���թ�@��+���`�y�����3��}��i�l#��-�9X�hFO�iF��'t��9��5nr��>��rXB2�
;�r=�1/P' �5æ��\��	p�þ�"���`������H��Ϧ(��YO�!�84�y��1t��<S8!�.|�46E�/G�KX��3�!���vBg�݆S��Sk�x�A2���O�!ɧ�]0�ը�@���bh����j8�� D�,�R�뭤��ԫ�e �
M����Ϊ�7���Q��꬜�2�v,X�E���mw,NR<�&��%�/��xrJm�9����r�q&z�pij��4�Z*�>�@�N��;rV���Î|,?�"m�dɎ6G��ő���j����o��.C����]�}Y�%ȍmQ�[b�"�Ǌ�(������j�-��>'�#|G�8�N�M\Y�2�Jͦ�*B���t��q��9)F�Q���TMp��L	�n��m��2xZ�r����Z��# 5Zw"S��)�q��+�؊=g�h�W��}Ub �'��~��za]���-桟�ӺD���l����!!he�O�6�u�C\��e�A�A9�{����E�W-2Q���������7T��Z�b��f�ت7u�c�Z>��qu~��3�a�(8�Ȁ�&��$}�u۲?��4�.h.�q�E�/�����m�5�A��A�4�0�=@DԩF(!�9���(Q��+�_�'o�1M.�Q��h�G�W&$�'�l�7�v�"$h!3��z�ڬO#�~�䁭u�4��y����X��\2��0kY��ւ�襧���4�%'�x�]R��z�`6C�;ϝZ�.{���y,Z
v���|H���MKTI�'��-��w�T;lZ��'����[�!��zv���&&��$و�+Άz�����F ��G{�n��lc��	駴��h3�Z�|�(Se�,��1� 7^f���u������ִ.�'l��`��|�C����=��1�V��]1�:�Pk�Љ��[dm��R"h?��/�EYϴ�A���.@�������C����m��;X-ܗ�)*r��濁3���8O�x��M����޶��:7���!%��tF7�xxc���tvV�q�ڀ�=J��)��d�r��X�sOϷ�)�p=̮��7u7K��ߟ��9)���YfG�y��E�]VY?q�y��:�����]¼�0���w���A��+u"�o��K��-��g�m�q��f��Xu�wXi����&�G	���u�_QI���+7~Fx��.|�va?DU�W������B�X�0Z�|�;5��,Ύ%�p�C�6����]U�Eҥ�����-"=�]6��J��kNC�?��A����H<%e���������͗a�����p`�po��9���:7|AK���};��-���Gyh�N�m��sI���)! ������/�PH�7��f̻�e�5bt#�18����a�-,����=���l���$2b���*��my+D-�lyf_�~ i�r9 �(���(��+���>��wjڈ����E�/�a�#Ԑ����(�N��?U�d^�7�A�;B�2��7]q�%0���h<S����`\߿��E�A{zTs~����k�ܰ��{�&!u&���mF�<��xAOa:�sB����;?�i���!9�%�H�2I��˓˓9~[���)���ϥ�&?����U�
�~]��Idq��k����� �� ����e�o��A�ᚎ��j/-Wk�3���͞k(���H+;����v��=љ�s�5C�AZ@�ą�������f��s�+ar[���0����E���(h��-)��;v5��	�}�Ŭ�D"eiqF���U=���)i�]�@Ί�H���;�r�2��wv��@��vw��x���\H���a�=���H2hג��eu2�Ge�-Q���+�%�y4{��W��s�IqB�q���7�q9���!H��d���?Ӓs�E�n�+�n�!q@�誖+��s�����ኼ�C�R�(���Z��BW��}�/PF2n�A!.�N��7���$'dQ���E�	�8�2LXn.N�/��m^�>��*�I�c�Q��Q^��bL��Yc.��Y
�/�k9CEi�'Z��s��	�%�|E���ZL9v�C��������>SG|��Тm`�)�l�巊+����ϺF3lw1�?3?��g�oDJ�]�	rH~� X*�ż�e��j��?�z�]����n�]8��[0:�@/ r�{���	2A��-�y.O����e��s�%��0�tģsG,d�|f�7u�KeF�e[Z���	P�VP�x2�!|f��k��H��zAMt���s���Z|������0;:�Ĕ��Z�"����P'���kI����ZJ:|9ihn�w��I{%�����߃�te[��񮨔������s1f`��cO�3^�iV�Ԥϓ�q2t�
�&��*��+�+���,~��f�L%�я��"Wc� >��b�0C�t|q�
�%A?��WG��^�R�ܷ�vh��=�h)a;i��bF��l$3ƹ~(�h��)�(?H�!n���;`�ċ�A�G8ܵZ0�k&/S.h�j�{\���iyS�֘K3�9F>��b���E�Y�Ɓѷ2��.��6��m�M�R��O[6�^ym�o'���V�4#��-.?\���@�W����i�n�S��,�)cQj�Xt�Z�_H'���\U	I�{j��r����<z�E��D�\�~o�:���!�8��Tqk�SY]��$ޛ�!,��`��FXSR��#a�� �]DL<g���K�x�U���\�3��G�ܣwԧ��d�Hř��	�$+�UEC��e�2�_��HY7B� �b_Cs1 ��p_��
��7O�v'+�U��dYs�^[�Gv<A�]�|�� �E�I�ވ���B96�;�g8�iq'�	$�? .�k,�u���Օ%h������n�����}'v�@�z\�<�f��%�x���3�3��f3�ƖCOgL��{�Ϯz�$S%��an��e��	�nԲAȑ�B�c�[ �"��u�\�����Fí� ;��o��+s�����?�<ѩQ�&ߑ/#�5y�:�(���~��:+�Ϸ^6S�u7�[�[���ݙ�5.���)w��侢N�ڹ/�C�|V��M!�PV�G�pM��${A�,`/�Ua�6��A��E�P�WGCiNF�J��C��I��f���gx�J��,�ZTC[='�<k:el�_�( ǵ@��N���׳$��)P��h�@�A��|���UGao�c@�l7J���c�6�Tۿ�����Ғ/Y�6���X���>'�( ������L�i�0j�������/����oQؗV�+�3)�sN׫p#����FPGy��5���K�觢7׼�0R�I"�w���f1nh5]2ܑ�L����&&Ȏ*����V@
��g"Ca��πӡ��LP���\�$˼`^#/�5���l�A��Rx��&��`��7��M�K�z��)Ke.���?�u��us�,�~�[d�Q�X�E�����nM�T>~���J�Ȩm�%V�'��Z	��Q>c�c ��N6�It}<�5t:������!�)�R�q̘�W[�@#�f��0�w����t��H�N�'ӎ?��B�.1�;�x�
��j/pl�5^���~�e�#�!M��4i$�0?NJ���塓Xq=��{�-���4����|�8^�	"n�Qڤ��i8[	���ɍ���L1��'|Ui�!�7!�3�yJ~����:��^8y�����-���a��G�0�������tY({�2��K�Zǲ�s<I1�"��A�{�>�a~9ᥭ���t-���Y��	X#�S��`���r O)�������@�0�.4��J�}Ld�r,��kT�?F��_C��2��|?u�s��Ţ|@<L���rÌ�Ⱥ?R�ζlh�tH�ĬPOUW��i����)f�	yW�^���o>]�0��_�wW�B~rÿW��xQK&�>0.�%""`�F�C�-4���x����h_���5�4��aq>�łc�G5�⌹%���-�9v ��pl�7�-5�����-#x	ao��^�tҥ����"6�`�� ��@e���{'���r2�&4/��|�w�:�	�}��b���Ӽ6Y�G}��n3�T�t�����V�~�i�T>����0�:��=� `��ha9�$��d����:IgΌ9��/��@>�p.3�xQ�8��<z��]��������ñ�u�}�>��+lڌsqY)VX�1�{&j��G�KX�]S�e>�����W$�IY 3�/�\~�'Xw�E�/��K�bv�V&y���r;�Fa�sp~C�:���P�2r�Ƙ��|�{O�
�R��x9�%����.������DF�����
,Unc�7��:Hdy�)Y������T	�e����8���?G�M .`�xg����a"˿J5�w jc�N �AXY�����~v�y�Ze�]�e�x0���\�(�!�/�2<�����f:�e����>�
����B���d�`gC�#��~,s�c�p%����^`Ș����a� ����Sc�qW3Ğ֐K�퉵�����+�O�4~��R0xw�(��N($l����7YrE�)D���Y�����![������ >i�ڼ3����}pm����;@0
��W�!�~ʭ��)kt�1��k��:����ʫtg+y��B� �lJ2-���0R��r{���<͐tu��Vg�(\-.Ja׵�a��$�}�XRuk��~��(|`�M{��',�]��Zi�xPg_��{EmmB�9I�H�\�튠~[�F��G��M|��9Jx�-�8i��nJ�s
��/�.Z(+��N��CU%�Qz��u��ғ�q���*�{��S��u��5�y+��B9��"����!�Ǘ�|k(�bm)�(�P�j��@=�(H�ޫ~��`7�gg���M@=A�ҧM�1	
0���'#bϦ�~h������	B�!�6�=��g�
޳%ҵj\��^���#26�އ���[��=�? ⬊N"W���4����V��4����_g��l��K�dE �
��Ѫ��5IO�ei���86=a�
���ba%(��e��.L��b��v�_�Ņ!hs�;�ؼ��ٖ�
m��6}`B�T��nZQ����+t
���%"|�?��
x���0�]dx���!�����݋h�G�m��Bar�R�s����o���zu������:�P���z�2��+8(��j#㝻AI\���ᭃ>$L���1�]�:�;�TW��^����=Dr|�O��WЀqUD���P��P雫�Vz�B!J�d���Hj����]^7�`�1_�z�Y����Wn���������$St1������S�D��,�0�ħ
xi��X,��]�m���}x%���|��&$�.�f�=塃��:1>L6�d��o����#�`�0�tT麖	����+� ?�������-X_��U:��҄6Gf/�
��V��:,�=A��g�A����{�ϦZ��)�u�	kj+����OV۩~�=�.�j�V�h�"�;�~\�[~�kvخ\���I����$T�׌����(�nM����N��j�k��y2r�}�T���=l���t=7c�Laq�ۑƚv��]���Up�C��M�l6m�����w3.��$ߞ��0gU]v��~}�U���� ��5�ݚ�̉W_U:E�c�} �Φp�"�*���G"��A.B$�Ǜ�]�\����>6�M�^r��e�ƽ����	��tX_-\�J�6�\����E]%���t��%������7D��<�y�(�g�=ak>=���B;U�;�yY���ॶ�(;2K���x�JUD-�4����CZr;�� /���r���{>�	���ôM_�\�T�Jv)%\�N����)���-����#�pO��ϩSUgV�vj��F^4���ϥG�S4�>��� A�7t@Ik�;u�s���n$�(�$v�4�X}�3~���m�U�Mfޝ3�"��ݒA��O:��?���W�B�K����r|F��Q�Za�j�(�	�o�2ei'�}-hx��~U���;�x�]�	�G�R+�@�z�Oh���[�>>�Bm��H�2�3���U�-��7��;DC�����N����7"����uO�ғ���pt��T�o�*@��N��!���t.�V[�sN�v> d�M�8�
?��P�\Ddve������p<V�N�G��-�|�d��±�k��2�ԧ�S��^����Z]s5,F����Y�_p�4���h��>�Xܥ'OZ��lV����V�V�mrv���[}�b�>��qX���4���BȣʥH�r!C�iKzO ����S�d�D<�O���������mS9P�\kQ��$�ɟ�i���	�(N�f9��ɵ�Y	{"�2hk��A��P����^�|�풃�S�K&���7��&��ƹ�wk�C;
��W�~��]��SZ�')�r��EY��7r�X��$x�T��qs�:�1&�ȳ�������������/ �BI	��%�P�L��|Y�����h��0���7��^F�>Z؋>�	^e��|�����B�r����/�F����R��+���wd��P��o9�8h���qj�ηmc��&2j/S0'���7�g���[J|Y�׏iw�a�'�A��+c�|:@ے���� ̳*ǻ<��\�D������:ȣ@^�b�S�[�5�[��#V+6x>�"�ǟ���;P����M�n]�"�煐]DS)��:;�����M/��ɐP5}a'^�����s3"�n�u�������p��5?|�e�i���-���q�	 >
7��
n�A�pb��^ϔ�j���@n�ʫv(r��e rP�,������s�>�X�����т�R���)����h<XYc���FS�����u�:U�Sr|z �����膸<�U�|�Śܯݧ�u�>l�OZx7��2���h8�K�L���Yx\M�
`�o�E�`\@��r��<3 `I3�X�BD6��Dzy��Ŕ������<��Q�f��u�b��~1�a�C>ꃱF��ꆹ����V��br1@��e���y]IF
��$�G:#���"n�ػf��_^ӎ��d&��tJ�#�׹~�F�6G����P
ri^�UΩrb�W������'<�V���
�*!l�^;�PO����+�[�E��{�tT��s8K*wꯍ��X�Pu��:@cX��Ug�;��ˠB���~�Z�O�J�8�%.�G�G��oFz�����I���g�50��}�Y�
 ��(��?����M��1�F3��á�_�8��B��n܍�ky����?�p5����*1כ�_"=L��^�������`_���\���b~�-���U��=��b��f����\��ڠ*�B/�����j�����J�0���j5������i����xB����:�${��0��V�/f;#v�-VBs�+SC��� ��X�b��#�X����!"��L��s�dd��9
�������7V5��ĤZt�7A4؝ �UwO@����ϕ!�߷$�l���i�:'&��k�I�K�/�*�$���SrO� @��{�[�2 GO�5�:L`ڿ�QNqN�������M�pZ��GU��{��vW�E/jw	��� R6�³X�h��D�H�&p�J5��MMCQ�Lż�pI%��->���{[ُz��mh#�g�ݶ���d��D��qWn�6���_"qK�4xk������B�mh`wF�N�P[��8��M�h��Fx�F��N�RnA�헁�v�)}8�ZiK���l	Q��-��ד�Ǜ���'�WP��An��h�G�ИQ�nv���<t��U��M՘tU��6���WکЦo�Ur�H�EqCy�����>�o+Q[���k�����x:V���'��t��	��u,��wO��i��z�-��/G�|%�ǘ�8�P>jnQ��^'�?��z7IE�
;2głж�Ћ3�(�?V��8-glh4f�&T	��9ql�,��y4�pqbA��&�ɝ�ø�E�z"�w���,��������v�c�3�`�aŇ��w�B�g�fi��2:k:~�1�6�w����*�5i���AUޝd�(���?�!Wd����˕3��#%��+7�WN��AK�>���gj�L͹I��ƦH��Cb�͆͆�V�K6B�+Kg��"ߊ�:���W��r��.'��F9D�i�ހS�bv]Q��!�]˫$�S�@Bs}�>�� T��Q�^qے�X�]��L0���>�v*��!]�`�s��ĮSMAv�� T��W��-\��F�"B���3x�?+�Q�6�\�+Ӻ�_Ym�Ƴ8��2�(Yў���++�w�R��(;�e�
����/�\n��w�࣓��}���vx�f��l���]���oO�'k41(TU��1���G�I��0��´XX�>W~��wz0C��g��H���PS_���w�i�(%�.���F�3�%|�Q�	(K�4bqx>���h��16��ʵX.�Wɲ�e�'�ի=��#moN"S���Nu�/Z}���?����^�H-���
f�lI�a���c�P�	v(�\M�-%E2�l���a*�b�3���	�|��?x��K��9��i��)F��B�P���Iv�ټ��ȷ�d:�٨#4F߁�q�A�t!g�O��Q.�bš�T(��Br�ڀ�{V���z�N!�w�����..Z�g�H�BCa;�V�? �4�Z~�'�6p0�"�V=-���ŝ!G><F�S��`�RG9�0jз1\��:�a����e�^���y���;ꖉ�t�v��@�OI����B����E��;�͏܈Ѭ˄6]�y砻kb�{�gx�l�����|h�I�!�R���.kn޼L���'Hϖ	/�sg8�A� �ZT/C�"�0�Cy�p��*|:���վ�p|�A���,�eT���@��DNh,J~�a��#�.2��O�;tH��rf4`��j��A�d��*�V=���|�.��A�( ��c�u=�z/H��d�R�������Y�?W��c�ȇ/f'�\!~f��rDO�/�������"����@�.�1��KD?�f��j��g��U�j1�G�1>2�'x�V�nf6�$9��,�HAlՃb��}�M�vdL��Rs�b�����ρ���8O
	6���"�x�Rh�N`V�:�>�$%�)"P&,��
�$�#�i���2yHi��Y0�8L@Cj�c��qC���\6���]X��KǤ?�����$x���AA�}�R%����)�6-�3Q��FE�>(�$ӟ�|�rfȆ�'�Xhd��Ճ{eW�K��.j~�%䲛ZX�ў��������k���A`��?�A|���ڴ��"���V��3�Ё�ܯ�6��ۅvr��W�����j�s��c��?5fv�t�5@��~�ph��f�@�]@���	�e!�Uj�*xF�&��;�ًK5���em��׬�Vq�1%��I��On/��,�I��?t,)_ڤڴ6±��� -lS3*��Ze�S�����ivGz0G:����$8�Dтq	�)IeP��8G���l�f�w&=�9n�n[�]F5>y�zKEN���>��C�8I�([{q�v��Ȓi�?:[Hy�)��Y\k�L���M���}aAB��X�%����}J}��P�.L����0��;ؖ�{L�^%�麎����86vY'æ���>�w���b����0u���)��N@�q{=:V�-�N�jIJ�����(�+�ǧf�a:����nV��3�xp7%��� �F�	K2�r�k7���E]nx�8���"�\8z��}��'��<W�� �km��80}�|�d��?�.Td�5(���J�v`���.;��߃2�k��[�O$\���l��n`��Wf;��� ���8Tє��xu��h�WR�RAa�Ȫ��d�]���k2�Ԁ�r���pOU�o����A���f�uvG�Wژ�,��t.� <�.��Cs�m8p�'��*��FAD�Jic-����}��`3I�꒲���zbL�f|��W�x9�d�J��mSuGݰ�rH�Wg�	=~�=�d6B�9k�M�-��}t���,-w��0
4.�V��:�;_ۛ��s+�lz(�=t�j1�hB��F��M{ʺ-[�1'��(����v�'����/��yu�윟8��?4�f���ۦP׿mN��+��|(HJMP��&��hsӾ��Ol���ほ`��C��q���.�sCa��%!}�� ���#tv�N���bB~�|����	�1�V�]�Qo(�"H��"祎To�K%��b 4�����U�ڃ�R��)�#�r�.O�^�M?��:�
�f-,O��*{�\6+��'�����g�EK��Ҋ������p��� iF�����Rms�AV<`���׫�F�*0��"�]{�93���C��m�Ge/�2���V^"� ����fέp���S�^��m3�B!Q0���ч�vR�BK�|�J�ӤNtM_�:�<�t٫�GR�ҭ���ϭ��g�A;`�2"ijmx���vi$!C$
�[ڧ�G5khO���0�J��#f0�����L�go���\�=5����:g�RF�~�NNs�~��G!�R��5D�7�E3#Lt~B�Prn�Df@��'��Mw���Ƽ.��x�8D�L��#��vݥ���av4ő
"%
-�Ǐ�KC�U�����h�R[~�7��Z��uu���?�ޙ{g�р��]��z+Ǘ�@�0fo�aStQx��㐁鉿*�}Ŷ��x?��z)����be^ۍ�d�ˋ[8:)'���)�� iߣ?�n���W���}��l�.&`%��[7��w8��OJw��֣sa�'����N������!^򿉶��_u�hK�9h]��+�w���9���Ý��?�>�����q�'IW��5#\�2v������ sdP���vF�Υ��pRU��I��Z�����~ݩ*�N�� �k���aP������YS�O���_6zd�g�û��HwH.�A��}N���N5���N6}���>a����]u�'h�r�ﻆ����V�$Y�s��"j�&_��=ec����_�<���'i�ҿ"�]Ь$��u�}9Vg	�y~�~U�a�ݔ�I�B�dlI�Lf��1D�գ��5@�6���vo)i���˛O<j��Y�<��o����֞wڣ^��߭�!R�-WT�x�ח?*������hj��sw�4d ��.R�^�v��	�����9G-���D��a���� ��/���{�KQ}��y�����(@j�����@H^%����������W�Gm
)+�,y�Rk%j�N��f�
~�x��O��N�W��%~`�-�gD����Y\��t?�a-j�d^؆��#`��WW�zͫT�B@>&rc�BXe�o� �TG����r�WD?�����_���	���y���&K�j1����ظ�Y�l��.����ұ�IFV펶9�,[dTUsQ���n�T9�xɐa�祽/���g�\�]��儹����C?�9���Z6=�XA|߫(Չ��(��8���v�+���?��C�����A��0!~��Ijl/e�=��D!�F2��+�S\5��ߒ�5�+L�(�y�@N��؃;�FoV�n���-*^�3qw0���a#���ŏ-�JH�GH٠�Ӻx��3���n6��\f�ɱ=K�����_�@�h#��)m������ت����������J��҅�ڹ�*��
�d^5��\K��x1�Α_��k2�`VN_v�x�o &%Kg�,����B����_��JJ�A�,n��mJc%s~l:�<��F����������C}d��O
�C㍵V��tB����,�-.q���}C�ƞ	�n��a^���<	`�3Ͽ+s�]5���&y4�0~��j��o�-��%Nz�:ɿU��M�d)~����ͮb�r#���hG��qU!4�L`��hZ�C��E@�������1!a����v�3\v0'�� 3&�@�LH�Hs^j]7���K'E�����&�Z��ql��
��n�H�YI���)k��WP�$�B8�_��Z��: R����BS�|�'G20D/-�Rϫ� �%�X��v�8m!�jāǋw�4<2Q���1�X�T�!�H��n2�dE�K��r�':@�����B��%�I6�����F�E�{�z����S��ˮ�C�ȒG_|�V�̪_��e��`������f����9r�Q��o��mo�Ytk��9����7$;��׻(�Jy&}��+H�n�d�NK��]O�p`���*�U�Y��^�?��a{A�M����p��,B���D�C�B�	v���t1���d �E��J�Z7@�7�0�`fҺV��a�T�kb	�<�\�t��������}��6cF���;A������/���+a?���@d�?��W5J7"�o�H���ᱺVb�E�ɴ�CZ�9`r]����Ȳ�u���6�HSk\զ���x���wX�ş��D�*G��gyc���x����uRH.�k�F	�Qō�0���k~ɹe2@���C}N��a	O#��Z:�f��`|q�9���ި
@��]�W�׊����S��ӽ{�_<AN�./&4��2���*:��&��Q�ŏhS�bW�b���%�ڈx�F�&�ӔV 9��*q�g���0��)<�� =aJ��ۺr�%�͢zR�f��Ɯe���m��y/����pr}�.?�f	��Ha�z�=�f.g��Թ�~�8?V��,]4}��P�Ջ�0R�@Jt�1���������i!�R5������T_R��:ٸ8�c�
�Ad�/���t\b�]P�!�Z��__�cj��ɰt�;�
&��5�g["�����CO�rtG��Q(��3<#F�cA�<��O��K��~�j�f��}��p�V���-�s<���jo�<�s�uj��zo�b�>�h�.&'�jv��k�������iD	G�7c�x-U�l6��Ȩ��CP
���c�RC�3��_�6��`��i��Q
��_��OL"r?❆|MT�Er����h��G9,�Q����CC[R�^xe�ͦ4�I��:�w�IĻOj޲m�!/_��P���q,���͕��~�I%Ƥ��Ǌy*1Cѐ�X���,�f���=�<|��_�.��,Kˇ��q�]�r��Č�U�6t��_p� S���BUYWJ��U�ƈQ�w�&��h�^*A��� A^|����O���E�w���7SQc�|Z�.��#�o@D��Iuh1�Gk���W���Yw%t�\,S1�����I�9-U�-�� �D�eܯ���4I8��q�&+�,ٚ��^ ��l�臰�9�'�^���>}!0+g[��}>u1��5���
1��A4�_���3u�oT��f���nTȍ�z]V���[�w�?�*��:��Ny%��Dd�N� �b�~�F����%�ϩ
�I�֍��P�K���/�o8������*����Nv'��6��_���j/0�[ >d����ua�ؐ���
5�/#H6�R��H)��v]{�O��]E˖v�̧l�SBt�?�0��sDK�Ez��*6�3�3#����찶KMxM`��=7eי�8����wqҟ{a�-�?;'Z�qI��"��g�M�3�ǉןL^���|��+���<M�2����Ŭ6�ˣfmi�+������Xm�B�*��=j7@�7W>��zl��ߒ��:y�����lN{�,������	hm��kA�.���{�N��$��%�hi�o���N�-V�Q��z��8`X�A�4Ra�Md�yz&����7P�Om���C�x5V�5A�ҥ��Jy��z#_4D�0�{~����e�+�5�|�T�֩�ߝ[���XOn�@o�!�1F_�9�%� 6B
tA�ws=�������=��������]�h�{�^(�ȩjN��4%��]��r�<`#^�@�^���̢�Q{����TH�:�\g���`j�
� �-5��a|,��<������* ��Zsƴ(���cz�Hۜ�x�Psk%MF���=Q?�צ��;x�(�D$#+��kA�$��.Q�����럣�"�^T�Oe��P�3�'4c�WM/A,.|��a���6k��q \ͣ|�Pn�!�!����X��մə���<U�D�1^=��:$9j}	�g1>jH�x{�Ӿ>аV��E�EN�A)�]@k�qA�*,�H�>gh�;���u@��3#6sy���N�tԿ��
UF���b�DW=xQ��e��;��Lؙ���)�(,��w��Ab���0���
Q��WN�SgRG�tT��\z���:aJ� ����Ks$�8p%�9��V	���%�8���d1�:Ԍ���ʚ�o�tn���vm8/V�Ș&�ih�Yl��	�A�ǰx`J��1��<җ��K#G�x��C�>�=���(��"��y}K��V��Zʾ�)�j��P'#����N�3'B�a_^�z��%K��D������5�OպDq3#]rx�0��2z��1L��nSa9�H����Y�cL�OX�jE�BN�F�W�kR�}�?J<��C�`@=*F�;g����	f���J�V�Ǻ���[�w_��V�oY�÷�c����5��['�X���9&���㤑��+�׷sc$��ntQq:vX49=�� ����~�z�=�)R*E�1ɋ��UIۖ\�Kp�t�|�������_��X�	�X��#Z��u$�t?�܋h�x��P:ݲ&�UE�t�+Պp�����v��whR-z+d@h`���bvı�S��*���������᝟m�מ��
�T, �V+���b����^ �G.&$�H7!��1��q���)�Z� ���p�Ϩjt���^2o���mc=g�*��qu&L�͗���zA����`�Qҷ&	eb�������ʰ��X�Z���0)�non��&��A!|���f�n��6U��A�h��h�6��}$�I���(Gאd?!V�8���/��ER���h�V��N�R���L��k��z'�O�O{��@��m��rB.��s�;Q7��'���O*��d��	���"�':��&Y��� 6���2�uNx��'}:�������_cK���:nҚEΘ�g\�Hz���_$��)^c�d�`�Yp{p
�.QK�-O>&��l������t1��A��#Ȝ���)���1�Y����aO�A�B�!�XudB��b.�r�B�2c���̅U ��4|�Tկ�Dǰ:�@���)^�4���_>e���:�[�}Ѿy��gd5�e0a&��	��U(���~�=Uf�/?$�򬊤"��pS�n�ґx�n[��^h��kK@�����j�DȈ�	��ж��J�}�땶�pa6������!w�~�����11���U���(�pʜ'။��+�:GFF*@�4��q�`]g�N��?��_���O�i#�
�w�5��2Y8��i^!��S�`o���^Y1)B�T�����N߆�R)Wϧ���V́��nN5�2#_�{��MVa`�o4l��:�:c�'��-�G�	���=�t��0yEI�nQ�EA(�<HpN5��@�A����(Ҳ��[�ч}�c_����i4�+�ݑM��� !E��X�^ �ҹ #2�2|������0�[Y!��sŴyyK
�\�T��v��0���E���'ϥ�A�,�W��;)��h����t�_HMӊY�T�N�(- ��v=��6��:7*4���ހb�><j���"���t�@��kp0�%gs$b�	Y͗�=�y㳛�QL�B�%�?zf8�E����?��V�����T8&��N��BW/�v�nG�'f��,�Wm(|�(��fpmcRف֓+�����Sڱ5�� ��'�7�݊f�K�(43� G��oک�~�w�-��z��xQjl�se)�� ���?�;������P���sRT2]���p��\6�6>�����4Z֤�y{��Q ߂��vC��J�!zks۔kB�����m�=�q��Y��A[o��9+y�!�񢼹�bFS�n���M�}M���m�`�g�sO��jy�m�m��SN[�JAY�h��b�[=#ݾ`H��z��6�;I	y��Tߨ�[7�ӯ����\�l_#}͊P�����_&©K���
h���<'��W��v����5�#�`~�ǐ@�c�PƖ �w��6Ԧݡ�}=�,O+���+�؁!�X��;Ѥ,H�ƺ�1v���%SQI*����1MKf�qy0�ּ	aF�J�L \�ؤ��
dE�x�J�q�9e��4�,y��廞`�F���n��h�;)��sa^?�3O[;&]��z^'p'q+���Z+����7���Mid�"�,�Х��H���TQr�.��_̇8�c634�7N�I�*	E�u���PFlZ�L꧃��.)�5��B�e��j{���Ȉ�ZѸ���%4��WAp����ķ��V��?�
+�$�P��ԝ�k0
/W�C�� B@����E�V�KuZSi��\w�"�u#�ĈW��Ƿ�	�4���1,x�_	�/�z�7r;�)���g�9���l�œm�b�;	Ys�I&a;��{��B�F��@V,P�;kv�T��� c��8Y $�)��70@u�Gr`q�7�>��������5$�r��GP׉yO�� �-;iKG�vqc��i���T�6֋]�%�A\rH?^�JHJ{N �
	�By�s2���nLk5#�j0�пl��a0�"���� ��b˞��X��{x����J�qS��+���-�x'(�{d��l���#�����2������݉c�ťsR�c	<�R�J����Р^�&�`�<-.y\�����D����n��؍�xKų�2��h�o�Nm#	�,��$o[e���?��	�Q�� ������<R�e���/A��I�rG���F�;��y�V��
��J8�����}�G�Lm�Y��HʊԖ�@��j���|^�0�\�Jn�qe��.'e��D/K��#;��.P=�sm8ʠ~�&�p䧏t��5>�Y;�=�律�~�?6�ҁ$X,�|y����i��'�ul����G���3��HjX~����`^]�3Z�O�|iF�},�=}Q~�
���1Ddd��h��Y�^�WcP�Bٔ���AZ��3�ě��#����5�9�3pn1�<��<N��d�h;
����[��a��ZVB�K��v�cO����K�}��0 ���#�4A��KWb�@�!�I���]�hS���J51�})��ǅvĭ�y�0�2�wlJ�2�FO�M�K٣���f����4�PO@�^"�i& <O�E2%j�N�}���}��Z��!�X���!\�'�N�!jO�K,D�nkl�"���,�>�֜��>m�=P�C1K�V�@�>��@��l��~y���6X��GEdRÔ� ��d����=�Q���̍W奷aR�0�l��̩l��H����h	���b�	%���vY�Vv&mr���ڨ[W��'�(r�c8�"\�_N�@)[g��p�B�}��:�X�@k�� m�l��)
�;��'��_j[]�AM�A��Ga���1n���#rp�:�I���-�:��3''{`��PV��m�&TX�w�9>x����<C�D��eR��|k����K�"����;�;LX���/2������v�t�B�e�֮�����玒��׍MC�Ǐ���7�^:���ը�	���9)��ra���á�=����4���k�/��KhCd�OB\^�f����Nt� uߞ*�����N�=�b�I.,5�:��a�1�z�i��H��ꉘঘ�g.�G\X ����P���;�fҌ�L�m�O�E�ډ߸�]	P��;�.��Jھ�ޚ��F|�~,�7�uN5���0й�tDRy��S`Y3F7v3<�X�Kx����x�R �
��g�f."� ��}V�5C������m�c�dU��@^z�m�R����EhZ����[� �f�)7^c��P�~�[4��z_ʴ�5�@,��'!5>^�Q��j����f�Op}2R�#�h�J�t=�(K`�a9[�}5(z�I͋*~��W684S3rU�Fo���aP`u�'�����Ɇ�{�k���Y:���!��][�d=Q]wXY���3�	��Ԩ�ɰ�!�"�Vj�	�^��ާ��Y)��9_�a;8Z��|f��ӂꃮ�m�/Ȟ�rV���5�5��X��rc���}������MQ��^�Q9�P�Rm��,0ĶH�d��k��w|�b0(쁝�D/�Mq����3l�[m�\�ܴ-h��;���+p���V��*�%���'E�_�i�U���#�Я�5�����8���H�� G�ԏ�LT*&�p��tX���+M��^`����ˍI*f�4k������\þ2�u��R9�TDNeɼ����_���elftr�1�J��}U��/�M�sL�7ut�&֏ �(A��TQA��TM������z��
ӵ9l�+��F"�.)���w����~��l\�q&�@�����uπ,%}�}��`�z�����:�C��C�ׁ�M^%�h���X������M,[��JN�}ؼ}�����^��M���?�z�P��0�ok%���y��jw}qP_�~�1vU��'���n�?2U���I&��C�:;�d���-�� �v1��
��ع�a�O�(b�_M3(1�r��scJ�Y k�%�_�o��ޑ��kΫ��ы�p�oͻ�<�'�.�f���I&��}�>x�Ɣ�T�����-�5��<�g4�%e.�O~��x��Xڞ�v ��?M�>^�O��@'��[o�H�h"�I��>����gs��a� ��[�.]\�Z!NS����x�bD�v���	���߿h��\����B�=}0R0��mD-H�4��?khހֆ)a)�}��*�tc�U)��$�:�8F�� ��%��>L(�d,Z��v��ł;:�؁.%�|��(Α	��z�KLm�})�U@��t�6��f�*�,`�6�HY��Thu��B��z�]��`h�ƾJ��O�sX�s�8��BG��}y�.Ӎ���(T���S_,�����C)������;$��6� �z6��b�E��(09s�;��.B����-�T�\�>癯>�g)ޯ�����\U~��gҍ��&rƹ#���g|�#3�c�w��|3���S�h`�"�G����@m/x7�$��U#�XK�N�L'�,Z&=�g�K��@�@4Z�k���Xˠ�ੈx�s��ѹ�W%�c���S~]q��z
�	~8��Sur��h��\^9�:�nrAt��7~٘�j�o$~���b>��_B_����PkZ��N�5�p2�]U%QH�%+�hZ��@�]��u�2г۹)C���!ءT�9E�@�.$�N�y�
F/f�U�iu�,9��q���r$۫��s��z�9;�+AɑU�]�uB���3�����8���|eM#�Ɓ	��sH.r�B�2�q����E��D��a��#��~"���?����e�NU��W��:�K}$F�+'��+��茆t��z��%�D7]흌3`�e+)�+�:a�(I���Zon߽�9閭+0��!yDT��Z��� N����|�}��7>q��n}�݉�R�zO�Ʃ�1������e����PN�B�)Q[�s��0H�bԧw�e�s.�DB;o]%󮀠Ȏ��}��U�9,2_�
�7?ߟ�����DD�8,��nD˦��n4r �P�X�h���w<��<��&'��]������~"�A��� �(�
�ï�-���@�0w��4�&1P�tcC��-p��@Y�("���N�u��t�'��R��"D�u_6f��^0���t�B�q���c��h$D|y��he��0��x�"t��B���@�.��J\�h4�}i�┹��)�9[^φ`����y\��mO�AD�Z����êys\Z�rP"��1�8IS���)�<S�� �_�
�-ɨO���iD�5�ep+��TC��L��{6]ԄL�* Jp&g���C�]2?�0=�3��Z(�[UUV��ѿ �����"��A�i�:j�!��[�-�T�8ޢ?Qh�W�o��y�SP� ��(xwUj��
+|O9L��s��#�J�IG� * <@q~]�[>N��$�H���:�[y����3O�X4��"cE���$u����J
|�^�_�Q��ο[q��1Z�no5?%9�5�pɅD�
��[X�x��L�2'��)��������<��]L����P�!��%�|[�ꬂ��Y���TOF�V�E�La:R[�攟(�>��!��'�#��5A<6��۫���ͮtY_�d�~�M�=�.�R�	������]����i!s�x��(�N�@:I�����m3�6�g��!֩^ya��GX�etV+��B��l�E�"�o|8B����J'�HFL�rH�l�#ON�R8�'��'f~�ꊔ�.1ʰ�w ����	��׶�I�>W�!�b�>��%fY�}��e���O{U���+?�_��#�k/��Z�P���Y��^������<`>�l�%�)��!�r��m���&T�f�0���6n�B� r���q���ۯ����\�/�Xó 6�w� ��Q^�F�x�����oe�P�����rtN�Jn��^��?�ʂ�$�F�Bi�ߞ!��cQPRb�"�B�иH\���0ԛ.�NLg>�zue�DL�fC�>�/��G^l��h����b����Qk�sY�6��i!�k"�8V����
����r�Uf���@<g:5�D�wA��й���;��ު��2�++B��Q=X,q�ۼO�[�^��#'8۠��w�/�H:�S)յ�C ;ؙh� -4y����|So�8E�6
_�ut�'YN2�]�9�e��$x�hp��#x5�y�~�D�㈖��^Jv@�­�Ϣ6�L:z9�^��,���*I�^�N��:�xݟR�>�e�#������`pLK��Zƈ�T>�O)�s�R�����UӤ����k�E�W��cT�9*�>�S�����̔RK�����7��FN��OtT�Y-�f��8:�ZS�k���� ���/�.��U���"�*�(R�Gz>����"	N2%-��L����E�e����