XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ċ����n��q<	�NF9����%���,���D�@�ڽe�p1;��Q��Epy�U��ϒ�z��dAX�ɥ�9�K*%[��/�׸�~*.t���6tvg��*@�=�H��+G��*O|�Vb'�1%���O�����S��*��:����:,�W3�		u��1J��İ�ɁX'���*Y�]��J�L���΢�jd7�^��dQJ�u�X�0{���nTz~�ݞ%f?�hր��1�y0vfO|�A�'��:T+����[��L~�:A:��`����������:�4b��꘰o���H�U�?f���)B��mW�A︄�S��A��j�7����HS�-�Es�X`�����B�#)X�h��3J��*Ao�f�Btw�9nZ�(:�2�0��1���Q���;��%���s�S��l�G��$���4ƛ���4B>��מɶ-�)'1�k�����P�u ��N��2����G�=�������Fq���Z��L�ޕ��O����Z�V�#O 8,�+i��R]i���K��"����l��Ȱ��D���ʬ"��x��M�,Q�+r��?A��cn�Ͱ2�#g�AT�`��Ҁ�W����Rf��P�'N�34D~d	?��9H�9Y�\�0��}������9�v�	���ş���OlS��.��iF\��>:�h��h.�t� �p�\� �4�~u����T�?�+���,�d7ϻ�:{���{���h�|j��������%eXlxVHYEB     400     1e0q?b9�i�ЈKw_�_H��(�3�.��OU#0tѢ+���<?�g�Ϧ{!)��/0�'K&�ۆ ^�����X��2�����.E��>f����oU8��-q���l͂O�G��AX�<Myx���:ၲZ8^1Q�(�_;��s�b��iX={��Py�m�"E�!�Y�3�O��T�Z�찏��$*T]�a��B�vj�Υ�*�Z��5>��?+qϟ�$�NV$��Y���EnBO0$�p�Al N6^7��e;Tl�΂f��Bیa���ͺ@wP�S!��
�j<�-=H�8j8�wt��v`���G4����)�����&^J 7���u81������m�bz�[�l���2K�m�N�Wi�lf�H��_V�ȷ�)��d�����%J���8��œ9r�w��޽9��E��>���}�����~�!&���|p8ۊ��-�k�B	Ʌ�) �������+�w�yI�C1B��C��6`C�XlxVHYEB     400     1f0�Pnup.7�ڒu�U|R�O/,��=;���F��e�$c��?;�o�`�����C�]�����씆v�'0 ��٢!ʝ�M������h`�Ύ��)�i�A�{t�u[K���yr���iu����I�'AH�(��œ�ĩ�P���">�;x�$o�P}�O��=��BbB9j�s2�`Nd���W�%�92z�]4B[��,��5y@j�R�i ��4CP��v�!�K���c�������wj&����V�}�>�i)����k�iPت�I�m�-#�4��p���#��jƬ�]("������鞸�=���!МoeJ79��Ԅ$�24+����֦���;	H ��a5qM��/�R�]����G.�Nf25=�䡨���Qh�5�~XlnI��Qi1��"w��]W*9��8���S�U��5�N�|��cJäf��'Y��Ih����	�7����q�Nk��w�{e�ѮK6�����7XlxVHYEB     400     1c0q���~��������d0��"pd����#Ѻ]v���l��9�:ixXE�K�n��C�{���ܰ�p����+'�'�'�'��+��>�ʹ���4ٟ_^�u�ҹϚι3�6rE�Uɲi���r�7��F�rr�o�!�d�yK�M�{b��� �_�Q��?C��9�)2㯯
��f��I�m,u5_+�f�B�;�z�4��kf�\`�O�RY��+�t�#U���&5�b�!�JΝ�'�l$-�)$�G�1�ħӋ��0B-�F��5hH�#3���Fen�����Q�&oQ���1R/p�eaPSN��-_}�D�PeV�B0�Ay�@K�D0�98�H<�	���F1÷+^�t�(���xF���1�E���d�w�%�� ��Z&�e�x�	�
tX����0�}&/���$�u�n��D�zRvQ/�
=�Q+����(XlxVHYEB     400     1d0�:QJ2`��Q#���(Ƣ!���dP-ʷ�WP}��xIN����}�3�nG~��<T�v���u�n�Q+)���!q{u���B�y?����f�)�8�������J��4D��U��V��AC�r9~.��+�yH��L�nM`3��	D��\�@�O�RHǇ�&��E�!�L�~@u�/���a�t��bi�i��z6o{I6�pD��4���{�f����F7���
��ĕ1�=�=���tY��jt�Ӧx5��j�ws$��ʈt�p��Oh�6_5d�Q�$������y�o�,�����bvS9I��\��h�ZCg��8[��Q0�X�*x54��cZ[�H٪����\�@�@�8g6?�ڍo�	�.�) %24*���l�]T+��T$�kRf��c�>��u���t��6q��s�$�	x*Z�V�J�p��A:I/o��|Z�A��@.#��`�XlxVHYEB     400     200iqYJY<4F4�,�~{,�f�密�r��O�b�;�Y�1��67V��k�`�ւ�<�&ߤ�4Q;��g3��wyp\~M .�q@QAp�
BŶf��@m�A�ķh<u���{��7ĄB_��w��$;�U��O剮�����w��c�Q-�iv����w����gN���t��(�i?2�^��)�r���pʓ��F=is:��䍹�0��䔡��\����_�V�^؄�P�Z�e@c�
̜K��+ǚ^�.�_E������ݣ����Qg3eO�M�+�)O�,#���X^�%Q��W��(���G�8�{5�},s��j�/Qt�`Fg�K��G.'��)��\W��;�T����K�׹az�^�An�kɆx��4���H�&آaf��~V����
�2e�r/3|Y�bc����^�Eb��p&������$�8��IY��;S�6���o��gF~m�ԟ���9��|��9��E�1`Nqc6�(r1����dP�������TXlxVHYEB     400     150��0�lp��!��h>\ �ȓ��O����Omf�u�{��%*?���wu0("�R#��1[��K�7�ce;?�e�:�z�&�#&��n�����W��n�&�!`ʖ���(�g^"x�,W��v�ca��	�^��-_T�9�^;��_��p,���+|S��+穋J�I�ꡀ������{�袙w���;�/�/g��`�_t^U
��@px�q7���n�b�f��X��|��}�z�E� ���ۤ5!Mh�}5�t���}c����6]��N�{x<i#�]F%��o�au���Eӵ��
`�F�y�b��F݁|�^���XlxVHYEB     400     170Iq��:�9�$B�ϾɽD�3��J�F@��M��7�0Ɠm�&�e�堊6���>Q�m��oL�o����ug!�K�_�g�[��l�\�n���<�]諝<��g��fn���iz�-�k�Ac��t��PP(h�g�S�����M��y��⩀xq�.��V��ACoc�]�@�ToX͔�	�Ց�(��Z0����^/�h�1d��70q8*O@+��;�� ��:���6~8mO�W���ʹ�rwN ��0^����%�^����
�yf.���؀si�jeJ�.��	���ٸ�5�ݱ\�}���7.��,���sC�o�PVN箫]s,^��Tv��hP�d�j�;�|��kXlxVHYEB     400     1d0���&�Z��v �����އ�P
����n�혙���Y�����p�ɒ$r���"�C��k0����ƈoȹ%V�#�}��c���V��B�����u�v��˦���9�����mGg�C�p�d�����(&�w�\k��}O��X�j�Cl�7Ȳ�;�ζTX�b�p�r��Гf/�F��->�]?��+�Y�TsHg�z�� �X%%81��
��#ZY��l����ha��D��l8�� P���m��)��s����Cd��6ꄵɒ�dT�d��C��O���]0M�p�u�LA�ޢ�[e���f�퓥Yg:D4�|��$7�Ŋy� �����ҥ�R�}��ؑ�?��xw��yv�S	�_cV�'�	� Q��n���!��U��*6����Bp�Ỡ�2V�$+�D$)�����2~@���	ݩddq[� #��vSDo/}�:� $HA'XlxVHYEB     400     190m��p��cc粑 �����ͨ�ȥ݁H1.u��]��?���aLd³����K�]�D��'�T�)|��s9��[����J�ہ����*Q_��"�8�b8��8{��v�bb#��웈'_վ��勿��ރ[X�f�.�Y�1��:�?r�fj��p#_�3�g`T�����)�����&2q5?�-�>ҭa�����-4ϩ3e�n?4�Mq�.|����t���1��7n�/�W���$�����5w��ѽ��I ̯�k��w��j��g�X��$8�Tnjξ'��v$��Ѽ��#��%�'D	1+�H!wT|�6Ĺ�c�ڟJ���
#���,�J8^��o�R�,�A���%��M.��P�k(ű�������/A�"�J;y�>��w�XlxVHYEB     400     190��Ŵ�b�?(�̌�f}tr9&%i7K<�u�g�FJN1j��$�<N�P������V�DJjl��[.Z�����9V��]����S��ӪB'G��jG��
�)�>��Se}=��!�Fu��n��9s��tL�#x�0G���`['���e�B�5���n�T8��.�]��䥂)gX�Z�x�#�l^Yh\���~�L�@��pS�?��mӧ��3STj��rX��/��(��*;U���{ȿ'�N�8^����=�OS���������3'~O�L�y��Q�j�/�'���E)�]���
�} }Ǖx�QD�J�^[T����F�V'# Sש-'u�k����f��N���͞���t#�l����3E�,��=XlxVHYEB     400     150*O�rLA�,�ZV�z�
�pW�Y�"�i��/�@��>_T:h~f�'u��*��T������pF�$��%��}��0��=Ax��d�qy��L�a>����3t����g�א�`�Y͛��!�U�wc�E4���� ���b�x?��+G7�ڸ����@��5@HA��Q��Ȧ�ѡ�`���l�S�>��X+P�%N��I�Էv�(���ߚ�~�ř���p�\�����_�*��F
K���ji*o���V���B�5FA[���X/[$����/����u�|މ3�tP� ���s�:ڦ�o����$�
7��~ˬ�qby[��XlxVHYEB     400     150f�>G�>�bs��UaѾݯ�Hw�Mu\�����Z�9QTh
���l|�9F�L�J�v��ҋ�?tM�@� p��z�D�"�q��vŗ|�x�'m'p�WX��P����;�6g��Ds���\}͎G{�P2�Hhf��~��r��x!0�&����7��2�Xxw��� �9����K|.-�����}rSC�Y�3bdYl.��≀�bQ���(����%5*��+ R�����)&����W/�Z��z�^��z��Mn��j� (9��$���F�H����C�=�k�´�>v�:j�'V&?�q� S�XR��(]"�ܴ��\�s�j��S��XlxVHYEB     400     1c0|6!��	M��2sƊ��.���� 
$X�Ξv���
Bc�(Zk��d�p�t����C�ZpPAIR����c�t\��kfe����2��r�H���*��9G]�6ɵ��qwі8\_7�O|g8�0�Y��;�9;��s'*�4�R_�[�%doA��c�@��k��Ì���A�^�d�;�E���f�{n�Uf�,��r_"X��=�/�5>-F`���m7���-/
l����F���ܪZ����\ɺ��
���d&^-숣Ct�<�HϺR�K�C�E�6����m����Պ^�@���LV(}��a�.���C�Ѷ����K0㦖3�Ͻ�g��p�r1��w�%����w��T8�S�.D�<����bE������oj�Jh�Z�y�� ~࿥�>�/2쪋��E[��i�6����֔�2"�\��~zQD{�J������XlxVHYEB     400     1c0F�-@uOox�m�������_mSS�;{g����=?��hx�f=�)�<vQ2W ��y���iZG��G�u�L!�a�I��B���1G Zg-��)m��n�%�55��]�φ6��*Q�5 �oK�"vz��Zz�����EQ�Cv,G�1k'�U�m��I�`}���ow�N²�7��)��WgD��Cn������E�������x�N�_�c�1+�0��[އ��l�]kZ�f\(��l7����Y0�c����Pkg�s�G
� ($�E�<>u��Ĺ�����Kr?O�>�����lr��k�"�5��_��&>�ߦ�m�����Zxh����Y�r�A8�#�S{�b,�VT�����{���(ޠ�*7�Kc`�a	Ij8�k�B'U�Xd�8Ǖ&��9�y"�_R�{1I0�:R8���&3F�#�$Fb]#���򵯱Z˓�XlxVHYEB     400     170�O�89:��7[':ˮ�aڦ2��sz ��+Z�������߻\`͍d��TF�~����5�芟P�FO9;�]�G�&��%d);К���?t���fz��7�0 �H�ɞ6����B�Gе�S�b���,���UFl��I6�Xua��F����(^'y�vh�*�+W\�>(	f�{�3qfNO����I7^��p���o��K���x�E���P� �&��^`K�ġ_C6����N���ۨTUG�+��h�T����1Ȧ+�@�%X�++�>u�د�rll��Ꮏ<%ˀ}k|�Mzx󲵗�g�G\t�ﳁ5��J��!�
ṙ��cz���;� A�L�S�k�m���%�1�twǢ��XlxVHYEB     400     200/�z�����`V�{|p�?]S�g!#��U�e�"&L�)�!h�U�o���#�־���-����L�~U4e��'~�[�k�Wp�N���yƊ�Z�iE��	]�:���JU�Q�dӈ��Q߳S�sR��;�)�w�o]hȶ�c�3�Z�c���,m%�`*�ڀ�k��r	@F����)��4�g���hIKѶ�/�������"���A[�ؠ�C+X]��+p穚�3� ��~�A��,�!EU�j�� L����Cv�.����icG�[�C)�V�dt��}i&�����U�j��>��e��8�J./��R���?#l�_����>��� lB�C�	&�)�̲^�c O�s!<#ږ��r%Խ����ܛM�܈~Y����6fLUS��')-��R*�5�v�`��/�λ��<-�
\;��3 kt_��_]t��ɀ�w���9�����~����5��n��i����P�I)���b��:;FF9���������^�xXlxVHYEB     400     210�",��!B�(-�&o"�2�!@e�z����G�nZX�>�vc�t���f�
�#P%��VJ�_�5�=� @X�V�ZQS��&�N�������o/u�@;3���0"-���Ӽ��y���#�w-�$���ݵ�C0ng%�Z6z��Q�^���y|_�i�͕I�NŚa�.���qlcx;�eJ	b���큃�m2�ܙY\�!^x�S���i!���yW���$�Wy��T�F:�7Ex�*��s��<U(z9x����(h�|�,�`�K49�l2��S�c�sz���|�LzԔpT�l�IpPc,"�H(�yPN`�~�-�0��Y/�Ί���	&���A5O�<�E������bO�|'���\���!>���C�&D�\Y�f4J�6�FǽxaY�mIy��d:>z}���^��!QF��i��)bD�t޴]�0%����Ʉ�#�5�
����;�I��Ll]z�ܭf̋ʵ�@�ad���x�oZ��������Ɠ���XlxVHYEB     400     1c0�q[:d���>h�0e��8����hsT)+�v;�-�Y�ۊ�a�&�����)Eq������O�7�<g�b��m����&�kSw��l̎�m�9���[�-��}��D�"�S�"�zy����tc��"��s{�	:J�j5#ʏ�4�F�m���^��<�1܆���w�T
�R�o�12#��y�Nl�n�WS��X�V��l383�o4�x
�8���pkG�ZqV�(�
;�|�^��Ph�n�Y����I�p5C���Eʧ	o�YCq��(�݉�##��H��X`�*x;xf��L>V�sa}R*�+Z ���a�~�N�y�Y
J����v��"����]�IM@W�����,
�N������+��V
��s������jj���!�SU�f��|����."�Y ��?iȓ�����Z	L��"<G�6����	@pp�7XlxVHYEB     400     160�z#`�5Id�]�x�Ba�t[�L'���쑗:R�3�"imȫ�T��<>c���T`v'������,�����lq�I��~�"�q�S<� ��?B��i�ׅl�,9�í˱���P<W��R�`'�s@��>l�Ǐ[vP2$��3�IQ��� �e촛���ZEQ���V�&]�~�]X�L����W�z���z����?='��q;f��ޔ��( \Ü�4I+����)�_��Y1H�,�;B�/W!v��׃��2Ց	��9�!vO.(g����n�[jþ������g��O-$���ގY�W��骢�U�%���"T.��XlxVHYEB     400     120C�?��Qe�������_���Q���el�t�r�Yb�F��u_�9�
����!d�'}%�c���B�Km�5,�+�R��Y�U�c� ��񍈍�������4c���4I=]�m�w������e��\o��<���� bh�ҾO(a#�Q-��J!�^�Eod�!�?���������Qm�*��0q���.V_���گ$�S�nw�&T<9G4A���D���e@kU�'�2]��{��h9�[�*Dh侵�_)�X+��AE*ظk�7)ˍe8�t0NXlxVHYEB     400     1607�C}$�F�-� �� 5�8���b�4�Vh�9�^��Qw�N����QA>�q�j�E�Ǜ��kCg�O��2�+������z|ɧ[&�"� c�7Ve�=�����7$u��~"�k���g���.�J?������mK:ܽ��/�
�c���l��ڻ����4�bB^Wግ�� ��H@kS�t|�C2<&�E����/�H]�=>�5S۫'�[,@F�ZPJ�����T�K�X!=��x��Á��U綵���s>ǺZM2�Q�C��Mй"#`K�!�썢��{FQ�˂L�w��cE��خ�ĜzFD�<ϦԈ�g_ԫ�xa.��"<!^	˰�σ�/�WF�eXlxVHYEB     400     160���������Kk�����+��m���6��i>��d�|�V	MLO�M{]:�s�Hh��)��)@i����+��jc��f�R���X~m����׵��8�'y�P�d>��(������k�~vǡHk����G�y��ز�H����JE�6m�9��!��zίԯ-��r���)+����mA='�"����q�gz�@�xL]��3�y����녺K5���7���jA�d��ˊ/v�*7�@m1v\�gj��C�`8I5��"t�H3bD¬�Q���1�hyMTv��(h�"������$������,EB���5��ua�A�a�j��\�QQ#�wQ��ғ&�(XlxVHYEB     400     200J��lS({G�}i����'�!b����N���!2Fkn	�_l�i+�� ��1Y��񗇡XA&J���7ʚƛgwV�M�4�E�6��<hjs���T&�ҟp�6GoN�\������t6�zJ+y��ݜ���|=�z�~�PqdnMx����X���:�X+c��n �X�XQ����1ph�(J�tz��j���s��~ul�	�U[�P���z0���$j(�X��0կ�}�a0j���h�'x�,y2�$R��}zu|8������_0Q(b��R��BA�tA��'��ͥ��
	�nYc].Ӣ 3�*�(2�"��MS9�*7}[
;,/ò'W�~���rq��&�n�����r�1�pe�����媧^��-����Z�+2��ڃ�J��^�g:���eM����!I�*��7�gHL���Ywģ��2\V�M�ni��bUNt^!p��D�u ��� Q�z��h�UPx#���"BW�g��U� r:�?��wQ��c�XlxVHYEB     400     1d0^e�P��Y�Þ�iز?�0����{HL:�8�7�dn�7r�&{�4�|O�V��J�8D�G(�ZPA�uM��+ ��=͸�<Yب���Z�������,ٙҲ�o?,)��o���j����Ʈ�J��I(��v�":5����������%8�:����,G������o��s �Q�zgC/� 	
��ZI߀�vM�m���\\�Ǭ>�bn�";r6+n*�H�C���J�t@��tEd����m^����&6n��D¼~.�[�Y��T�'x�2�@i��8#/�b*�� -T�v͈	��ӕS�j�<h�����^{ym���3E�7� 4+��2����c�'H��@T��|g'�B��v%y�2�)6�����9���^����"g-@�)�W?�/a���9%E��s�������٫��a/�ɣ�֕C�v$� ����@4�x5!R�DXlxVHYEB     400     1c0��C[�����Ӛ?��F��f5a�/# �����N(dc閺Y\';o�����X��{h�2�1��r��ٻ,�:��\�L;0��_;N
F�\,* �@��4�`�M�=�C�@f��;�8+~9t|�qҔ �p}O*}���6��1Z&~"$���XX�
��.z(dd��np���d��r۷"�e|�y*;R%!�=2��z����ͱ
���ۜ4���ǡ?\���^����z����.
'8H�M*�\��C^��2 )���T�#�t/$�Hr%�E�##�%��=����g��|�7�@����@%s%�ef1C��mQ�\�����$'=���n�Xb�2G������3�;��_�k����Cz�����9y���-�X?���˵;�3���59�@�Z`�[vm�i�^��u�ݿ=l
�XlxVHYEB      42      50�4#��g�X:`�r��H�������BK[`C���:�"���')�� ��ߋ�;M�FE���n���ĭ����4C		����