`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
M3XyT/ynG6I4Ck1Zu9rpefnR/G6iPbWRXYFzLKXaMvYcRHn2Ukmh+4prSLW+Qh1wRyG4YEvSLjzh
5hGGyQKJH54ziOwTu/Xw/QfGOzOzCet1BIZpKhJnmgEUqIQj/uolKgkD3/rWGEZVdHVcDmXNWjIG
RwdyR3D+j07glZSf0/yL0I8hXkFTq/lvzbUv+fGhl5fOKTfPjrC9zWUPqFZMItPZTLYOAntAwRrK
WLuLrviTRavvn8Zu8dqdtJ2bXmFie5cnE1vEPKNMjIQcj9yi4HcuIBs0kui/8CmT69yH9IISt1CX
x5xM3ddovO9j1iBX8UKQQsPVpQyiEDlVx+bOuhAQ45VgeLvnpRYlBLPLh2fzQ4o4KT7dUN+Nnqyn
wHcyZVhJhYlgi5ajVIxBd1flXpBb9A3xc4mWWHUkbcAyr1A2DO8/mqjs2o9iqH6kDXAuZ/hWOQMk
HKzAAJN/JnnbeRtKWJ/9gdGMNnUsGTQbJolf51bJ4CXQ2RLmPO6tHsk/SUnnup16lk9jb/V825zo
jcwkEVl12E1PJ4+KzpbGbQ14MikJyNIvLEDzagRIAet5KcZEnUfrOxy7Ic0rleszSl5EXtGUrY/Z
SPonBYaRIXC2Rqgb+sbZV+HBCfArDbCjqs1JAuHEuVTqT58brzuD6RLV88bRiFtk6UE61/Jk9vRA
7DODKkPHDl1JHodPUqKpG2N/h5yeAO1CH9nc3gHXZvB9F63WH0oFSN9EEHpl9ZOSIKO6E8r/OflI
rqINYAcfMcEv1zx9eofVmLP+EJ0vjLCMXaaigjkwi/7aaOlDdElNxZmejoHgRmfspi3H7TUpLtWg
QgN65bcRhPax25Nnq9gcG7NAQoQ5pID0bpkWfNbiaVAWrrCSNJXk/Hy7FcxX2O66qLpGBfaEh5Rg
Puvu0gmUFfEJFWfxTHB5RFYvmbnFhDERSMLELnNH3vpaTdwjQQ4HRrPMI2Y6A9Cc7R7fBDBCBAsC
INWgRJUDq+2sAdmIU7XXgxi8PBIGCIVI/eERs1QC2vYii4gQTH6gzVdcD7L1f19lYv6xArCgp4el
GAfGeEdiSdqg3U1lwDNFZI1+CC1k4Tb4ym2BckJlo1toBMNbc42qc7Nkb14MgFfC35RmqC5t5Cd8
AtWds7alJ7dJSoE6jJrpC+EFO6bC9DaQz7lgQ2ZgcRBA0CFbtpSrETcDB7HlwsqemvdMZjAZe+Mw
thzswxAWGdEjWGYYdAfOGNdxftreVe5I7+KkEacJ3SNsX0o0f4jPea/22im1IBvQ5rggzpA0dexa
9pZzWBa7fZyPZZoLfvf3cyNZEN7KAc/ijUfIbkDTkUIi6UmDNvN9UIVDNhDCFpE+skOuwkA63/I9
4762pmaukD59OPxZnVwMQwOw5xAuR8VVNfieiCoYEsIWhUyUCjw5nwBvahVvALiW8nsX6x42qIyw
WpwDtqJIKWhl1w3xfUMQiUySNC+ceK6tlwTVw65+3Cpvi+O9VN+5s0t4cEOoVJLM809+RXmrsE/I
ftYpWenjL0qk9k5F4JYk6T9hR/Wikl7HqsgrtFTOd2j8GEvg5tclj+B/LGHHXcBIsjAUFXg/ru/e
GJW3+QUQ7J082nluN7fI1r203y/i0laWe6MrQ8WbGp8N5psEXvNe94mEr74J4jEJeYMhUdZI4d/0
vJQxPvxnRE/f++q2sc6P5yQNF7z4CPzhN17QeC0WXY7NoUrb2k4YPI0p0aX2ymOtMrHrwA4gLady
J5GCnePFOqSvWADcIUf4VXEFVzU4fpr3gs1AIymZvagS2mN9dh19JBo1KuQ4KvGiWxt/bVe04G/o
ekX/OMyWcJEo0ULzakypnyM/gSnUYC793AZw6b/SdoRcTmCy51lc2olqCQB+Brfi0ljOJtGI16xM
qGWNq/wPUg8wUc2os80eUf0E3kRFzxn/YnQUgDp9WKXHmOtIWk/dX+hI7ZejS1Ve89Vx32OpSlLH
tT6KVRiSEuF0r76hgkpMb1G0tHOTvhkjb9suHw/N4tlSQNsfE8UEGx0dHuJEKHKbEfpgcOIMnedD
aM3wEWJ1tNJf2y3plEvYDyXr5zQGpypRXoJdf5ABVFA9du6hYe55IFte1oDjsWjvdV08ISXA/Isu
K2lC04oxgKwrVoJVz0fMTLW46dZRQCr+bqBr25aLFhKbT/QTxT6rjCP4CeZASzRAWVHmP5Bq5h6G
fk1Yb6Zk/WQgzCM6MKO4FIGNzMf9n/xYfPV3VCJupca0jGAIDKRymunZtEbyPFBXy/SG1n/mgZ8m
uOKlWWDQEJJPKOARCZsJL99FMEMWGKAPydQvlswbqjRi0Lv9SPOobT3gX/6rEmRwm2nAQas2+O8M
6Z1Li9wx2XWCqlimvBC3jjMjxEkbVWwU6FJg8RVG9eOkomLHxvRb56Y5J4cnQWlqqJMIwveaDnRE
FncO8MLLZ5ALaWjO3vdcz/iSlJLjmLmxHdVjws3SXbHKDA9w3i5clTCAzmhjv5Z9+FpQo/o97a6q
+eTcMitYP/z0isPD9asASHEKxMn68O3m4B7lnBo0KC8zxX7Mvna8r6x2V+em4ZYAgSf6+Q6oYomn
omnjaDS+cE/BGqSauMSS7M2bwhYk9XE2KfgpciQ7jOxOOiSaTJJowJTc4VK96mGBowTr4tMWlBQ9
KN8qPzIrbkAcdQPXBk3HgHV4Rf4fK6dH9K/FmB7El6xsuojyM9egWxffypEyXb+hsmUqyglnfvSF
STM/ZTOcMwVVcXH1sa+Wsiyv2xBOGRhqjzkWtoMxqnz6XH1LDX+9TGD3/vDHjFzpA2gIBfDeGfZZ
9+ypRQECPwZknRRWNtuzkXej5Djl+dcBBEBVhwkiVNTnbj77rmanvVPi0FSW43Sw2Basba+NskxR
IdvxW2oidr9DryhiQ9gXvnckNchdHILnKYW8Kf4EssCzdzJRsfcNj08rUffDOqILDta9WytCN1S/
FuhQedKbW2HRAxIWbHQmk/YiWwcmSl//1NLxutuEGeWyt1L4zrDi2B8+J+F0Ucg/q/6Jmahd1TsC
0NwPPqx8UuIspuNdaRl9MqdXkl7LHhLLqYHoTxmjmfMlvX7JmSTsmrpqATCcbHKsys6miiYDmXBY
NfsIZ/0oTixmJIVr3zesAWE0QWTqgrwxDWamUnpvkbzY3fIkh7S6gUlsPjBtOOfMrKfZ8wp9S2s+
xMQvpfb5fMHj7mV9+JjD8bCGw04MRMiyRnr0wetl2OjhLN14kq+g4mYLSKR0ZMqxOS3W6Kt8AxGj
/Roo5DLr4/KeYewdNQ4rRK3dcZgMKKRLzbvBugkNrGJAlfYuoERPOiqTXeRL6EHPmnSxfmlZnq1t
jIgDiJGw0wfFW9cg28KOIT/KPsMUJIk4VOXNQeD6gmtT8GdzADOa/WarWABMDtgdNC+ICjVrFKqs
Gbk5hofzMhPy1+CpWgh3hGWSbmaOjefPboTjvGfaz14RoDHezkO3QnbzYLh7FonLG+jX7Ziao6te
CWSb1V26nwQg9OsGeopRKCvllr7f3v5ZW7y2COGk8YabUwVaXMSm2G8A+XmtMHZqQYiJ5VPJGV2S
hKi2QyPwu3v986gMceAqz5OBBHLJZ59v149JayC3E2537aEJGe4xRgELuFF0h8TUQxGtkhyhgksz
BPHzi9H+GGltrBFCckAkaprUS8To5Y/O9JjgF1mCFNN0CHqWbexfSBUuABf3PFG2NBX40MimTFMA
FPQPZ1q3ovb95eaoTcbZVmr7lcQ8/yXQRSILzNiPX4r/cfrzDsGdpmLlnk7ngpTKhbaSSAdTkNub
oMpcjelgwp1FuxXkI0jivKlYUwjkFMKFbQw01lJDSELQezkDKmKlgunmsRSyHDa5bXhh1y51btdV
q4ZTcc22uUfIMf0V0WEZy0uikTM3NQsXlXQNxPf+j9ad5VCZJjejtRazLLVcbEKr8hWAUY7X7Fu3
rMTCXrPeQpZkmngA4CDty8ppXOic16FQ3Rt/FGTAU/uXK3VhtzSIdFXROkYpZwtlYvW5Ll4TJZYM
n/LZE3QAEejVkoOOjg6XQn7ZVHoF9WO45ACVF1sUZPxuMTqMKL6kGF5ewJtf8V9bmSHle/v4ESaS
rTqDsFNaiNQ1tXtDxNTqkDNbw8cTg1byTXJUUNH8hV401PRre2l/AVwAJoXbnacKptuvuMGHpt9B
ZaheNSgxihklRQ5v0KGabtyDN84XYS+s89IIuc/dSFmnSc/mk4oKGT/p5GseG9DqLBVAevIP+ymr
qUsf/xtMfO1Flc7xdYOMqkbMVmp6ZwbrW9AhJdsNUEWMQ44XDoSkMmJ1W/T7tGP1W0f6UOxIvqMp
R/R/UcDt2fFYDQZCGR0EHei+4iuluvh345uE/+QqitIsGnJw2TJ9uoTdqgMsuzzEdz0BSwbQmB3o
k0ZDnF+ZrCqMNs9ukXhXRixNjsuDZCT1RR0b0AmSjC3eGtWhkQzQwcFivoNofqqmMGoQ0j0BrW53
V+WiH4B3pYS/NL0iifvSMoHOcTR0pEHgbe0mXxMGcnJT7BR/wJdhlo8w87hJq9rO6xVjFJJYZWzp
85q9Ke+0kjpKe7nASDLFHtjhL/vxyA7i7V/Rdya/KLHstQYxQpsHKbkgN1C1zuhfigFoogGscobA
MvLub6QGMVkFOn6I+jzBJxXH3T6EzPn9uFLkg7VqKsSxnWeY39QtiFRrxaN2AEYbIHMISlGaQtSH
OhhPUiXL386Qqtnz3q5qyOli82d2pX3lYbccH5Pmy6kDst6glWSHwth2JiupIuXMToLu3iNNFJew
T6o0TF40beDaKfwfEMqLbAl20/qvDgUjtguZERlnYXm/rBTsquNW9u3iZwt7wgZn7JVy9gZDnI4f
b8Nq6mUSvZDGQ8MUS06+DgMsPdowTu2PjX2t4w5unGvCIGE5G6qoFc4SvUe4HRHewTy1envKoZJy
LGn2sSQYDd2BPXdFNcfdwCYs3Tw5QwCTo1teMqfV5M5+wydC6NhepGMmhu/oOuuyirOrSECjXSTk
4PBm+mGRHxyH7p8rdVUks1SzI8sBFOObljzOw7PkRSQrWbWML4RmwDJWjoknxgmjXBmsh/coB7QJ
36EvfOWXfJepWsbF7j2NlnsdiFlRGA6b9Ce+pnXUWD6PC026Q6msaPUGu+Qy5l97vf0AU1+GdQFa
RMZHaYrsJitoYcmTUaXiMWvoN05sWNS3WM6uT6A/FETGl8Xx+fqyrQUvCLU9Vl/uthOvajyBHzZV
5wsz5z6LGlW/pbVXIt7HtRSikBmWxs3/XRwvbsp4lmf6YajA4oj6zWe943u5OVFPKXRWPlKX9oPC
QkhT749wzV/4LWIDShRLGZ70fDCFybEkZ3so5qiGi/kMKv4gumdqh4/NIwzCkG8yJubOP/M625X8
6bavZMyrcq4G/m8pbMxPO4gpCg0EqJ/sboQrR498kAf7PfEU9Z/XsfUMus0U3g4VVkHePtmH5gEz
PaW17/X5FKia/RHelXzAbtb1DVjeiS0xMvugcDUK2V7Aoiud43BIuTRUawSjh/oVJslDm1cR6H3W
TD+W2vt6MVSFvrKxZOfsqzymbb5FBCxxILxpGmxaTe8mBEX70Us5EnmjyXI0YCBPvbQ3j+NeyKuc
Ma8BsYYMDGwVikdagJmIUlHcDBELcRL9Reo8AfA9GIXc4INfR0btunddmf57OA9rGYGK2gslxweT
Tt60DvjBGXI4czGDjVYDZMvhg6NI/4VWUbWfaycTTKapq2OD0MF+6VWyFtfPnIWAbueHRMqEhd5n
iUXRQIvgscFd1N00vLkooNF2aCIVW3HDAUcZj+mMGJgZKmn43mEEiS/Ua+ZbszOXTRDEFh0QwuWJ
wAbfyorTv+AjQpq2h9VmtTufb9cpsMWR6dGPbwUEvdkfjMRBn3ShHuEL0K/92QsLOZgCHqb4IUvl
GZU+tBWHeVTXI+to/24QMrf2kumwoJnN8KlmfxQ/3ENhDjaBTPTJT53DgwGqy8ERZlOqMpXDfviY
oiSa9DRC1+KiDrVS3/4N+yfQK8Zi3cpcxH/VfUXeb5KE2uhHTWeRn3yxiYxewFhbYHQskWby5mOA
lZzHbYWRqfWrbTtdFvu1iuqfSSN+zBiTolqdnWMndr72vuKxdSnnIqzFnRh7c2YtfJ1s/J90Tvv9
8Dq9Mp8h40zsCT86ZzBr7PC4dOsseO9y1n95669AoYkhCKtwGczkJWogb+pZlGUpyuSC5a3uBEcB
U+bmdIoBft3Bk7TVGHyB982WxTLNgTqCpx+I+G5yutY+rapa9XPM7WRvLBYJ76sxhVyKdfzkSvUj
ErpawHmgeRU60/dghb2HClio1FpfZJlng9gryEyJ/PV4jHE4hNSlhn07fq7ucysjvsDvBYz2xxas
WauMXBPt6ldbYoKh+VQhPckv9DcdU2ir1hKIkuGwBQIYTiWKtr3GCfxJWmEPmXnjmMpUEJrkm302
FfsyTvo8f5aAXzr6v6LRuvlA6g3HDwuE5+uZu7feOaLYDp1DVl9OwfTPPJr0BC+sqK+ozGvRrVWc
DLHKEIvi3kmCw1IbkLvXeUUlNb6t9h29+aeWQ4M15eXE32fCsrankZETrKYvNBRLj5O2ZtPQ9oZM
sFTxIektDaYUk9JW1rYzNzq7Ehi1Y4EoBvgcKNVRyElr+I0jQrLRtiY98YxfZMkcV+EVtt0yUu7t
Qux+dILD1JMRxivN3PR4a/+i9mMZQE9nxwzKn11noRuccKnan6l96k2ewt0Du5pZFP2SqHRM/6YN
JhrSDZJq+22sOujkmI513vNGRncwhyJkuUhlmE5MZwHbzwSGr2+W0HIqY8vQ3AYMNl2/mfe/zyiv
uYVWIdPQkwxFWr1pXIq4Xqhm6X5zu8dE1kVQCqfiBcJMs2s73GMlGo45VeR+dgJDN14aDyhPZnLo
zkjxKfZ3M4+13IC9dewP6zG960kgUOb/2Umq3QsN5j+8I9SqRphHjchsYSVw6AM25wySPfA15P9n
xiwqo/agg+deuYqO1r79g96Q0P0T86ThqJwPXrqe043kfRXe29SmWHW/t4CnNtbfp19xnziV+3+2
Nc1DhzpF5uhLTNNXY0kkbLq8Rq32GoD4u597B9g18t4WHhS7xTNNzJYQsE97sOzLt48p9e+Qs0EG
HqigXp01bpmcksVlTdLOCvD7LD13v0+6+AAamwjnyTp3K68XgEDqmVSKlazdxGMAVsz7ZRz7k+34
bippzZMygX9GSOBpj4nKSgRFag24V1yXWGwxlqaBbD1NMV4hzzdlzW9LuGoT43ebvFzA3w49ZMqO
0Q/4+fLeYdpi/4zCtzz3aY13b1A6frcNDmaNFA25ftj6ciOQPlj9xpy1uGwlxUSAAOh6TuFRZjRr
4fDdBkj5vqsfMzU2czTCRCDntAYDbTZv5S7tOA3nmaeHBLKGG6kqdd89hgEXqqHsv1t2QrHPdfKV
DK8iaO5UoZdMlwrrg3zXFJQ54xxVQitn9g+02ASNQfA9Z30MAGENG+TJw6yatr60CrKD0mVZps10
1iafuSMmYqEKaz7k2kHZYBKmDQtpsQAvEvtE1nfEgBkcHGQCbJKEW9eNSO2l+Tqy8c/vxiVFVcyX
dkkFdGpi8ZlZwRJgybj48OzWgyId/v4Y+n05GfcdQXT/kuXodmcpUEUh3g1SpypmG1XG+DpDV8DR
KVhlhvlVmW3VL6xyp1QGNQEdv+YW7wtTE08Zc61Tcdo6/iAIUSIEeBVzBSq7Ptgsd5vVrBgu5v95
jBKUKYetCVX31qMREYQWtzDXrcrE/BTqk27FBSSzEH+quSUjRhdtqiNdngfHGS8erbnldYYd1Rms
0jO+5tqEBy0L8SJGBrTCPZkAIquaToVR6AKK3RxYoN7gCsKq0rrxRzbMSeEd8/tU3fbVD8aZlQxD
JaCrPRjgyGnO3nG/kknA07VoT8Qby/fUAoRq9E+rB1ppzeWeLsPtXhkO0+mbsHQ7c+VLwM4rKmKV
cbn8hWmzw/GIforLbGfvjlgP5y8bmVEbVuUkw69Z/Ktr1LWJoDYey4nM3W0fDpXbY01/peLskyxd
YvecPkzVPRo4zw1DeAHLoJtRDDpwBWqPsen4Rc8MnWG4ATwxwBOjvnrsO3BK8Tm2t5NMLPKTVfcV
nctB0S4L/C5hLQHsrQlpTn9Sf+BPfBG+0ABtdYrU0yavhmuj1ccesN8+6mt7kSfI15fpJzuBoTT+
lYHfsahXCZro9AUSuSObYMJREH10NC3TDJeknTVlpiLIJa1EbHM7I8BR4ELGGS+EhmwDrT0Sffv8
acm7cULribmkZq3e9ZsSV5iYqxd2Vl/amK0t0jbJslEmxqaefAfRkaNcNRx5gsZCSu3JEqHeBsms
gStYtas4wW7wAKkaCsWKMl7BAFMdOpYSj/XOhGZLEOCN5ukHe0j8g+nWfBegiJ36+AIDwC5vgR/e
XLiTkyaJH/cjpA/+XQSun0x0PD6pCALfggsQrpN6xLiy9AUr8pMTla3PCt1nyC3V0HP25N9YtLNP
yzOuecwdhq6uPV1co+SKz3AhhF+mEHhkCrbmte0eYXsMPmIXVp0Qo0ksuky7JD9GERgMrMNYrVnc
1c15ubclkqzGOUK4qJkgaYnBqLnEVbb6E6N+KMxq+oVJru/C1Q57qAlpHc8KPsjB2cDoWK3qsviK
UilbQtZVKTvctup56+YYfFtd79ihZBNSn2E0y9cLmU674LUPqOewjotOyU27Z5t/wnO4m3N+aUdA
9uE0VtLbhkoxL3R0/5FV6XVof6ZUfJnR1AjvWhqB8nEJ1JtiuFZkJxqesZG/ZDyY2BQT6f0BNZ4m
ux15Tde3pbbXMfXM0Xtx0ECKqli9gN4sXLkRSJ4+eBMQdhwWKc/KuBJ6//8sd5PW6NgTaypxIjkA
Eccu7nhGdYdYLYYtQMSOFJRAip/TMTQ0ef2k8V2ULkU0RPMix2OtJRjN8thyhBxZV6YhyJ+WnOnJ
j29hjkic6UlL9UFaYjXnR+00lwzhwzh0BBAmAJYgd5hKLzgFoRFUbR6ga7mboXpzWJG/OyshUIY8
Il2cu9SHhmoCZuMzqQAnMEnH2Jhd5xm+OATeKkKc7bxvSTdI2njkv2/s8+zeWtZbn9mwloYtg+Bh
F3vOsOlMvXpKGz6CcrlLGyNUg0JZmMfeVuPwblHh6BCao6dmhT5EF/c+z6y02yU29loE9u0IUx+Y
6hTpJ3+cXPnQDSunlVlMCIgaE5NG5deVJ56jE0Xbc6zSZ1gmh8Ad4zQhGjKJbdXaG5jVgS6NrOw4
5Ydi9nL1ReETDRAA7hoXyx4zQUU3zK+Q82vHZkg0ahOZ72iZp69qR/XlCKo3Z07qpXnfNFWvaxi/
3sX9NoNluATaYtvca3F9cE3RAACku90UbzWVVmrUPFCDDq16ZcxwUCU+4QhzSCarNgSEe4urUWQO
pM2Mh0NfJyeyaHjy4SVZcn+5kLkATiKFSIAQoRLVaPNAQh0mZ+D7ioMM/7kT60nc3/46HNU6d6eK
xJSlIBOzXBn4BnW6aIL5EjwbRsz4fWpzo7hJPgYaCoQtyltNCFH6kH+JlkysggyeBQaN6yq0CvYG
y/HGpDxox1NgkNJvSsUXWrEXNUhHR3LIb/miRR35M5ntnz0zEREYSgJg+IB1U61bsekB24kMal3k
st8Gyj7IkGJ9Bssfi4Ocr+eIBSe7uhAELBI/WyUNXQtKmxQF0tWGNEr6HvzzW5PBR0ppzr0v5EH5
bShkCEKQ4WW6wJC6dQI7ol/Uyvf93Af4GwxBSCknhYYSUk4dQy/3YmCk8ofNHgpz5NPz/qbHnN1X
Lp4TKD63UyzVEX46rUJMtQrHPiRMgZ4bOMWzR1aFH2FHIySnJhLUr5B0VBTDLsFdIk2/eDGn0VZe
gzM6uGiDi/aIS/lB1BknBs71QFlU29sX7oNjl4+TuyE0LzjxrvuEouKsf/C/tWCBMpJWsUMS0i5x
ZqVjfdMHq450VMKd72/gM3fmYu/eP8XzYvHktR8O40xSQ8wCbTJo2gLWuDeVDpFPIWSLhqKpsRUw
gs4iYq1wXDfwi7SkIDf6evwqGJEfUSvImrDygPZZfi5rq4OsFWeebUW7Btu0zz/SX5/x0SUG7JxE
zbe41nguao/vwg3yibU9/vk5HFm+6coao8u/7ekqKBp/uOLd42vAXcJEahOPkBbohK0lhUEFmybp
JuEdvivYGQMVvrn925kZxr5xu1EIL8na9FBhFofw1PAce4uyHEJVpNdoEsZ0fdSv4jkY5esUQX78
6uKNPTQepnX+/B0DaCLhqqMpQV4/yvzzngTlYXdMjI8+8dQxrrryTqMFbV7b0tu2a7BlDT+PduI2
Pt9Usud8SZBqhLVATwsDeCPfH+71Ys77VK1MyLPKesKByZkQqCf6n2FUZJI3eZHye0kD1h9mBcWg
WD5fPv45QZwPX/N/cqmmDPZ4Z4y4xpmlBOavOaTNHd3zTKt26/Jb4skIUXp3BibnFzQjqW5A+jlT
XSliz+RGqxezy++W3jJDXkWNoitAHdc0Yr8+zFiHWq3JVc1FcfNX9uce6WOtIraEL1e8iINuUOyD
AYKrsKmBs5a9qOo1RRNa3xH6ZKtvcCuoeDyseoz+Q2Bx5XAjqBOy/00WfVMMGokbDnqkSns2Vr3k
sba0x1LklpjfRclZyO0MiUwzvttZEsdo+ymbCRDZyPfgDSQGRKSxgd9li8h4anRi+a2wyN/r7Nw2
1xyujD2CeRNLIN8gWFPHkqjLduelc7L1aHVOllUTyn/Wh+R4SgiKi2D4R0ME8oOgpFbOkT5vaRqL
MvP8oy3laBHQHpd8+6uVd8tAvVbr+L7O/CWYUvQsjqVkHGU7PULZTVz7YCXMpcVlNo8x3NUji30r
jj+6Qh+heKxvp2ewMjtLsteCPwOdDtaljlEygMxNizuYITH+qfZ9uDlnPbCOWV9BbhzO4YLfqRe/
SCzKWN8vDX0u9qVjqcKCRpXH/COwzODO8nct7mLQxZU48DVhv+IDdinxuCsJmaZBtCURf/3xq30T
dzYiJfp4OPVrZI3VTYo2HYG8U2hBCBNosttcPPZOBVRekcldQL/WYuQsSp9GKZwZxpT1iIoe7gCc
13XSmaZ4PvQxyRXopRoUOKd52+XB6DBCT1igPolzT9ysktfsLC/NcEXJCQyqKrx5HbwJlNdqkGMn
/F0hVvBJ6FB04ZgdY4voGh3qtWlY
`protect end_protected
