`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 100176)
`protect data_block
/80mKLS2nh9UUBikn8H0CEObJMyEi0OTgrwD/qUZMN9cONGeoWiFdspwjYWRAotVTfa2p/HC4mQq
rEnDTGnaPEZwRxKn8qP6SbTmyTX3oXmEnkw4uNHRhJJHCwXcXLiKrvUmSbRKOziVn5wSxCsjkmAK
qdivvGHmMDe+mq4IgQmFLTyXxVNL4lmcOx+6IIjBkfomUMw66xgyKpZxgFYQer/rygGvzltCw9WW
wmkNjt2r+HBBEmxPgC07ICGu5keQpjbblbDD8VDFoCQNXXFajzYfmGlp4NRAU13iE4VHHyhUV02O
nV+0f2ySKXw86hhN7fdv+qmnjmKlAVu4JJdNUSAdZSTivroY/vQmOEGsaq3qi4dRGDHharthqxyA
NgiGEUR9BC+Ko5colIcsBjrPN85thbtUXgGTwCGPqEEmBPl7ytLFQFhSKcKXz8MET8VVE+x8l5DF
s4mr4LLW0ll0ECk7oZXpR+5LpLsj+mIvvG0jbTTyr0fVtPd1ycPpZDuGmzr5f9WD8GplCFmYVqKO
4oh+xw38KAtXVIfFAeEOBaK7PaLNz2uZrtOE+msqKB00oW85AdqjtNUW41DRkUnSwmvcnZER40xd
85tjfcAXM9VSFGwAkm+wmDxsjIa4ogeeS4cCBDWz3debOpYW3fHL/NB3YXVFUDYH0S/MOwnfyzkG
MNCAHJdiYiBs78EuGVN7FweXlsYEkbwUnDwErJ6cdmj+C7xldxhnjA3/HdmdwloED4DHXbYsqBau
haJaEVfJFUwIOOeJmnnkkl3+3Ho+CjIdVwNNj0YzcFI2G5KtVHeI20UODk1N9KB0GBoSgnmI4GjB
Z+iCil+AjwJndcIeZ4e7xW33KRHuhZZkQN69g0XK2NN4RtBeSMLUIHLCtvKvlVu8phC87ZUavutr
F51Vhoj1ZgYEOaiQYYFgmvrZDJA3lq56CcekdGzXtBxoMJrL8oqeVJ6Ep2GrM/kIKOh2Kji/i4ZQ
Peh28V2cBTyss51RgAa1h1pU0uivz1WHIfpoaCMh8lVCNrJ5e1or8CLwt+uX/MKxXAKKS4crtMyE
iahXRFXdqRG6imuOiohr5lS03lvbnzjJH054dfUQqTiU+39J6ElEKhpdFb/L0U+gfBS4gMuD4lYJ
/l/k7nia5Pf5sxSklcGqSH0bS9JqX/A3DunUfLjspt2wT3+DrV71Zuu3+cg0v7ieQfW1+g5V3bJf
6G5jYeginh53gaaWMdFJXwVQy/MOCysu+AM2kN2pbSeCxXu20bW/2HCsQ7rqiO9JluOdmQ9hxsEi
1Dvcw1ch8ea2Wpoqx9GeaoeDQXQdTLU57/S+7EGbtkZ0DJhlkBrisGF9q0cZEOoaVso52gWtnRsv
k/sPlSOWc91/GuRJvBlU5Z7xigtfqqa/78EWHSUk8ITQlPiWjLNBWSaSAtOwrBFP45AnVpiLRLQY
DeymhuiAKw1oDxYy5oGo/ql2NogipZT+KX3sFIKpQnc59MFjSBouONHE3eXdYOfKtkbi1whoLw8Y
DPveZ8ataf2+lPLQMrIILqlxOnzs8FSFFuMMDYFttAna+N1wWHgIwk6n0bhthqyCIF6o5oH9TUTf
TdS3nXc/ld44ZC+vnhioQo+qPT8vzBPM28Cuba66FWcyPPdmjO2fwr/wRvzCtfOoO2lztZbNcmsy
go2BZdl0ohh4RUYN26kEzORD93OD3zzAxxniscItoHk5ERQfr3OnkUEtNUK55wfffymLIaN6BLro
B3r1zm7aGIzrbmwxqDqM3UNQL2m8Trl9lBMD3q/3YNCqrjzyfzunGvXRU1JAQccIKotUMjhnkXWJ
k2Fa0M/hpjnrBTvTxXz+WaOm8uKG5eMdRM2vcQn7O+LyZyQHdpi2ZjauAsV1946JviYu73TwU+BI
C1+AX2KdTcC26RlLbijQOOlYOsZ5Oy7094AZNE4x8xMCVIF7gmN++alOPecp/uvQ1ZHr6BqutyXy
IHrHslo9x7ahTevVX7yQsDLOEqXyVGORyJ5UYKBAZuE/hie7JGG0PZ0tUHtDRJSCWtstkdY99em5
Dog58/ZWAQ8CgQn7AUhAHXaYEg8waKv5wOehN4fYUALeYolw3SvRanYgxp2TiDkhT9W7t+gtKBD7
QRv5ZsZAzjc8ndt8WFVyF+iCmPO8DPECE1+8oP5Hojz0d8jMvhFT/c2h6r/LhU0ymbo2RkeS4CEj
UkWPINVJlMxF3prFIqttkrFIIHOBo/qxecaw3fxP5kAlNoNZgHbBnJRguMudkIzscqkDFCOpxKHS
slQiW3rHoAMX3yi++Ru2mn9DcD45x9C3Dskyfw5Zu8JZp9B23JRDBSABzYafs1+P0Y0mWSS0xER4
d99ZqnWflFsvLlw3bADEgQPWtMbmMHTZlqrASPbqBKQ+wWL2DhMcTotj/e0gGZyD0sMtFW4mJcvQ
lRYXUivCSXXFumFtHjRbanLUdN7Sbk9qkaCtPHjSmMuYtS2wJghQ/YBgcu42J1n/Wk5gNtKjCbJc
4RuP5xQuRr/Qk3dEp/iAjJdjEfUiHvX/zu1kK7svyh2zjMhZPAVCaIeHXBhbQr6eOf92RqdG/hwQ
U1+JgeeUFUG+GZ4I8vDdKHBsTq3PiPzDHbdhOQBWwkZGGBt2+BkX8yMGk91t2Q9c/MCEInSQmXCL
NGnOVsUA6WZtj35Jukvi8a4pPzG2t7ddS3PO/GX1X8VZ9r5h/x/vnOd2XD8xE6KuSWxtJZ9ZaKUA
v17BFMzFALHsRgzs13eZd5PKjY7jZ6IW9aVqn7pjyvRnKSyBI/grLsLhg9w9GqGUtEavKdBmKQm3
R0FK33Yb+Udk2og0RvutK7Un8xIv+WhADtwTWVhigLPOsv0P+bCw6McJ3I6BiM04PAiwfMfDBvlg
F7m/gCr7X/OAndr4mdtnuVcuWEET9bddxcOsx7lB5+ruNzlQg4Dsvvx31WmRhaBmXxTC7s3IX3sn
sQ1yfLdwOs3Ouj6iy0jEI6ECpCIHs41y8maollk5PzufOylegreVPiEgTpfZW5W7YYMvoq3gN88w
TXbgPNnXWLliGb5brEjAoqAPWNk9dpETlnatMeb8HlLF6WoK6Sh3n/jj65L1WWTL8fuFwuIbpk76
9JNna29m0rhmrzF+sxHQCQU71dvA+wL9dIA7UxOzrRry1LVJO7YEo2SVB5Y0XD2jK/pnvXeu8gb/
U7VW2f7lZO2w9yyzYAiZOuzesPZXCeAvI5pBM4v2vrqr5T6L/0hUYqZ80p7fXjHHy3DiaZtHwNoV
b/XhP9M9EVvmwv094bOWvYdZg1QzRn+aDBALuDdNnrGxL/HW+Yk6r6ZTG4dXks7GDgLlxpZIyZDK
+kbZdxUjmpfuaOPELAFjTKXN7CT8VtnHQ1mCgkXBG9YMgAGQlf1RUu2HIVzaNsbCyaahTeSAdNCK
md8kBWq7km8eITm+juVl693Br5+QsbGQZuxxsapIe3b9Y8BnP11q9Lbhilcr1lNtlRaATh0uF6+4
za+rgSHHGwmbBthssWy7bJBOrPQvfhL+XAP4CsTmQhnmDeNVv1pM8lvXbd86MH+hlPWn4sLsxAB6
QnGYLXCqip+bxzT3vAMit6mKpMz2Q97qI1IPQDY5jdBT0k1DZ3eVoDxE6F+fnFiTBBCJH2464ol/
yZuJIhdHC/TTsA64BsSU4pjtM71XSp72GqOu7GasvNrQTnp+Cl2F9tYzYK8exvMFUezDSHt0qLVv
oWXsfqHWqMYYQzyOAwP2Cpxk54S3tVOe4M85LCL96tdbs/YGn5Hqvvpm5bI2sUAz0s+A+oIcJBxh
/nHYDk1efz6NhMU5xUtG1Ck7yXzELfGx24y1c874ZjgyUztAK1KBY/HpGeAj3pjjzx7vyn+0AXQ8
jh/pYmdt9xXyk5r5ym7Gh4OC+5iSDTfyhsw+wNOdnJqrloMpARXbGBKhgjmjLgaUGke0ViNKOZyx
bQ8qzl7oMANTNq0WdSDgAffBv+t1k1+U2ZCqFsA2Qn/trRxUpEjUCm4jrBvA58lQkwRpKEraBjrT
2wtwhw9WlSPEASE/ITQR3ZqIpQ+J0HkCA0U2fidwBROrWEkl4EV7OIe5IZjQ5ZBjRaQ+1X0gjkxA
UcAuAc0z9RERBhc0A5V/+AgUuujjtRwGhDLWo5VJSUOeThAftC7lmowyA9N7JTZqbBwrC+2NAOu0
L440kxIID7vEbrWAAglgXBtw0qaE10rhyz/lM2leT4GRJ6FWkarszi6N8Bmd44HGdCl7hnHURw7Z
R/pMABXnnVwDmQAACcx9hpiWUAtvoux7XFuszqfAyhWxS/YbGwsMMx0/Ue7+AEfp8MqOoD+5Lnli
CQpPSDXbk3b0thf6a1q8HPP2m4fvZviQlvquia/7GrfO+SDLzcNBYrVSbnm+A9nSROt0xWiY1E5j
6dei6YoHzoisateYmJGhPlgD/B3EqHVLgWXRNB/Zarru60p1eLnBoGV4yzgQFP/oydEZVCRdSd19
gX1r+11oSMCiYjE86znMfGKLQDmqXhzpLJE3nBXPWyqT7Z8PC4yvTa5YMHqtfCG0/KplwXXcJt30
drJU2pRFJZ5lZf9fpo96mbk7kA9CaraEhzVQ7kxS84iqjoDhvVGOgImUxM8wUA5NXc9hDda1sdz4
p62kGNhI3hxnuDvHipA6SFEnMywViokdb1e34qms9yhxoQPY/lqYcf9KSGLrMHRnVfCcmy4422Um
cFn7w4aInYokeRkyyqxKlNPOueRcY8y314o1NQqG5ysTkhIDlyAPM0WIL2DayeKot6mVVDdsYH0X
oSTMeERWtvle4rl7MlSAhcZpqyyb2JgYMftWkOya1rYutp6VgsUV7mD9DKrPlkPsB9i5r0pZuKhT
kvZkekmdystbzMemujeLvu6HejxDfgKK4lkIzHTPjjOWVeLvSV1MTSR2f+tLXn345Hvf8N61ssdr
cKWd1HghlPVmAiOj2t0X05ABMbXiURjJ1lACk42hZlcSLuxR1rj/VmWg+Gwf85ZqyDcfzo6nlEDm
vfyVOLGEd6pohioRh9W06B0eleRP07R5LBNUjWMI7Yf9PdsX9pbwD+4c4flySudLwMuJcYhH6iYC
gEurv3BR/HGkqjmeHEvHQMNdFtwbtaW+T3OcKAUHnR4ynQHKBOA9JaMk8QaYsc0WoxijTfMzHkXA
p02a0neyDZZanL00GcPXl1AHqj5MA4mODOEcDp3tjYqwa9aoM/mCbHfIjat0EnQH0lZaSABS8pL4
ee7a8fk/pjGWC/Bnhn6nxoJBHAXMyuH5Orhv0y63S/pElAv6TNbGkT05jEujuzy7vei8Y6tkypK9
6shm+Jp7FyZ1SwPCCyu0YOL4v4eWl+INYR+9zsO9sG1i6OUWfRf+Gwl7NB0RGGlcsTa7eluvssCa
HMGcLSCbfYGTetLwgIajDCFyJ8B/bqjX6vT1hjo2+Jf6gE1lwucd5hW3rqh2Q0/8JwwWAJvChOVd
PPqHk5DX1OqriG74rY4Har80dgNv1I6DFbe5vNaMI27okU0C3Wp9t/b9reh8ueMTLckz8kNEnTQP
nWBivZ+shil3ghtaQbUb1UqECbcTQUDztQtzL0/SiNGsIKp3jXwiKNFSRy65PsLrkH/xx08cgbVZ
kCIXhLcsjq+gDjI27ZzdYXNQhl7mqg8hbmt0zmVzgYpCqzRFnY483GK4AesoCxaCHJygfStEqnn0
pJ2Jpa01MxUNZCgvjn2432KDxNikO8aHl9yD6S0DZmMd/OVr4HGyRCZpeZPhGe8NWNkHFfF+tVSg
TCbQB+XQ4wJ7bJHJHD+p9FqBb192lcn+OlKvzIR0PAxghLa/9HbEs2McXXFEDf6YuZz6Tem4Auqi
Yk2RX+WlbBKEFMgRWQe4oKEKQdxo0F1cPetnAb/2crFHnz3nSdBT9FQB0/POhgRgbCbVfURO4qZg
8wRfDp+94y2W8ZOGIHzIYtXaRmRWTnzhyQHE1SyvlGXuSt2IV8obGQ0WEER+lEp7GLRak3iX17yf
GlYUAft30h+/MNZC7JcDIwQRirgBMT/D3hHdUT9DPniuLOIrBlsks/RZW6NZ0lO5lKMfCUkirK2R
kSLaI0rSX0OSuLdAIO5tIeFqLv8tJZE4XSAB4Hy8tNDoBZOh2uvYEl2XfMSM2LBhpjQUKOZRbMUe
IDdiFogXrSnI8Ou8TCHnewz0mpZxTNsJZ162ckhpPz2kjCVoabTY8uun87xxA4WqUPH94kNw0G8/
eZwpGQ82N9lUYOHUjCBoVNJsYh2v9Z6gIyPh32LqhkZtwZOT6dG/QE0QrfNCQVfIp9F937zGH5XT
ff0lc/k3DRLzb6r5w9Y5P25FsREgzlnvn9VvhDGRZQRT9qaTe5zsCa1IHVMAdjtbfIA809cUiGuy
CCxrM9XYnVvPWvdta1i4oXxWPbB1hc/ghH2ffmMdhQSm2x/vK7lygZrTUtV+DHcO5PS5fjLdjdLM
EsQTRRHrJ+OrTR4vuySv/73TnBbOwv6CYNxKMhl9GufsqJ5UswkZPU2yBlK226b4OXqr+EvbwSUu
NWla8hEyGRUKZq1pXjO+qvH5XRaE17jmtXIgGkm8cFjAQ/grlyB2sKURxxE1bb3rA4Exh0CMRtDa
m70IMTCbV533jZYVVtgffddRh1kDufU+QuECjQYf32JBaQP18AUVoh6nAmRQ/pPM2rpNw2HnsmHJ
kPMuZ49WBMQOHTEEqE5Ajuw/cBQIPmthdb6FKfKM298DH84HXHgWUz3VafiSp9BV2x2jKp+gMLg9
YWjANj26vR2AvR+AKsyiGhdy4rj25+uLxfOJbJ6bJ+8ZjAaU11qwxH3pagGotsQyt1RrOivKdj0q
H07gnKF325UTZx7IxbWzwU3jVz1OxE8T6P9GmjFpLJP7xCC7r2J6aNt2H3LiUALTK7BLHxNbn8jv
XBVTa479iXZNqbGbORyc8IZut2wea24tnAdEk1bR20/V0DCa39odPS/Mk8Yb5Us6oewbTq5Lagig
m8d1ndX9k3Mb2c+OMNiloORZ2ybECefsXYzt4tEWFyPdeyaKmXfQpwar5mSJ3odlZt0asG525+Qr
pDPfEG/U2inemBS7OWZit0iHStQ8mRo9dFWbqtAqukfx8Tyxb3bqOHQZMpSAQ3uhrbTalsNxBnhP
KMPvk3Wy1TDUsxPvZgXbU5iE+EIVmAsy4b5scoklgqOX/Z7MrGVh/fd0FqlAwGmOupt8ohuIPpUF
DXUltX+0O3SXKdaMuVwwYm2DDqzObCwU+rtQ+OhbJ7t/jxACclE66L09s+JZzEQVLFqd81Vr8hDR
HbonSDZE5dLP0VWDAnvWsqlCILKx8SulzuwO1yiTIHO8GXOYiEU2XHyRsQBZvNHqvMn8+XCgQucO
iibwjE+mT/Wqf4xiGszliTYsBKBxUJ6UaFqczUrCjeFwh5wdAv7hHE1G0Uicc27bKADuoAX+for6
7+Cm+iJDRh/cxtH80MkcS/JkX5e3RxeMiTLkg0hBkUoypzu1+YsFQqE2rzPdf3hE3A6BQSeNzE5Q
Gi5ARTx8eGtYgRFue3IrYihwdKDjPINX97IxShWSdzgz1WSgiz68kygqaEG0GA2BPGDLG8fKqBIO
gtkofoyhIdwHN9EJQrtZYmiU4LetQx2C/e7KC8N3yWjDmIKsgXWrsgeQVuQryaaUXunFZrdN78cy
jtdTqAvL8DcHUT0Zi/emd0jANwo0q5OxFzXkjKQe4VMXZ++BR9ZMAPyaCx6qbglDYOztT3r4w2Xp
xufZd0LlvQCeJrZAVj9m1UufWTyxRWzIFTyDr+f32ZGGHj3hM6jbcepWjrjgUCAaEWXxMzA81Hyf
gL8aNmMp/JhtJfCsmxtMlUqZLRNzKWXVrTCAt4zM3F3PoG+Xshc6Uy3f84H085KoiQbFlcWPH613
71pvlbHcP7pWPJBnGD4BKuBkOdcURGdIfvWTejMXsXy7bn9xixMVuh4fH7dzZYSwmRhZFJ+muWxG
8qP4Jc+MxVu4VgvaGqju1Gb8GBmg7LkXzfgDPz79ZfMW2CJ1cAnyQsBZheKJFLNSr2p+xJg9fFqQ
IE0KOTipl9gF9WLN0++3xtRW0f5ApYnb0TTHguOXmig68Dbi4JCDiA3PC8rfNTsxEhNXNLFm/dyF
g8FCRCLDpJOr3YH8bwTWGQTOasPvRukgx73jkXbxzKRB/ZBtRBObaTZ14HR4uB+k11A9kZFNZQvl
osHRLkqBwWxCq3/F74Dvxm5pd07mhw4ijZJ+LIFVHU19k6KdjDr8PND5TKvVUZuOsC7/S3KWPfAf
ByqUjbAiwEp4etUGDopNK1RuHKB9+T0AOQ9vj+zsl5Pm+S+lnDMTniRCHXr3egcXVefAFNmX4pL9
pwkndYZycW6Bxp98nlBFCAl2ZdAgsoMPhKCm8ttSbN09hD2MRRp0y0crGMnp/hx8/9rVgdyzPsIv
HL3iX2g74a4p9kIotkCxExBB1EbLV6YgDE7TCsFjYJbEZCg2zeDli2w5JQyd31H2nySs5CoxFoRv
MFG3nF6aGmoLks6T9P6nRdL7Z16hWKobMjqQpPjtfH/dvU/8l7BJgJiRZdam4QX8ceNjBM4JCnPQ
J5iib82JGCKxprcNtUzAF5IFFkl6TyDhOVLaex35RsZwoL29IZpfZce73SLkgOakwZ8ezO/m8cZt
vBzN6HtfICSVIKylt196nK57WabV/jD/0y3FWlTzJXHynFJEkoEPr7n0TQUWgD1tUvo6P5Cvez7r
PkoKUfvHkEKoalRuKf6Js7ZN4KcqXDvzj1yJ/DnMMLQK+1QEzyAynrGGletjLZkXWV+tjkTR+czX
qiTguSFoo2VpUK80aAdstKM4uc4ojYmE9g7ulmPua63B/oQg8SJaGV8uQ1Shq6FjZjJnl7FOfDNg
As+zWe5H00xnq1BA3/vPVfjS/xEVeFVfDzdMistrqJl6w5hKnBK44XzUxe2gPHS5zX3F6Cli6rur
99qev3qkVCUuDzC4VCkev3i4EKVKdso5V+Gm0BQ1hTLHEJMnIDt/g1rQQwGiREILL9AHhAWLHCdm
CoP20LlG5oCciM40556ByKynaB6cqvZOaa7YDABnmhNG70FVIbabIay31sj0qTE83MLipI44RkM1
kK34FIi2EvXmxT71dghJEiC6VJcrVvltscXtB1CzkSu22gYkUl9XuqvjTBLAxfvYqk8ZOgtAX1WB
vB946/YejLLNiHbfWntgyRpbowqYi8jmAIfB37azLR8AiqZ/pVdoH0wsHs5hkKsct1TN7GVf9+9M
HAibyfYxFMoUylAFFu4ArWtcwDm6oU888Sp+Qs9YKITjfL7MpQ+gFiCH+68Wg0NNtPzgX9Tq3625
XzJARYkkIFDnyG92PP5DkHD3FCp7CH5wUnLT6UWVEmeQ/sd50sZ26iOfphFpxWvx7HOSPgZIetsX
oBYtZw1ZTTybuZs5etunZSlQveqZ8clOXyyF/g8djFuPVqxAlGu4e7IGGPWX97ziFoatlurjKGVb
Rsd5Et+Pqu7KdhfcVg3W0t7GAYrK490J4A3Lm5f1CrYaAl1q7c1o5ZFM5NuRG7ZBqb0wXKZNRJ3+
/E7pzfJDpdVuvHtcOJZIYwDklNnVdSCEHLt4u1jjAPqB7UbmE+LwmDE43YMhI+IVCTZVbghNPYCC
VlwlNctukVpHsA0tjALYxxr0ofiKMCwBgc5vJHwa3VfyDXV9mj6/BjZUStgS+rdLM5GAhWhwsXiU
8CIrwZZU14gWnkYHTBdvWTi2fLaJLbulqOyAoPNUi5X59B+r5JMjky+vbJ9iPx3i7CiA/J93PAIS
+Ok1wMBM9s/vWRrssj6HQj0Wt0UNfq08P8oqmInPfo+G2FQjsYdOcBUPLn3zokMj+//HnD1tyjyI
4zjLiDyprFebIe91o1fnzqMdL45sj0Yu8pAEWoOhrVHwFDx9Dq92kYTDWjFUMUYkuqidKfKhwoUz
7KoKkKbwfjJQ2aFMQILKc5kk4mTi+ZTl4nCq1mShfUQTeGoDlm8h08CRLZw98WZLnI6faHPumKZq
VULBPIybi0pzzZ8dYpMKW/VUm1SxVc++0TEGnRlwuuDSM1EN7X6JHWVn4Lcxeh3LxG2goFsKmkUg
tu/jv8SDb4duNzZmb7iTrG6ih/x1nmvocw24YVsvf8TeYs9G/W0Do4GV3vgxTYY4ip1z/8rZ57PN
/k/xQdphH7iecmA7wtWkGfOVA+BgXywRLlHw81S0iqGKUhC3XCnpgP/KbVk2YKB68yzP6djmG4Po
qsFLCBdrMGOjt0SiQz1qw49ubJGLdBQ2f/wqbAjGIIUeZ7h3ulFk0KMU5nXRUH7f5M3sGMbkmqNB
TCXjnrv4Fjg+OElqj2EnNcEjxJLfCVbc01TXltkmz1uvOh8IW8BI38lVuvZYU0QkratwakiKlgqm
KWJd87ulHX4i8Bx2QuC3fhAcyBpA57aMT9QIPUM+KrnfTxnEVQKORp3rDblrWv9z+aeTDRCoGyvg
Ze0YwVEsoA5/GjhfShJ9kxObNLpsu3nbFSXImhwavweBKKjAa14tFjCydPqYPOWjD76gpm9Oqj5n
jGN+BsruwoOeW7GPPrhKF3EN47B/jcD93trK58rGj6v8yhe+fR0NHt0oeKTqy3VVo4ffjG1NIiYQ
Aw26gf8s9SipAR4xCAVmKB6/0felhm9hBX6Gik7yQ5WYKIo7Iw9dHdYu3ovLGUZGe93FEtlTeHgH
DFCGieg2bqtHhbDBCnGIKrz7ZsHWrcw+bQdIpI6XIQ2g9/puLvnz70X+3uCBwnhCQs1WMDnOXOJ3
rsgKVyKCBhFeceKG4iAgS/ehBoLoRg2UnU4SKVMZUlEOS4+kTpuLoZ9yIAPm6zU7kkqZbOFOZp40
b2yHakg7JL+qLmRqpmzzRhLbIif//z/cDYhFf1U+1QDBmm1NLiojHNJ4VKHTnx3NrvEbJKvRAhkS
jaL9iyFBlg/PnIUeQuCCDHREJvyi8aFUhbUHoNdfR6fumSPuL6gUEDqOmPaUjP93gqSgHLZanF+2
03WdKAoL8cW0+7ayEDWNtevKcuNkKGIHH/F0Egsh11kHgu7ghjUcKVZor8AkcZZI89WfSGmdK7dx
NmOgDsVMNA367QKo5Rr3l5g2qKiijKsQ+qu2Enog1atlWjlzwk/zChykQlwFtx4CIManZP8ReE9q
EQKb7AL1juk0inhJC07H1duxE5WC8vO/VjWF+WQuHa1aCGIlXjc5RUZkcY2XgiPef7bmJ5nuuLx2
zLd12wfv5e0VcdF3M3hsFa4FfBGwNVFsXHltqnTO2KA09mPmg+Nh2agW2TfKJ2lXep6Y6VruC7FV
XalDrxV2c4UkyMVqXaxAOaTerLErwov473XBysAzAlixkeAvw3A5ToiYW07VsEUL36o6fp/4uEtP
nQf/CDk9RhfqA5ERE7oeyOcg4a0L80cOOJArBg/viOuEl1e33bryE5Z2bZYfmgI5KDsxfbqgzUiW
P1xQgWW4aFXR88NI/mUTLKbsN5vEK6gRrrxaAzKtZeRh7C/Oh+oX11wQg6Ezfg58KrHkdiqn0y7e
pzxGfv/DiA2oMhYOb848xP/G7MhGRuz76rg3EZhvEltB0NnbXV4maJ/f8ucf9wYbr5PxeS+UB0nB
Bl97LLDC1hzBD0Ngp68BKO7ZmZDEprsJTi4qXgoHvd6Q+Hryw1ytMtcqN9VtGpz0duMKSx0Q1Asr
hQsgDDYhDFCjFbT4SQeuk9LO3vi2sKZKHRNsPGPLsopfjELYMw1qc4ZxgmNoS9Iu+jUzuSf6YGGF
fyGhbPS8vjNGHVajyjdY3/0zKxaQq/4DFzAB5n9LPZ+mM/2KCvVdlqI+WbaEIgdabqvRMPTJY1jU
S11/gHmqC5y+r3Oyk8y/Q7haVRp/HBUy5pzfVw/k8as71VTep6G48PjIRvklN7lJKfTG92qab5H7
cRuhgkbnP9QjFgmPJ0MoYst0kb+SviWby3mB0QZ3LgCVSOqv27mwuLLBynkkWqi9gLt6lomVljIE
rZvr0sF6ByuQL6IyoXDkTBBQwlx3TfA1OkG/9j076m2R9Dem2wfVS2MFH8Jv8Af0qgrjQ3aW4gAD
DdLwElQu9fy/NrMKnW6euZmhP5OJyDatVgK9+sHPe1ObRG+VO/A10h/hcpM7odvBVgMQ3Tk5rQLp
0s+KfO09aa0XxtHFQ/4j5eKBmzpkKp66SU93kRORmDboTc1Ocm7zXrN0kP5Pc8G+XWQamvR3t150
zP3l0GakNNqxyixBXKVkuOWub+5sGqLp0zKZl8KhTD9vOi/eajb7kWtBpohWxV0NTHyui4e1ofIx
Z7gYAgsIOWwxNqjZDZbwQGXRAxWm74wd7H5Mo7M66B4gEBl3DUXdvQdlSD96+cga6//96dUI12iW
PuP80EaUAbFEYW2tiM4+Ttebv426h/ZnZoth/Yf9pVvQQV6q+qL2pVyE4nwCouYW5SI1Nn1O7fZf
6QiqsCy9eGBtvlcjaXCl5AsROAMPs027AWlZaX+05GGdOgEY+7Z5LISzAVeCGKbjqJ8cvkU92j97
ikO4wlTRsBnGKzva9lK6AthIZ46OvSC7FCCgufzZcrfNGRfDehRvZRcJUIf2IYHykY0RIRRbeswz
+Ee2d69Mjv5eL6WE9tSn6m0cQF6hh6xuLk4MxC4ye9f7S73MSEj+C3lBVw6cvngJqcra7VQi0Xti
tr0MRL3pG9dVQo62TrjqcGKyN5ueC1pDoQjhhnJeVjzcD+77hc/QcKLYwysR65OAEHtYvbmZbu24
xphIYhgFhkRV3ld9hVpJ7J1kcW1Xoak229uuTx8H0MjzvXFtuiWa4zWQ/lU/s0jWyshrI0ML8jqP
vTzUxeQV/O6/CYjvbtv5agVcMFpfXY4i1OAqp0vz5thM0reXOsyPVu2Y3GTdTYaYgCx+h7dnjmdJ
cOHGDuIoVepnf+Xn4ZtiKWvR8pDKJayC0Oo7LT0JhhBLNxN8HaZjAb0cEOwwIR9yD3KEE9CvpXiX
Eek0lpBESQdXz7gxWxko/ADwzD9zUFTHUBL/wREkfUeS8Z0cJ0JcMrPzIOh8912UNSs+fo/p3OPf
g/c0AUWClRraU12uv9fNGY9eQ96dGNi+Bl6g93NTdaJDYAFJIJZYVynlDoiJpuQsnkk/Eq0Mkbiz
otnCuXStdJxChox8rspbAp51GlLvgScVFfOaDJs+hmEEfSrPEYdJCoCITjh4IxSg5Hs2wFwMqFBt
B7bTH2G2jjz1acYmm+0pb31dz1x67g5MPw7smL75mkBlf60BEg656bbnacMIggVmp5nWhTftFvSN
pFA/MMllmaINTvbwnJw/WyLBIEDisVwaHmG25jy7mkUrGQQ7LANSz6KBkgGRZdz7UUXwDvBniJPj
EBqqQLXIXRYTGfqje3v1HZO1G4+6KEypxuAKngS//8ppiFsGcVcKiRyTlYOhRGGKwnnvlqlU915f
hJsCivK/lNguRoHb/g3dfsnyXfoeaxmowDflAexuMdfLIs2nR8Xucjbg+ynxFAkvz1bHCUA7XoZd
IvBqCuvAywpbO2cPaxEbt8GDfFiNIeQs926qEBkoqYoHzjYBdl/77ply1DOvDMe1gJVpQbKsZBub
TajOJaNNJlsDqgn9KCyepDoem+ElqGWLIYkJ3TRAiihERg3JxgrPXLNO9BtfYiSwMhuytSZ4SOlL
I1Fg4hIrkF9kZsgQFmLNSe9Zl5rZX1HY4Toyde2H8QgjxwSxKkE4eyl7ncX5QKXCmVl5uCDSFlkA
yTNCPFYVWde2fMlPcRsqHBxooy74Yh7/OKaimXRkcw/8XdDdPE6kcvgoX/1EJ7qSgxUIVYRmH07s
ka4pxB+4iSac46WC1eMAUuDX3vuFMH2BDLoNMdIexmw+yIdhvWYQnmMP7YdIzVPyT4kcIt4FtEe9
0lZP3T5WVZWqGV/TUPKozfpeS5uTgBkr8NWbKnehYOvVN17qZLjGzUp2hiX7JC4n3MAKo/KSGln4
NTpSzy/HUZ4qIxXEwGqUoHItCDq/7z+yVeV/USDaaMC3+/nphZgPT958rjWFKzShgpXqPOUtv3rL
iscxwkXrzt90hNkUdRukuOC3gC483b10e5X52kb253thzSB6lH7UZXgA9T9ZliZ1SAEwlul4yJRI
3pjGMcT9vl8saAJ141yM1wXb+jMAPKTkrxGedhrN5iIKeY5DpzdhX1gu51Hvmf7eUg6ZzDWDMNXM
+BDppNi6lPLqKaqylbVQs1HepslxgplIiCagVA6SKvDfqQixoL9qlU50fi6MZz9xkF4IKWucG/+Y
4BxH+T4okuaG35D5nP37S0eQO+LSXvtyKyWxL4XDoDgqDKlw0gC4Gb3eG968/i38RJsgwWMWjjSj
hGbF9wcdOGS5N30nSEWcTYtCLPVrrlFTSIKCCMLk0qk4wlbyrzsH+I/T4gQ2Aumdx/o1/spEgqCM
m4IxtBbnIwzPXUAJlvhEAj2m96dY3Qr95OWYLPn2D/Uz5faB6v/b2i9Tlp1FOL6c5E9JJm12lJsc
tZN+Ga1CdpH0K4HeXz8vUYe7tlYKtNczzw2L6K5MuduILw/sOiOadZ1XPU3CiRlxvLBlqRTech/Y
0MW+yZiys5skZShdsHvXWg4lKGJKVH/rh/DS1OCLFiMT7KocydGutqPj+TrDMPdv/YOs3ketjDH0
LPCYvGsy6VWmjubyA/ejUyECMKbS8AFR2RsdU+2sJO9wypaj3/a7g3zlR33Rijb3p5gETiwzdT2w
g3OllM9LHLJIr3rDl0YHHZXDDx+PbQ+AHcNfybK8wjm59dPDUOXgzHXNp/XlGpGQVJJM23GgCT9k
Jn4FEAO3pzUV5qVSlzwFb9aoUhZlz19QUx1/j/mjA1B3ppkkhGY+ppIb7fTUNry+DDv4utc3bTYf
m+XGmx6Ao0K2eaz+p5ihwpd/gr6+tEocUlb1hpbeiIA7alOciQAqOzf3UPlNyn7Ug6ItZMUCkBcA
caBnUlfY8jw4tYmcNDAFKdXSGoQ8mzPmqoJ2Ne2wBxanmrqq2ym0MAqAT9CGdbxiERk+RW6RiB67
CSxHJpP76vdwM0P9++rxqtjcftM/OsYeKXiRWNMuBjwSZtBbKWTqCvW9YsCeUfoIIZ3iFHtY+V65
/3Gj2fyDAgXj9fE3gVlxk3Y2HdE0JepncMsMhVzfYLm3Zt8fgf+93Weu5h9l3jCGM4KMU31lUKq6
BfYzoNitiGH50A5/5I5Bun91aE2qnSwUwSDSdfb5jKDTKDBCnidi/Yf91xqACKeMLphe/EdaKp6C
kxdnih1G2SB7mEUvzh1oeVjPbQeIkVsESgALZ2YRqytIZx885rNUUu6xfNnC/lIYUu3I9t0sLKBy
cM5f/ExEtqRLuEDj9nKr5kGEiMGwzt+cIE02vrM6Z/D8blCdFKuFLbdDR01uw81x2wnWT+6kPl6F
ib72N/aRybqsN1oiWWxNRig7Iis5TXdMs4+a19mOYRjldtPnyvhQHVPPxWZAajaf5yc+REsX3GX/
htTRxD+FgKRyOaaIatd0ZMwgBtYWHwOy03kwfrfkUi3B5l3UM1TY3xuM0ZCTcQ0O9thQF0syveZn
OD2raO7vR0H2cmbucRgeWjl6H3OwBhkDTgK/CYgr9qqClMdcEnmGiYFBlSvbO+ZEzYt7mw1hkh5o
ztQG8U3+XXSXkjvRjxLh81ERXslekDlprwxYJAk3Jhdlhzyo3kzpv/S6bBfxOU3rbTCEBqdWJVe2
WMN2Lpn+txf4doGw8cvgbrH9Qi1IQfUO7I9Zx2852mnJHZHsRnG+U2HDyTQ3HlJSxAIs0hslvQLt
pyp1uSJRXSCX7UpIGwUu1/RzQy8TgsnP0LrfHtBTv/SIJ2zhiFekKSfA/mU6sTXpKVMpDj1kzPmH
pI97NwFUfl+I00nkxwm0CoAPgRcV1PWYwZjkEI2/S+rjjdinhaYn33/psRSEg0AFD2xFNWbHuuhX
88aMcQiS+bbk5YGXy6tgDTw1F9y9k5voIUh9JCdoG9LzuCVPQfU1e3gMp17Y7lnxxqVaqFp22dRS
ybhYso8yoWvOPqJj+ey7UgHfot840+IhX6mjJXVhldBGIq6Wwlr0VWqWIKc4oWB79nfdG5Ilt1fw
2A82/FjvX3QbJmS27iptBswPExtM5VOK0aqal4bBLtubnV2+nU+aIiiSPXybDzzPRq+DVYVKD2ZL
WLE3IOlSRGf7sOZfQXQS2zIobAAtnqqtYjIU0prrB3yq7pNOMdYentgmhabrLT8PSyAw9iamwvJ8
yYHrThVZnNsrS2h5KpuKpsvR45PE+SXh2Kb4KqXvjFi3A+UdtNLfOFAPpyTEe7GnySt3s1Kbokzn
IMMgp5az2IuFb+mPAdVHN3UsOW6seRNeSsyFy4ef2MiXLFBF97maxzptnVzw3dCzSwvTEPOYizq2
y88rmFPIcNczf6H+Q99PvvPNarU1XqqZhqRfTlsVSOVuHA+tzm0eRJO62jOG07jHUp3+4VuQfxbZ
k/XQDIrqxXnYmpjqbF8KB/bKetrJcE++kLfybLTnVJslzPUYC/NYzmlHHDpIi1KJeJlYz/mn3Ynr
xvsY0ReUQnVtTSVtDcPXOQ5weygCz33Qg+W7PzbloTB+ook1TldcMiZCNG88DyEnUpUGP+K/1yrq
DuELmfp6sUFS3mxMgTuOObEgaqyFmMdkMt4mzPI7ctXkUc7vst/vlu8HFGDsLkrd6HFJHWK7KYpL
vz1gnenJfHjzzUyICcoIPC4lWLkpxGemhBDc9TtIYcM9fwS43wu5ge6O8o/ccdJOkhzQzeoEjiZr
lyEr8ATeeCIIq44Vz4WVhFD0DZtgTd2/Cnlwp3Jw2DQyCDOLz/kCT5l3JPPbV10FcKg8LWYud2le
oU69Srd/TpSddNCGXxrtBQQNBmFiGXykiUEP3vemuQ5+eg+Vwxd09K0fpCCV6aFza1phQW7xQpOC
os7D4AMtPomdrQDvaSYtaVypbNx0bU2phXkr2ubDxlxvfrbBOg2THD5SJHMel43D7u7fyCvkz4r9
b0EewupO4vmjXuP9KvSTkZnBwY3M2O6gyvfC7ko7cYaZCKvKsePVhnNPzgmHAr3t7TREezmx+yBM
1XFpIhkxKI6Ohgn+3f6yvfAI9NaoT5DSvtcbzdVSJw5CGVl3eFOFbl8OSU454SdBfFwjbH7/ZgCX
inUlSalhecU3neLX5/106Wwtav4VwZKF/QZ6SbWS7UwaTbTDiiFuGQevK0cO0/AbL/cNG8As7Ud9
DXil+nb/yWoSxpudlQxgg+GtNuyKsoaSlMqT1Y6IVsc6EAUMBIdDUN0GCxZgeNJ5SUMD6mM6Ivi+
hDSgydf/lyWDkXTztQ2kyO275mK+kQY/tiJYHsy0QH8EQ12qKtq6Vf+Hjpq0bBhDXUQAS5y4UQfe
sKHz5f1iW0b/6xM36QJ5izsqAO2XZXYdGjm4F4Vb7mFjrVO2ED5gEBH/Hkx2v1RlOiXttOFmG/VE
5YMaPJNr71tLjXQHZwjWbf4pxBSAI3/3smHh6LXmzfjmbK9L4zGR8KuMqGev/jQsu5C7qwyx7ZHm
aUEJenLN6ltvupa+q3MhWxTPsGz3uxckZethv7o+vB7fwQEZ//DWnM8tVmIytUIwNMgrmL/K1FDJ
RNdOBJ4Rasxb9DSg4Tc/M9TBuxnOwvYEVtWfFNT4KPhmwZr9N2f6BLhmJSHMPn5EfdGeaQGtsOZk
/XVSd+A2e6IgZBWBhcL27wgU86IDV3Uvb6+cvUH7p1WMCC2R2hieNPy0KQQb1A16vqGRmXYfScIC
EZZ1oIGnlkuQUfk0g61ual2Hx1vQMMkQRYxRu6Psv1NGDnVWqn0CKmj06X2UaojJOi2XvFa1hObS
xT+eJK+BBPuxQx8iJEDXK+k2i1hV3V2wDiKHv8toFJUWgR9QKiBt5Z5xB8BJxl5PM6q7Wvii35Ww
+fPSi/ina38uEPAeLPoqRsMF56RLIuvd7fnqX8Ir+01yC0RqnIVSkpaIn0E8RwZ8cIo5JLjMRIoB
VhRHqJncfuFJSPds8DU7ahhBK3sG4Qz8BJaNhGY0EauNO91CeQq62DDXCRLQOw9zCvsTSZfG8T6V
Qofuz2HCC1O5at8s+5U5bZtp7nRHw+3obA9+dxQfqaveo2WiFqhfasno1//ygFkB+6IiP7XqAezZ
iqKPG6BY9JLCO2Wt5Ugv6bjY3Ar1ST98FO02aTec0JN7FZZuCQQYrhx6s9s1kgSeaM4kajFiqOgQ
jSAbbBwf6/RzCq0/lavRWG+Q327n1HvccIOAfw1w7ilPTCw8233kCiJT5J3ewLv6QKj+gUfhSZa7
Q5peV2qZWKbfnpU1uFNYM7OWOtgY0WwH9v/MO3xv8ASbIp6PfCK2hRTe6wRnzrM7Z/DiosB8xNTq
S+Dzw7LqJlGhd4ZFMDxsau4paCVPVQ2iHCpAgWbbPyPvesoOHVmcVuRCjvU5hXGs1Bfkw6npzYiw
lv5faUejIWAZI3q2apy25pUDh2CVhhFjeg9+TtwJwCj6MaMc5ALRO9GEX8W813FqGueplvU3ZhsG
yZmVOIc7C+V4T/kM3DoSX7fD8SgMhN/3h89dYvRwY5d3tTAxbOuHEpimLCu2SIbgGrcNyM9v/spA
nDJNiL3wcGcMBCyp8MBnZFOLgyLELlhF7ijS4M6xDkYk5LlzMyIS06aXVh9iHFL+q1ZtuKHZwwTN
KtZP5LQl3mh9vg98ThEZ2Kv2WDAWD7jWj77qQpneCw9dSl7EFEXwS4vqyxpXXCQBUbLzv5JkmiLR
PdPQRIge7PrAFb4YABHvxIyscfmHq1o4rSNpycvNBgWpVj0rHOjKNeqVXePGOuHXno8w73iaxt8Q
PCCg3cEbMaropLhP0neZ9XuOj6wyVLQKhHLNGEXc1rpXMOTc2Ytc2gQ+dSuyfTZ7DM85Sy+DQH4g
xYXFekJeHWs9dnk4At9Me2vLb8cQuil6Hg01symyQyJ/a6SQCdbQ7+q4p/zydqQm1K1ni6qYNBg9
iS2u+pSkcScJDnolvBPTV5vWSTUpuQ1EXIo7W6JiBGniYGc8vev3Kjv/nsrbzcLL0arWzNHCqtLy
IyYjD/85/iI3v6r02vvG3Ymz+6v099BMlYYoVKcKkcyHBr1mKEa1KzREyjj+06WMyUEhA5y5hkvB
Y1jG3i4JCvoLSbCjqXOGLnblZ1BdmcNZLV+kVaCJnzK+ZTe3IBKvm7PBNl8n6BzZc0DyDc7hPrO3
OyJaOpiFapYXFvxWlUhWIsGYBf5d1UnDI3f8+xE0Gcy1Audt1GD2XnjqUGewuZGSEzn+hN0doAO0
BXgwDiaRm2YS2Z4FqxtvXb73KzJ4X5sLKPAFf1WDMKdpUNmv2WL+ytwmaNBF0akmS9zdIZqpziKu
1xjC2/EHhLmGnyZDqvttPjaCtvv31YMdRQNcxfvNOFz2eK6NhKFbcOgCMGCcioJPn2US7n2kGZ60
ZWWBSKscantRxiTRdFc89MztlC7w6KIOcGRm5ZsPjMqZB6oMlFUn709NN/Z84jKZMw/ZHJ1CwC8H
LDU1txbAiqwGOdnkkNIMj6Vjpn5azEzLDDKs2y3P2XwedDfb9JCgNfYYgVTMu4Zh0Azjd/QRViBN
PmDcLuA9v7y/wkNy1rvn3kksibkl2tTzGD7fplSq9/6rPN7FHimHTaoIiuEB/Ov/b7DttSlFlNkQ
7DaTsT6zd+6LmTn9XHNvjKzZv9SfjMBDufQxSx8Urgn8mO9CytSgQr9X1mKLyp1zFaHflIwy/5R+
5o96TXQZvLj2+J92waUoJeMay6guxD6UuD5jbIRpC407YMa3uv7As0ZvsmcuurSW4pk340oFv1NT
ZMAApYrBQeR9bpjG6/dGs3Y8iMsxCn3+QLB0iHjbvYV7Ea5I8Bj8D5YpqPzlc8fQMi1fB31GUfsJ
A1Vj1gfDouJ6O8iBobWWb8wflufLeK5cw+o9B7IJzfg6zSN6lYuMOpa7EPiDxtkSD9mB2iNXuuTS
xE83qJviB7+m5oQkwoYg2V1GYeQV7fKtziND/uYLLIkD+I8DZ8ZFBECwl21qvOs9mank/CC+KCFR
CqOQTPP3y5p+9VrBwvu7y62U7+2xrCVbxX2VANv/lK0wPglM1/g8KXG+Lv+nzBvcPjvVWKO93KeM
a8Aj/D1BHwdKSrI1CYuIrbFX9KsjgFEMu3BVn5BxBQRBuF8271nOHfXNFwz8e1VwqNOSMQSbafqL
lqOLLta3Wumprka4I8VwJkothOjOtFQpaiavEL+TKOydvIX1weo/7xq8dX7joqrKccJK5Y3QVZ64
3VElVFB3VQvjkXqQoujzzpvLBMA2Decum1p73f9kcyfkfovWgur8L92LF7Xfa21BBJVFogH+PIjd
UNpWF8CYyfAUs30gfJP+Wozx/ygaLW08TzUma8+S5jhjg0HfscbVItS/Pmw/yb/TaoDA+29otomU
eKMkYeSp1cuPmgiqnUOflrhvk7oCO+Gd5el7BzzfeGHx1sY/utTyah+CPQHpwX1uf3ewaMiXa+/W
986FeWlLrn7HPwNWz/CVXqAa6OnotV/UGLIu7c3HBjdne2fq8VUIGoiAaMtRs9dvWwB9mwl6BU7z
HKu0D7zAnWO+CdX44Zl3d0fVhsfz/dRtIqPDYzwu7mv7rb2CJrpvICjA4RTvuKad19kVCO+fPASM
md4ZL5fWfEcVEeqYu9+MtAuCNyfKl/4b2iRqFLbpoj3Ysdhvz50qZYUZxVwJa4DmhUzZ7ChEjeKP
hywQF2kQlEZgVHeXiH0S+JIqzMeX8OyCfnwCWir0A/kfe3sgzlEreXicQIW/zKcjmcuEAL2WK1OD
bzkuvvqzRAmXLymGsbVHXCKvdNQGSQvrq6spe57nDgaTOaXzaY5nbB4y/pmpYraylNSHadvSy8Ob
J5wuIBlUBUvJqaWywlgRIuK43PwgO9bT3R9kQIc7SYyvWxgjiQan28bSX75UiQY/LePSlGQn8du0
3EoIOMO7OEFgWvjScIvEiT68DWA5Jw5BdyaH1KD2dHvAsZcqWzpTe3s5JSejYb1CAczM2DVS0XOt
Rp02hpGd451IfjfE3y/R8L1x1C59Fcz58PDqUdlNQSzJ3OC3b7PahmCCH7oUkRMKUvto/JJocIpC
+YpnzA3Ba9RKD4H5b0Wy1mEoAJ6mSvIzjLEN4Yf1Kp5rK8n4UX+Fjo7xYu48v0KAHW8Vt0j1x7Jo
b5U8qwyXOpNhwq3UmOm8vRPasMHOQDKDFrmCOjFbRU41REvnm5jAgQPpn9MNwucR8hhFgwXG5egD
tcle9VQMrzUkecm2+pDeRO6IWPB+qWE8gmJKaf1h1WuLI/zwLXJtruEl6qC7B6csD7vRx1ZFMOew
gshrlx1H+LLxCM4aDMapDwdcka7PgWfuKdkDXD/DLsc9UR6cMU5MljoG/MmDVvl2I8Cvd8wXiuml
su9icTcOd9NdV5ucOFElzIZmDOMcTzn65udo5+AQk//L2LRUlVZK9W30v1pIClVNaqfVptLYOdpB
+Cqz/8oK+LNEzKDsx6/D3thuozClmPw62MrGyRmETDYVf1T2n/TjNjUX938OM5h4h8Qf4eRyROI3
3FjV75Ge75VH6zflggUep5vqoeB3ZcY5GjQlyb+SIQ/bMM9KaYM3YdeO3w69E9U7MvwwfP+7lrBV
cY+RuP/kQfYCwXoXaEDxsJD2PRA7Wnuc8ecJwQU4uGrCbkcyr7DGCaMSvnUQ58ohW0z0w2WdL3dI
sPHr3B8KzNh3f5K0ecXhrXDOiw4D7yQwot2oKMCntHJe/OZsjy/3rlwX5RwXKTBVh2tgkfYU65Wv
xVpr3MkVhfD0hk8odOI8iR18zr6wEOwxdtUtjJmUihRQB+rPfC3YPaOBO1cLlc/WnFiPiYEji1iM
iD5hKV/a+a/gIRQuu2bhJIk37x4BCB9MuCAXSZUib0yeM6VQSqzAC+p+deDFJ0x6EsYgsA+8AFaF
IjoPftMq0m2ohJRLH3qiAmijT3zjsKJgAhjWVsfAzuLvu4uh7L9fDZ0bRRzNvtzIlt91wABRGqdp
eea9quZphm2RF7i5f4f3C+sA1RFCAMkbtqqEsZS5D5rtJH4tLU/rxPhrMLZWQKTj9H54DbIfe4NA
DbcowWYtedxmrv29Xtf8/V/MB6Ga2tV83V82q7xfp4HCY95ONZijLUJBB7slboBBgliI9mb5uPLf
8/RJcTZ0Vs9h4w+00rpIABJwEDkKTXIigMbPCj9DKfzrwI2jY2AjpHJFNRwciadzBuBDDEKKMG6G
szGM2VTb2R6xVUTl+/3UKbQb1ewXGFhxBRsJXCFeLTSylpTUAQLN4oagy2hDMN/eSvXVLXSfVl3X
i7PGPfp+9ZkI5cYLqdZhXtKpHhx90L3x+PENv1hay8W0ais6iuohGsTscBeEAX42fu6rdhsALKAZ
er/mkJz0yDAaWay3nuT1J4YlYL5hK/9+OSVXlcGlWsd9w8jn481y38MX0+GmtKBEUqrUXjyHA0pl
WFJvEKZYP7VsA9hTHCtfKkDKqg2Ffz+f6CLcArMbMI0wEeWh5t1sed9BINAbg5kILr0xyDpeWeia
KJsGUacrfQF/U3o5wi7DLmHx97J649RX9a6QR0kcS6Xsz8Kwl9yXACcJgxAfcS0C21RPU44eDaip
58oiy/4trsTiAK+IIvlQ2Ttrd7ruysiCEd5GxxGlluIl1rCIh4ZsAL65+bv2boVVojbtm1udJX3t
/cDV2IRbJ4/oL8pqSY7x7ksQzL5L5J7TDwRPtMsNxydrPh26wJwxK9RxAtNe4DK+yPPhGlGpST3U
jIrPM2rwAA7+in5fFAdCzvGB6EHc7irtZg6e53uLZJKK05lB2UNErQ91lpoJON8L83o6as8PfGCS
Odvxroj3YXAC8OH2JBod4T5IIHHfrPeI+1JQrFau0iClPhfXtFr8ZNPd7r/6IWTHfikfznGTRskH
34Hxy61R6I422cWq3rfUQtzVJ6MYTzAoP2FANgg6n/aSb7068USBIblv5RoNvM+5WRkmSVVjM7UJ
GPIXuoR3qPQhsHYVoFgU5g3lI+NVic9KNwqEWTpnSA8DG1T5qtTaKO5vJ4ZYN9/8KmgK+Vewg6T/
pHU6lI4Hw7nOAUFWNno5dUuvX+NeysBZCpZSRkyo3bFZluRr4B6prsS1aZAs6wZYfIvd8pG90+/E
wz38pI35rD3XfsLdHx1chA7Vizge70/SLL3DTjljFGkq0vyGfl5Q8J08HzNwGn/P/s8BAFOWmO9V
v7p/7sczzriVx587YLcoonytNwoVG39uOXqUZmiUIE/dqiWMtxIx6kFh6QBXEuCQDskqn4Zjr3g/
Cc3/rhzUX0gJqHdrc8bQ1THB+PrTlJkfH/32fSXpIo5IR5btfFUPmpQA14hYEDbR+7yocGVzYRMU
7S35FSfVqFR5lMGk4aYoYEAzsr6rqGuDkkSeQ8VULlkPj1Y4sNFhLI9M2UqAj5RaEGdQbWGLGF4+
kvTkqvf+DoRsiAT2HEsl4ubq81sE/F8+/Hfnn9pmydJxJgzbmupn3iDc++IrbQQ6HWHSwBQww+QG
v75utYqCMasUjthT2TS3LQb33CUrkKsss06+o7DM9jw4vDG7PKBcPq0HF/uCxSB/1m8Tn9oeM/vo
2XkRKiNC83/TZ8CGyMEq46ISuIGGBOeYHxCZq9bKJYC7ypX4mDzRd5/lSgPSrkZxhCRkMgxJB6/0
b+RGEJEDDkDsZTLBp8G0NY2HyJL5QTtUkLwb9EhM1giPZSzDb3/oorkF1g503uzyKLCemdV8ruWC
7lWFKAZL3k5SA5q6bSVzPczzKRX7fTg2+Y0WWlQmNk1a2JtC2uRbLtRwb1Di0xfbueJ62Vl7LiYs
p96IfEEZMiIbWwr0fp87SVKkOwmdQ7idV/58OE2b6UiVaYYNFvbTiEibBCccwKVpIehbSXGMpaHg
Hs4hb7OV76qxtK33mUEAGTkrXTKGaVnvhrnqINYxP5a69pu6+xCD3KUB6nTrHBacDNW+LAGC27/x
XXdJe2+6u9E+6IRkDQR+oOaEBA628I9yte5ngJf7yFeTY52ZHrsf1wyqt6UDmOWQGwlYug5IRV/L
PcFslqo3VkPHvUdh6s/zu5PjZwXrDhLnSHoZjDevpV7AmdG1lX/xnLEV3415pE0FDs9MxCCETW8V
4A9IsP5k9gg4iwFg9e7ZqDqh5BuZ7anXPa65aF6xOgUiXSw7QfQ2j2vyb6n3ECDMaCRvKHfu3fZT
DTafFel3rZQH+BV7WYG806TvH12NN112oJZ3NT7FT5mATUwGuPXasuFq71VPCbPMTEzLFKQ+42TW
E+d4oVRqpTO6eGcSBbVW8MhK3qj7b/6yCyVl3z6Ccs14VCE7l3og6RMExgdiRlhO/eZba7toeIHA
JMEVp4snyGhFl/JUyIM4buacbQfF9ZrES/m+bWZCpKBkzjmc0rFaiyMUnfoOctVK6cC2LBHrvQ9G
DRjD72LPoJWkpmp4sdC8ZJwF6O84iysWIfjSb8SHQLUA/P/OBOmzeG8aRaAqrkXCoiahbIV+cMHv
sc8+qE/SOLG9BThF3ylAn0JRiSjZPUqjxuS29DtCwYvuQCv3fkRRz2JbWuZwQjm649fKB80CytJD
HCRTA8voAE4UWwOUqGX18dz6SjlHFSSE0eSUAFluD0fxZmGrlg31H+XGHf0ptMaVAr4ZWh4xayQS
8T0HGE9faxMlFlvBKUi7JWHl/lfzUQrBeCDwd5qRp1Qv0z9YoYvpIneE/xHedrpz0tATavyOk0NA
I8FOKZRdRdPIdwVTXW4NQRrGX5dsMSPSU13b3j40MzA4Ca9rng3WpE75LxvDTFMiIYx66WuyPG8x
y1Dq8OrSvkuCvcShAqjXYjjzowHCN7ObqC7eB7iq0gaXvvydqB4KwWBeewZ5E0X3q6q/Wgdca+kr
fa/wjWLJi+vaVMm6jN/TQs+NXBX2ytCrYAhqxGZYk6Vhtf5KxVPBxYykv2/rU2r8bqm3qKVfL6yG
zIanHO7kjXR9L++P8q8W0KBe6uysbwzqtx5irWUEcoPobYIxsHZbn0oETFrGTnLIFXSU3BxuaeQs
mopzb+M3h7XligLc2vLd30nrEo3+0czjt0QfOBDIZcyChlwaURm0bCadhi5YRQfGAJ9i4/82xFkb
TzCYUDKYScE/8uFQf9Y42W2Wlo45ghIGaQMWkk54tB146/qJvXnJg3xYOLjYB/haaE2DH/737c+f
2oIq/vwt1jpBMR1rcn477LNKGIHvNEPhI30AuqeVcF2F7HggtaFoED2ihuzYofQIWarbdAbgnk83
Bwfde2dVRBdqp8ABU07WoFlVtGj/yyTdSg01R3RpTx6QjCpnx4wmx/o9DWWDbBZhaCmiiC9s0G6B
qTOZ6Ip4kgswsNgHPAYijFdRwEYlJcbiHRCs7oGer8eGz6IrCbgB726iZeEkU4k3y1RpTImikFi7
m/kENBLaPFMCCCZL8/7dm4yn5Ogc6Fra4ktb6kb9G5yNijCb/A8kx+x3QU0sD6sknDaC4HBhR5GB
GyijtYb2zCTvnhqGzuRE/T7HMT3uOdUkSZB5FCgZSY90672taHx1MNnGpAXv6sikvh9LS7BrIykO
/rkldmwCYkZ0f+MlU7m0GRSA+rijAy06E+a0XIdFYNJ14xaZ2iaM1QwQmSZRXZw3C6lAQh8o5dXW
YSHU35R5VQgo98hwCp0LD5V74g0dozt76pTOEtgL8R78/dfAMt++memYOsY7QmjIxG3Ao6/RhDYv
eZLCXVsNkiPfz2Yrytx0m7kzLfyYJMb6vKRTaYZIZCH4yIhIgOioF2y1SqFINg7RB0E+opstv+/V
CY5cvajMlQ23nkTC2wukBcxSuN0IRuHNMTYWxU9jDA6ektaqC4fGNJ0Sty3cvj7KhXcW67LFnY6V
xaZwqMdQnvbEtqwi/Esk7ZZpNUVlnw0mEZj95M0tvpRUYFNP0VNnB96nUAjzKTUlHE+H6C1AYtx0
I4UMoTqr8+KFEkOo9fmEGlwWA+SVkiP1AiAq6+TpnwRimU2KXn43bPiUF1UWVXuP8igbNeOo3bNs
g9lgPlbGZNuMhSmJrRkWFqfT36nhLaIXmARYkNQeC8/hh5XIfUFQeKjCbmkYJVNHcBD0v1/9fJpL
nrTpkBueE2rQMAwY7e8zYGU+hevO50bz6pMWRPqNF2TrHKEpEwtwL10NKQEORt3cwq3e8zsiOcLh
yNqZcbGYcEZVgwsDWdIZaz6sQtqrSPJ2QRo05Upk6J8e4YmNZDy8mjitZBUvkDWQaSEFMFjRmk+g
va2lT6i/EPyS0MbZkbuJdQKLITIeLgsUKveLeYNsWKHfaEu9Qp0pIvADBcq+kpWz5nMfpcD+rrxQ
/hnUiAlAlDvbrtoF06VUdYulCFgkn0f4MFGrKUE2hLqA3w36ARBSXYBIrnjpuKVdQ0yqZVeVsI4P
huGE9eYoYejGeTiIUTru7Cj96eieGe0txjqnUB3P4hzpCS0+icKsoiLKlJWFT3KByPYAjn7BU5pE
PhnqPXLmgQMSIcoQwsug8Gbe2qBaTT8pPzgj8KuO897PGPJiZrmKLztmzyrL3biW8KN9J1Z4lQjt
fPacwyphMTcpXGV5S445Q/N2SUWXJcYsRih0+dJbP8e2n5TD5yNxlawpaetHevHlFrX/2Onu3u5/
eHTa3DbA1jwGXGaKhGnbonBkKU5J6GsAKQBj/iShQvHHBMGyaY+a3AQSlA3oY9c7XQp4Ky6EHGUd
ji3OjYoA23Uvt+d+kYfPztSN12HXvAYUwMYwLLJUCfEdYFLaAZwUx1JUAMYZt+fLS6Nll51wAIcg
j3zxSdeTKC3WsR5S1fpD4nDKgF0047dc/icG7IB/qMRe3atb6vZ5q0hHsCl6lvYnA8Q421kZZCHN
IeqJQxPrDNOid/ygY2AcnJ4Gl1fQVK7kygMJsKZ/uWxroFY6YCJmM1MRBL2v2o6A3D5caDDheRr4
CErxYTZRdNC8lJ6Y7JFjLdhkyxfYsi92SoCxZ4m1Kxoe50aF2068e6IrvnCmkQsakymLYOtkPikb
j+Ec1p7aBeDFQ0Cs4fgEmrObxTC0WdSuyFPMi9fVLvZiLYujzf9ZwLublgr8cRbtOR6wrYPrecRC
0EshN54WX8tbC3m+dlwPYG/GKiugYMeeV+yEGYWyfufBe28VQswfjsPZ1ZgXW6GrNJDC8kViD0Pc
WVazUcyd31vENb1gw9rxLqlporc15HUtdXqXmz+s/g01DA8lWw84JoKJXEMNfeqppja0+AU4Yctf
C6ZAk2gBnGR9k7XCp0QlO828xLFfYPinmzjGd9kFQnOKUzgp2AsaiK9v2u0OQhmgUbzmJOq/Exao
7jb2e4wF8thMeSWFEo4DCDX1mPKyJgv9a3aGJ9gtNrOYN+nQCZDC2zqwtgegKh0g6rUuqk1wkUwZ
iJz9Tu+PP7YuGyANZ9EuG18LhNqDusAljl6NTZQATzC5A1Fv4aUHkc2prwS2lvwc8Qn24haX5Wat
DWjf/po6k2Wsyb5z0kV96aDwsTrUnf63NhYYLygdZs/DK3jAcMR3e3PfZhOobUsEsuchSJb+GF/8
fQJpMpxYDeu6ApK2X0Rwbxbp+wrbNTFDpGz0SNwISWq9rpsA2N3bIxHJ4fdwcD1Bjhft4VR06U4u
fcyUwIl3B8nNp7hLixUZYyUkN12DOFtE1yzHOayD7HqHeyFHyokiyz4n1LL54X+PaovenSqwArI/
zKN62DKARjtc9FeZYAQanqV0gId2/65KPqvu+EhTR7H525iDx5rldQuTxwrnpB+Yz8QIQdxW5IMI
LHi7pG6ePxh3v2/nHl5OFmiD4tTKbBc81kBGf8edijgVT+7kx/lv/8ymS5h6lUKXVpO5y6Iw/Ga/
+WXjYMQUh/KCpJKsNRb7+mgYd96iCNvfO02ZmlyvAeJHKDO1ojRdcr5NfvqMrkTQjCP89nlrlc5+
PmvLzaAcw88cuGlawOEEgwCUmef29zecN2oowun8bJEVR56vTAtyArUNOSl7agRecdwdoJHZnYll
9qWVB5I1X9mwmxLESvAVUytxsx+U0igZKIp0pP1bpfLRCZ+kRL1RYDvp8+JB5gluf+YCOEnwSwPH
/FaiHS2hMWsBdt0p+Pr36FRhzEtS2B69KpfmjLIvEVBCPNYV1oV2fFtgyUAhpMVhV3aYg9IHVC5S
7gM56aBP7wxOsJuQg/1hSRP1tD0Abp1A0QV108m50nBX0JPpMNdn7x78tcmqJ3EXzOOeH1bJkoay
k4AtkBOxgIzlxkR17HQ2/fo+QjmLzUoKdr3XPmzopTjZc+g9TQ2FLwR1jHdqkgh+WUyCaif8Oxfk
92/KJSdBYDoteTxm9FzFviklYqlJfvhpzTWauBrirN63X4JiDIIJ5lEF3jVri7/AJCLCzr4Ih+OG
h8680y1p5ZNDDpsOV9E38OBcDAVRzGjGMMuSpFQ5n4CdQ1/ZmgQICaddsQsy7DmWKY/cg27aVtkA
taSuk5GlxZ2gcvFbcyHGBN55KDhQZfef6ggmFL/q3JUITtDBqh+TxqWRWvJAPUif1dKCFWWYhaFB
xokj8FI75S3sH3aimllYl8OYalErOdFZGvSWVTSlzuY5l7DKTP265XW8cfebWtvD9OFsddMI7A3D
6FfWYdnPAG42xp3k35qRE1ZS/tS84rK62+bOmC0MIwe6Ecz63UI9GEj9cIsItuv3/PVaw0LKKRGG
Xs+SIq61A8lNJ2Zs1mI7AqwdmSUDNeSiOaKmeRLNA/dLZzz7IRbnyt9KLWEr3HeexFMfBs+YZnTS
v46zJoEQ0HKAsTN+gcu2lrAHQGVGXX8DeQah1DNFWPU4BdV3uZh2KKVfp70fX6/gKclvvmlDJYMI
v0T5KFqKrk8kMt8hddBZIBSUq7GmkvZYuFwbCEYcbtVq+7ARHQsuDSsHXxcJmiELo0RW81YzBS68
ibZo8p6EyGMS6wNPec9/u1/xE/HtgTcUj7JORgKp/A5x+8fBISUYc1mCY8o2UKKRgHYSNV8G9/m2
0e39XMUErPv3D+PIlO2BVkJ5CfIwxHzu02DmeF9xfSDVYjslFldMj8fPCgQ2uq0NMmsVS94djF6o
eIlLpXU+LgpeBNr/gHbsT3iQKzL4E39vaPtWVKqImKjoxtz5izFeNJzQZmkU2WPsaiTexk5gHwkH
/2URcYS5izgTF7joK1qE/xlmKEa/RwkZn++pxwOnyDSr1o1VOIMFS2vgGgYNSeEtF2qMWqTuKUOu
fzHarYMSLkRdHjqCzinzDOw9mXyT7Ukrdvx8OzTnTXZSiKjCY8sEUzsPK6VAMMeS6zaEVenkXJTG
6z5y8fccTsXymxiuK89jAw0Oe0m8Pk/3dyGZqwVwaqCaVcadt3Ndg34HvhqozFRmcd7NLVdzyF/0
b9i8+NG338MBDmExTjSbtUoi1ype3/zkYxIGi5P7k4yOvYHaImV8ZkOmzVGrANPGaAinE4YUvFlT
zq7VyBK5sNq/AtymgwUJejh2T31GA03Ho9VLwo699vRywzDliB8eUag9rfSjSnLiA4RVo8CjWIyS
WkbegC4ymL5q1ico6bpUMBusaxTBmiQxaga5YkPgs2Qh6deucxOMr1MRj/Jg0Yct+Uo8ZSvUZLFb
cQ5XCRxx1TKr2xVptoEMlM6LEUu3SFNZ/zkHiGpaaIlML/ympUBW+7gOHwnwPbKs5yEBpaQii1B+
3Vbdg9QOHqtgAInmWQfo2RiYHuKyMSPdQ+ynyGaIbmq9p/QJKnIw/GI357PqFInnzMv21P6yTCQY
9B+bu4hvqoUZIo8tDCTGgPBn7eRpNzPPa9l+wuJRFJZekZwS5bQWKAmlSLLKHi+CMm39ZYur8szO
GDN0eEwvIJvTyGpnrcqiFQMsuHXBM1aI2xdLQWqzDPT4FGBhH+MqSS3G65f+2uUXwMQlS4u4Sm//
ZPMoBRbMpC1cYNKzvWgGKKqC2s6t23f3o+d2Jkp8ZQVLy+1hARSwbfzcEQ27vNWXydxDXQGkZ/Br
CWHK24j01Wdkj7ueefLNmBmGpA2I/pHWjQun2/9e5Gddd+jJYw72JbILuxBQ2iOKrmm1I30uYcrP
ME4iuCRbr6pm9g5UXV3x6awaL5avH9/R+YKGyUe9KBvXw0fV9g9/v/CR51x+/UvQBxou7CJsawPQ
SWM7JvXyr6QX11JhX3ZUXMK8ZCUGdiMxTX0DBNrKO8JIR2H/BcpqVE9Kxtrz5nhZWa3cI+RYOiKh
slTHSj8YN0eD7wGxn+d2AlnQuTw4ctWajELgJdTKW2X6otwdclXazFqz/fH2I/2rZMB9FohjlBBe
T+AiwL/BcsMZCP1vbJW3wnC8ihf0lQFqbN8YZtmwjw/MGFzvJ2cml5Es6/sw0y1u6B4wpynnELe8
dFuLMD4/NtaxuH8ii69XwP3uzOyxPIfnkun9mg+t9nzHU341ug2j0lzpPn82Lh8xLgFYC1tJWjS8
hyaERf/rWiPA+cFFhLGZdHaTyNR6xGjF9l96Y3pV6h4mJvDWFQwYmljSuwqJKpwRc5CyyIzyes3T
ZeEu9yqKa+8cRnpTrtc5WMPOPSi6OK/Qyr7s4hnV/OhBtyBUCNcVVUc9zw8JvJDpxG/MVi4tB5K5
xkzY87yYsaeIs0FcRdLS9YDRLvOyYEyyR+Btp9V/xv1Cno951KsTflQWdmj83sapr4CuqtIZBr5D
MST6CPutKtkcTLjZeAzd2SwZvJ+XAQpw/yLzxd3ufKzh0U8K2nCof7CCwBHjDR0SAMiXG8nOSWqM
9y9I+auRGXR55snIV+ou3i1a4QybKVR39Lgf/GT6e+1+0tKCSWeOiStTu0fBohqjCsjnCgA99+JC
RJ6s3KM6e0dkGobRbuLcGlaEJgoh1H7OpZqYjOtDf0U+QADQSy6LV3ygrjpW2z+Z9kfAgeYfskqk
3qHCXZ5CWolN2e9tbJ9kGgb7mfB/tnSbYI7eTsNIxBZzTsLBg+TtBtmeKNGWmVjJBrWB9GEMmtjl
+wHg4lmkDYtH9NqVftN34uo0Js4qblFc2krICOqqHUbYEM0/Lxt9ldB8OPs8l7l3ZaJcZvY/MvSs
XJpD4HdijgAwTIJkuBDsjRycI4nsbLB+pJPtPhgYA/4uAK1NZa4O/IjZWhnqCaKPqFY4yMoNSC5f
XT4R6ztUYP31tXBy7l8hAeiBEIQsljz3l+cbVm94eBhHY88+IvdtSXwh5+Jf/oCdHtG0YKC97t56
jokpjcV9sC8g0uJD36zY9vj7L4mxJl64/JFSRz9Cg5tnKRHupMb+mGOjyPP3+5hEn6LMr2ZOYjAZ
qa5mQMmo3Z/xG0/LSwh2P9Q9wOsgtYEN89KUXSTledGoNN5HSg49+kHtRlFzE/5Wf9FvNsFO5BuV
Xlw6tUNaiSA+lq4xBH4j2KSQUJfWNzuQk0ECakjmFPy4IxSTHyHXNvBgQgkCFLmVHvWQ7Rm3tx+y
he9Z0jCTH7ecRWwz2s3TFSlccDRSrfFXnkXWcKKLC0J1ZN/04ducM1vQ4bLfWuM7jHUX0N/cf2u2
3L+Acr66EjHN/mmGHDhBKlQO0ckmxRNzxZETmK9zaIzn4T8PkWjFEkPO/g9up10250l5HG0/eR1h
nvyba17zFcpmhLLXgX4vTCaHzAtvwaTgHTtcsJgV6qHbmORMfTzEXQKNIP+w0vhsGFLeZFCIen2n
OvsE1mANcOi0OmEqpi7CaANHT+mUJs/e24DiFN7tclwOec5I7iKRdhtA2b4QDgkdS2oK5mFjr1Xu
o2iUxz5q2H0Hvf2dzkskxVo8BKGUoYSEtWb/qlMJ+EXQWd7XZR7x7JrGcm9r0FSz9XCnfQeHWd2+
G1cJRb5JGbzBleg40it9RXrt5E+7mtWFuraSABxBdlJQic7Oqdy7G6VWjAa5Iwhv/u2/AXpXYox2
OHeaSF2GHlyLB+tdiYfag/UToFHIAEuAM1ODXigTN1sNAlgVfH8Mfoi8fbv2Y7NJdQGSdCa6HomW
dm99yeBF0Ytm27J0U3zKqiWP1+uJMVIrioqU56fmRAtch6KqVd2l/MvfXR9AVLmz4ReZTsj4KSXQ
anWbWgXA9PAq8uBjU2vV0nPNw5wj5iyW7B8JKZbrn5adRgcTxY69M0z4EICUwdDLZVjljprhUJBL
lm5sCvda+ejNNlfbilRRROUkyM4YVIp7/xxK8JrioBTkugh2Ls/SkRBP8rXNVsRJ7KnQ/jP5UGaT
xsqpGe3RXx8SqUqftRxAvQ8nduHUHf+cQWIPQ/z9hn/mOADluszSxE46xj7mlGdlc8g/myyZo/vX
MuzIjne2Akvgia15Vshp1CK4eUB0uWFVcg/CPcnohwquMnnrfQdgDOYI01UcpjbLixnBuK/tpZEQ
eyh0JYBZpHBwxHSuuIssNxUZ8FMJHBKUkEqF+MzPtNEjviMLYrHgcyQ3qIM+qzppNC8/QACtyUR8
hh3TTKifCFspjIGPvRzc5cFDpeWVVSd7nkXkdqKIMpZw0Nk4fedouMSAmqvVHuljcjMci6ucoXzE
EDWEcPGVpw/Vhfk2W7RB+2vi3H+VAVr4LsnRXPwq9FtkehmlN2rMucP1BuzxJRZoGC/JjI1oYWC3
pttJbegKUKfGgL9ljkj5UlVOkFBPmnF5tRr5s88wwl7268fsTLq+UGsnAB8ktOVBVKJ1vgdLkJQl
m/Av1U/t/nOHsXeE+c5ceUXIce83W9oByg2G65fsLT38VRNAASws8Hh3Djfk4xBJdr1fRZTI1tNS
u9AyoNQ+JzxHYfFx5WEA7F8wQeCreT3vk/4J8ByA3jYu+2AnZWq4YOUje339iNG8tZvm/qO/SSkJ
IUSAYw7ddb0dElNLmRTTdWTk/wbQ9ZVDDSCbakEFpnwL0cHVSZ4Ly3MtNSyb9gNL7qBtAPuh7dM6
8BTgPQtUCc65HIl5EK+OMkQIx7yV12h2LKLflEhD6aX8wwLFRhELKS3x4UM7zx7+bbWrrVo/J/oE
6l0d/dSS9yUkQ5MAWu7SZm8aThf7cuZZLzfrB2O5FZBsDL2cGlA/LvPjvW3odnJA7escGOtlvyVe
OZ9LTxItUQr7upYi4l/qLwmWps9cL02q39JVjxq0wMzVQyvXramOa4KQnpeS1/xAN9tJ4msyUwkB
EY02UROaju9y2WXUcNZJUa3jyMcUeynBQ44fEOTfmGay5MgIgT3wkDAbGqZbrpigqHOcMAgd8bno
B9Wn1cz5fnq1Fm/dvaDHEFTxjJ3lWAhbeydSJg7UAR6R+35yN574TCK3qaq/hha55tHrx/Q2N0ez
j/VACjlkkwlGLindECzocvTTWRIT37AMNxcOlj/bnOvME6fln3SkV75tvNOWv4QQWccvBYw0EFYf
3nTqxCJjxR1e/mC9PtqLkmy4l7NmruhrAMVoPtMJ3UZ4Kl8E2L8uKfwqWuk0KtLTcWI4RaN1unyE
egMsPng1B4ffoUcEYU2p/7Ug9wXXwHSayqfrKUMYks/7iy6vqAvyPj+2MjAXLTYlKMi4zRM0kgfz
UIUgx4LsXbMnokAdeWvyjQ4hQy+qpsJToqe1zvx2CxPEWTvSAa8utEBaWmK5Gh8jsYstsZZUcCtn
Bqu3icKQoi7O9chcLVo/rvD4vZKYUPcoIWpjvq4RpnLE+UGWiIcUnZIwTxO0R1jBOC/w0p3ImSmT
RNmaavcgnPfNhas1kbk3FSCJ5jOOOr5G7c8D47BorCyNParqPcwspBiFwcBGM6X0d65z9G3N+zkL
4QoNYSMnVIoHdQ6XttG94sJR8qvM8rWko75jU8+VvogTavQdrg8F6TuBmJoh6deovjV2HIMQVS5q
enM/ENJHRiyZMsjcV0t7YZwXVInsf3heZdaNkrtifW9friuuNPt5hIaA4X+AhQ0Z7GrCRs8F+WVr
SzodY2W0dNctjpkooyASvMUutNj7VchBNhWAQmRvGryaTtG7XvME8MajIKH3TvRKIDDHVBoDljb+
s53aZfYp/QQZ4fJY30bMgNpIcTs5cDMJ04B1eJ22z3SIw/PzD0tuobJKJpXjjPbxLwk6bYaVJfWA
I4lrz+HEtM2/vqM58pn3aY2G7Kg5e+hqfiW3H0X8hpYeYqdPYVoXi3Fu3/jrsiCktWl6eU3Xh0YA
wkTX/zLQIVxwFYpl3B/yYvoS1fbCXd8QmXvnVMPlYzbhoofcSbSCKGkPo71LmXz228Z9e67aVwcy
uslQswTKncDK21z3YJp186RLl5AevEi7Sb4q63/H1IVQOrL2mLt/LvUeUGtXeH2NvbV/zQLDp+KY
2N2ETFAlWlEP75e1cF0ci3YA9cTCyfRW16SxnHMizVEfqRomh+FyrJChcviUiPPzb9osYundwFJv
iMFTAZehpZaNAdBWJ5XdyoyyM8U3rrT/UgdwyHHi5T8S9N1kR31FGdQDkspMjtyFIVIlCtk+l9g0
VJJk36Dc7q+Y7/SJ511kpzSr8iM7OsrIuiTyOjqIomg25PiIZPtHZhpQpKUWp8M0agWHOKOYiJ72
zEjDMnFLUE99VVppCl5cQarc4azzPCSUXD85msrEYicrwQLM8xtc4vMLV05FTA7KGthQOFsn1oTV
E9IvkbmH/73SaodHKkORgp7NhGKfte07K+834y0itj8/1fGW3K7cLG+N9Jga13+/DcjhO5smHEL4
PoMwcUO4QIK4ukB4/BaQLFxIbyYJ3KJsBkRYnfqAyc4g8S1qBB+hb8UuwDcbyqEky2iFeNlM0OoR
QCkVdOfpA++UTEGIjmA9rcg3r9j0WtN6pNeOvUH08SkMDozUu3G53js1YxpbnWHlyjp1JdBAG6w+
FllhMz0TdBkiOBR5I61g1w1rvYlCJ/UA2J2xsWoVx8UEXcSmob2bOOnRUwizIE0vWDfSrXm20okM
9ghTC3nMp89JdFipV52/rkUKEXZ1DAqngcD8fkifI39X+uxPrcIxgqMOTSemvUybXzKwJSfjeqmh
VdtkCcjATGyNOC/3d4219frVeNWNRVMTIexykkF39dDYk++dWe8zAMrHrLKelvkcDPS77nX0ZEiO
mcN3wvYQnHg5XAKhtnhGcs6YgIntv2/KL5LkesyScl6/F5dLvzE7tHPmsO9+6nt0iJCQwp1JlxVD
BflSXQevI/SqwAJ3tMHvuKd9BM91hcLluv0p/TWx3GF6vo2DvCyxXfklTUNgcGk7B5QOw1cltnfg
WMXxXdUEFFCol9U9XLBCg0hogI8A8QGmLO9eO2zeou3CsblCM2UrrHle09rYBKaKmPNlKK0pGj3H
C65V9VwZcOWh0S7C7QymuCCzZErI9RNbI7ihRuOOdqja+cWPwSOrcDwThIkoPr5o9NcrYMqk9yRc
BJZ2GCdbRT/0OBA1EsA5EIwQ8We7cV++4uWK89QxCtaKwBydj8U+7g4I206hX0RceOaSmFdM2xLi
VmZhRhC4b87AurxZKAo8fZk2NBEF4KO7r9aqO0VPBeXNnVEBqrrqmB5DQlIw2q4y3Jhy63SDzqMy
FkpsA3zQq+ejYrW0nBYWg/zH8qg6/Bv/VSnjy646Jg5k0S27jf+U/z4pDCmOlUO08WVzoL8/3veb
c8mh75NXjJRv5YXiop3rUg3o0Sfif1Uu0KpQkeTwheH5B5UI58yZwbEa70RAY39G8MvPfImax60j
x+YUzWtbvzD2v7LVXyyhXnrVdK0quM1iNF9uqNLLMMhYg4c8gIBRcxQTwmRdji5e25qX7yksqPqn
bjr4/Sk4JjUJEHbfzSPMVVz+Y611qb2cACmqGOoItZqL5o0uISho/DjDvgE3ffbHPE0KvhmNwatl
2V0c2iqLjnGFUigbrJHbR6FIA7P+yZpSTRB9nnoaxDFOyc0Wa4v8pjUlI9zUnrsDM6YTZxqUWd8R
h/M8ynm14Eg6Xv0kYWNZ3BWYApHp0KeNHtcna4KL1Q7yeCj/NRPqjkhiRGn8VnqmawjZVh7R9V1R
P5XbANk4DOBYPdefaTTT05tcrg6bCMvqlFImXjFNcAd3s3FJ/eoKwyd3PiJ/VmqBpN3zJ4mPWdAU
TWhTeKsDhtAByrWW5qG5MSNubb+i4ERHOGJxk+sYGxcJf2Vpy4zIU99NF0czXsAdxEfzbW10MSdT
OAyiAfMjnYjppMJr/EbHiagN0kk9ROqcG3aUblPmXd8OMaBfXceEo5JjV9ldMRYfB0CCUCT9rdP+
LCCnDjtv78y79dNAXZRA7y3oE4VG+zbl20jUMAS9Aqm1W11aO8AI4DKR4NBR60zAZUJl3DFUsH3P
pzPWwX1QWcWjYzv3bTdS5oTlOyQ+0l1l8Pfd7vLKuM42QJRKQhjv5FdYlb8lLblBAQbE4iaXE9wZ
+WBz8vToYkZ7rX2m79YzjjCx1ncirikgTezHJO1WsVYKP9uWrFu1bLkzSL0EBOdy3PRCWGPYXQ49
WN62IaCdpnsDR1N/8yaCAk9X+B7xnOiRvMiHJuiHoJEtd0jqxgX3hnwDKtsU+7iNGQ/lh+Ldn4kc
rJpzWa9L71GYRCgDSILlpTZuMvi0kWdNVF1+VYapZxIQIKpA4ZceHI+YidA3G8qu1EU6wfXcRnE6
dKvWWqHwjH9TppEkDp+uFXwwtXZJmUSj/5snIYvMUs/I6dcyma8HQGfGLaV7cb4Fh9czHuabJpi0
jKlOQqXwYhb4R9n2Hj8ACDch0sb14KXyWQJWxfa5eE5n2aiJgY1sjHFHj8lW8kwlyVKWqgce3Jsd
eceTrxUVJb1sSuwEFJ9dfaxNGNOf+ekUWdbYaO6JVa75spPt+kbo1VJw/M41gVzif7GWvamUYEMT
HCTsv2OD29+OySxnb5YPpiCT/lpxjGR+0RuS29CkItYlxaOGXfGC6AW1E6ENf7PvmMbxwRoEBE99
FjmISK9Ycd581XPPHvkakM9wzu7k278FQNqiIQDCLvPxJqeooBw3jEwfL0dm528P78S/js0ZEE6q
Ih18iwUvnzkMOGdbO6hT3VHVeWf7MmU+t4pW4g8GAEZ7rxVnvVyIcAQtxnY2FUi1t19/J9YPLbHH
U2i7eE8cDM80Ok8Erf7d2F70pEiIMLLVKJEvL2yFOOH3byDUoT7ItNrok6gVV/dy1sScIXszjmcw
Gxhz0+foixw3W5MUtTegsweGPY6FFZMpyDxpuBaqi81YLkMBRtTxJHdYDmpkgq9MNDds3IvouPk5
ptM4klZpX8VEWFZqnBo6ucpaGBxHaBypyt4JLyaE4NEr95642RaAUpY5DAGTniAhhR4Z0C/oJMt5
3n8Ma7+S9HmVzzE2H4uv+N/r+HcXJIFXnU6ex3pOYkSwLG4dbLM08NYVr2VGlK++1iIuLVKvFxJM
7QniGydgF/wfcSFvB3Vxm1Y3ylAVzLavirlsGoBXLok9wVEvyFpBtTb1O3zBkkQ2BSMQH+gf1xSu
TlETWHk6TCJNuiMQoyOGvN52ZuD+l9w4RE7Pkveu0uROmeROrZnI6P26R0JZk273G00WNbVhZOBT
H6UNtNVFPGmaU8fgCwXrCaz9L0vLREV/rHgVGe5RcwUfm+UWg30SiuHiI6hMZaak2vhSYvqUj+OH
ffmZDkL6EsYkg8NQw7zHiAJJpOcPVULR726eqPtIJLIdUZFKEr+fSZkx4Tyt0QTJntjFTvzIGXr9
fzg/yglRW0J/29RMw0+gfWjsQtVcaacmyE4a/yySkGRZcoa68dA6h8b+Gp5l02NfgvjEpRyd9vDd
VUaXd0Wzk3RDel5fepSkSppeunaDF6SjwEOZ8P4hMUCrb/8JKUwTkIMCTHhVL+zGDg84vLfLl130
fGhDMDphpD7M7XB8bMHEhom6tSv5j4C9hOw9rP6hqLlNyEI4T6YM9o9aAwSyWFOgiwfgMlcKNee8
PZdddToi8thW8zSe8m1RbmssCALEExNBu7j/hDepTVcAZdFVZJRuBkhaZEgzNajX2c5Wvm7I1d1s
OBDLivTOp/LMXqHa1U4ulP9l2XDm0Nga0xOQVH3yZjKJ8LbrRI8Ym5pVVVfdwRxfFSByMqpf4PLO
q4P8PFwJYhFGxCgzyXZ+gYuPh9b+cyWjEiyAKiSjXWzauOFDL1HuILytc3+1pn17yGkliLr0zdOh
8k65N9u88qM1wmYBZH5l+9qdTfXJDdC01yMBootXdEqAl9aOEz6T04g5zamDQCejTRQZcD7HD/mO
4kYL3deSMW7G2qVNZD9UtOPjIPsgINIjmtESESiQe1pNymKCU7bjdmiZ6xgoYA8GLehVCRUxTLps
HQBp2jnwuBS7i1XOmJ68kB8fiXq60EnNMysALYcKKGhRWkuVlIQoM8p2A6G0FGzsIKeQX28Vr1LW
PVRpN85w6Uo5DXltle28oJKlHiWHKOb3mlA2Ph7bkIo4sZFPkYMLATA4kiMISClvqhFwSvp1fUmk
lK+QvABlO/OSTNHIM3PTmu0Xq/O4Px8hcyd48oGCF5gqRaKkbNtsw7GxbUdpsR5wXLkHWm6OWsyh
X2CA62WLBSUtKX7uhAIDL2OX/z0oL7fWX14FrRVsfvyqe6bd5J1io0/xy4lW+/9khwXo3pRnJniD
WqPlmzyTCqGrlwVDDQW22BxjGghwwjM2Cqj8NFf4mNzwWcKImmyH3gVbvQ7kAzcMlYSI3aJ12b9J
mNAb6jAmpQLobC0+7Ia3cd1Xe2fCXkPZgDFjbCOPb9ASO9bOPvAgH18zsyEDzOhRaDKZDxN9VZWI
OeBL7ObV8w+JkICbSAdwJ5HWruaX4gvIG5WpRJGMHO3ju/p+iPg7/+NnBigrqy3qlOd5dLQZRJIe
zYpEc5Gmg7letLivboln9cvtJolthAhBSgABgMq0DoOl2s2SISUvOwIPJhr5u9hQDvWe3nOsbB8q
xtfwwI1Bhj1rWBGsAkQXL2lSeuvi+mIwqnslkn/uqZdyOHssKZqxecCuvOp2AfrMhHrnF6n6FzPG
2+U77oa9qaXb2UHaZG/saYzccss3bVxHoH3GilBTSdVxfPcDr65npmoSsvw2EN47oPgWrG1kacnm
8FUOygA3fpIcptn6Higi5CLYShBBDA0HeSOUaj7QNmb5kG/RnDDlT+MYfyBj17ylihHxncknfUW5
dNS+Jk+vmycbfY3DHG6A+ohO3u2h17q0aVofrlg6xmBtjJE9Qp7uFQw9gK2/2QOQ0MI9uH/5Nq0M
FwDv8Gsg9Dl8x9eoBbVu5aseQwz1IZ4F2bbo6Uch13Gie6q6Tg3pkvHi87meZYZFrJDABMr+Aq5Y
WLVFPfBCU6en6UO00h9WmWgi8ICrU0lw5R6/efckOvVw1aMJAdCBfXzG8J1ZEhgk7ZP0oSfW+cR8
8S7kJztOi9+fdhDXMNEw7/Gj9RhSmkegDULvPQkncqZvbWa5ruYF8niYwwDY9UbuWmpXtbEd9asA
Aoq27/pR/lBuJGBdxwLY049lE3TBefHfb/MYd+vJn49Ct+nuxuPV4pn05UdkrHlbxfX+CGk3PCLx
NWbaqWUZJZnYSVdQaF+xBY2eH7psGVKbrRMIGMq/PxxhqYYWC2oYDhMikpSt4wnHVY+cOGxa413u
w2GQfrutLgD+z6HKqp9aW3eRmsmktoMq6LQVhzumQXi4Gr1oHMfSJi7EM4perUYtGQlaAQsQFvKT
fJ5PoMT6oJGwPAntOOml8pwMafxx3sGSY5nKE1g1Yg3L3i9M2jPPkJr5USQIIyXVsAkpNxhxCi0C
/8Y6jH35Hixb5wq/xmcRByEfae4mBfE/D2TCz2xG7K7EY6aDiiAAuz9VVZl/PPP9HHJ/ePWN8UNx
//Z/3ZvK5q7o83KvFF8hFA6YW9A17ddDzCoQtbJE4NHYrbX6C3CnvbTXCEN6OS/NixHRhcmVMjk+
pFl2EPDyeXOCP5gDH+6XA09wdIWI68AGoO21Da0uExrK6YjzdMda/9efZs/933GR0EQaPWTCszfn
jR0dNXfbZZQCOAO9hvgzdbNtnBYd27Yy9Az5rouS432mbrHNOKY9ycFLvy0AawJnQvZCSTg4Xq5k
SehJ/pfa+iG0ky5LWaq4HoAt+7dtUg9o0Bm72s0rXrqC2H0MJ3vOvjm3BJ46F5EPvz71YnwPHTx2
PAuvLzokGOQp44vM5XqPT81r7aHDcHJwdLl+XZmYbqilRvfgalecMdcXno9niT+Vc25WV4YSdwjg
97fMUP2w4ltFd9434yjZlJooJdMB8vsCiQpwUeTeJAywqfQx+n6t6MCTsJmF488CIhev/sunu8Kh
73AnmsWlYZZhRcSbnap+iBCdMfotbIg/GKSRCEoKmoKVS+O6oN8UzaTfRwdLO1jg5b3JsVjlQOZe
75CBZmA2OXnBkteitafpKl0Tmmuq8vw3n0Tcs6hTcBkx5KslTx6n+MdClRxtjdPLtEpA1f97soWv
tXGBdA5LBO/yn2CAJX60H5B4Ofmib8L08e8NEhr1uCM3u4SaA4FEFhCqfwZmYUhzga8IFYmUv6XB
8JauGkito4o8U+EV809vzXDkw4R9QTYkWlsZ8hf0+q65ulXIdmoKT2kmQpFugaEZTIcnRkGhRSEX
OkmpJoubks1S0Uj/E0O8hrROR9neCBzZ1fjle7WbY9o65MMoJ0mxd0zYQp4naKG9XWmNbwkJrz7N
IznPqZmZUs2GSFGEOLoNBVhn6LLDW4PeXAntdNFILHbm974mDfcEiuH6GDuvBxwWK6tZ+jtLJtEA
9JfPBeVyaUdao9yyNdSg+OJJRWla0uU/GvfC2Mgaie+Z6VcAvd5frqJo+Ljj0r2QB2gaN4n5uTWJ
30fxFgpaT1NWizmKiWB1HOOk3O+EhwAKymbf08ONwlCjEItEmSddhCNsf1D2WqlQrTJc9YTNbAZ1
dub9rz9QlNw3509PGTrbkbDUw8c38yS0f+BeIiUHcPOy2giMopKyGCKbd/b388rLbhETHKSIcUxZ
f71Eas/LNfLBoN3uUYmy/i1uZ/R763vdXCv5dkre+g/GOHm9sghOK7u/+0/d2mEQ/GuLmbhFcDrD
0rJN6v5r51SetbpXedJ4Xrkf/GuSsL7XiLW93gi6oyWv+jq2H4agKzyJI4PNJxFO234PSvvlv1fd
ZC1b6kEo8rL5vvwP9G88HDpVhoJnFlEoYf/BN90akwRqXUFwIsv620kAEouLtyFhTx4a1Vp8kl0i
DQ6/pg1ZV2kzblTOAG/J+JJe+7wb8qAFw8+kBfomCvDX+hcmN504WMBY0gPY5dQZ+5zKNFo1oZxj
DRvrDVnRPirLCcLZbucXuEpJJTZuAeVxJoGrGKTUeV1ELNJPEzJ9aZuRkaPCNhbPR1G88ROXSS5p
iRoYfkASX/twChFp7qEWJdBovme/M7yNUAiXYEcZxhN0VmHlomCNXZrVjjoTUUfP/qj3+4zdTTUO
b9b0Puye+Tzk92HiQz43FhCAEdM6JbOveRNZw6Yfj9W+0LmG3YyoKFcKJtexSHca/J59YQ1EBpPd
AmNJeBRpXqAnsQO97Vn/XMrU0V9PAKB56fz51/TrZ8td5u66ogsfKjDMT7cEbjgkpi32kNaaQ28m
D/RgVa1dXxA+aZ8tw7iR/3ncc+ejrhh3Rh9UTF6XedJy1W6jRTa7bXN90JbAR/t9A0t5aRhbRhL8
GHHcFSsFZSo5UdHQxKOD0FDiO3UZlftCrWc+TPLzobyO7RGEKNyGT7V0AiW4E/xidC6eHj66kGCa
1zX0g18hidvGmLbcTNqHVtbmoCDr+8MsBHltrstiu/LV50ZQgtNy0wC1ac+L5Toxe2atKk6ksT+c
XCxcRdEwy5fpm+7xu+zwu073R1ypfZ+QELwSelAa6atcWoPbriNDWv1XpwhVW5GEp6dvL1HlSo8J
5yCdorlwkvSOLZq/9gjW4AU/vt2l1i0UjYrQP8M/wLyEgUO12AudIVavpO6xbNYtjFxxRiL70VwF
yOIp7SF1orwuNJAX45f/m13GktCunfpaKIn1PAMcubYNdhABNRmfCJohqxsT9zakpv/mr1OvjrWU
NwCywk93xiiFYJw1J/NRChXQanlu01+dDLjbBZpA9q0lAkerwG5L2hfrXxE2zOvoldacRSFPjTb5
dWbETuz8isIx7PklZH3YK2xfR/Jp6T0klt6X1dvDNqxp4xTQh1h8c1IgEjxtoSoUKWngYZV09Sc5
r+3hFmUaBTjL6NsUUsBRJq1BkBFm6JYZASpq41iDB+iCARK+dJbX/bScyeGLT9gaGNpW/CvZYRaK
9TtxKSgr7H/o3vlSuUd0QhcjGzqvLs7SmZfxF3U287/+KL3oj7Da0o5F5nXMIriXZstjlDTnV4q3
oSvZUZWfHjizpG1hXW6aXjNX608twbyJ1p/5GiTyI+vKgHciOkA6xwxoHqmHgFU0ltYLCmaw35hu
W2ZUnuwy7Cn1AXeZhLhlbCNOuT/kPMt0yOL4QbGK0FaZh0rpQMSq4bkmgYqvl3du5zryX1qhsvnn
RjKGsdn7t0m69oBnBwawYcRijNMp5ysYLjKvS4kMmhoEMpH8gkrZm3re7FsdL4z6G9oHfSZC18oy
m07Xz+jN17stT29jLY6xJOvZt2mdkSZLeJEg+YX5tDvOmhk2rD5kSYsdrNAiWqCUerWHyNaD6KV3
QGrrT9F5/SBFalZZnFYUoEY0yIMkC1R5sA7pwF6wgcWOVGSUT5mlhUbD2V0+Ylt5tj53MajRBiW0
HtkHnO1MJR8CZMvXrWjtO3B9l2YAQVvnBVE/gsT5C4LSFBiZyoOLaNXU/sq0Vo3QLqSQhZMXEDdQ
4zMcqxoXwsgtm54pI+4929vz+gGVGSx/Yji5pLlvP+UQMkGXtxfmF7UFwf//XKBDPPhl8iz8gP/2
S5TBQtgNFXV4g11x3gsJl8JqulK4etgoTTmDrvugaJTBNXjcSPP3C3Zj29bPiEGrA3s5bv5WQSap
vkvWC+bDQSBLLobStYemhgw1G9zmoOQiZeibFTxWkEXW7OhnMpcwuRFfFo/JHhiW99kNlttioc5V
otkVgWDRnlGcSkYroymi2BPt3BloPbV2XmVg3Qfdc91xqRGB975ojhaKP1WTpA1q10embLG0iNiW
GbAMNBCPXbkzjBGIVfa41GrsiGw3Za6U1JxVBUkNYmD1CtIHmgwn6CV9gR7jKspUUFD6fM1Igjc4
5t1FBKWvMnCkvqMvAsuJIWNz8/w5pZOiw7KrPBSNA/8BfhbYaqV629qaQu7Rh6YFlf/ffjQJlSyP
XozO+r51Ov+IrjYuZQ0C28ouV56sXykFtGGSypoYIun2XaVu5od2ta7MCpYUcFQJLpa1NsVRrh+a
dS9HL0FUrXs5JbqBzxZ03CJ9j+oF01ilXdF4dmRqidsz8fKKPvD0TCAvH6G4yakXSrsLAQiYOF2W
fXhEYjOFtn6HWUaxeQxnRUdL/6PRLUWBQVEsBXyo0cU1rNKIZOdWAysM35XSpKOuKXjX9ss4sTO8
hdMAwBUGs6CAn0SFbBk7FmkRjIIWkHxEKHNiKe6HJlWzgCPRKgaf+CxNx1K+NIBaDYlJUkJw9nWC
wwitXKm2S31qe/fxK6s01eiLFo6FJISNEow+5RWBjBP9nbxah9yjoyFSqRC+XmWdVaNT915GO7NH
whIBqFGQwDtoCOXUl2W8QeG7MwEfoAJ4LAztBQ8EQaGqCp37VnFo95pB+mgqfD0sdG56V2tT9D4J
Di967NRSjKw3jaA8P7jQHkLNLYS+O03Z+vkSlU1ghq8URSP++nMO6kFKjS5/Wmm/0OuWUx+Pqxvt
FtYO6GMp/3dczcd2PXWYk2m+u9wqYIr+AT0XlZYpYGqeccrNarJ7lEqheXZJs2n0zLo5PzjpLvtn
FCz/N6X2q5dnbubjc3+eWPB1mpia8rfKqYmwgbybQZCq4FOTi7sCmjJ8zU1iB+KZD6woqfhzLSOk
41Nz5XzJDSDEYw/nVRtRcMRljgOj+ZaXUCerV1NhH8z4kKAAnClY6F6S78D/+8plJeimVP0OV1oL
uzb9jqjp8AwNehKKEGic3L4i5DkfrkcFV8ARrq24O5KrBes5pmMoAK4K47yMLQ3rWHXQ0o/+l0FC
Wc5EGyaKFdr1XUaExz6BLY/rsFQufxpRnFT3OiTeUZ/euIidUj2D40ozyRRPdzcQ4Bz++dH+sllt
RHXSo6Eh0kbE15O0ASV5nj7HJbrjTc2akyfcfFcWcKiD1Lee+t8U+ePpBn1dagCHYj0G5U9m+XyT
TiQLhZnTZmObaT4HFmlfiRmnA66CGanM+pHRM37v4s81mMKz3/a5Vuuqxo46Eb5sln9I4WKAkvC9
2tI0jp3XReQO6qpqmkg4OUaGKWDDXJ4AZrdGW+8l8X3iV40H0FzLRtLBYl1t2lsBjlZdWBbJ1F83
Oe7pa4755YKt9PYaMTv34zlFcS812fgeGYdxUvR5ojjera/eV9eL45T5ZG5Dxg5XDv7Ji9Iobje6
nRudbQx5lpVnWb8TH67vgc7CQ5z6Mg7MZFYc898xyyDKfhLDkKksNkZIY0+gkAH+7dDjxlYmCyt6
t7kcIc/8YyEWetw07wyCuhN00+tf1XhDFrlruu9OUyWm0JGriN1nFpivM74DbqFW07Bqv6ZJMqfi
Bcth27ylx9CIorZY2itVyQkMFy5GW3KOLWfZDhnRV2T3ONNEykaW7LeEKcz1j4u3D7TvPz3mddlg
T2T3qPaeT0h2oh+O06beN2XcWzGjskelq2Giw+w0kzq5r0tTHpG6eDnwrHuYEVV5JsyCli8yPkG6
KUTrD+eZQBsRGKyRWTnNGcNu2bV3rF/kgdtU42z7lt37CeWFg91ABHs0uL7LYlXbAypHWDGadI0L
aENcw7FC06irUmO/Im7DKlDG3yNR/eW1l2CDOYlFnhu8ql4y8YT8oN9eGhi2gOyD/mLwuTUVriFf
ht6USm9fmQoxW/hRCMkud5VAj6+UJJ9H0sUTk6x+aQQ/Sp1xSeBprPQBHkWJKYo/NQnmk+hLPRZg
xiwxChps9hrcON+fNdXrrEFXfxfFVaps6rwstC4KVc2JJ5DiARtIupHgojMmcnWwzSWbRKZBA3nJ
4WMiNzNpQJE38KjO8TiUhPhl0OJiy6IlR4cPfH3Uc6TxCWIDp5HEOO6rbnh5iAeTfqt7Atr8rfWO
/H7sTzbj9UsLEqXjb676miGnvSmbQ1zTPFZbCltcj9xGA5VX0YHP8zCPegdaHC2LDJr8EJnQAJly
TUPVbYR4ZsMBuhDhaY69kSIg9zjILSnQAti2pGwZzDsOto12QhxOpeWzcf+24qQ2Zu7VckxA5iwt
/5UN41Ebwm5SnmF2zILrTQu4J3haVSqnJ4Mx+6tEWWj9Zo0sdLTA9tOdM5YqpP/6/AUZR1nWJHfL
eojcXwukpqzHVeptBRk3+2LIMUi7e+8q8HoVT/nPNrsLa+EXkM7EeY3ai8V4Ndsxkcl9WAd1iKvM
GC4sa8MmU7JlqeXgTsK85z/3RAKva/W4IagtbU01L035GfaLBIVp/AgEYSVuA1qUa0bxrCkCQq+P
I+aUopXoalsCPk6UU4EtEtT3ghHt8mU2bQ3bM8KhZeGnqaxxAJV3FAgpiNXpKHsR9lxRZ0+OxFti
S6xjai1tcaOl/v9gVRE7ne/5Jw4OOLshkRvc+cNz4fWMqTqTz2L7N7tvXupMgHnOlKtrEg8vPEvo
od5TsOmZfXvOces08pR1sYfIWsMOCb9D7ypr57ZahPTn6h0NdEM/2VyrDdWYd0WnaIbumwEt9/Gu
oJSqDZsKqrojtcMxfh54I8boPL8mB6uw5M7YCFfHDHgrLe95VnqUs18l4fcKC3MnIxAv8wJSxZuJ
RfA6cRUQq7yBSFjs0zXcw5rK85Hh33N73XNLGXTiKngcLNhhT8UDdYTxfSlV5eR6ZEqJ4zA8WImg
HTJH4vHYnDKMyv375QeB6fK1J0bVWwoL21NL+N6rXtot2cI3zMsjqXZExxBZW+PgW8MEWO2yymCP
d9hpKS6aEH4v6x3bSsDyjqU+i97PyjkIyjt8bBCf0V3jnHSuTuveIk8UWrpov0WJeXDvvxz71gXd
OYg9j9KqcoxiSh2xPlOS5uBnRAAo7Zlgvf8mbkIL6LZGL7z17SUvZA1FcKzI0+5kssNptrBVE2L5
PeZjwEwaTXQHP17dyHTmi5e3Jz1iif3qnHGfV9PqkHn5ejYCVc2mfD+vl5Wwij+K4M0/0Ybw/Hfj
W/8MxAXFmcgXjHS0anaGr3pAHD0lMk9Huf1Sr/0gmdDgerSNQNso60g9vUHgrbBce7SafZ6nzGO6
tY7bMy7yKeBdl25tjaJht5wT9TGmfbur/4oSouAU5KyQzaoq5KTLgo6WLTtLYa/5IPOIJAPQRzMd
4wR2SLeogMQhWIfK595qScYcjvEEIKp7FU00EmK47IAAbKZ7260bjpDXvVIqVguQgr+EkcQNWBZS
5pZn9HSHAHKoLNsgFkU2sZwvWYjNeaywnVADnhHM9ijCDUN0ynaNhoxeRuWxe1GejiDuZLYRj9Ny
G10SEZ1CLREXhIZTB9iX6EwAZnLMbW1qUEPTLH1HHH64RE752E8h02GnNTM7G8N6SbXBozK9r8lS
vK+ebYlnueHCseZQ3wgVgsnl89is9PEcOvRKxP7Jw+DKaXZ8GTLu8efW4EHDtL0soJk7rywACHqv
4rC1DqHtIHRh7pytvDiRNI979ME984+AxLU4tR+0R1j8wHlaDStKuczIpExibMUTv8tLx88/uLHJ
xWs9gGVGbW538le3U9rGCnpubhZa1ulNpxL8lXSO+MKtD5czM4WDIGx6y7L7C22eMED+ziOrUzoY
hLNRGzSrGO00ld4WxIt1dlsz51YK8tFa5kvWR7t1JQj7pz9jj9uR34DvVXy2VBlZUFWMMtwKr51J
9vugJCCAqvRm+ZmbLPfEqVUsRPyR/8m98eghOd67qAYu3ExrcsTPO3YAF7WKq3u8F3IxVglhEgU9
3MvCtMFLBqT2oNlC+D+30JUfI1UnABnnO7BcxpZ18DETcc8T6ztNMitRO3wgb8eTHK5RbZtxPkut
lq4Mtd9u+abWkqRBydMR56dKClT338jnDv3pew/CZDuTb9osrI6RiqAHJR2B8e6Nx4vM1/fU9xY6
whJj3M69b/Gi1oZGvxFK6ESFLOZZ3E0RK1vyYVy/SWUx+dUqQpgnm3DBxT10dxHHwn3vEZUCe9n8
7fqugSBdzT8a8KlX9EG3Oobyp2/bNbNU7azdotUPsMGjNPtmc+dccVMNA57IBM4A9R3ruibgMC57
+bh2KmOua9Rza560Esc+Pduk2LsIavU1jamuiP3LHDwo0DYBjWiAkXN7VpgmUNm+TewOmY89NPes
Ih0jUVIa64kDbvo3cO1i1UD45hlXvVoLg2KPXbF4Lsn15BvqPOYoSAPW1NheOWPCX40nUSkQJQqO
AdxJ4xHzHo5Alxu1OJS34l+Hg0e3O8CCGc9KqCUXft/2R+S8lEgMQtM2gG0uhokvMiPtL0PsT5t2
7apmz8CCTjSziEkjFM6jkYyB0VLEqX2sUqwo3fX0nCZQRkFTBAgRAhBBJgic+iyALZRvtQepUZqP
NxmLfXj9TIKR57w71IiWrMhKzaRDaGDOiZdhCtGsMtHqBY4azybS5V0f+QMKNSjsW1TysKrLqak+
2myJ/ShjjBdYMWFaljorH03ZWCKTzUR353A4kXqk26ia6h06JhpDL04391PFzBF0RZ1TdVX8I9/M
h6rpjcpVhmCLYiKdmKmWuWIuWGa9+TSbOkFmXIHiko8UYHVqZ/o/Ors7hetEAZ2Xyf4xRtpIRKBm
+ahqTlPCWywiiL9xfGQc5JdbOwzoVko4Fah0qSvk9b92m5qUEesF2ebsRNtZ5YxulIbDLYgcud2Y
ZL6tBm0hbyXKuw3tJCEBwp9N++RT+d/WQ2zh+CcQP93l8OKSbTESi8KczSgYZBKkzWjINPU3xjN0
GQC10SvxT2eJKxeKDDL2h1DMiIuLcX2sKdQBtRsdFNh3TW8J+RwtJfJHc9+QiGKscffWFMJYWQkH
3Lo4PQy02kUFRyzxblu/Xz6xiNR0OPAhtJ5Z8c27dhxxQRrbBrDd5K2JOlD89xB78dI8/QjBONim
J+Rqa13ut8Ov36hu7njExtfoHvUKsmYAJiHwTppgleHnIjK7wBBqg8HATSDg+Mv3HctBs4mwy5ab
EmXzuZCJaybk5v6qbIiflJGYKwsfZ1kBStJqn0EuEwV/+qN/Z/B8Ini5WObFkQzsMJcZaQvWblte
Z+1t9YdUNaT7Vr9QB7SON/ylrkhWUT0H0loS2o3AK0NDVq1yv1K4EEU8/BXe/oFkTJRrvR6wIJ1F
yMA+cv1s2NpBt3JaMl9boy6/WzqjDPYTxHzIMg6rBP8GPPWbSs80NJI6GDi4EN98sH02ZnSWd0Mu
uc+RFZOQFxIHtgIjMvUIrGyLdko/YqcdTZTTwfnoSO9IfuD69EDE6xyvJoBGCnEcKucDGF2A6Dh2
fB1dqEIGENbo68F4ojGP/DmfDbZ/Z7QcwWVNC2Psr7U3WQH838ThMkmJDH6klUvUIak+Zw6ixlCf
3eL45y2b+wlJcJpd5FdSr99BlSFBl254vMR1oGyHGaOKL26HPFX48n1hxB2XaH7YifpSN5eyOkpL
4adBj7keC/KihtyOaNBYaSSqlPo9BMYWLSpSoHxSToT46riMvLphmjgrgdxWxH5TqUTBIRp2GLmY
/w/C7ZhyJ9LJ3gToX1ozjNT96QpId+E+mYsnwwMIWQFr4vP6Q3olr8Uos1+lPXk1KJOWJDnCuyg1
tNqFU+qrrWJCQCp0frje5QAP3fd/C3hvjHCqi1AHUhFtwtjs7Dsl77QdwSL/tIhLIwsg1D65oL7T
87iTiQRiwQaTwg/WNETlAwj2zrUE9ikKi1k7EOJqgxLTLWJonTCmu9cZ4QaQgygutodTjSnG7tK2
IydHvM2ozUykJaO/B2Ec9VYWdLUOtQoymHX1r8yAgl6pcP+oMkFvmKcQRYjbmVahyOtxbA/eoGuV
hLXNMtTvKCJG/BnLkGZfTb8Mbr5u+xgos3/eloEdgowlKzcYiMGpOmVwtI0nPcHxCnofeXFXGTCs
hmW2znDwlxadGZcDJSRLcaejRYSHBhsp8F0GoAIYygumC4uPKBcm0ZGyoGZytSEWb18DlSP/Dw3K
wLO25yeY7secbSb6bwbFWNr7H16qRBe250h6jaa7A/DcNY2X30NwErHHInsu7eOEcIqHHOzhqFte
7vxZPhz2R7oUIxJtH4CsU6n6fNb2kWNqj8cQZgK3AIARAvdjcnIKs1eSOwB2a0giSKprUKubfMc4
MTt5byygxDkUkccFDnIqgA7P0NWQMPH0imaxF+WrCFqRIVYIWctS9U7rtnDzdu65Pn58CE6gNAaj
yb0xGygy8plI+3lJmuQI0ZVXrqZqr64UDMXsLO9Bj+2hN56oQjWEiPZ592LWXefAQgN88BTfO9ey
BFvvqM5y9ztIH2c7ZmMg+W7z80GJqAevJpr6s1Trt9wxrB0pdVmBelHPjN22KAoiuleOvBqQkyAr
C10tByb8UxVFb3TchHVGvc4i6TX0xBdQBqdzIBD00pX5EAG50dwHubu0TYlPECPr7HXLrggfaJCu
UwAliAGxUDIvfLjcBub3bDldIQqHpe2jAofxB8ML6uA9RsXqfvtkwarrf98I0i1j3jIAr/afSdZo
gWQx44IHu5q+5xRJg2l1b/l/kUk06Dp/dhY0qtHJuSKiObofLqeYwm/zLMLzMO53M4+ZyzyhhKqN
1xKnyqotkyuJ8wut/zB7GBuizW7m24DujDfWfmAPW5TdQXjMb0HwteMy6B/K+E9Yp9bSaHsLhr+f
GEgWWpZNadGminxPwEG6LH0feYgbrxxLjNBZKR5rXHZbAWqjh4qLyQpE2oV2yi2mD4IghITFA1Gg
4kvRNRmWYKu7heG0DWGaD8Wo/OiJGShcj9JDAmCTF1E6odTtqCHPQUcwK5Ufx8i0wCs4CMOBwwIJ
hYMMIlGzim3bX6JDfD0SHMQgWoQqhvNx8kRL12nebR+YB6LV1jk9UG8MYbuesLLK+AhuUk6d3RYd
VWddIMnzMdL14GtjSaMAUe7qzxivWDAnAOccCfHY2r+077hlTOUmUahg9eib7jNIGA5eBNQN83kc
C1d7u4cPuS/jS6hTyMjsmgH5VeWWylRJ9HkK+nsUi8+V7b4ygTXq2whpRihJZRtu7+7hQEq3GnAA
mmuI33yxDfRSUZhSFB0IXCTY0/j29KTVP0c+sXGlmwhb2Ob65ClZ/sd4UqXKwYldbVYf6/Bltxe6
gmro5YOmz2dB+3/0MXbw6YirkVpR9pZ+ecil5GmKzDCVSMSTl0WUtv2cj4l66O4H/NdO9/I/9Slr
YpA4pXY58SLdVVO5c+YL7VSZftKJ3MqhkpV6xRWHykkXEWOyJPYmEfhckfY6xzgSzvf2ndIyJB6O
UmZKGXSK2Y5fWpKJU/wLl2NT8jUQvqbZg5jn8TLuL2RU7De25XjFbjJrJPlVpVnCX6Y/kK/tr0XW
GLKVsDPrUgnSwDuSBC20CBuYbIWVaT1JB9r13xLUcnlIKT/CLXpMLyb/MNEvoluOgXhYdyunHsU+
pxVkcyFSb317SkYV5ZMnTXhFTFbcshdcDvwMVyHukfKCcYkJ5pFznQCYQ8NF5gHFJgTl7Exqn3eB
Zo08pRE0X2HIClikucFE2VF7HDL/axSyoqgD7EB9hnzhcCP7SgQa/qCWeGafFwK6X3hSZnZNAJAX
QXYgw7OAewy35ncXJLwhQb7YjvsjQK9zvRnyvNWAAH2MnPM8wepLgSNm74Sv8JTaoqkrGI2aMXK1
HknmVfZ6pMhp9b9yZsWq3GPXy2v0Ri8RLwiR8uisFDYWor2s6qO2kR1HYxzY915AdiADg40CF6Af
8eivHCB2het3sWHK9B6aG70t1Bg/rQnfREyFVaD8Ev38HtjWkv/HQUIxX577oWoqgDTW2Hh8qg3f
ZblL2xuAVffcaMHZGip1xNmkGagdqZtJclkykHKF13ExC702t/f7NdhisaHLS44HHnUZZKxQFJU3
q5GF7LAN8t+Btnih0Gi8mfcLRuIi7F7qORZC1lY1gUv8VseqxEQEyyr/qVIXJ8CJ6uhFTGuS4m2b
SOt9xOYSEEvikmmkfyjVs3FdFxZ99bBTlt1GwfGuDKVdhvPvGFpkNqyXt6fU5RUMnCvp9uHapHlv
0b2TdZZuDbk385b+/GFobEe8URKDOMS5YjZugZjnAmwk7Yrv/AIn7Jrnqwr7L59hn9Yh35cylnyt
1nYXE/9BiBVG/wQ0kBRy1KhCw43o/Z19aipSO35XYTxW84GlERu+fHDaWKqjnCpJLir3swHK43Uq
I5BirqsV70ID7mpdwmxGGerd+p+WpbcjYvY0B5ApXLJTiohR3UYlGabNjTktDMVl00aPFxBw9l1I
jmooEQaT22UmVdS185rFFuLVfDFzzfiTeZLeyEGSPVssFkpeSK9f/1VboBDZZ5rJCW327Ah2ZiPG
4OWYRrIhxn88Flxwyn4a+sk7YTv1VyYBRA2q91Pkw3ekDduRe6Wf9J+Ysj4rYFQJUc72SgWiiLjS
vsfA09VKo3kNhzgnMr6f0ZjqaV6xOoiNKNOoG7mOcj/uzuVVqDI1jJ/MXhT9YX+vC/IHSKJbQixq
k3FnBufukBUosAB6kSAhBY66CHJK4q0UNeIJetwvDTW8o/lxtX7P4b0MpXGKD0jJGiw1UcdC1rxm
obY6PqtOZBQDZEXMQKg0CQ8Sg1LG0ih7bSUpnKgHRxC8bKnOuCzLgETqvy7Htxhs0tozlRUWEgFQ
z3HCqgMFnCl7JkQSFoawJjDmW/cenZ/lo3v9ipi7cfVaoCTnMCtm9nNr8x4vQOcqW5n9wiP37tcH
uPX8yuQHrqotyes/H1sefLXovLFErIGkIhocR3Na83kMtTJGBgtgHnrSqftDY9JASajPezZ7lNiY
5FnxfDeiY0o+dAVUtJjuhqylQ4Y+15x9i9axAIcjOIUJDP41CQjUPufjbuJDIEZ341fMiWKWSfYD
Nw3uZfz7pXbKG1+swmacRD+zRUDh3B3i9QeEbd8t7gKLkfi5N4tSDO0Grn3/4uuPbBSxSu9E9ZQx
GVr0ct7XYidWm08qVIxarfoc9CqLItGCrL+iqrWA2ZWx/ljs5lgdWX9jZ+y0z/iRUz0ubbwcmkrw
IbjJnFKqCDw3jKQozmnkrDq06aMonY+niNlgNJ4x8mdWXH772/84YD4FoceEnV6Gj7IVeKbdSR56
AP8gRl/5ro+8yPFxIjE/GMO/GuTG7DQPWdVo0Ei4j+h1V0fn9BYrAU5VGv60TwTenec5VC1HvW9d
/TdP3TO+Hwz5cpT9OQRwV8WFcfibSEGCBZC50OTPoUk3iJSHgMF/VL/ZfZJ6CO7NQUYQkqAa/NOF
atLSgqHSH0yZFJMV3B0h/a1FrkML89VmTUgP5lA6HYRoAMDRkTSlxZw8HZJoWa1fLSrBdqSUzc9o
5Xa3TLLarzBfwbDqVRbxLJeUueNcfxnbvrepi9n2TFF8S/DNoNC9Z36JPn5qgFiIG+CeBA89nuWj
JYtcZdAM6MTpyYTSI+l27VARgja04Rg5M7+XhX2TVNUHrWvwPYk7qwq9GJubUgjvohtn7jmrKYv1
DaEbFpidY/C6yjDK1I5u7HUat8vzjX74h221CLuhHhCFj0lG9VJGK265g0HncjgTHnkSJKpxjFLA
WEERTT5GdcuBW7AN05/1Z/h9BCPsEwpelNmg3KgJB+PsFDYCvstkEsq2ieB1OoyTw1wtaCsrbwBu
aVCmh/diiT5b0o39RANt1McU2DyyodtahvCoLcLHkIeVe96txcrliCG/iLqdUUBVc9LzuNaP9+CP
ihp1F008MKj8WTB77Fs7PufXOqp56zARJs9tyyEqHya17wn7ya7iigrzrj8p2654adA+QSSFI2xj
EsH//GRhGtH4Ql18H98unrIB66AdmAskiQjhGuKc5k1aXgtxfYwaUqVhoXv000lhzJlPtp+URsKb
+WTicXIq/EEuEZsxUfUkpMGon+6Xl0YcVK5m+hqHF8Gc23G2xYk0i4FGcJCQ21A+40XXqXZfYhIx
V2rxcJ3TKOzCyqmF+XWo89Gbo80IY0QlAjrnx+ceDANo8VDolbIHs96a4v2iBlw6/QkyyDpE74hu
SoSaUEQYAksqNGtYx7MJ9UEizqGjtKljX0/aRgEPdqRRLhVLfsmyfQ6IbTIAQe9apKjSstfGK2jV
3Eql/Fu3LWyQVI8H/arAyUfftbSKzuK5KZ/i8uRkvUmmlZ339QHYyXjabQLOetwTKXdBYgNXP78I
WCGECap5oBrjuTJPol8ncQr3/zMb86J5sRcG1kiGs0nvFObWFXnhICS2cjRoQntqOM0UsIx8fdH7
PrEjsqqu8Ms5JVtJ06JRPY5uc7U3CHZDPkLRSmWHlQfJfQZQGP9JB7bUEZEUn3Oeu9x8XFLfE9+v
mgRsW9dyDkwE+Wlja9rf1w0D6YrWaPAtc5H5nwBjrNTi5OC7O1hjn+TVCBpFpBW9h053ke7+HrGB
fik7pjt9DDI13SXfZ7Doi6rz3tfJ/4RoAav8vrisXZbmJTeYxWvWqp72ki5NlFG1c5yutKnZ0Pck
/4HgFR/mnln6addxArird13Oa6L1/qhffgKSaulTe4Sn99gq0D8e4Sb/KgvbQdI0NAD9sNJ/2556
TtCtJb8Bh/TZujlyeC1/42IgKKSKCqPIF79sM2swHKfCvw6hFqN2OQeFJwYJs0hM3nftv2g+bJUB
R+V+OYaJkNVirQU3loOPIszf+VGGTlKZDbRKj6rlO7GYy55SYXkrkeuLlIrY9Ja1REmsUxALIPm6
pLgd2eurz55CXjQhTMd+L3GSS/44dQwRUTHgx6hzDoroEaH4YUjU5PEqZrGEy+H9MUtcxSc5f2O3
9mIncIiobzsJb+a+7oxdMSIs29iklkc7ZYafJuRo6EYdV82WxSGi7qqDAcFd15QiEI29UQNN24Mb
U+f/cTj5GPtj9GtiUX7IZMmJSvy9UkknCIiJY/3+R9W+8bZNpoE8QFYgwtYehwRogd4FhlnUVfXg
RC7p7+TaGDJYJhygeih7CSCGboJlWLm/tsn/GTBREf7jbpx5XT1IcBGLFS2vzpyc412LwW7rzXPh
8yiJaAEnX2uUCH5gfWuoqKqsTCCD7qQTCslPcUgoSVYIjRvd7xh3q7SmHlX4kfNHY2jxrmr11ZrT
Iu8PDv4X28go91pYLvVQmDsAGeHWPiLK75o062vFfK9J6MqXdD+m1PysysVTotVgHLT6DNz78AhA
3tsk8E8ac4DGCU/cHNXtdcUiHF2JUvaH1VJQoEeIuCWj4WI+m1Ch4R5S9mUEQE/PaJiZzQqGed0W
Kn1eQ+iYq8SFWmvSnAG19IzwmkqP5HpVu2vdrGD0e8POBQVqjpb0wT3rkXPU70c+uzUXVs/TMfQu
T40qknIKfgXrZ+epkzURomrbqUQPoZuH7E9wYMqwwlIePYuJhD2dgVf25CFmLrC4YZ3B83xatY5w
1fWzMbf+USP+5SN/wEtJ/d9DDmRAjX8+ihIxKKBCp/oOCsyn/hejWBTSOf62LQfM5cPZxAEsa4Dy
27iwlBf0VDaHPGgmvaVpInf1241G0MOnSeewHw3bamXjZvujFENCIisQ7Siehg1KQFCK4A3hrIHG
4lXd17K7dbkrhPdsQg8kUNDReC3cSiOKGloZkLPgkSbZnJczasUSSJFpJzlEahsSRowDTNXFULov
iQhrs+m+8MYTmmmC6666MD/UxsGQS/PtRXUygBW8W8Dzdlzx8weh95oYBIQNniJwWsyMiTyeBW22
MT4GSIs291mdKJ9gNF20IryOuP5Af3Agy8fw5Ieh24SbZXdIFxjESC9Fazg+H+8BBAz1/FC6JAId
BXNbDgus0nek9ppYwbLW23DXj3Z/KPzQsFrlTsxYVqwnOKxPG4Y1qPbOg8HFqeJ08UHpX9BrJ5YF
HI9QxiZKc8gvTdD55yVpaZyX0S4cs8zt/S2C2de7xo/D5Jzh4uvXPagEgzSROmc2hBsaMVCppDjr
TPoxlN/DvFc1aWHXLu5x9MwNouhB3aunafGsRIyzdbg3lHIULyjv7e66tarIHLLT3YoJgeUwOU6/
16sLeHcyMa6zdAAldSZKmDzVZ+ILL+tOdV5OoVVreftIARlWGb37yWaR5ni/OhEJWLd7p7zbIsFX
uUxu4/xWz57VySkoSatpN/hOyB2DgEkBbPLeMom3V2SqmgRddbdFNhBZbWNrWBoy5Km2fEi56nCD
L6T5McIC3y2Sd/QVrxK5Qj5U3canzG39w/KIo0LqA09c3G0jxC9OeK8qd2IY/pq/hLfcq5QzPl5p
N1Hx0sgzNsifrPw2WOE8S0TF6XjDJwh1LFU2QAgc4OUuSVqDCFDkpBLBTkMtPtzXGIwd7EW/stTZ
Q8tXyFV1oJtwuNnmGdu4ECtZ+nw68PvRrcQrUrR7PoX2wa8bsuq+bS40TujarSN96TmFPhQJMnTs
oBKppkl383j1kH+qZYs5XnWXsRBp9AGz8wlvYvXXw6ci2o3j3CmeiNbKu83M8h29xUN04U4Znkte
aciML2ffonzcHqapOGkuNyVSSbVRjKH/wqr+gJPvgmVDhXa0+QhM2WpDSKM7w9b3eAa9dt1mRf38
7hIEHl7d7Jnjco+CSArqJU/UDu0OHGp5pIXDflPJ+dAIolgU74HN15GB2dqYEIC4eLIx39jrYiyZ
pssvl8H4DuobkPU2vg2Lvbg2Y/VulcNjgqVAKTR3YMMgmFmP1TWAxzyjXa2I+YtKBqkCuw1DOdxG
8lxLQc2b9V1cPfRwDNpzVNoDuVSjbwHzHg9SsJ3m81xgZ7DVQRpEYjU9+OT9paRBqyK+HLyGR65k
ukLgei221bhj5fOYjK/THf9+yiNrIhMwl9mP2CUklUn5M6k3seJtjxYX+y+KDBAE4UNbIkDyJZFH
ZKV//zwhPM5zEqW4FLv88Aovn2islTx3nDQqOWeKbZemtfbGe+PAMt0L1twcJMhvI4hTEv4PaT1g
AIrFea2bXELJw65dlF7EcWK0F9Iv7jT+wdrlj4vscV8eLa0BpckhT4TSRvNIfWUUqq/tIH5+Av2M
Qac4DKSzDbfM46MVQB4LY5KyDWtG2QAi8appCI3A3EQxRRbxhhJuFhrHpyuolTTR5RQALz5DsDrK
jlilhkAA6y7U0ttGbK0MDFgd2l4nkNfj93zD+x1BG8pea4gk4FFH6YaxDh1sO3fMPy4NfFRXtJS/
uVA0JdUb362+8yx2KHr73j9ZQKY8+Gnf7xh+SvuRDYHglUrpyFzxNkcFtvmYr4pUCG3U5hjjeLPT
hevdsc6/GPa0J9koIscvy6XiUlVae6ZOI6aMnV6gEC5Wl81Sng4+PwjwoR+hkfnhbyJmH6Yjnh1E
PyB6Y7ShM+P4XSZzJkMtE/LwdFDGxS0MNp+baKg5paVtAmZzbzl6SWeQ/+mPQI5jtFJrrna+905C
XDTV3OvUrn5o4vRKSP9eK1tCaZ1gt5ndo9Zv4zlc4KB2Rax5sUTGbUaSAtwVn41TvXPZKAoIhiHX
vYTcRYW4J2suVLbKW6jbNjwlMg26rlnZ5L04RU/wBk0V5RrtQqTKN1vo/rU6OCF8+vYZ3z3yB0T2
LmYQPJUhpUtMJXw1sU06qOeyCFmPqIiIuvobhzUHWZCZ+jqUkVYt7AeKl34xYJej+tj9zBzbEbQc
vhPhg4d5P6mynXm+w/hIBEaAabo9lwKuRv2k7L62UmkRKv7M9FWW6Mry1sPL1WAuf/azFIrZ1HV0
EGyV5kTkVggoXUXnVMe9prpUFQrO37DfsZ0qQYKnTEvmPYKthVeWHtQaVGIPX7sSZa9NJJe9mpZC
vsG2xzu4hrQ/bxklhVd4RiAuk4vBq8w3vnckHMSXV+i2A53HpMJohvyZXDHX/Z0T5grgdcIvJ9VR
RDSiRu48HeEaGL6W8UYLotAp69CJesV9rIWYwEJkVLVQX7mSIFUsttwsAv5ZWW7KM3G5RujC1Y7V
DeEGbXvJMK/7PdQ1G61G57Sbr4PwZ30REyvlU5Kgkf5CyuuRl4I/SUxEuqAxkLa6xLZ6V+5Io71g
PU+6R9eJkggv4duhIyt4jSeh517fxxqvgylDUa9vEc+jhU8yX3TrX01L3itrqWVXlxU1S+FQwrPZ
YOtMOhgicqBA/y6lHFpp3YC0JO8hntCMHeVhB7KqcF5PbiWT6mpRQl+jksun3evOXdi7phT3Q529
6K+qCXFlqWFBwc/tCD+RTPYLNOCplfuoNGwJLg7RJpE1JFeEwn06CuIg2wvVj7LVfBpLMgYqtvuu
cr/Mwk8AQQg4r+Qmb5lOO8rQuGs256m315D3r2n0TWYvEi/598zzWY4dGRMUUTZmNr/KPXl+Nm1n
gAgppwKyeZlphzX7BquiUu0efoBvi8CxBrjMokZBD7ziGoAseMY2DnTvBN/Sk+yxv0Q+hkHY9Wre
zykzUAMJMX6/Be8x/AvB+mB6kCRMqqHD006JsjF5PnfXDrV9rkRh8SaNcFhJYjoK2zZh5d4FGwJv
SR0p8KknsZ5UlmJ3XGuQvdm1aN1ghdwGuDdkbRXSzhepUsd8cSvyNmlona8dW7UEDpHxr8MbUP4+
uT/A/pjXbdyXsyFdqVS+b862a9sHYzGDFVaJN7xWJRLaGvwlU3z5YPfSHZluOLB40kOjzYu8Sqon
nvBHncuAg8Owuy+HlmNZ8ggmNF7KZMCOsEFrG789jX/jxG98RmwjhhiqNZcoc/oyMG/kS0eVv5QN
YPHD3hB3v4EHmfHkp9/UhYD+r18hMp4hsRX1lJc8argAOYOxzLPLes9vqwSY+KBfaiJU0pBem9Kz
3R3EzZ4JhktRrYRvY7FzCoSoZJ42N33Fw7zEgwMK4ng6unb7nToGCsSUVK907RAElgnbBGYKg+wj
kac8gWgsm0llAAOvXhQ5WyRvafUEmDuqx22LJrARNaF6Grl8tAQXkx8ltnAgz0K7uVyhroUMbBFb
Q2Fd6bBgJG8xyY1hWcX8NI0egZBexX8sVxXpXa+Wm2nJs57kFaPyKN5mu79GbLaPtlRLCukNg0Vt
ZfNqLMCgQ60FbBBYITI43FXLBk2/gO6uNacpktSifyQUASa9l0GGuyWRK04JuK4/bhjvqSs+KMw7
hcVud8gdzwA3zytpamw6y6EEqsRmB5kwjEsLzTrw1nG2imdIB63xJBMrYRhyC6GeUX6SFs6KnUSm
8pIcGei8F6FNeuN+Bx5xV05oPWcJcj31Vx5rW0K2OAyHdQpiOPzdnRkUiwNs0mAsotEjH5x3IMLv
GtItRt/EYcSmSZ6O5DgU3hQlwUVjRZ11vhVSivKoye/DjjxoRvn6x7wCgD/a+8KFHumYKpOFKbW8
prpTDlvpbJ4uXVgu1GO3Frwd92XrrGiU4bpPBJLQzaVKJQ8q6egFcag9Sdlvuc+MVuoFHFXM0nfN
dpNwl6l23oMJRVWGCXnaxdvWVBpC1UgYmW2+HMg7DNjGZL5Xl95YAuM/qJBOl0j4cZQ8BTmh6GOT
XHhuNrtFkSyYfmkwwnLbSikqKHjGAbJn5fciXnfqDHaMvsAsuLi7Y9VhfFpiy9SO3QEF61+cteT9
V+uFm7UVt6xozLe7Gg9Skb0c8Rp3DM1Ob9vrHJsmDFwikyCaLgBQp9f1cEVWCc8atiRoJu4p8ZEd
VDE0WaomWsI6U3ZHNjf5UCSN7kGEaYdHCfg55cmlpD/5n/oy4jI4vevdFfdktCWgJKBViGvZI4FD
dbRpM6DpyFf84mt7HF9OaxFs1CSymDWmfs8I0mbDaEH2QMhzSX1vMrRjAqvu9c0WhA3p4cqkvcCw
y8zxPNY1OP11+o3+XbZDgedrXwGh8utzqhY9WVlXYUqvBJ88/QPps9WMn8GavhiL/E7YFsrjfTdQ
bzwYTLbbN42LibwO1HBTgZOva82P4pTcCi7s1h+AYv9HWYPxbdgu9zeCn4rRqlSWJDYOeKQYOR5c
n4cDLDD2p5rOv7mI6MUzc/mFWd5p0vFRIkmQxiKPMipoIMBtc+k0SMK56LymLD64OgJybOhz7BHw
07FYoVrZtm2m8aw81RbDof6pTk63jHEcQ7eQxzyfBSQ0BZPHvE2ntnHjIsxSlk0T4W9iR31sBZUD
muGg40+TeffqnBHv0n0Lh4Us1KXH4zHrY7Dx+9Uj/NY3KktS92prELRFe9b7y0sNbw7Sb4vFP5gM
p/ycBO+/TSeQqlkA/fQrB3e2SaeM51317P3Je4v4Eb9E1Ru4A4didKRh0515r7z9fu6Qk+HaDHTs
uZt9B+5q+TP7bLkquyBau1RDASZK4Oc6xYMa8Vc9XU/1JPxqtZBOOyWrlO18tAA8pEoMJD3BZ2xo
s0sTNOeVF10MryyfahtqYOKUp1QitcT4GajtnVD6Iij7rr5zEu8xMVGv4m0OgLNSYTMtOX0nd70R
cJIUY5sFcDUVT63sKFQcGWbRON7TAG5Br10sX89G4jAuhCDNzfG0C8ndDEP6HWnokd3MXD4zH5Kg
9n/Cmy93tP5U1cGVrKA5YeXZIDERAVo9WDk0mpE7oOkPaIAaXXkr63YakJkmkt6vgNXALIBhURQz
JfJjFIYrZonzRbc9DknRihFkORLVawvIqoFIxRjl5toGqTQAbTL4uPiZit/V9W/WUjTXDDcOMiOl
wGLoX4yjqvT+Am9q4qstzNLwV7v4SD06VXHJSxw8DuI5AQCXg9KMMX9slEl8nDHJEakHBhAdSs4c
43HYAZ6NUtmXQZHgOp5WFnx/+jcIFLlUKFYTfUIv1K8N8qEsxrJw8GhOS2LlZbQwXPdM5p/nIGfE
C7L5cA+o1bRFdDdwnlK54tPFSIcyZt8PR/00lco/bLeLy+3YbdbdFxSsAYs/x7Bj1k4qguH/L+mA
jEd2/OmY1ncSFAt4XKZ7pClPzFZNV2TNCVJXdFSspx8C5s08iyer3s+5bBai8G3IRkqi+JaN2NJL
gj+Umc+gBEW6sdtYxs8qUOnyXK3J8pHQ/N9c5egXMUc5W2c7a8HU3UfM3HFdbybmLhczHN0CtndU
uSHUyYBgSoGZTww4eA8sAmDVTyk/5kteIsm+saa+PSrxfxCpIjri+v2Pqji1jNZQaUrf1xY2GUCQ
ojcc2A5sDbwMgvfsppnLAY13kkrD4XMBmYiFUbzzB/9DYk+zpG+F/MP4FJETzBEEMcnCnGc4R1Uq
Eq9hv/uRqE8MDbqQVPZ9BvPMkxL3K/9yjZ0HnrCFcbya+B/IorufbP4VSljMXVjhJVtyNr3I0kMU
cmd9xlRZ2IQBwjS80KbMHdvtNYx+SsApICY4YGqUGXRlrxS9X74eR7kwc3zQAW8od46x6/tSJOtA
uZpHoYAiXX2/4bybfh18HunqbRkYzlB9CsOQ9+a6jd92WIVjN8Ren/O3JLIaNr97pDlZ0QxwRkC4
hGjqBQqRJLEunbGmp4hZz4IhP6SWkb3qiH/j15bxr6xVl36gVGJI3Nj8GgUSOqnazZJtjJdLxH7r
jnQQNo18HnxGIr6XbmDVhlsp3+eARsGSZOjj1LWAg6E3MFdkL1DuXuXir4zEC8LrX9mvdy0GiaBU
M1RdUUoILQFKFJGhv1IJnEu48m16Pi4GPn2A+A0bW4voM/bmwomsIyLHoJvuqdGOlgkqNZ1hhzVL
FTvv3kT4dlfXnr3J4KAmOq/LfRS496ZrFJ/crKCiKeBHIWcjN8gTlhve6udpbc2vdYDYVp/FkbZr
rV9j0JhbP9RLbJYwPeGws+ZPWsANWGE6PujJGWUESK7sCfQ2r6F8PiHt+bodUgSf6uql/BX1L38b
RXrXfDc0hWXohDm2H4lDCfhUid0GslhQhRwG4fBdDw9bScOlKF7RuJs8gU4RwjapKpMdq5UFTP47
Zhg72vKSD2DF09mrV8vDQ5aN+pwLOfeeqBF0nAxQKINTZTJBWmn2LT9veAxDbV18iZHrce27OfDC
qX+4b+fZZP7I8PkD+/Meylb7OWpvXOEMOM45Zi52IVQ4XLKBvohHTr1L+P4UwUD8tLSQWGXbuKcH
6FPcj/mPunlptusjWOJJZ3J0u71EnEy9V71qtnI61Zd8uXDNUXE5O0Yq7Rm0WlZxJFAFmH/hjYlW
KYOKY6S1DOoeLnj1S2DDc1FV3G0ix81CBbXC7K59SMYwloM6X9fPOqxPYGwzWyJaHymsAEioXV3F
9l9N0VM8sszluKbkY28AP9lGehq0SDAgV5+PyL9X92I2iPZAttA+2aSxpmCon/mSih9Yt8Ck8ta+
b8H2v3KbtuZ1f1TObfszRbjjkAzj9S9TS9BNYklT5sZer6jLV9fEHrmLP1MgH4HWknhcVqgYP1gh
Mj9bgrMujdgxKy20QYcFFTpyWA9TgFuzxeKDnhcEBvZ/2Id2ZQUD3+vYlnKwIO2hdzeIhQgfQE3y
WT/nLqvb03iCGm3WD0oAxqB+f6D7POSyUJz+/+Lpxqd8XvpddwZJoUjQlXYegKKewsT4rv7JZqm6
pRpCODSE8Db5AyzFgoy+xkraiQEahcPOzOcrbTbdK0vtHljU8teCt6ELcHH7aSDHPW3B358RI6OZ
OUwiQAyCeiTBTo8CJxKLWo/465T7uqv8mfZZwZIh4KJibmr6hoOMTN8kWqP8aovjHWVZ3t81DKLj
wRhsR0vB/bRiQR/vIf2FbJRrqqaUYIfOd3nXfVDn56oRw1w8V44aF5ngPvGlwLzQDX0iK8OJ5MNJ
DoriCJAiE3cJEWeDn8zKpzMH27q0vL05Cy2yRwu79t/QkC18IyFiLKBlbsZt+/T2D/AJtt3WsTfY
s8YMIaeDRROBkDZ0XS7SLMS7ET8tN7twembzfIvZIE32uRDcZHKp4gTcaRRiDiQihbAuYqPq7Tz5
QYRziNPHlMCTVtWVAinpVvviYVEuxbo7IeO+3R2kZ2mxo/ZIkiuRyzBt8UTPVewoYT2hKioZRSbW
abGHWMdbWkuYe3QIVyAL3b+Tqbk+lwCkHqGkVE/ZLLkeM7Riz9ihaOWN9t4E0NwuO8QZhFcvKup6
1+dqJJgc8aLnQ2hkzeWN9oQytiF1yRfxHSSPHYUqgpMVuvQ3vCtEA4CelC+BKAV0fkk4R5uWcm7n
p1CU3eAx1Yr/UxC/OFImshOfEDNSC5wLFTfxqiWTBBVR/MGJAkIgDym2Z2Pq2Wd4g8qjJYjenvaI
SX0vqlyxyI7KEgBPaed7x4oPr1CyeGsXQVKk4BLMFBAxeADPIh8/0NINvoIHPe2Sa2dwkm7ES/xw
cJrfDz3IS9CMNr81MezSnyhSvhAYoBDVT3eF0NpvrSCiize2i4hX1Z2bnm8i9byy2WFG1DF9s7RO
4CDBodZDxoOAODv7RU4jtEH0PxWcbyTu+JWQF4A8wsrgFYpyj3iFxOmxfea6dJvvR59mbalgYpIy
hRJaP55dORZJ5/mPI2NujTo6jF3n84C9ACzAxvDeRwxyKXOcDuxghWaSPmQszqSEV1ruZ+mlsDSr
3vuwgNWzePqZ90I6yHGXVx4WdKeKUjL05HehcICKbbrKkGS6HVbTgfLuxT66QAQ7zf0XzK4r9EkS
VMR4hbnJX8YGJ8mzEz0huuxuLz+YM1SXSw0MspzKOgNWEv3Q6WjVWqd9aY4dkK2VUByzG4a1G73r
svk6IESlmjTh5jAs9ogYgmFoGhMojfcO9rYw85r/bcAHfw/dStBd0bUhTSXBSCcqmtmja38aZ1Pu
mZmWwGgJCgJaUo07NOskhzPsPZde3AtMWVtO5s+Hx8OltaouXtoDZp8CZLrmn3h2CDAIHxnCzXW0
CmJYtlsc/NDjr4qdmBpYIdx9UJ+LyKk4hld1YbiqtWF79TtS6eKlXL70CA1MeaazaBjS4i7FxYc1
gFCKrLtDVqFgOoBfuyNFYsakxJmEIQIjpkd3l1yp5VYagDY9mmmK7Ve4u/OmSAmSiCJtizjz/2S6
c7duTUM2NkqDEGyKP6nxFdz7RbCIDzKB83k8/bylxb7mlUl+Oz1ZVuGaHTVQLv7ZhmNsTT1jHpYM
R3hgnr8mFkVvKcuFkTIcbD4d9wZVfANHrxtfjnWrG3+of990ib/gbm9Rp7PDUvuNAAA38dh4Aw+e
FbtB2mpOHztDAr55xAQ+D7iaNkRvYFZeMHxJ18XmzzXCAnuM8zPbPHgc9Ee+ZyIBo3DDVDpzNzxr
VxjSI8kOqMsTOKCbE6SqMzvA166xuTuwUs7FX2SQkLj+X4utrvjriXFJ4Z6ed08MyWtLSGsh/YJk
/v/ysr2b6FqJE9ZqDk7fJEVRq0meEqzg11kQQK9a0vzDIhqs5vR25fctVRaD5IoTsNfp4FWfBCcS
qB2uTvMlresdxeO/lL2k5Z19pSELi96oNOJaYc1jAJEOEmKTACROnbNFyraXV60GK/RMcwEOd9/v
DKwt2mlpifYd38CxzIdDBQ2N0CjQFRcaeFTPmVg8GP3FkIt9HrcRauSnaEevROixGirABxVi1mhI
2vC5uWR2Pphvsn00AVBFp72WA+OEJu/FPD5f3OvjJBgslnl0UbrulBfuGn6vhd46XUUoCrAEZ13L
fiUWcuGyKE8bGHQVjQ6IA5wPOAAxYjuQPACG50EAtdVMNHUQY/TscMqcZQ0treoRgeCLxMIB971z
iPXbF2qZPLUSj4UpW7fXtx78vPXndeLVb8l02U0Av0cFV4BHV0wf88DHRpyDOeZ5UvXiXjbfk7j/
wT83kdfecMT/l3p/o7jLKWDT5WwiBnOsupEia+m+3JBYoSKO84NJkp4+qdJygB+P8HSzz9rZ/7pQ
8pwo4vc+GeyFTbHgHbFfWPX7m3Whs2FQaUKFf/ZsuZyKVHDA6NKsqulGx1UK2qC/PCn1yemprJcA
bAIfLyy1/FBfVEIXKRKX21LU20tTm+1rwo98JiUZvE8J72JQ4d0tD3CNUqwSmkD1+iyrrIpa9wh6
KfsvUoqj2ObUeQQXgU3njJhDJMrrsXlMMxI+oABv+5bmMKZ2RrLyPPsccRYQYk0xsJiK5EuPGC8F
ll/lzEIhpO0yLofjMnXpgVl3D5YSWE5H8J3/9VT9vkd0YhfPJyce9OQFZht+zbZ5ZnjWflEH19y7
cJ8VnyRqaKuFsn20ywvGcJmF+DCIRfLxyx+QzSUO5iWFEd/2v9Vsb1B7OlouLGTV0BIJ622RnofE
FkVk+0kt/+a2Xq5Jxb/x/RUU5VU2hYx8FP4X0xVwLQTKWD6ZEFUDJrtoFX8Xej+JsXsCkumbl1qO
tGq8iiZCijzM+UHr1tAZ7QAVanx3lBtl8/chH1sxDbivuk5vx01IoXYILaqhfDehvcIUh4pNuuku
0JzkDVJfd70d4oxcV/KUNgCmfSTUyGVeyxQ7FKnJbZDwv4NpnLEBl9ybjvqGWYiBblje0HTZo9rs
q/U4nkqxmFnZU9XgEfJ+16yYhvUGhTecO1JpZinju5b4ODhN2BKsAbt+AjU1DQ3pgvYVHBFCxK+c
AQsqmtDds002PX8Q4n8WtfeQvMhOpWuUFZw/5FP3I0BG7dQ8HFMaEOtdtfwr4EKLS64hGG/FkNUw
pypvxPK941E7ltaB4a0ucJeB1gmfs5v97dx3lxWhnqIHFicCfdgXBZNJZHJaa/4tVMJiQhqJ4/0a
8nsw/278r5AzzaeJQbOmXl9DDnmhp6Y25vCvKkpQeIXo0RtjNkml4aujIaGw8U+eu6EH3k8VxOXB
1EkEzWTpxAlxUtgu+4mpLVrnygDkF+hnhsk2UMGuCSqZddggam6bGwYe48NXWVqMnn80tUXFBJLY
RU0ctSfqFepNWDS/8S3wRjAKbYhgS4jb5gyUtALuAmyc7/QZROWyDVP8UsNdYw3daiLQCtDO6s7K
S02yTGhsuf5dfSjkoBhWWakfglS5Q+X0sR0dKe6R601L5CBKOIundDtTrPsYZW2wdAJJBEPjytat
mQar0hlDNIMhqgmNqjkyPWYcLOFNr14MtVbv+yIQejr+ykjw71ma4cflPNBGjMAdLWe/0E60iVhn
3rZWqPInX/c84ybGFtxs7oWWmZ7vSecz01ohBgCwSWz0H4NF1clLtv9gknfhMf//J2cV7wIBNzJt
SD7LVhQFr8f6gyyYb4PdxiyshBDHf0wOMgFNkyFX3G+bpmXHiyDdkFryIAXMVWw27s/UdBAu3CcD
QK0tb08osRcbA+/h74U3h8P+lQCq3tN+zNUMUTbHXaOQldoUtfOLmca1NXy9hK2xI/iicb7oS1qT
WnmwYEQht0SoDxZw/3yZ6vQ+AvX4w0KHtXzCoJoh8PD0R0NR/2h9NJHipx8L25hBAS4QIxn13o+m
iHPgxGBrgUrGZ2SHr5aPTzzZ2G+k0DXHTRXzB7Qk+5XyTUeVl2WraZxr/gHWWbOFWEnSPT7FewnE
PN3j8yvKJx9l7P3Oivfl6ofz5S3hBhXt/z7UPnO82+VgYG3i3xpLJ0iVVJAemzhmSuZ0xr6toP90
MMuANiNZsxSAUauAxD45W9KZKRXGT8FQV+KU5O6QChG6L4+unjcYs1ZKnJRYe27BgMlOWSDvZji9
ex66Ut6giAVl9IYVH3kwp0QNcmlAL/BhQTaP4i4PMZwXvn5jwO0ZKwiTg2bQSPTUJjK6s5aFxoCq
njjfWtyEdil8aXdnihhuwldRgMhWoCTIZhIkLTRItrTm2wqvUTxzzzvo26s0LSA418XUKiXYgCEI
sylQ5DVbCyavtg/vqE8yPKtOkRSMCY4ln+2504tBHoNuobnoAnzj55tqDNY00kEF9jFjb9dLGvhw
cuHh2Pse4B/VuRmH0qPpH0t+j/gsL4p0cQTu8Zioc2EuFl+jhDkUo4YRcmcybYcHrIPlS1MnRZkY
+LuJ7swZsX2y7G1ZvGaiSnlXdSTm/6zF9f0pbAjgMl51IlpW5/SDS48L+iS6tg+eGgsBYIFRgIPX
08DtpnLDIkLM4yeM0VfG1dDZVXltHOQYkvnAZpADmVpk0sXht5VNSL0FTZiEPyyeOQnfwJMGmVJP
5xCo/TuXOp/WBlL8wMb5mCSKTgH5MzB/bAKryECa3gUh1P9oWns26/BcyQ8uM8fTPrucyRMJsVJ/
4r8+9jtSMM4SSBwCYvhVljLHgwPARAtG3LUfwXLVCqeOuNaGMMMFhg2LNgmNhdmr4ZuE1nf/n9CQ
sz11CPD/rRSK90LDxl53KB42NgD0NAf7yDdQUegp2F3CdLIsT0uoyPvqmCDYaxWjRSZf+ZQYkk9y
v+nn6qjborw5/fGhF9Mv1CBZfseunhN+RHVMJ+js/7pCqrMytnAofzvi3ZOXw4R82WWKo522LBgY
rUtndUK+xfF+qNX+X1KHjxUplhbHFMlXnQDF1MWdaFjEDcdEyO9t5y3/l4O8DJLPjPNZADPL2ALj
sgNxhfV1nIhEoj52jPSDOYrZsAM9Dl+3DquormBlCSqILR1g757jk1y7zYmh+yG6RGhAUE1bOo2O
ZVb8e0FCiMYZAgBBNBoP3g65Hqq+t2RtQ8dK1mKU/tvtkAv89JCabfb428HgbJ+yEKHBlQXJjwCJ
diqx/fE4VNfiWinb89zBDRmvrvgqDo2/coIhFVD88vvavlWEwGcS3L6YNn6TPuBgEgdGvC0lV1yG
GhANqO4Ikj4yjxAPUl5pu/znULWuON7WMyVx2G9soKf1PPrKZ3yPKj7jTc+/mApdyJkSOGHKTol9
f8CzZIew8Be27O3Bg88GBisZ3h1cqhgvxPb6kFs55Cgn2phLAqV5rB8CZT/sv1tgxNdv6/cPiLjX
30jvYT5afrmic8CSCuNGuIoMHeMACL5xZvO+asA4sBZDkreuDL6aERFfC4LUjTtacpc4aZOIIJSF
a3huBG6W+cfMncwjpDgzjv6+HHLRU14bQFctDIDgjPnaAii/KGXbTo2Ei6CtOKDeDGBW7UDPfVDr
OsmKviSBCn8/tyYgXtte1ik8pz3piU4YEnIgFDouz7+NE52dEnwtslxMzJZ5QIDYKTAgS2TqjBER
OBa9LN67YUUuR94AdJsIKzevjLQC3usQwQqhmPcAHPQrwFDfNsARe1v9++nkasGwFspxK0mpDmZ2
Rr1on/U0WgsQoAQPbosXRC4l/wiRaJF5YFZ/u7rpA6C6oo7rgBfa21ALaQUEv0lbN7gAed99VeSz
sStl6m9E+vB7RU5hYw9ITFpdfuObjs8Kuocb3Kx8OaG1cg3Vo6Pp6WLgKZfL2MsgUgkWEosqEikS
Qqyhgmrx7siS4DI7eiYjPqQCcVU8ygtWIgTLwtSTuK8lPRFp923PCFXD9sMkz7UG+S3X/ALjEAl1
Uug+XGRpRKmucCW1U+/obryemwzFZ9cjmX30/zUU45I7DFa7zr8FadWKvlOPXNIRWDWpocrEjtnX
gQ2bQGpyD8neT7a3X4OnW/D7bIJEFAz3XwX5qcEt/fkDWqKOgsesDEwmkmGA7NXIwhZvZyeUKLOZ
wK8zecg3w1i0ogkvurDQaAj07S0cmoFL+QuTt3eGsWEiz/grBZ/jD1bWFhf7F0Y8VuC/J/7GQMC7
f3sUfmInIRYXpp35P7oby6W+Y/hUUmggIjCh14bGiZuEcZ+O/0guL02zHMRI8gjR4ZT64Lz/nwHo
G3lFGEeQyB+J2FlxMezdNRg1kjNDBKYhGQrXVD0HTqbvROH4jUBTegQAsoJjPIMZHtxp3EZVmIVC
xCuN/6TN0+Wz0HlsQqJ8xywidZt5IBTE16mOTED+xrKs3lGlUWtsd9WMqI7dnZckRGjcFTcN19WU
vBiKeeQzROOABbtOI2yyOKIZsrqH5tqJpSY33gKzeQbEYJvgU2XYDFqrZ6XC0DB6tgnL5vVBhmbD
iI17k4btDM63O+V29yW+s5wn5YjOMy1QyUuwA3thREndwql00A8nzXusX/c6TRNk35OCBgbVFovd
p2iEFwW5qfQtQknRWptgq+9yB86U/SmSpA6iNy9aYtAaHFrqbrGsNE+158gcRtBWU+yjv0FJktT8
087ZLaQvyGEtKvQ+aRxCVfVtnvei1cNv8yF+9SJo8QfTkmM1xkC5zEqsbVJjE2h0uLO0qe+l9cvZ
yxbcu8NCaXdg95nv4Zu0M2xxsQmapshSwgOlX7hKRGT5cu/dmhluYhX2FHAfVg52tSP6Rep0rxb7
jSZ4f78BAs8XFcB00QRWw9HHo9RMBbxHOwf1jS5qUoIQqhtU4YkAuIse9mJvOAh5Gd1ZtmZ3NSrv
Xo1K3R/VBvKTCcexmEWPCEx4XcOy9J/6Lz+QJEUcbo3zGmSj+4YGW/5Mpok2QH7KKnJswuM/Cd2w
24iAa/AhE8j1x2InPA9siseHbn6LUYv4vNcd/kzWq8QqxG6KpaSIg81hwR0r/VgPhboNwFOVauAZ
eR/1i7oGYkemTrL5Jak8WkZPydGjXWvqSU2kp6E+V/Vyv6tqFvZ2gL/zOJSWXHr3OxqIyKFvfk02
4s6a2ixJzSOt4gnrrV0v3e2kAOO4rco7dfkvKK1AexK6fVOCofIpzEgdtDXiXBVbZa1MrDqPnl+o
eblDhXBIjiP5mJlXZnR9+VnrXW80DoPrLum3P0o26dV5kPebllVj/2BvUB3ZoTmIgDgY34sYj8/a
X9bn8Wp2LgDWxi2Y69zDY2iGtkphG9AqPeGzDdYKj1wTaFKixW46j+P9s9ZfCgo/T8+3oHmclZ4e
3G+GZ0QWU9LCroNr8/FAijDWumcho/tQyY5SJtJb5xtAdlDIs/J6hljMdZs3uNbz9+YNiLwBuKvN
bsHXhinAIxmD9Rf0cVzCK3qns07FzWuCvR7n546dlSIt5qhwS2YcNwTCLy9hY5y0qXWkdYjD2Fks
99K9kCUfv5r0QB+QaWrd+3xYcI24enmhWOkoOM1Dfap+3Owb0OHl3+othA6G8WT3vBymxFyoE/TA
5XpbA1fQV1O7oPLbGEbavpoagl1dUbz1QE+jayL7lhGlGFv0x+J3Hw+mQA0IKWo/DseJk6IOyXYB
I7sFd2UXiGcsYq8uAp4N0jmawhYUZFuUz+VLlUBzo6pD4gRraY9dXMgXQI90M6d+m4y341RZbWJL
JkzsEFupQR0VLo2aTUUhR7vxoEgcokaLAnFaGK0X+ZyztptxxXXfe8fAGwT4yu7PYFildykWeE1t
Pygpjtm+7GdAhujXsPlwGw12uhv9fStGPhB3W9NboS3964xdnKKBXdgRN0C8Feo59J25h4KmIjdW
TG+Pxo5Ht/mihwJDH2IFW6NNygRuMT7M5V2PX/Ul0i4ihsmOuT4xnyzm0p3jE6ljZrnrXyvhyHY+
feMWRz8VSXDZE80+EijikmL25n6L+VmX9MiNz7LyW97U1RzYbZiJtcIaqXnCjCAWI/crKikGk4Da
uZ57JK7eCEZ7TFPVsVJ0EK61zYDg7syERg33589bnttscbTEeMGvLO5HDPYB4O0es7MViGUnHtjJ
PrPS7DYaTRdWNvUtrZ3AazF3jwF937uE3ve9yIqu7Asa25eunXlA+1wqzevpUHevQkupLQW7DvJk
17uTT4GIVjxRoFTfQRzcFm2Y5jaodLpSmi0rMZHd9RNa4L7JhSTIYKTqNj6gS49KEPgB1fTobol2
BdIajTCR7qQoJUXQxtwj6wW1MzNzSYBHnI9fuFngHD5H/UE7bBwr2VdqkFcqP18VQkEBXEeJvSfy
kOcUO/DlFJBYeD4lkgnVoT+JkOEjGJl209gi/VkA0OgSVNPOzADdcuGm9GzcMrcU27EfZLYzU7h6
jVUbhOFpQxb3ZezKCoDGW16YJ65qlIwx2cH4idlJWMfQ+hcu4qkEUmUiRcUkLj+70MDaYtl1WFBg
ITXvpVsE7p3Mh4hohrhQhTJTUidpveKkzNJmis7BxcFKCtiw9kmrgFVmxJmpUgBMCRebBoKNf/+G
hP1IUhhzeGtoMgnx9IstiNNzCyrEmM2yN7qLNjBdYRb7ykJWwpfYpOk+hJ2fXdIUmjG0JyJFVSQZ
yDc3dzSsPwosJ4BSOm2RNWQJkXig6mAiQMO7hib8Ve4n36v5cHCjTr4XQIrWWGE9QhGeM6bCEPMT
8T0VGesC+5RqOgKR2w8lXhw0Kr4BcgHTJFmUJiTl4kf6v2+KHYOo5vOgxW9A3SsyD8zFw4N9KtHD
bXzM43UAgjbql9Rs+TlSnWCKcITFLezwZOllUrt20UdPM30sjKSlQZ39ianK2ATXA+DkrI1IbzYf
gvB4znKUMYpUV4MMdslpl4tpnfq4pYyEzC0+6bpOmCQcVFLHOaYu+EUMD3W9JR3ToSU/WEIZul64
/bFrY5vzzrlJzVv3K6feE2cEovPZSg0YYO5pSxegAO2Ajd7g5RiZbRLLoiZOg8yAz+VvfODJSI7d
xhJ3WZaMr6epOWk90UCE9ZMPeOnPlsTXYUBlpWNtJ2t1Oldr0xB4y0nTOJammDQOqrHt7yKYm5aV
2R6ZUZY90rrB3omttZ/GwNWD42Vhp9FUL6FaKLvl69Jo+T2btahUmonOOjdYQKoWTPKbp4HumPGs
PlRYZ/zXvxR4d0xuPuykSGfGGIJBR0Eqp+iQczsYHBjD6e8MjCk9qPx8UBInm3r0p0LsdKH+yKvO
/F9ntx+iWIr8dlPy7FNix5mgmXG+SLRNuj7kL7Dc+CmaE45EaeA5PN9ym6zYw5iDA0V26ff3Z2Tx
w6BeeyxK2Ok0Zh4hEQrxAxkvfjmwzFlU8pAi+w+wErvwlWrLMrKhlNowfdeMcTpnj+Rois9m4AtO
bKLB53xFHG1yieho3ofx3lEUfgN3/Ji5abFfnHuZz5AkRRpO21EGwL9hqrqSJUg5SF1Hp2KmNHPv
h1GXPCnCruhiLJzuRc3kaRtt4LMW+jnH9s4x2Wfw28bF3npjMdS+BYN/UKVSnAIYmFdGjknH2Myx
8yKHkfajayk3k75BkuuC0/xgWFfXjiOTK8x/aGHQCi5mXAANEcSIZtHgq10Qgn/SkKv2kRDVUwDj
pWaPFQgjjWrYlAHwIckObQsPi9XQa9VVxPfCH+7WSAOA5/CMPj3fX/ckE07jbKvREfK7Fj1mba0J
vB0FFOC72sBCKu26dtlW10KDGTT0Evpz7fkP7rcRZ0yOIO7sXed2Jkl8c3bqSb9eYvz9lZu1Bsrs
1QzfYzwZGsvJhhXgXF6F9bPfT2RLWY6BML8jVj4PpfX4TL9xHfqZUDwkYWaekX+cpQvdm32Lvmww
qaSDI9nd+FWqJSVzi9flA5KdpPmSEHLlO7VCdvKXrWE2bPvbsFkzuH5OpEiUhzjiAWFSOwiK0Foi
UaudIY/xDhLjc/6U1MX5bON6IgXSeLQMXPcujWf/4KnJzAzS9gvzPln22NGsRh1Zo67mldukIDEC
WwydAVSxQHgwvQlh58gdyvV2k2wwQ0lnz3zyq4j/E4bOmAUeurSNtW+H08AsBtMGmPcnJgJYjhoO
HTVCjBbgF4y3aInXnFD49Lj4IZuiuJcjgVBU8SxMvlIHtODEXu9SdEjWVfim1G78OqY4XiZduhvY
oQ7NBGkyPgVQ1ncOaVpNje4pk7VoDPm4y0QmMmPfNOQ0kQ2SZVZoWtL/3uJm1Kad7t/dgLdAHd0B
/FvRcHn5Pr0ghP/XzWGVe92M3/YTroJUkd+r7yfgvz1n8mAOSuWg2m+ggOfYlT3C5JbVPoV/EJLC
T23PO0Wx4eTrPcuDGIK3RdNC4S8JRZ9E+QtU0IQad2Y5QVRHR5JUB1BBGzEe/7YE21HrQjOVBTIF
uSuznwyLEL4/0QPd9joDCOaJBkqhPCcbLRPbXjMx/8KtMoWRZ7a2MR1WE9dDzUf7fnGJL3B8rIeC
7UCHofWADJU5WO+mSOsO3bz5ASvBTIdX3b1Z7wxDsRI7FtMZO0X14awIu1oBUqYXKqfK6nnVIF+A
L3p9SUbGm5QaVPn8+ghmdvdceMgIX7D1SWroXRSm88R0RqFQJY1hmHb9j5drxAnDC0KE7oRR9qc3
0Az7psoMRy+qwQD9AQSf/SnqriHOKrXUZ2Hc82aJY/nZUi860hejYBPegvyigTxcnQYQDVTLrNZ3
HUD55loZ/n42w1rqHS2K8uUb3WlX8Q6LbsthwdZJ6aLR+ZnTh4yfWMnRIf09gLmDuzAePIavyOZv
aMnw/7FQdeNh2dn/Zhkw32ZcayF+Usl8Ht4qu4TMKBg5EBvyUuQTwF9XUpNXikGlNtS0H8RKoYZs
H9qEO6Avw2Mlg1ELNjWoluiZae4XJXR2oyWdzmHb1D1n4r2RJVPFtRHzxAFWEgd3QwAY4TDqdhnK
lZ5vLt9BUG0w/BHYQ2aNfEeb1IaIWBmeSWAHoj50KOJle0ocd0AlfhbgZGOlq3gDs74WkKdHeU4G
xsXbDwA5WP5+ubzi4mTHz/ORMymuO7AS06Wmj0DTvWrDd2IZfJ83ikySCvcKynAVMxCjiEfRpj+K
GC3YKz4IB2x1w1o4hvg9SJsKYNwbHU6j0+WAUC03wDa3K+V3U7Vwz570krSkpJvNhnCK2HJhccFt
6AKcTW9zsTWWznMe/uWNem0gUVEy/eW24ZPTxJI5Co3CfQb24kkUI5YvRKxOVpLGAy4c/DplEuZi
ODrun5bSIXps2ESHs2KAd2TXbHjGX7RCGzeYV7EM7SUIGDe6sOfgZBYFhrA0r5LwA4AZ6V93LTaU
wXOLjqdOS4J4rZyrW2My/sxzgciMd7Fez5ESsOY2ogQ99nkTcyzBxe3b1+qHGLd/C3i7nSVLuhCh
l2R5QrkS+ENrr6htcgINeDl7CzavLap8tuXxbEu8uV9UMcZguPMya9IVjj4TfKiXqHNATDn/TFRB
4gD7jhpegcHzbW5mPpnlHEBBv2umKHToUyA2U0e/jsqqbjFI/yx+MJx+40pf6qZJ4sBakpVEv4AP
mHDxdzpQNaE2LC9R8qX4vIwaLghXEbibXj5OnrzapIkGTgY/KYJbsyziLWuQGJcbh5MwA0yABKB7
vTyG2gE6SvPmMxUJmY5RdNYW0x86R8iXbWg1qKcLhikfnYzDGkyjtkysaOWW7FCls3hL0pZ9rFop
jSFYUwq4SG/aVPHftpNMb6hF4LHPeMq6X3f1xfqLvch1fSlXLAO7aTcsP3zHAd2b42QFLV10Hgnk
J30o+v8PJJAxzvNA/0j9jXw2oisqQXctLufKnPX6aeogdxn16V5m4yZdIO1mjggmrskUGNlJbYkQ
kUz7KQ6Gh7V9CPm76ReypWJr4enSDCKrXWSLSVKZRpkqXx7lcNucKEAv3PaQfpprzjJC+j7osVly
GR6CmVqPMA0tlLi1Qua8r2BQcYQcXNtjhqcfc2yzq+dvAnXvxMwKdswvmKzk6iQum2EZ5Z7bHYE9
cGzThwuP0o5lyc4P8rO/ASvO95jnX5PXAmtVX4bhm7M+4jZutORsDBOdUUBNlUiJLQKizTHFG0hr
wcz4jzhiPIEFg6Gx7pbBsi6HiP9zr3K3tXXwsl1qTm5fMMIrh5tVCJ67Zf7zNreoBS8IfYaRBy1C
j4Y3TXtShkk8JTz5eu8xDCbeHPS2JEyfdh82L3aP7IaO9cOt42WLBOSDhz/70/qqhcD8XhPVm6Kq
IZliRrTt7X/8BOLywIxTLHIijHtC5db9EWIhWy9rMfp9biUWFF3QznhNu7jvcNlNZE7VbfvitWq4
aAYAUtvhgpNg3YRSHKtIdaCctZ0ZgUHqIM9HWKmAABTzuhCdon/BGfCWwqsioxZWu5PPQ45ldBqn
m3gEa/otqIcL9KtPaKWnfZJkxrtL7g05jfLI5ECr0+9kQU848MMPHvGMg5co5xHgNoi9pdi7vkkE
UYkjVAxQYC/jxHPWQrquKxTfGpsKCcY0501/Ps2WJu6aqKhDTny9Wo8nr4P/Ccs7/EKwYItsKM2R
h+hxmGuu1v+AYSIok5W8Uj+yxcm/aeWzvCFYiDMcYH/+CFv0qQcWSdfQU4GSDkDtr+9VQRZ5fXXz
oKgNLamLuI9GVuHsEfnuGXeG+8TtuqYKk4W8IsULVKAcDdIz74U29OEkwAZKfPYt02T5QlqsHO67
K+Whx14wx7Hl/uiDGhrqYe1YOxZIsYiSEvqc4M/iMf48it34yUOZLmgy3/ozUcWcznQl+4rFLFSE
mPhMzxwSLsFHZxT8QWfXDDS0hYA8dk4GX5XEpqUgFQGTHe/lR5RlPhEwYrVZw7zjZdWpeyImRd2c
YVlLdZTHJxf5qXDGkhDSobOqK//20i2goy4X269fN3+KI0a5y9n4jqEsTYErhtX9vkcD0fmiiZ0D
bgBDcNlrM/cmeiIicAULkNUQXJwhf1RCyWrD/uOjsdyZi+QjqzK+tcrTrTAnRW3UCRzpnB8K/GFc
EjSyQ/OWtBpDv2fNI91f1a3wNX/nIC7V7Y37FSltxCcEmeybHf2VGt4fBMlxdB4Gheq90VKBiSfK
17Cv/DRTLwlSa2OFhmJLy9XFXizviqK52B0WRLEwT2dx/3QdjpUWcGUEXA+AevlIQOtFdtjTf37e
/BWM3NSoCrXNAiRPVkh3Zirt9HFQm26eo4P/1poG/3GRNQcWfrv28CsygDQn+Twi1WOSBII2RqrO
PKOqKs6KUKVRMzLT3hBbLK9ey0SLt4f6hGl5sxiHfP9nIiuTWq7cHOpoqAMrPujwTy07aiC9LlM8
J/oxm4Jt0EzisU7U6AANuBJp/hnhW09doTimb159uObjkn4cu72MedR9ztpIOyfcpFuM0R/GyjOM
linpZn2b9qh4c7ehXWFCrR1r5RmqThr29r03nZB0Xveps7tPXymitxDOWXXxWwV5NCzh3EsGkbM1
n9CSSmQUsY5BWkqsgrB10sUpVkpuz78ToyR+4W+X85bhl/qipyVs2ZKf8aefWKxKtDTamXxMUVmk
0UMG0gVOySi1qkHz25FdP6SFvdfU+ZzwTRsIQ1B+wB+1+RnyHhL0cCJole5QYvMecd2DciAP4Swp
+Ix+LchnYLpo3HPsjji+lCW60ikBciIa2tekvD2b9dPXiMpwpiSMBT1IG6Am+dTDpDnGZxpmuHN5
XERmE0meZ3z7qNVyMlprr1K7wnD12UjF2fYhyecXcWmuJWLs7O0qDw1t6WNM7ufcvK6arywJfjc2
0raZH9TsGLeiVcENevdUMGxFN027rh1mEQ9MJi9P31WhX54IQvJFxOY8LMybOICuZS8mpy0h6uIH
nH+zID5u7GjuRxY9QgoeiFfCG891uJWVmJ7YE8iiT+WRxz+zxsEwBQaMNoKBJTTxai4JX9O2n7H9
KGcvX+WVyhXsOxiTqWy3gjZm8DyM4MmIaT/sB3OZrDviVv9H36LKpa5h9OMiQdUy2VRgghJIeaf6
6Ka4DMBqBcWBJ6bjvCup9PmshQmFQniAzl3ZPR9Ia+C042+RdYhv/488qyFinE1B4t3Z6Ht5WXXI
J//8D6+J5iZoW7h9QXdnzAJA5Nzdy82Ig+1fnwhcXO90YshSuvfGM+WfSg0PAEbi+H17yRoaEgX/
zzKILumB6saT6YLBZSEcUhTr5LLBdqScZTMSwGXDP6MI4ytcC+TsuFvkd90kgCgakF9RuJYZHeUM
dsUQPgWBITERNmAJDyyjgsvEBKSjRoO7O/bIVrk+RiEzyVC9C4cYvTDLi+gRXH0nw6+qqbEd37NA
TrRr1BJXYOjbtt5JWC5lYM0nHd+hys/U+soOf3zn5ecDrahJ7khtgkucaqOfKNZijG4ZYU3g0KPq
HVAncKrOLY3czgYzyWmBzyM9aBREWyfNeNdpEyXcZGaIH6CLECsGSqztfpg93zJznz25EMHNnDw4
IpqtK5z2WN3oq82XNwjH+oIkjqzjJLPhiZg7PBdx7HvlPHcZV2c/Lv6bJOQOzZfk814IKjuKwG0W
5V3IRNsAzcglZYfM3WL7T439VDuDaO4wSGUGEP+mKad99IAmEMYoJsRyPbmTBFEbMcW2VePceOXa
gQqoJIMfcpnbPQO8bul4NbgnelQ5mYSFvG8inQN/4Gb3GFcw+GoOv1mFD4CTjdmYBdCn5imWQdS9
dyimaYueB1CSmidkNt6X8WmTtpYwQR4dvw819cRlCFatH/gjun8HP2VI41A2+bNqISweB3tBX1ET
LnJzDAbYi6iLXfoIKmW8yk2ntCGaUQtLVF/QldHUYYDn6CVcBGl3tFN2mx1RbcavPSGeoFre6t4z
1dWcWAIKsJtRYBkhSfYi0M/RiYm7ppY30pjB1asp7MmYrDPa2AYQgChpErf0vjilYLOYsVoAwiQp
8iASvYqkyanMLJMr8XFd+LjhfzgCOqvdEAIvxyLRUmLAND+0CHIus2duJSGJRJDcIVvXELKI0/Qq
7zMGOPufsUTCmxWyTIC1Gv1zJ+YwIFa89GMefwV3PTy+QyYEq0LGE0HnZO9ICmkyXIN3AB4RtEwk
+hNc7PDY0S8el2QksffIKWVHyUd5vmOe5YXK7rOd6EV0JaSF6QlAW2xHqkWmmb4R2G+sQgWm/91M
42bg+28doUQ5oQDor9aBmrpCh607QLc1TeZfUpDQ7V4jqX9GgCP6Z3HVAwSaXMMT4P1JcGnbPCU7
JC9Q7vSM+z1S1znRqShjjmevxjb5qqiiKxxnybTgOUMWf+yKHg2JX32aWhOxtvDBM7qbheqE72rA
cEswlmQRkq8GakKGCUNLeGSzKGXzcYbOp6DWNPsg6IT1QcU06jr2ElYIw2VwXwuhMa5gWNq8xz8+
qpV9a/cLsnWaTJy7c29nQHpHFR6DvRJqkEtJt2ZcWhMxBKoqXAiLVhD3uZGc3M3iWm6EnoTRO2JI
crLlDWMTJB4r3iu41c8Y1csPQ59Cy7JEC+O20ym0xAzAjH4zWubG9luGKTcErCdC/GP6F+aukFmm
nw8+3tly2vsSeUd9d/fLyGS+G03ivQ0snSW3VuMjHBmQ6ccgxltZnEIb63dkZ8wxjtpN4q247eWL
OD/J/FxJf8Qtxvj7A/YjaRzn4UNvjRqAVMnzzZ60eSMYVLdZcpRYMk6gsFE26Mt2s3kFemfH98q6
BsXRTuXLH71JzuHrjGQExRnDZGR+hC0IM2Ax824mMEju5dS94Z3LQOEu5iQhtT2jbPGh3I9hgVER
9TF1lMvZfjH3IYnVudDWXvVZL+SGx9qZ8MTlqPtWgVt45qS5mK9ewFVTiVrgIpODAtWrmY1Bxz3O
n6i0+1lYD4E9Ndc0iqpIf5LkwPnL2DKpaX2vlSJCY9Rk6scvdfOqd2enNGxlvnzf2sihR7ThptxH
TubRk6gp6f7y671Yudo+XG+ey85so8THjFwNHY1BI6OqXebdtfB13K812VAsIllDEdbqWymPS+WY
I3zWTRs5HPdIMRokFqlsvO3+szfGxDLXYZyn3M9PRE7rZ3f4su0ZVTFjyAVHIDWmg7mdAaGSCiGU
D6m51O6xT8lXdEKMPkNo5NrjxBnaVbyAxb9rSbXr+oJqtIGpxq0OsGN2mplX09HgLlCoYGkp7wp3
n62cdTPofg2l87MvDkGuiTeTLyf4vyfwoXxmWR5bN68lhm/gFMVDh6bzPOt61TyPW+ZIEMvuu7Lh
zoiUNIaGr4w0dGgFCPsU8vux+gy37YHZcloMFmNFYFHNhq42iead6crO0NzlRm6Be2YtQlQHEiha
/Nsj5JQM+zdNyh7GD4iSTpecdhrJynp0iJkdCAUiNlUa8R82D7aj/yQdIdl+HEMYTPFNwWi8C7qc
ifFpnNjaZWlwaXa058ZjTjw9DO3ZkFnz215HDJWGyAn9PACNfgFeIBNCCfgVDBxkvw+sGG+mhxF0
XYY2fTazvFv2OTUZhS5cQcCJ7tgJiXDInVbD0K1kEvbLAt3+6YRARQP+nWLl1UCekZ95IathGMEv
/tHCJNNBcLiFKR11ZJi0I6Z9mLwPcIGHXp4V55EwjhdnEqNKQ9HLqSoEeW5K5gnqJdqRt0MCoZrA
Dq2prkLdpeHMO2B8SeAH1Bf3P+e+yxlOLAAWTX0eTSeDvsRKKZ3zMx1ZnXpu52HPccTK1MUCz4N/
cdCqB3+LucVhbVbTCqaY3r0IcXXpED2cRWs7G93Pkb9+iHvAK9luVHsHM2kUoJ42QEeponwyDD+z
ht9D4GzdhL6vyXQCJFzzWLQPjb6D4vBye5h4/fGAsOTb25nBrQtpgJBf8uV5Nq+14zYPn+BO6qTX
bHr8ijaxva2EaHU9op7uoQSY9nnhR7Xe/425UqE8IoZmUhOaFH6FzYZlwcUFnx9m95QBvrZCLX0c
JgFQX37SuZUZQwFD9MEa7h+zIOEQjjABAMpvWw2E76C/2FiT2bRDwhbKUuIESrMs2IBUVZPpwnMN
PGjGgzB3BXSUpMPa4OvD19LpTyKR1hdWnXvkNEaFlQYeQ/Pw/te5yqd3leu5kNDAJWCOGOYLlrzZ
DFBjH/EXsD1e0NSG3kKcKhfc5+ab94sZD+qElLmW9xdC1OgSa20nP3MfmdJwyfRJsOA3qKPGD7Gn
ggLwZB1UvegQlGRWwQaZzgMzgS0kqTw4iXbX11tac8aV/WpvQWoszRO9w3Dgq/WwrK+Q8hy96MwO
6ffFtgiU8NrKZBNgWOQcwq6QO/Iciw30s4b5ieF0NVMYh4X4XIYCbbGct3gfBPhLl8l1a7Dl/h3j
N0e1sYp2xk8AZPyVcwcIK8ZMuYY5rYmkmVATm+x37Slz0pjN7lXWbcSRDmfIXgpUpbcOFKwY08BB
vhzlKodfpfgVZJYDACl4GiKXxCxSABUBjrOR/AiXE9VLlOOV3bcL8oSso3AjRblT6Nkt6Xu9nYKM
GG26vgzgPoKUuEi+R+sX3XHepkjiVWK1WNrhsfAV69+NmnFkiyBUwVdH8V/pEhK3DL8YxrULIAxB
Pe0NWqViYBGOB3NAY7PsBIOkp6ytw1byzZw4HNzc3Ym3sEY8uOdEndMSXZrmAntdCt/bmyMdljb6
iD6CF6rGdO4JoOq+L8+3dLJDqjBcyVMNLGxhaFday8JthL69pfVnEfXQ30y/Ii0EcmsObw8cd8gk
zByd7fK/s2FWqLeQxdSBTbBVCGC3ryrNUWKQOtnS/MDl0x+jWcqCBut8sy20Wt2VnoqClL5i2Q3E
Yc+3bDcCOAEUKEB0s3gBmLYUGhd4iFRuqZTEfdd+Sv48ceSwQN2aYoD7AZYAYyedTVZQc9S/JGdz
tnSqnIsW5397/5glV/OInUYdUaKxvaiRKJ+nWg1B/28+7G1Lf5bI4dzKE264m9DSb7u8J93vI+2I
Aq3R2FDgCYYsWZtU2e1K5GgLx4xV3y1XPDP6zGs0Lnz7/plVNQPvfCNnDLhM96aATUAsaVZ9vBwl
1W6E5uLDiEay+kiai0uVNfMeiG4CVXsOLt9G8zlyIp4ZrmdTCFgWG1Cqms+skUxmFJ95yunOYJda
xpiAh0b3v5XEGug+zMGhGHIPhMUSLgba0FQFSd+Qj3TG3h4FwHx64P3b3QVoddZMZHCukBEZW54E
aGB1CHJjhRytwNO1WVkGuaQuR5GhsPiDXVDXBCYYEe9dGv4GCNOeXYd+gcjh5MJfgbtXpV++Wo7R
RNpBAUNc0FEwG9xg2UtCiLm459Xd63M6Vi++Vre/KPS1BSkrI60X8P64uZ/KVQW6mZ9NhX4qMcoP
E7P4tDAMyz9BBI85Cvn9KvPlxBO1sZIJv1uGo7/mR8r7FacCrbE8q191tOOsExpPUSp2IOXcC/qZ
5zoM2GA9kk4sisjXol+T+IUCBOEQAEC9J3/KsRyJmPdvCfNYTO4MOvVqBZvPRX9+lvfRKlxDvdKp
l8YWGyDeeo5hThCifG6mtqe1+d0xa7UClj7tHrzjluYxnqy/bFLudN2BMNYOGAOEsX00JmcLrH++
5DXmPbf52n+yO4q205ucDr0WfA0iUbuuiYsVr0BF09wpWZqkI5ZqcLoOR/d3gzoN3RLlyzxSI8X1
DLz2f89zRUgDzQCItDHto43EM9CcJMG6moXCMIPRtLBqE114rfD+ZVIFeLk9+jKM2CaNgLEBaxth
6v9xWyhyleP5TI2Pl3YdLU2aHk4XwChqQP5IscKGSXjaV3/XseQp4JTYFemtqruPQRrQHH+47fkM
KutR11US59aCvD6Rs1WidOhROeRq2kUQoXCz47BdMhEgRR9FlmhdFYDJrBaL9YGfmJ68yKrXtlKO
sE3O7zcZiaC1ziWAQD9pWAec45FX4GRXc6RJxTB/pdUNU2WeBQiVx02XkjvSSclVb6Xqccdhyont
7c5UF2BMZB+86UjN5t+xu6Jl9/rKb2ir0SV7mpEiPzwXxGvokVYWoRZyk5hMH+JSrUKMJuOef293
HNczfdxbENwK8IjjwZmUP11Lj9pzf1qD/9sbXwbgWiwypapJmKk0LmSicwuNttrceBgal9NwFG6y
mOe7eQLbw3RgN61qirJJo5XH8Lz0k9qm3ZUYUjyFsMDvxY6RosK176+QtpPiww4w57Z9ocnm/FWl
+cCKwoNo8RVOxZ3jh/805C2Hyter6U6hT8qM4lkfrtAsu0jTHYwXxpElHQj8MsnoE18eae9jiaqk
Eg5DOhfe+hEzPMbVCgShUHaJqJQry2WOoPBXUfQ94SG7j2tiLOlyOK+ZGBRtQxToJ9z59mKp0EUQ
Gys9XtBaaWkIVeMb9rNoC5f4/tVuOt3WjfSDrpDrNTr3rMezyOxLOgzJPWI27QZMhykecglsD1Ue
kQDiJpQQGHlRh8zZla06W2/gzEAPqQCXVDZtXOBRWGdKUUcV5JYvTsc3DzhfnYAeP/Y/cQ37QuR2
Lqh1NInGLyG13IaVDgOp/nmV1BWRjzjZwjGlMvtdOnfRRT4nl7wMOVcRXiRPLSpRxYeaASbQDUuS
HT6Mra1AOF2DjSMFgm2GkEe0sVq3Y/8CMMdxmfiR39EPnpUNLTOEoARoHIGnqkFCnoSb8tG40hx/
1zTiEYyO5jrOZi3WyROzFeDIbJBiCWGqv7vIPEcVf0DVisCrYWCbcI1dE3SIxzXGwnIMVqV/3RoD
Epzi1BLMFkgFG2O3iijRq+quOo5VNxBYE+RRl034vxSIn6q9HN5AJOxPXsmUupeWACwcdwmjx6Fk
j8j+0IDWILsSeQUl+LIovYnqzlaCza5rvAf4yS47emMXBUw6o/C6osoe4lhmUPjlIlEAlOz0Z+Mp
HtgEZtNFinIIDKKT3Dc63R1cuIMoTCAay5QpuFg44aIc8PMss1vUSSjZup21jReo1WCp616wav/Y
cTPQ6hpPdnlYh1gpphbReZER8nplFFCQOOrQkJJMD2853D76GvdTvc4FBJNqrsKq69NCRYhr4frc
/3MtRYmFKY/D+KXYIRwSPOikVRmeHymJim0GnPQYjeGgw1CuecroCq0K1eRgSLOsvDKqcgvbEejr
uoYUjls+V1ZkZoU7k6bDmizLUTJJDxmwEwo+LGafTiOI0h/hv6aImXwmK43KTSrXKNg4LDRscQ1L
Hfl7IKRz63t54IhwZGxa3FaxulIqR1kpv621FjzI5plUw2vQuhlw2k8YX2qKS4ZLPXFnXX6Lr/bU
QxwuKzpgBrUsYJ95Un5cyto5AGevNq1ouYfHLfNjTccfcUW9MaDdjJIu2HrqF0TLjQWZxwfWtMGq
Fe/ac3d0dQUeetHQBmzJEVI5M0V9nIFoMTIfftA36/+ka89a0kYaGgTb8wkPTbg+XVF+L6oEdSOO
qpoGSubzbhlbLf56H8x+wCc6mOhFYCypjywe86OOGVFGkjsEEcJHJVzNcAwE2cJAZ2wGoFEryNu1
HDRxG3+ZskDk8duqxGlmIFqu0ETySdJ4IIl0Zyb6hAOC0pExtvfJ+veTQkhSLEIJbMKDt6FY1fIV
Mts8sRHnMp+GGVxVs2tT5OYSyQ0EDlf8lBAZiU5N7pnLnCKaCN+dYlorcy37DfiOkwpSbHY+2+ZT
g4ja6ZTw6e37doRjqPV6tdvbwdDL71LpOLeNPsGr4SPGBvgqE65mAPnSJLglPsGXS6O6q6Sh+Fsr
57DgkrjLierjyn3r7ddAjGDpBvOMN3Zk4AV4CM7gnS99QmS8Myn/IQTaY06O2569JLzsUyd3W4n9
cDQnmWBCivA8LH+X22eWacFWb8tljoCXbMHBFXrcrxWUEFX8qbG5GgYKVarhm/j3JVeZE86QHIUB
YGtzbpCP0/ae/y445zuLhpUcQlcSFfLDy8FR8qEhBvCxeP+E+KKVUPmrvSWiJCfKX1i1cGSDtif8
RfxBZ3XqbJtXNxReY0zSNxXZPCMMboAllYDvQTqhYJ7jfre1Kt/NHOg4RHL3WqNBWHkQG91G2hhl
IHOSFV1E5fp15J18T1zAUBEbp3tg9AlhGjqQdQgHAfHF/4ZN+jm3HyTX1TZLdH2UOtqOSTr+Cfjb
rxCl1R0HMVZiww4cft+eXlX6i1hfXqpTj7qi8iBw0P454uceIdW+fcLWSouii+Mdo58qO/ofEmy6
UPr8G48HJaQCknwQh5nstu8gCRGEPnZTWmaWnWo3iV6tRKdw+Dt5dDti3yuRhbKEjFdNDtt55Dpp
2JnpBYKwJyWa7Xr6mhXZMSfgy79MG2yccggheKQwe3ScSc+7hOLUfgg9NFa+UuB0L68ChKDMDHSe
TYucBw4EHFbO+tM9cdh2lsxFAySkS5TxcLqygDoOmvCGrAwjT8AqH5X05R+46dOADQTRvAB9tfpp
tFUjL56kIPfNX2zLDz+Luw7y0/hUbKoGq9bGAlbooIk8Y2JKVtdd7Kiu1n9X+08veF1G+lN5KZnv
M61uctX/vLqrn5vXcfFO4tf8+s5tNjrqlf/k42IurcbReZx7BLmvqLGEqaI0xFWebwCyOcOKEyFk
i27rZG/Jg1c346fr1VB5VB7UBFaA/+FnyoEGRhZ8SJ0cfxJRMLH/FwgkoJzr0aApPo8Zi+nafCfY
qCVmZHJu4zOS5BGGviOul1FgZOXls7t70l+8sJONZlEwwGzNwZ+rcYQzdI2JM2jQ4zrSZx+Zglqw
nf46nUUExU7IA42Gna2t4ua1LrMnl4VsLUEroScjrJAygQ0p3M/K1FBlONTRSocLVxyoEx4HaL0I
Y1SI9NvrouyWvIwXZv2Lt+AxK68EK3ndrFMDWO3QK7Xp2V2cHOs205Jit6zYXZy71CUjAL+cwqOj
owO01oaTj6SxNPo29bgewQKDxttKZYsyk3ZZRPF/dXqdCOOrGY9TXkedFdOQq+T6gSwhh7Ep2bbA
McxyhxW+QOBOjnNRJomwmDfQU8tsC4hLPKTLQkG/5drs5H8N4jR5ML4xSA0BBx1TC2uOwDbFu/9q
H0a9DTFEjyKYE/ijFUuEZQ3hUWL4659xROWXuRXdw4KhXnK5n3kNcBAaKXEWIraSVk81Dq4qsLLr
KTp8YtB+MMnLBfWk3ZmBh5jtx1mIppgq4STCXd1sELQkLJstIX4qzZBUWeI8COkNlU+N/A1fVI7w
ZugoJwZZ6u/Fak6uwTCqhCwBH13Th2UCPdpjMPxxhtV0ywUzyaLCu9SlWJI1sJvjLFBIZCxQ2GdH
7yHdO3R1FS33ZSuO+HU0t2DRDxw1+ZIx5iqs7+YkZIuHLIfU8OL+2CUGeI3uC9aGXsI5XEjUEWYn
sY04wUzCPTDtRCftR+4oJLD5wpp2qQNn42gYIBSTuPQClCoOF+LHiobIZkkwukuq5WdRCX7xrXcm
0ZYf3ztA8XQx7+rS+/TcqyTMnxrQ2An6jHgFpEiYYOrCyGTeaciqH8Oag/89No7GC3MGsxN/Qm9R
X8yyEg7+nxnQkFPQ8bpIXse/lzbsOPjPwKBMbAhM56VD0hh+Q3VbbNIbtZdbMGnrzFaJD0W7FjCn
B3tj7f5hk+LYghPlw1AVYk3dzQSxiiihKrsZgim/J+xH2eLnCUyUgfCmjd3sVqcRAbLGe+JtKioa
jlAptzs+eg6WdSiTgleOam8Y2UxNKjjA6mcOqYzE97uxHExyr2AqYvIWGoYNARiDFV4wJE3953m7
PaH6BSZgVsR+xi8cNOzP/TEg9MJdjDTDEOYv1hlYDT+rks77AH1+93jui99MLipQ0QqJmcVxXcZP
nMwj/koLc7MRv1ReCnT6iFlrzNmuXz30oRMlyza6p5RK7YzJd7tmEFg6+1Jq5b1H+ZSsuh32gsTs
0x5FK+Ipy1ZKuE/kP/ydbbJNcldDadZsXDJ7IMhThS7g5c+jPub260e0vOENCm/VEgK2EtkyK+Bj
YdmegNWrcxyn53fVngRNAlwDX6Zbd2tjdhJJc8xDZ6h1IIW7Db/yxf9jxDK0w9Mjo/hJYqJ0DAZQ
eZJsr/6WDlmfB2Td0MmJ6nP9CHX5PAdQwOzfV1u39UaMYA8OBTvV4TeIjYkaqDEBCcglXomUyKh6
81INANS0LI2xjKLtj5YD4FdgNqwdoFwmFvtYmfhSfQBZIrkV7OtCzbRtAtBRxqHuzKoMa+6qnGt/
LEcHyOTRPcK/AEC+j0FU561gi0i0JFlTSMLdZ2XjSX1JY3rPNwVipJAh/jnQ0eJI7WFvaZa5B2D3
8p0I6WgZQtSOJSHLxw/iC23GGvo+XQXViUGwNhsZ3JT873PfRWPW9HAewFJSCSqjxUvoQa9sABlf
5ViuH9O04MZnmXCC7C38yXYp1ftPp2tCT7wHhvr0lvdvQxKVBLAxQ2dR25zXquSGal0Oo1wWMBJQ
98tFqDkwzZjFzfYJcmNHLahVlrDB6djIjirNTEzljACCebLWcRxMtId3V1/pMOvDlOpJWsWR91dI
bbVtQQmcfRLDEXm9g8BB9pPtV0ysH/YEChhrTjHdELU+0a04spa+a3+Q4mXQ8K4fRQLLb2XVC0YF
Ogj07wnNef8Hor10ueMsFF+eSPlcZSx1+LPnKkogsPLiiyxD1juW7z427eDfJverOu8bCSSPrNtE
WvH6S+KFFxHfUl1STjV74B4f0nxlY9ozEp6S0+zDyDo3excHNQVpKX4LPF/koWs1PXrREe1TZbLX
M5S9zObWRVZB0KRqqOnc1+VAt3uZw9Zcs7YmbZaXDCoVbWB2c8OKsxipCRAHLhNg6CU4NZLPLmSM
iXdjSAOk7IBPWBtdT3z/2JtavUp7am/h8hcQTZrSLxt72dQXkZ3GuyZ9OO/KbN7D09poWbsY6+Xj
T3lcT026hqoK76qfpzrJqeosxOB2LLyA/97pgcQA7X0y4YbAmHqkOELXBfT3++ivIF2kSEvqxz0W
TlKNluUq2Tk9B1eZ4AYwKSuUa6Kcg3DXi20lWAzsz6lUWGrZR3xYoi7yQKGDJp33nN9pQRRQNQXn
e6C8akxfslnYorEbfCTlWWqXgveJnNPULh/DelUdFsbRyIeVZ+O/S9Z4c1VzgTOrEC91gQxHvVSH
x5xfL8cSvtK581Mo3ANY3ewerLCcyxXoBK88iV9UyzReRHnP06MyhxMaPQqi//vwtNcMg/u1qew0
dQPGWmAAS2WxH65yDggeVd2eTr7+b3oHtFGYQJu3La1T8ZTxF/DVDzjtqbKZ74MJE1umYcOj0jjl
E8/yXGItS8I5mVOp7Zq56cgx5U7m/HveMJcZdNA+QqrAwm83M4kZMnW0U1OzGWNtRp7sAPPF8H4E
6UP7SpO7AimeGPJmai3iVoB4PjDIK3wkvySSqfXiso2CwGj3/Vo7ezra9COXFSTL1wpxzYsxytHL
D9FiycrOba2HWiqUwLFG4owB7OdmEmTId4A6hH5Bqd48pkw9xcY2PtO2407KQAYRjSRa+mEQDx1d
G78vd7XEsKIhHQfav1xM/eSYYKm2LEDDfSvxycuASi3ijpQ3RfpVj99RMkJzGgfa37go3f4W7SuD
isNmfrtgWUJdYKbrN9zsVGRRGK0RTVOwhBUVYJyKrwrk5QyoOSeUCb93QY7Eba3Z7CzRsLNvM/UU
xC1pqOkeNO2S8rZ/kkrTOqfyPPyH4Ly+s/kbpruHwXF24CXHpE31oD0/l1WOpm5/wrlIqvsdICnY
pbFa885qoMosTqSIhlNCKYRGXZYHGYnbX9mSewk+XN1qTw8T6M3uecCEmYHzXgjg9NVHMWQCuxF2
wH48AnJpbO05pZceczoXcHhuyNXUYbvZetg4mEoG5I0kmznXJ2zszgPOgS8GAzn4HaRoGWzyA8S2
EldgqWnqSPFDO8wxbUFzWeJNv2a7FZvXuOYml5VvVEaeyL7UV7aa07n+zJALHsQyBIEqxN7XxFFj
z+0LwakumiUBB2HNtB44SgHQVYQP0tFJLRtL+9572Eaik5Va/Mo9OXDD+9c74n/J61Atli+AFV2e
VwkQtyZq8vYqTMUPS0WLRzjAIta6dk03Asfl5Z9cUf3vmaAWMvq3sAdbp/HEO0ISfyRtj+Ea1wk7
tmoPtYNWpXEz22DPqjItm5a1cUPgwTcV+qOF5137OcYEP5xVnrXMLi4uKRcfLBXrGxzaMfmw1IUk
egnIfN0RTQOgrrauRy8njNfFpOLqsCEh5pwHJn9zrUs5hyc/g4W1ROGo01g8oEBWQmCAuTyqOivD
f3J3dvMRZ9rIaVJ2K6F7k+DQwK0ZNSBUZIWlpqvKDeFJxMCrNL8htI/qXh5ZPN+8c8OdGU0extHD
8dLfgXAfQd5rT9z+biIn414RArdRxVwooPhimdC/O7jXaUWwBumPRdNORFnlUgYn+LfqLsuOBvae
gF8ZZ05lVDfHaXHlzcZKA6kAnKinT4Pmv2fTWUiPk7C3g+Lw+de/65Cd8peG7eyCrFCD4tbhwvzj
i0+CEXLR8vgNklxj5+kCHIA++lh6Zfd0d09wxRbVehjCmDeUwC/iYLMv9WdsVJGK0bTAywk2Nzxf
lAYGzL3zOGm7p+TdLi7ObzXhlYNnsVkbWx/1QPs9gtFEiK4AHlPN4eFa/O1yuP91EX7qEBONOA0n
z1KJ+8DDbaH5X4uDugh54zy10Gk79uU46VtkjcqSzfYsXbu0qkvO9P3nO4qYurBBR98YBjq99Qh3
H3LzKGyuk9kZl11bD2DZzFzykf367RfafU9V75FRjFv2OWX5lsPuSmbY6N6DBuTWJJeKKhOyFWfu
4fzm5p6wLzK0gIXT3GTKNm7InNfmFn1h2+lc/FF7/Qq0+Fh6IQ2KwgdQUyER5N3WPfrI9vJIQcec
tKdJhMUddlwwMg1lousgn43f5b11LFBHQS7VQq7dxgFD6DYMLcGkTJRjaOJ03NJvtYP8bac6oYGk
0wQ3JTh6+L4dzQcFlYRIqz6NDwkJe90ohLeFdHa/Oo1o52IWxPichGJPcVP0gRh7D39K6XKMexkH
toMZER8ZWOnwsxvioXrc7oajgtre8uSjYnjwD3cD63exeVATAWigC3ppZTX3myd271s+YLfP13I0
48BMrxqhc6bcWgcNwLtsNEp5k5yq7OUwhJW8IIPOzaBcfQOYd9eBhYEFzLNfe5hzkOXDQDXQrNuY
bKAyvFu7ZM2QKM7KpaaGcr91HRoXrwFx5ITYURUizI0gMd9Jrvzjx9m7iUeT340eK9bjgn01U/lc
OAIwrhEVt2iymy4/CyRxVL7ucLM5FWfjLhLWEySs5l1XKR5BBKut0LlrM0gxHyMBybXQpfHzkIFk
tecGM5nvDh3fB759XFoO1a1JmtF960z8F3mnX2Wp1DbtcnyxjiIsX1U46hsTr2VwjxvDEYfDO+7L
XNJsv5NpNsEQI9vIJ93FBFgXlWAIpCJMjQ00+1CbiZLwRFwXYV1pvi4EaZ1PAUrrsUjE+vdRO000
AUc2d0IApYQyo09ouGgNzSDkvT29LT4dbvN5TvWg26bY0RSZeBnpmJB55a/w4GZcN3UUt5XScdey
52/tq2Prk8mhypC9oXVIDeBz6zKEaOPbxNz77sH2GnzKypb64neEdht8eOXQEeu/xEqx4ZDMNdqN
DY6obDle6w+qx2NcooM8qUYd5XGt1DVaSCH2IkfZBMrNIowskIqF8FCa6HugtxDVVVlJGKyGpuI3
xQgCNCJnDKcP7bYp9ZaIRrXUC/ZDH7BHXjqc863uFy2Li7lXtNzjMJ9aMARwVEwFqStNOAFKI7EO
jtNMhi/CMGu0ELZcaik145q46b2UDKjwTniq5pwt9PTbnCDTNXCjhrC6tYl+NYz/UcgQfv4oWjW1
pGJn0qpPHIiQXnrlntWqkCH64yf4knxxiptjmLQ/uGbkILJC3jMheHKX+aWM9MFghpbybCR/fn8a
0Krk1ZzadBIrsrXTSTnXCzuQvdHTVlmrAR8foToA6V5OIqe9GzLV8VoIXaigO72PhPX1sSaB4bpE
w9DylFAxBLED55aBdNL6JTagCvMvuXSvK1Ay/SUKL7UTyWdUWiRmT7VEUgZpsIOQJ4qvB9o4jsDc
h5HioZ6x/BcIpwIN/zXa/W0AJ7xdXWPPNo3fjx8sDxt9HvkM5LqkV+/0sf1Z1w4HBKP+JBbeBOXQ
QKrQ17KruK+3RqMvR5WhNl/r8b0+cNw/ESWAqXQvW68Bct97JmKDmuPntUBG/3w99h+i4ux1aP3m
uWXxSEKQDru132fkh5/NCxmzhSAvH5Zo0TkgGwzY2vohEyv5zrwv8rcOJ9CJC65N/FgrMC5c4rZq
DVt10R5OxUSd9kUNnUgM1nBZk+MZ1ATBheEvToB/bDSD7fvmA4yo9V+8L+CzSBmb5WgxLthYMUpI
7nZfc+lXBKaE7LDv0EqNLS/v1t2Dg0iGSkxQm5XBS4SGCt6VvWJA7Re6kiQ1N/RuVkBqtCLO9QIr
i7ZAX+6W0XwVy7DaXUmTJ2z/0aZYpB6PPNJmL0D1VwEq/viqHcrJueKysKYSj97y5l1U+pV0SLNo
bYFhj/ry9AaeE3FL4SHXhEzX4JPXctFo0os0ThDf7fAXAxb7/+uMyugxLcZgQTLUsgzNlnt+4eIL
DixSLSC9QL9zP2OErVViLX2Dc4VdktdjZWde+kGJsIZNmlp68vyMrD3C+wR3iGU7FGDFAnTQ9rMb
cagSeZDtkov5TPxZhkj84Mq8C0dGJ04qOaZanoi3oDmOOgG4AAB2zcbSQ2RjoK72Z2eUtVw+ikUk
UvrWr8M2K6DCab9ek1SNaRIMbICejtz7pKlhO7EhI7QVboFVR50VCt0H/4mYtllDTmIoQ1xIMndG
0ID7fgBSMptxIVZ3JF8AYCZ39LgN4HUoojz7gr9numqkd6oLwnKAWJpVq8tM9TSPff8mbCYAhCvv
AbjkpmGZgvEojNMyHU3gOee6bqovq/btbisbmQXL2fnVTlKcdE0K1q3J/Lu71dmEddvAjrZWw1yE
fbXVuxR79Zye9e5KrVkGnrzwVHysO0kVUKazkQnZ+G9K0ZiFjn2q9U/nYNc3WTzoUFYrlVvUyALi
7B7ni+EcSGLQVA9xuj9N4DcZC33KPczEhs72LJjicvhROsP1P/3vZMT5yegSaQF+sL4ECuMwE69T
4HvXmnJvz6X+uzmHeeYTzMq8jLNt3fAUW7rF48X1BbOL+Whp/EBJn+3IXs6+YNh6wJXH2w0n11TT
hJqC6bDXTyZinPCWsYEFTi3wzCRb3K0LGYSxTON56DnS2/eT75LiJF45rLY/q8GQYggcDhB9Sl78
evDF31kJXYvYs26PFu4iAYZ3Ulp1eSKcleJ0KG5nje1bVAqHufiAmG/9A/Qu70y2jKADQykhZCjf
+Z9oLoQHiLwIP1piS6VLlueml7uKqZzys8QdbbldkDRlikBefkFoDeb5yfnjibkKPLd5MVHmIq/u
8KnT4TftDYiVRq4uVzsngWFiOarc8Gu7Mj59Rh615oG3tg53Ck5Nkq60f915m5Ir0mxL2D2YXq+m
8pbEDEOQMcfzQwXAU1JmwYm6EWBzmGG9NhFwiGdUF+wfHhxOhfyY0YIo2AD7D9C5c8Nd9LcqxNMI
6VYJaLLiqpFe1+svv8IB0x9ekBzgB9e3isGBOffCj3CFNXujnx+AQe+TBlrKCQGjjTX/VP9lE2P1
TJaD73ki16KScGW+eIm9m+XieQ38JdpiYc6xCeS3ZoAqghPgGmv978/rcboIVmgXcUREcPdySeLP
3U1qkj9/4cSJJWk2vKaLhPnea93fsEc4sBfMT79DMUeI4xBrUUjCIz7PKNpnoXlu1VIb8NQSTS4m
5rx/R0EFYhITB5FvI3R5diz/+N5FQxXnuIC7erA/8gDG/DU3yqmLh8tmrmEszM3kp0gbE4WIFsIl
KTVYXJ5V7KegqiHO1yTQYm7ITrLP88LTwDR6IR8BPoFMdOOvuD93ew/+/IG9U141xCrCka5Newib
oCAIldHqA3V2yvwUAlDNU6FoZUd/B0ha2SbLcxEEKilDWsvip9tlNd1BDZUtRAH8ZhiYMgUu94oE
NRqg7Ph7EYk0uDgNjhibJXf9aiImEeqd5eZn4lETlLz/PG+7r1QZXTci28r/FUQAOU9pn7bI2RSl
MesYmVBFBLXxEAA+TmQsKQKyOX8g5lFn5xTRePde0cD2dyZDtZarCdYzEe6pQsBzoK5sZzJ5rEuu
q/IRkH+cuLjxq2j5C8BE5TGfm7Lt0BUOUMwKaWzclWUUc39tHoIcPEOmjQFXrgEWekF4N5US9QVy
vEdhlyJzHD3/7YXVwqXYjEwNwDpzWihyMbhohvN/t7Otm2xEN0O3KVlG1NaH14Cu5wXb1dF8q+Vy
VVy3TMUnbXyXSZRQlT3FCSHzBte/oKRa0ChKHGtO3wYLIW89DgTxztgIBW4NnqKk12079zF8VxYY
OieJCB6aleD1yeobsr57t9EdubpxeYJsuHqevUNXYEPPEyQ/ULF1uMClFBsrcnEwEUt6QwW3R1Gg
ETAWvJjNx/svXc3GEGG9J8ZWxXyVehaUQ3hpilZvcHt+SI7hkYrErEa8ZyhhMiGwLkOeybodjX6S
PTrnUY7KmpDjm6T5yhaHtihiw9klLihop3e9vymtSSp+ayX1+UOCTh2a1HAFq1tPk26fLE+dDLL7
5pGlCq5ngzCWDginuftlqxQjZVgS4PFv9CVohjBX/nJAJT+36HG5O/wOkh9DXoyrtfaAV1N1uHOp
MJBlqX3wty3gBly2hD2wiGrKi5gCwZDtjL3DnAGbbrO59aS/w0etmIy0XIeLBHk4WBKl3PW3C3tD
zQARhtyMTUOWjxEXbHno4NevEENNslCLRBoES/8vP2IpK7OShnQ7XZozajgKLePDRBOyklPXHRNR
4wGtgqsbyCxc4KegW/UBdHVTCRxWki3ZXaGalDoG+QwfJzRoJxAwgun7tSFxeEi9xTptNCzO33Ex
1qJYhWlVOqha5TVMym2LRnL2ahIfThqBnenplZa+fqDp8FLytgBvfHCpgsIu0UX2ORM4dU0t/utV
rg0A2/HpACBPB798NHF0kJeyja6g/OtSk+Iqi79sF0XBcMgPt0kXmGiGk2xOTLHPjkeNnuJBxLeS
4NQ1HySBtF4g+yODVCtPykQA03J9GC4LoBnxSyl2F0ZHVqwYrqxg4qFYz9VPOexcz7uZJqBqcv5p
xPw4T26fK77z7iVEIQZ2/z1z8gibI9CHcMMlavzzDpop9Byhn7ArbGEUxf76dhK1xtDW/umq1Zf7
3a6OZGDrqlTAfFImJiJktMTq3lp/TtIpIHS6xFwckt3NaJpbGOG62N2/W4RSB+s+Tlf/gYoPobaf
GWIO6dKPXd4Yp4ZZ0J/4mGggH63C6xWm5IoDFOxyGUEEqcOVao05mdA1WejrBkWZQsisZCBzUM1D
RlaJK9+fx99OIqDHGT+pX4X1f6rThxn6hRMwX3nuc/pjopELnBf4M5Dxh8NGv11ef0q4+HYnGEJ/
kGkChPKcdXzoBpWHWM5n4jzb8FEo5r8+qL6oXJ4UKZZjhCpDp+mWigBKaJcLO0B9V5LIpHc8s/Uu
2vi8NPffM429b640JCOuTp53wtU/TC6IFFWxboV5qPKtoLTTcgjF0dtRJkSgLwGRH0gPRN25afDa
nwvLSM1hXL9iG7p/1hBDEFHNzcWCBY6umy6qjJc4U5oPvtmC6WFfcAGp26UYyAALIE1tFSoxQPay
2TYYvJ1T02nXAObkeA6eW3a+b/uhbSsHwvXtKRDFEulONLbTN5dk1nj7HZRSkFRVcqBjnR5jLTao
EYVlvdequXbhnY1dizKBhHufsSyTq5qmozWBifcfKEOiVyx4GGOMaZTDn9VoAil+lJ+4wnw6CC4M
aozlvHAR06+kpt5YZSF3cPyuvr4Bb8pseHl87oHiCO8kzHBCN7skG2It6UphNs5RHzBj1/1NXMmV
tecnj9RfkpkBYwMRPOJx316RyfoyzFkxP/cK0fHin2giCoN6qfqCr2gH9fm68tjK245E3dSrQABA
yjsxdvGODlwpsj/om/IK59n2KBrzZ1ccuunAVD5KavMqHiLMeBeRoj08HAZCNU3vSoExYi552En7
Ydc2WVTDHF64rFuX/do3OdcmsGga/3E8eUuVEh+Ii7PXgkQXCalUMA2ueUi9FvVCdLc/n2RZ4wTR
dWaJ5Wy2EILV/Z+25XhVIqyKI8f83alnlgBVETS2zN6FUvGcc77rluRKalUwJhtuE0v4LEVl1N4R
VSxlAk4eEwQkULfY+KcZv1qO0ZG1ubEVmteEqedl8uKzo0amGXv+iABwxHfnW6x3zMJ2EMDS4+9X
mChB2GvR0Me5U2Fk3zJx8XracYFOOs13G8DUrheAbVxlXVgCq+uPLv+6p3vtzA8nfesGIqn9EyKH
TJMx8Ka+4rFTohGkmWaq+5IQarP5f3Mjw3MrUTwGYBm7SEU+stSawqzilUeAmFVSSHqofYS/UgWa
M+UhlvCTuojLahvoqxW9ZwggLqqm6MzIQASrbIJbA/VVV06yeyjpV7kSCKPn3Jmhzr9UZyZsN7ub
vBFqEoL4wjOAj00wE19b12Kf8ePf6ZoT8qvvop4v8GdfRybAEkIAhaXC0Yo1xx48GRGJoQR61OMM
wErKS8Uebq2RanSuuWLrBxFyQ7S+N6zqpvezlSHUIc+6E7FIXioo/cH7qbIkq3pTNvHUL30Y393B
zKjE8jaWi5i1yorAOLv1RIn9LTslVnZF3mDHC6BX4tQIm/yYUnAOhuAjZevoK3tLTXca2DY2JXiU
59KKZKUqt/ijdq0oazoE6v5xc51n09WbPKrr2d6pi62lZPKI2gCthGxEE+JuMLmjH6BEyxW7VXiv
8K4OM9fUi1O5ABgq1L+xFw9YRGD9iUudHtB549FRXwV4IUC4Dt3cfjp8KHORVaXC6nsFdFFZCBkJ
BKhjPrChrZ0rycJUORlblf5wVb7cZwR7jBXf/+syxPuUPFW7PldJnnpT5w1Nj5EdAIXyA25A5sMy
Mp73EifRYv7/wbePrWW44uTkc5uzEopA4P37UISNxMoRMlSBk/H6y8P+kjwHz/BpFe66XEEGu/9x
Ukwa5V50CPI9NnnwOO1RVLBEl3/n29Tf8SepsDexA+XV/F4B30WMWRDopmvc5MYaDj7j00m33Go5
l7AlFskTztQ17qM5LCZvlIsT8uoVtF6ipuT5h5yP9Uo28/WVEvx2kdVYyjT/+RIXGXG/zcxAomWj
NZ/io0FqpKaIOwyHuEDjaBVATkQsf0vbFfctrP8vndtqNAbviKr2drPbf7/0eK23QSGHbnfPR0vl
5Q3sI/zow9M5PFGR/OpIttYe0YLC/Lm/ByIxe0Auw+4xb+Q67t0MQOiWasmXBMrL7wXngajSYA4O
QONND9qyqajUptxX/vuI1ihfNgEYG/O6WdNiTzW0opvNN++qHsBFMrnkiOgtqX50M4v6q9jgNZv+
gEF521rnlcCZO5G01mkSMLoRRSGQph28W4cB+DZp/WFR1XZexFq+mgFrYRLlSgjLtv3Hhge4yczc
OoP3itJLTOSZq+YjK6pnXiiNG7w9fxHIExeXT53Kx/ceolQiPjhKpY6bZoV2+bTaYSCLoa15Nkpm
1z4IMxvSSS5iNy11aYYBEuPkDhPaL7JH9Ber0k+BvrqhyKzQIbMKhWnLPHsMQ0CbqHKuz6O/BNPE
vYp5B/LIOKctDEYv9Vfmgbhn8QDgSSUWxSyC1OPhmY7AWi2TEAg9xMplMdNxVrS76aPa4IQ4iqyV
o8LEtipAcfxrsGwQYzZOfSPwQPMiDTMjf0VhHulEykq3OtsCDe//Z0YIOgs/02leEZxHqzzBtxdl
fX9dq9RswcgfLvOqtPkzORBIBuM/clEGPI5PGj1tdDYxGH+j9DdIsF2eD+C9K4PBzrV+YzAwHpwz
fcaeefpHEc/yhr0ppNpuwApeolVNoiNmj1tFun8WPikgTE1gD42dhKVOqwg6mkgR8cX34Ks+NQqp
VLhwluYqoio9fCDRHjeSJWUohtHOXULCG/OBo+lxLJlEISZElEMAkAcZ2sE599G7rgLBVwxxAd+M
X42ymoKzFOIMgbZV/n6MkoNcrZWW6YOfNqZaXoH189w5fGoebMOq1eO+3AuL3sdckns1bMKBl7HJ
grq4JDVY8kLFZHoz9r14aiK9K/7P473TV4oqtim9lAarCQEr12neT667uj5RoGBEKUOVVKFQMi0P
3x3LrjVxa3peXM/P8ahPgwb2YtPuqOLnI1jGFZiM1f2RhrJI/2VYgBcOMLMtLlpA5LFjcbGWOqHo
wyly1+k6gYPN136gl3j5/q2W5qqLbnsWnS27MuHT+D9H+1CCnIpzQlhGg3devH6CjjKzMiAZZM2N
PEoqWATW8z3st/V/47pwkthr96lHJkI+q87duFTmdM9fdhNw7Fr7jVT00Om9jz9v1By7Jd3896t4
WV4Dpmz0F9Kjx8OfwdnBCcsNzi95Ar2u0rsy9J8w2YylfWE5RKJt/SPuHv2m5JPGhvS73unZG4Xx
kWDaRS5x6ptDmZoKkuCpbOHD1p8OJi4QkmlD2qm6L84Zqw6Wf56cfYIC9bnhUovRGSHggta5PROk
lIe/xfDjILQZtRfuybTVhrQ7MbUK2p73PBd9q5v3MZfEvhb8r4QMTROqb+1wk1ytGAbgK4cXwjhF
bBBq25dQiv3fx0rv+gSyzrhCRvw0+JViy+tDzkbts3OpuWi7Fc6EH3A3O5Tx6/rMshxkfM5fMzu0
VEe93CtDBmjuFzyiWy0OzJYdsIVRkmrt85ArLhDyMpnnSJRpYOmgueApsvLg4y0O+m34SIfZdgOk
/6AZFppp2+yA3kQsXOHHBNmo+8D/SOFg8/t6zgdJEhrCouy4hhXQO0o7ZvYN/YQtxkLaY+rZDncl
7N6Nso5xFXA9NbtBUa71a3kV8q3pONeYjHT2dzDmUjk35hmBlzQQtSDqW5IExfZqJmKOpGQnKjdr
03uTe4q/T0T9aEmjRXHL0LtXHpCH+XHDNmx/Rum+5vciz1hCWm4hQkVLYdBIrrjmqk4p7nBkWe2a
zn9sAFc+wdZ5Hx6rVLqqwMKkn1PtXg4UTkfvIHWocu77ysQmRTmMAYLEjW9eU2kQcjwoGJXf8pvp
gBqEp78TysQwnP13V8HhmN7SfUbY2fitqiWA5bRZ9JxIN8wJea2TXNvETy5/XETGxfOYPTXe9Qj1
IJPG50p5UeUBZxJHd85ujO054n/sK0CCRL8KFTIh7gbo655IIT8cLvszVELtMp9vKce4TDgOX8QQ
Rq7z6Wsx3o0AdGoIhdIG+neMge/lgG3EpBQzh5hnL5dcnfQhEfkQxkaHdXouF3TyaKlTCSUnCPzP
EHZKVs40BPNmBjpvEOhoPIh4ADzS4uSAzgzKKF9AFSD+ImaOJ9aqiTuMGavNInkL6ixbbbJO3CRY
2eu6VZqkac9DL5GYZBlxVDi2ltuyIs/clmCDKEbK5LKcpihpooIdCMrpbmykg17LI9YUDcTlVx5V
ebbtWl5cEZAgwfwgUetTjOx55T+1iCJgOUMxFedTT9Sz/9S1apnQ33SnJA7y4k4xyvIwgpN9ZGYk
uGHE6CWw1fqMcZJ8lEEo2EYW0gYb4gN4vB2bSUsk6rwIxbLWHisx3HhBVJvBZE0Hzg3FRMNBMcie
SbkJHAOVYauFotDElUWMIKNhX7P9a4BaDkTWsU18fspGOwb6pUeL037ufoLW8ISOjEUAWDbfaUqk
qvq8YPtkuDjMvpIbsolWn0c5BZ+Kjgaljn5ObBdmpCvYcASI8bDbcmiStOPwA63J1dis7B3WpJJU
U9gFaTnX/saOVRmxkLJDalCoMwS89wsZ3FC4ofIk1KdZ+P+WaqiQLRR5Pb3p9w277Uy/cuLuLQBo
CW8sbYxrmnrYytjEiu2rDx+L2aD1hYI7aoS0EDIZeVVwX7KXrdMI+CIlRrd8O3+zBLNjkurSS/tZ
1/a7T8/BSe27Ucz8K4Uv+Ds2Xjo/Mob1w4qF3GGcXtLLSW1lSs3dVtrheUnEDpbuLY5i3dEu/Njt
onsd6DCSkljvs3QznWJDV73Z/AzseM/7vnvuibDRF3FXpffEMAaotFUuJEDKI1p+n+jeGupUI9UD
9Cm6UQIeE4iHf46frqa41ryv0WnZOTGEADbhQR9zJZ0Tqpwqg5WbM3g64sE6dzCd3X+auk7AOhry
g3GC5KaLcMkmOoNenxzUV8ZbBnSu4FnZCfUK5vPjEJbCs0FF87SUo2uODGRxFQiwKmXoTSpL/sOp
eFs2mjQFdqeo4I+raR8CNXOqfMQYHSUFuc+LHMCLBBw03VzQhmxQbyAwZx8lK+GU5NS87QPa5tjs
ff/oXLiKceMjazdH1TOt1k8O0wgn1Kb0bfHF+1NppFTwCNeOzvapTe9IYpg191HjfNXwkuEx8uDC
BdRflsAbxxVayYPg1dwWTb0dokehOOhMnKTc/+IAOFF5K0lgYbstes6fO5op+UdFJxEA/LNr2JKm
SJOlWmAI8inBcIfoMUzv1pAXxAWGy/eNs6Gwi0+zyeYnH3T8Ks9WhMK1WQbP25MStXnQE9BCn8oy
coZHZnoiNzzG9OkgmmTK9Lsc5HE0qSRJUBUUVXdtV24w4BIu4P3IDLp6osOHe/4G2svCRJQUEHYZ
1fXbe06MaR+PR1esPUdr7qmYznsujUUOPxSB7DG9TtE8ODzL0vEIyX0P5LZYbdyR4jPYdTYnvw5h
TrSCNNdsxpeUrFL+Vbzrqqa/WP7+omIGG2Oc19NiA37SBfBqQVShsivX0tSFSY15nlTtbmR7i53Q
afh0qgBOKA/6+kyI1PgzIo8un3qFA/wqfkrp07B6+D3oFO/gTsdGa1ha5AAKzlMTugdVII+2eECH
iegBPxwh4qsHV9AcSVRmdmXCATin007zuUpMcatPYsip9kTNNAaTw08b+aR5R8cL5zGs7I2mUhFI
DBnv0k4fDqxK0V9yK4kKP2Wn27qMrWgVdfzRmjRvtSCOIuvvnR+Rko/VWrlUqEko/f4CYsrwj4k2
Qwz350nk+tMRvtQRY1YbzgItqMSrrA21cBceC8MDNX07AYzx1v2jYAg4F5W6vv8vJpWoFmbPihQh
QjxEfADxNEOeUsx0BvxkpYBY/S2GNYtrZ/XrgzUxgBoZMQxXIvhGkLLMi2Hrq46F2yu0NSg9eq4B
w/8lRjWqjB7gwdowb8PqaXS2lSdpWC0qYMbeEXEAyj2TMTNrVGztDoaNAzAk8DzTqDtWrxs+do7A
sStsXyDNYmAeXkjQiTiNeKpoicz7kpFaI2QmWnqfxICAnotfgu8dziDRnhzIN+7jbaBAiV9AXIED
8YxM3cD/E3FZcmvxQ3Xh9EFwShuXMujxcQ4Rd8xqSoQqQF8jukYS+zkK4D/Vq5az1M1nP2y6i3dK
gchVNdY6twxHfivFwCdzuRsPNCIKtEGoWNqndk3OzsSBAIW9sZmveGr/t4Ot+cn+Ohae9IBVUsHA
9vt2LpgWwXuunvi3+pLi+IxgWIzdikso18hhNHIO3pb65yYIYZvzq6cLMfRTcG+k0Gn9pRCdKVWd
rhlawxrGsH2zKw0t09NR2LNwlZJnVDZ411S3YZEXcBEZtA9MtLthKcLywlJFX9TsBpr8QQHPQXUc
iZDI63BcVI6A7R8Hx++EGmYNJsfLBHw4T6U6hOVPawfiZZyBGDAyGO3m150mbTTBT0T6cF5gMczN
HcCfQBaTMBcj9a6ALCu9ydNsI0OyIUXe93926t6DUAPYT/Dj8+YPSgha150OjfXc3beEgaMohki2
rq+Vt7Tg5Yi+hgdf7MlGBTuU2ZvZ16uWu7Y6PLbL9O1rCwuqmnz5Bt978IVaJTroFZROniXJ/QJL
NLPcFK3JGjf6St8AmEeQpqoq0SXcai9dgxh4gbZ8PODsZCrm0IMkEBqLnYes8qKYVXDKbvoeg/hl
yVBow4zozCCmLJtGfs57MGaixv/S4qF7aCM0KC40DdqSQiBD+aiJwsefdtCFhwAwMsHQVETp9TZc
eDkTF0w7GPYQkO+TMKPaGsOVDm0+zTfSj14HKsxV+kxqdPODNUBinQx3rhBtxGvq99Gt7NWTTC2w
pT3H0aCKJVbtvYbGP0bum53fEcZ7pq2RfUHahHomyiPCNA4c4euuKm3ujcTDbho5LQDfGGgg2sg1
P5YHg97p7pjm9OH5tybyTbyY47/9APys8hMwqOvy87Aifsxoi63bw+mfQaXhHghD5d+uLz4DbUen
Oo8tKo00KEZvL1NrV0S4NqeLZ9c3C5CsAkBKgy2tjv/1v/Yyh6iCq5ImJ19FPVtMNSkToVI8GTei
eOh78pJZbYv70Hgrtix/PhOq+SJgM2ng8WQSiPat/mvkiAtz8JmzUsxr7UXs/SX3KSzGeFzgGVIz
1dnmLaejFJDGI2koIn8C/3WLSlaXE1IZlkQrWFoWJmUaS489iei53V+tCHwCmvFu82GdawXT7zgi
RSPPOQRDGa7zwN05XMBYdZfvi1aveYd3KkOS86qXEYQxSgAFbkPgxLJwRUYxQe4A+w+pOEc9G4Y4
Dl+UcjJowvQJi5YuMeuLN5PBcxMYcDniQtqTg+iurBjtxbB0lom3RutW0yB+J5hQqDL1lj7j1I9S
63p/Hv30cYa2XYIpLO7faFCQms7scJmTb8u59U1z3J9GH6f55EHzDHZLkGfyqqdKx8o9TFXYq/F2
s8od4Zqpv7ScP10Mgkg1ksPGISEFZR8uJWwKJITFb3DweJEEJAyL/7kuPZyZSEOj75JCcpCMQuIG
XWylCjrW3tWi3kP0O6eLXf3T59uTwprFxWmezLQL/lzFQN/f9S6k+kNL+8hyD1DdnqAEYP46KVDk
1B427Frmj0jhSUxq5GmMrLPpG6+8a9BDVkR04IXsNy/exUco9d70BrBW3PNeexkdoDWBO96N+Ymt
UStYtMtomebhHahiVYy71c8qh7X4NAjPCWMwhS09FNxItYnKC+7xtA9pKPH6XYePwAA/HoXBsYVe
R895YPFRAfZRYC4zZAKSAK2jzhn98lOF3NIcfX31v9eXglOTC92RpxYELBzvfIqliJw9iZcRogNH
6gbGjiBM1489vGunQtLi7jrnJdosbVD8Wf8TxTUWM6asbZZVhQO6a8tzi4MSZ7lLrzykJqbJBwGE
sTliB2sZMQd0aVzYgFkrxQ4IcL8jQfbKBAL/I4Lla7m5TZqSfeT812l5mwoxkZBneT7cByAse3Wk
VUhpVqKWUL+U7jf2Ger3fMN3Yjk6HAezncNXFIkyiLQBGGo1A3eJbYC+JQv2k+TcDgvAAM7leQch
+FOGVRuuSeeN1HyY4eViNayzU5Qb+c0u4yymuCP3JNCsmJs07J8FBaYa10qEQy3zTH/Z4n1dpCSA
EH4qd9F46YXJcXeuT2zgyoGQusvWwNCDG154Edjc0+KoFDJXY5YzZKgkJussdQhnP8awpNFII5sn
Eg8PHpJQtEn35V7C62P3w+/HX+ATBfgB+jN9cp2mjK+8cwhFRQ/eLmApQRE/+BVXskSv06pJzZkt
7Mf4cAr+htZXTe+QIoM2bcEOvfv7MnpurOmK3wzoY308Ai5lW7SaUG5pHhi7n7nF5GT0/MqTF5mM
hujOH3nkJNNJZEu3B4DNzMqkTRWRgYkpY14jnzgG+q5PH4854ZJ1b3YpFwML3Xb71hk2Qp21b+Er
kv5cXQQJwh5YsHIbrrKu2yqo+oCT8TIVVwGFZM0G/XIht4gPszgzcCoGxpEge+0nQfWCb/9iM71H
nsBIpJE3Dk0breQg0GN8/d3iP63b8xZ5Y0TPM8LyJ8629xaF1P4SsCDKBPbVtt7qMtuj6CIFY0e8
0ZPteUs65A0F9arbeq4HldZzMcFxvK4FuwIKnzsmx8pN03wVjTHeR3yPPiRN2WLRvhsIll28ctF4
G6TfON8jW6XVCMhMfuGYlJ1NtfHbuTPXlS1NWMOqbd3sbqTxBoodxFyGgNFq2NVpMBZFFVQdTikO
CTRHM+iqjClfHLohoDk7Plr7xWqrGhiAbdyTK99z+Y/UEjfXTLIcHzaRc8eLjHl+gFp0dDMDEYNy
jsVfq9ps40a64+AF9r/yrBSV6uwc5uJMFQCe2mVn/bfCI5iMjc6CWHchQ/sbF6FBuchcok7TxeTb
++QR5Vpje5dAKp42LwSKnCxnwWQhcAvUv6t4Xq2JyzLEep5Fl9QuuN/av5k5ZYrDz0GaAgvR3EO7
4fy3kmvfXsD4ZA7vgEiqz995x3pquQAltwk/QwpQmB75c4Ny1Dh+uGFkn5RA3wuY6XnY9yXdBvPi
cOZoNZ7/hlff6DGOqNp8liPC4N2S2ytHnSF1ZVQsqZ0RY3jvLI9mYzhsLrEk3LwcjPXlvsavUmAL
SN1W/cRed8LJBD871UJtL2P6lAC9nQUOfFUIq/mHQ7O5vmAmYJ7Tb1anmsSQdcxZmY0lELo6tI0z
Wdl2xs9UauJcLmzYalAsP47mkd3MOCLsF3q7R0UqxgLjvULRwQ4uFgBIU390jG3Jhy3agIiLydMb
vOkNBVo/vFC7v00Sjhc2wTuqJP2jPbILFUKT/TYSztWvkwmUujWUY6hcuxLDxEYUCK1gureK0Mp2
DETbDE57XfZfdGGseI3pUQMI60nD7vpyqxuZpJof1xrxJLFAxeXHIopsFwjXRMUu48TJlioV3xty
QoppR16XiZxQtPkXJ9+DNdE41dk71WXxV6USXqVcRfRpoCbnTMQfRKwrpPb9hHWjAmYUjP9qx0Tk
JNf02EsBEQabwypxLuMJcKGn2BWH5YOCq85kXuaqtB882letcd36YF5n7JxixSWzl/emSXtdBwTe
ds4Pqa/jUnzy7JKQMq8WitTn/mplNViOchhSK2b47vYlu/mdNhtOOEi7RnUVdZCh6miergAeu9lq
GNCHEIauQYK8nS8ZMmsI3/0fDbTRlM1zFlj3IK+/OHH1aAh58QAGAnS7qp6EpZIl9y8e4kC/LPeu
h6/0wT1+7FlK7rUk31J7fqxmDvDaT+tk8aDjCCbzuBmOUwYSZJu1rq70GAXindJtPpF3TfqsQTpi
UYbxlhc8+gy8v86MGMcOBt8+GZbeBlYeE4ZBIbVzmpmf25Zq7vcX2gM3SB01c9HJcswP4PMTmx5Z
3vcKzHP33wfaVh9zMEYmRxi+2s3sRbjviSZlSNhD+YNJNB+gqBcxOhP2NmVuZfpf+KUmZRLFRFCd
d6BXGFTXo1mmoWOEQampxf9Xv4QKP1JgVatsNAjn+SItnWjzKnvYTviCCx8wDKDX3ZSIYi389abA
mOgxlaXmYUff9S8H73KFjEJ3EHuvo24c3Md+jlHthQLtCYZUSQFgmjETcLAmGRIRO3u6kRnHm17n
52yoznzEMpRgKzfcHxAuPoR0UpuUNeryU6piEsskdQ49/unASDV3lneGJm6lUrzWN1EvKW4/Sk3+
TnbT3tHcT/Va1LZZ+0924Pwol9dF29SuHfdOiA4N+xCjUC4g6AGhwsTVUwctASM1LewCu7typlZv
OhretoWstVwIhjJ060q6iFM3ZPzkOM6CrjfNPBiHh+cCerMDU081oOarLRG4SuWjia3oIbzvwpC7
kcxJhP8RQT9tiEMQEewht3+OWC6ts46YYhn9b7k42B7uitBGSuGTL1erSdI1f+KSt8XZ8iq+f4Er
IMFXUFhivl0KiT3zt5jfueMyV1l8mzd0EwXwpbA2aJSnqi8EugWjUBe+Se4jFqrjmEuFC1nUwJGc
NYxOJP1UCsgTMklQwKDQOw75CSznNHlYBMU/SNoLtCcjKvyg/Q7dXCJwJw2XezcBeGSubTiEnOtd
BBJTpS34A8+lRK7AVDnB07lo+cwnh6IGDPpPQ0T4XVyFsgaJ7HpIHbVP1ZkuzJ6dibtzq/58s+m6
C7pl9BzYVhqakKagUFGzUspthh4y69jmQNY5mj6SXSNHRwtcM10faegpCJ0fRWS7506KvnaPvU98
fEemgOCrz1ge73RDSeHwXWPr8jbNoTRfpqgup2yLToPmInRC9x8rIHuhOQOlNTtpyrIQKZd9nSt4
oZLbaTOHKuSxyuT7DcGzE0vRU+dnyclMW9FH7b4x0uhCasqlUhLJXQ3Y61iSuZDO4nKasAt7YM4k
kqY/nmnHyg1pb0Geu04GsGEiIWmoUdV6xW5GKbtkApApfWTAa44YROGmL19dC1HBToaTPr2BROFT
zsvxtFyvpQxgzg01LBD+m2HGL8AlMPxKwVunlfkPwv8jK0AyWfcjZyrxyNIlO9yfcYYLsgkVBFSy
COTEovY/Jq/N6Al9po5Z81wLpdMphpc2/vkGgacxf3EOGirQfbEPpcbcZ+uQw9ZOTgfNwkASlkSc
JdS9EoOe58mR49bc5mlIB/0nnsbLRGI8XwiBGMymfBAJDYF//Q4Z2WQbtCtqhy5TKcmENA/MKn/h
ZVkVLD4HvjZShPw7BRekqjBIJiY5tFwi8DsBk7GvANoHFksEUDM0xKmZDeImW29ipuZpJoSyS8yJ
TWeEgJ0/un6xKtojdovW6BsEnydAqEBCUP8nRQ87lwIp0+5bXKFSlPFB1jgDsyY+FoaZct7MMH0G
zWOb/0qykqEJsOFA870cHJAW/IQmWcngZ2Q+ynsTXKeMBIuPnrsmpENB66CnPxUO3Wz9OrDBnKxr
cNCgSyrAVM5h8JA95Sr3DTRaVmpHzGS3DpSTPTCLBOXpNU8ECcEBC5MFg1LKvuWJ6PVGg9KDOXxQ
GQTbBiw/KJcO3GC1IPmugKROPkSDk5D7CFm9ZQET51cPwH3FaYWtLjeWQxy10YZYG8j8RwLsBnK6
5vrNKuC/E7B1lHNpfPHZaZRugAMkQ/64sFEEYSL94XMzUt9FRbBe06amtbudTnVDXPnRanMfhOeR
68CYfO9k3D0+n6uhxZZSlnyqKiNUJC8q6CSHzJlnnk1MtcygcAyEy5Ef2DwMqJg4+2MF9dJds36+
XG/ew7mXdP6XRswbRi+zCLk9IAtlnn8qet47MSbCIBB6yfgGbvTKGAHMC+xYALygRS32t4/IhE8t
x7DxGowhy/XHQps66Qw5JgnuLEKhk+xgX/gNue2Ui+gawCXtLEZCaHm90QwrPvJWF9rF6p3fvrG1
EpzicYjsz2sWAHKfT26Iq5mNmbdOY2E2ZbDhon10yoeE/W085KYtObY0BYvMe6bP66sN5T+WgJ0W
dgJPiKGNZ6hOc5o3vJT6o9lze5DHZhgoFykJyX8819jr7nQcPqDR4Np/IPMqknNXqKGNn/rNeaff
i4AvnxRRKHjmtE3j8nZLadaccJzLBdmtb4+yMZW8LWAGAWmxJ3gh1Ip4gFlHyIkPnLEZ/Qxn3Y1n
WYKsL2iuRf2evY3YcXlqXx5gifiF5WV+5nKyZ+9c5tXYramI+iP94OhyqNrV1xGYIw8fZAikMpxX
ct3FEg7zff9CIRGATev5PjB5zA13r0W+Oh6GY7qGjb/DJavtzVtBUEPJksFaqm+L03iHiYQ4GFAH
5CaFUnYCIrMDnn4PmuSK30lxPZAcG224MRQhWIIso9HPkNEAcXyH27OlNny1fmHgADb95uZ/LKGu
17NaIBiJkzasRcy5XBVGtg2Sigb7xDGbqYcZWaFrVaBkg30h2jmJo/S4AqU1p9yRxCQ3R1KnxCCr
CQdylyULG1wtGyxGSdvclc5NRFlWRyku5mVVK4Drywnvpx2uI/45A3ZySEMSL2EdqGYYPtGNNJDj
HmUdBz5azJ/FZQF25rbcx7nwaWdWSVPwr2udSepWi5uy32EskntqBHAWkd+iJtApnNT5DvkAYJ2l
e6uMu3Vl7QYQSMYXKdaltFySSinn33+y9vFjVHc/XXDjtPsKjQ9q0y/0C5S66GD7gIaWdb0wOC02
713nkz7fJJ5r9sA1bd4PGaTW2dpf83OfPW7bYYjB0X7vU9GUc8c8YBahuG7n2t6sGfQ/LRyy/UfZ
9NWzE7RCG/W8zhRxT4a8rNJwNPh2smeLF01/gVpqC3JwNxtQh2h0EcwBak4QdINsnMPz5+9qz4sB
N5uR4ZE+Buql3awnNh8LDKHOj00VX9Ul6choWPV6gyZRsrqP6y1bqd9sWkx7V/7bcd5TUn2ZTwRa
Q1drW8glCu5KnojThCuI+tMJ1gZmuv+o+8QhajNnhDwWzfVF7heNfAkmL1+TGZZ9X/shmUAmSN3G
LTvGySA7/b4Pichn+Rf7Lu3szQU13kAXPljgwxJiryxuSQQOR1DPLByEiZp7YHNejalLkubbnqds
uJm8dvFe9k1O98XkeFg/ZllqBP2OU/Pw64YkkaIeT3HfyiYODk6oWh8qqtXu0a5wT3ZfC05CloDU
941vOT4ubKBDnWrfCQLde9S9q1LbTuXRiJQQ0RxhBvH4GQVS+kjZCM7+Y6CMTFV/CHWLsC5h96/y
hcA6M9/Tp2i/klppDbjTFgU9bTfEE15+KlClenNzLEpCgUmwB/VhRXQmq2k3oOI7UJq7cwjxk0GX
JdGYIOJ0DuM44EpXU43Fioz0z3m2VHAtVqFz7BUb7FenLc/jpvOJkf/iaallgIM4SkVeQh3V+0U4
Hh2qIGKgrde/DIpiIIuL1fK0jmUeRlIRtphUZgw4igIr8eu0KvbRJnAvNh9JDosEdbW8a5ZUtouI
rW+bx+WrIKTZW6+3/chP90psoe/Kp2R+NevAwnQ1RNQUp3ldd1xnrPL2buo7897Rx7eJkv6lcjGR
5r7AO8UHhRsU+9FQazsY+59WXJsaRCBy4ElQNghgxkPKTqbm9/xGook7V91dWnroPn2IEk98orZR
WHDO2opa0GSI64rGxyUMlTrcWSqqea2U75eNw92cKsdohumsthWhpIaVKDXcvglC5noOOXGNDmbP
AQ/dQPfWugb7oboadPJ6twVGf+DkitIsssM0vAvZfM5PRKRGOUKM2mO5RfrTMvzj2grxgQPjyFQP
U8JvOIhsAtUogMX9pLmCKVaJPlHb9k2j6GpeHVWRjffWRXCgxQr+Vqfvix3ZZQe4+gCH2n/oCwAm
JjBcgKffjChIjKZsoWJ5kL3TTTWq3saLGYdMIX4R9wcg9GMMZp/rJX9U5o3cZ+1EeRWNGcKx//JN
MO+NgCzGmGgRgCFuKOwFvozCfrF2oxLZ8WN68+vlAIWgNKgqbX/jYkhQSyDfQ9b/5Rm98pap5i2n
cZheEmOgf8V6O5CuIUhook750fkLZj1Cx0o0XiK/DbIGySOBHFKWq24zyLZ4Fy+hbxAPVHroJ36g
9eIj9FgRMSEmrQnuIk3hTE3gq8S+hfNPB1QGkIe5Qpz/H1MoNGfIpSk1//smMy0BMLFaqyVoaBFv
cRjUnEH3lkKtCIpT0WaTVeNDMEpxKxwmLvgjb+1+pJ4u36zTc6VPiZYgasOJbM+C+OFdiUXSLxwn
z/FJUe/Ki76om4bIM+BJcJHojI2q0r/UCOw+PI8ZyQFmiLS9ZK++Qz19vFAIiRtPl9w9C1yBcoPX
BzmXYowpTCdXr7P/yWZBmEddZ3LYl7aqZGE7py7kHUn5JS7M4eTuJC00brQbjNCskqZeM4fBhdQg
7a5gFfq6ZjxB6NHkc60j4DCRoYGh+EloynPK6MiXhh2rsHnkGcCV+XA/CmrBZPtYOcRdSG9aeLb7
EXg7wTAIeOKZfFGh6wa9sChTeLmSu29zph1dyUawmEKa3NnUcucZSw2/KWQAzSIt+CXrLe9U+xRc
7bdYwo9Rsl9aMWFJHNgT9JY9pmEZPElsFTaRpY8JL4tGgiQp/2c+SFWRIwXGmGD07aNXkpCZ6GZ+
yV8cvmnwRZqpXFHw29STgXD1CSEsQYb4Y+ZCxpSM76P2kjMsxtC3qZVuSdyGJdui4DB+r7uy5P0Q
3k1MvfEaVylAJw+lpYI0qknQvOLOaukc5NuN0uF4ubadU/DBUdh+PNWCeKWpKUdN4NzlD6Sswstv
al2r3lE8CsNcZBzk3U+GUUDD/X/iipqohkw/9y0t1UGJiPbGyeYTCfSihkTjaoWrMxA4eHf38RFJ
OXjBUmaxWmgitpLKtqzEhzpdcjMGXxi9G75t0YXuQnSLSLEKCMj9QF8m2EmjKeWH4uoShg5f1dc6
Kc/rezImHj/gFyaIbrrhon+/KapTG7LZQukVvB/I+V1JIGwIDqBhIxMK3jZLoMQv7Xb0uGm0FSLl
9vFV7YEcSN3UgBAObCvtI8bmlJcakCfaijOCrTCUvZdXJbY+xqBfHSuGklVGoNoJ0GhQQKRANJK0
JFpR7AIZaFUBize1z+2voSW4DJuV6iI1ICUhtBWifl0AvK7cuilqfNjnw7v0Mq5222x8BxOnyyGY
4mDZ17D6EdjR3Mis5euG0KdFYdfjeT2c3PyI7QdFGv5g/23XZ8la/TZCuSOIyWVP4Hm0/aNh1t+4
Nqtj5p7l2PUaq0PXz87XRE6sKrJCz4u7+mOXLNbuOA3P/C660DlcPrvcod5g8E0pI5IFCfbVJ+9J
NYMvLz+pIQmZ/oGRVVp7Pzjl3UM29KcEzER54eVOpVBB85Kh95EqKqRCnOOcM+bnZT++J9311M4N
sDBm3ygCBKsOWkMJHN1fMK1SwP+0nv6l2gJqUcnBNioLM9kAsflWycIxnRFIPxKMXAKpYt56iIRK
tN+MM6k/W/wrVi6phofPic/xEY4tWGcNgLeZqnqyyorYOSN/baMzpF4dUQqCSmJRUIif44PTLDZI
GNHEe82Bm2XEro9t6Vb7v+OqmDa5ooNs6gI3981/k09lm7pBmohuoEu6hLwECJqpYCMEs1X6l7S/
P6A/e1ywfj77Qg/7Rsfht4ynZIkl2eQtwfaxIGCZdCuEKSQVQsCkoi/4Knf5UUGIqkPTGtpno/Sv
rODK1nX+7OCisVkMeIlFXNG4pBd67kPA4euAKtcruqG42fGLVPb5msHTzpeEgPYsAwdX/UQuB88H
TNDP73yiwo2EjkSeuarU4OSoAZ+T5etY+cVGXLiUP1lgmD449tHGdutZNDAVPyz/h4d//qdCMtXX
gpMQiDENt6f55GaO3GGeiDxojvx5EH95eH4lOv+UfrbIxcwSS/KvKnGQee3Wk4HhPvmI+wtT451B
fUTr75N1gel5KRMcDsf6dYdAPuMwOKAmb+W1yuW8m2COouBjSjTyZIRb/RsZET+H2jSxu/x3TyAK
p72Yw5coV1t/znw8gjkx46prFAqT3Gn0NOBhrNDeSvwa0YxenZ+HGilaBvdsuKVQ8VuB8ihChlr0
L9RVRIiG6zgYl1DcQ5uJyU9VpbYoXmPHOuqoDYIeA85MlYL4bga2g86BguKhrnXijjuEiMOCUl96
BldRNkztyJCfOzBqwQI3x2hXftkHNTkX3jCJ9Bm+uKOo3K1PKc2Rx07C7/FYfj4bozavlGTBOahy
6r4CZrMggdrQ2i8N4dztTh9QqQIcZo1eFBiFOLmQgMcYVwb437lU1C8dxevo5YjHd4+DEqLiov0L
9popMcVmlzp0nLvblthUeg/YLvmIKtmOOUxaU6838JUOKyUyl1eIE6zMOuZd6irxNy5m0cVazz4s
kEIzPO5S4Y9711iMBM+ooM/dLglSyitOaz/ZeklnK/SkzKSUA0/HKIE1kxmlwqQ+MAS1EwGZM5iW
x7Ih/mWO5CmIFdP+ZErzYAno50EfBe92sbzefv/4i/AHKn0o0JSMj469nboZN4Yh7sobAevxH4sN
EkSW/8sSq+ePmtPVhPmpfUgIX5QjeBPj7JZEDbncH3ZhHsQYC+b9+J94TF+CsOc2oaEYrjhOFqfx
C/29yYt+MZZFWsAJRVQfi4/z7T/Fu7ESKpMJJhGv0IsKMhR5qm0mpoMImc7exQ8TUjosFguhMJVx
o93QpYMe5Sv06a+UL1JxAs9CKnviNFq58OgfmH5bHisD0cEYVKMr+pQAVrN5vYkiQTQ1Njlt/7VK
42qhKbjw1bbgfFDTWuJ6n+QRiF4cA9xRHEkjNqQamflzumh2n86SMCi/FNyr9A0xWfXRUGc70iOD
ttDOtv7Tvbgpi8RE8UslA3rJ43+2xhFatYCQBH0po7ZIYqp9KCd+GVl46gLWcgWpwsxe3pqX+3iV
nD6eqMCq9dcTGUbzs7AMqTRmE5sfXbZvR8t+xkWBPpFjHeYZpfflNUBgBU4GYDfVkHdCx9UVW3+9
HChBfW+S1zn0behxlvSzQKS1JvlIQ1H/KZ6jNXfDA9FkRE5f6f1+kSrByrjYaba5Kd0PZLKp1zjD
ehMxpcaGdsyMYB+Ig2EnhrrJUQQIVsaCwwKY2UxZNHYP3CxNXTtb9hTe7fgOgBasszve1q7sVCZm
Wr09ksybQvBXjMh1FC8JPiAby9zE+U8M9w63FlFeWt8WCwq7RHX8fxwz5mrj70BofDsZvzU1SBuI
dJwxdqX/tT5YSfNitvBDEn3tpc7QeGp4KhmfMHipt7qxjKkSsadR9A3YLuFmp+xiSuY1penj1aEe
ld4Br3l4Qy76XOkLnHHwU2BmoJsjKU5AYOQ137p32dnRf0f4zp8FUldzdupu86KaCC6PuhuFwrKw
XhT6AkS8D50DTleI13Aqs68hzm4Z7vSHAejr+jyCe54z7y7O/2pAbsYhIVk7/FEYm4nXU3hHDYwP
5xzdbH2/YsJzqe2UTNJq1icbstHFgZNV8XSSE5ryUEVuLOEvZG4to7WgiTAgA9mvLXZoSTFkad65
DrpZsWYlLiDjvf1ldw/zYhx9C8gAglZi8iul2kyTFetsAxfU1RXw0+hQ2Vn158zw15oUpMKgMN1M
wHRVBcB84rMrnE5CRuStj4YMoPV/JIaovyaphsUPsvIgyRB23Oiu+S0e9ZQU8qkuGg1wRdhVsKd+
3bwRhdjyBbwFkpF//BPVEp4u8ApM32U1hjBKzaFC2kKg+88s1drSMsCw9bTGolTuBM5aBfaQ+oEx
HDGHr4gxROTZBgPE8Gh/aNO0wXpiHxQFHbazt02X6fKpQOmWX1llSZBtlXWxwi+hEqw7jWg4tyV2
JQJZNTP1As/u/6oIEinhEHU8phLcUINZv2XD930xGfW4jvq4I+OVsNV17PJ4ATachVKACh84olHL
HVw4hbA2GUV5VpHwLBy4AuwJNzxYe2Iwbe8RxcskpYz0tApFnrc3cOiy1Q58FeIPlDk2eF85J/MA
EfPSl/+ZCtD3BTQfb7UC6oxR7eFnyowAoFvc+96qZNg3me8JhTeWhISDNDRiNrruydGLmIk+lFiH
scd+QuWSZ7ImbJ7OkCR7SBZtb+kBxW+mihjlTYUOl78CDmqtwiI7BPSn/1bHbDZVj0eM1WBydBnx
wts1gkARARIGRdOBFz++LCCZdv1fJ203xYYiCe08e8BHJsp9h9ROA806YG0tAQ7jhYJ0py8aFfl2
C1/VeByE5s4agLJcfSdIaHpXs83L8xtg/m2uQOFN3S1IYvkJNEUKymxbEDmepsPOOgZJP6/HQo3V
yVEir9Q2WIhZ0rKhIrGbZV/GzOx2eT9wPXJuWJi5lCODYGigVmZWgk1iARXU5ffmO9yffi+tWYW1
8thJJAN6LPdMEgPnnOFHRteGL1zhezptzrYF0zyeCCUG4ohZjLDcDxfXrTk+LRwf4uq51VCFNnJZ
66erW/vYNmzePP9L97hKsr0b4D0aeEHM/8h67D7st2ginH8ZOIRS8z13jODJk+uyM9ZQU9++kbdR
JHgs/0ffasiVl+cLZzTrI4SHKcn9yo0bjt8SndBRr/m5DouzLdWq+B4AFX8sMXlvxp/ZGDkqq/A8
Ev0oFo6mp/sGQ71mBtFwxJwISIzykZh3Hzp7DgCcx1HTPsYt644hp55Ww8C/DDnP1MgJcA0FkK/1
MV4AwZ8EWjxi2vBFs5d5HQDQZl/0Xaio/Gm0Ca75zQwqUAJoOiM4gaYmWrusn5lPtFdTNdv9NEIc
/745myTSC4MYJKOtC0zmzpR/CWrNVLO71vxpfyPE0ZNGuuBbbjkUK5kGNOdKIPish3zyDsvNnNYj
RVJc6eEWGskVMv4wVaIKA+nCd2uBqR7Pq3AIrOl7lI3Xugik/GVy6tw/M5obi0RFMuY/S6BV8b0a
w/jO13lioRbfWr45haOYYhEvkziLAMi/gtJf0/jxIq8J8o9Mhy8Zea3xI2yVeLTBik4lwVdy0H+1
3W+sXTXzInvRlM9e0qOxDMui7D5zI/EmUjMRM1Bht3T0Byo25qgBeJUMuWn/YXoCfEZi+zo0mqEc
4i/DvAOycyaIKYD7Sj+LifdswAlHALmtXyHGuL3IlTzAWhJNEC3OWJL/t3kyyahgSenp0ZEw61ZM
G/iI1LrvTENK6uxyp/oPR/P8PITCFATrVF8PKjmA2VQuCnzU03Dqaq+qVrT3L9Pzx5SHvarSDvV8
mHOIDccGvBHslsOw6oF9zc6upqPw2X/Ng3VDefW2W6jINo33q5ybaI41+NMXBOGCg48h5RAo3vMY
jirOsDh2XG5gUC0RuDLYAWU7gt0VWSKBBITneGOaJh3ZVi8KGAQD99DCrqMrk3U6ZyOITIgAYA+t
nDPvVi4c3L7/n3b85uz1xx7P50NL5abdRTG6giqJo8XtV66GXbAeHSg3bsGvuIp7UWmAk7mVGArS
PT+rUV2VothX0CORb3BFJi5xHExuwOdDGhXVQ/ntMXpz82xvcc5h1dshpLGXopUMt+yn6tP7eVuF
UKrm+PfUBlw3Amx+3m1YIuX4HKQ5Nq1TI8ksFjekqmZhZxiM6IDlhjSVbLFcbMBnVBStOI6x5L2s
2GV+1ZhAlbPvK90QSM158L44We+u+KgAC7sBMcNOjp9jotfMxl/CTgQP0N4D77BAETh6Tex7mROv
BFOtOExZ+7L1GeTfGavPtum3+MzdI7YlGby00jAVB3BvlZtaV0q9e36iQSDOYoQjHutgFh7KKwZs
EPzF0TQQwaQiNfTd5/NvdMcSYB2m2mwUk6+mY+7fN/8K695hQuVLwt0KlkaG2ZEAg2rQ41FXXNoF
avs642Bow4by9rs0Nk1f01ZNKZ49qe2ydvyXNPvUXvY+Jyz/9rQxvlTmoR8wobslpYNx3jSJykgI
a20+Laa6ePuB/QntLdlR0cCLzQwmsfSf6/qEBC5F9MeulNtGI31MAnA7OXL3DJsbQP+xfbRbiVob
EB6dUorU/eEKzAoAZEDM+9ek+VfSB7fk+iyyCg3BJQszPUmSp2JeCP0pG23Z83IaZqFtKRWFCKIm
IbqbkO81E7gnozOh8yXgXEmvj648ylRK6kaVfk38VCfoxS4vfcKxWIqDwaQK3Qf8r1QhVoUmDiZn
3CeMaoX8c3+rmlTV51eMEt5BpcCWHhE4olJabOLq+gIn0/1nuHq53Gj0HSnfN3Kyg0QAUClqn5Fk
Yu6mlOXy8Hg1O4ZV/13zSUPSTIHsFcertIcXfaCtqqA7EzKPtK3rcB1OxJQEot2ifw9MevTgek/H
lcz2sWB6TV/hP7pcEKjoFvDdwhUYI3csKFC8ujMp0v2YPBCGwZv51ohllXfET19tade285guUsAY
p49UdlYvvNIJzdSzbNU5QO1i9KOcyMgsUqU3O3Zk5Yx+8kpBcdxGjJLdL8EfZAgIg7W8JqVWpgdo
iXQkKQ68xBCHYHiLXat3bgVDTyuHFPdpXYaJruM2EzZ2JxX96A3UfUcdh55Shjc7tVVFFhz04RCu
qiEe1VSVTeMs7X0w9rfgM0CE1cMPxnwuGH1fh84Je7CpYlOfhzxOK8R4kTzITsemMHUX/fjw7aL0
MeKQNzSmfheoK4geXtW+n2W8OisB+aa0iaOdNM0if9JJMlAZUUJlfccV1ltYoZ1Feu+DDv4mPQ83
5g1L25O2QSOzLBrv7UsDEWCqmPX7k6rnPjpLghN72RPHd08l7itQZHr+zYuIqTYPlU5H07LrI0fX
Gb9zDZ76eNf/7CtnYpDQm1d+e4YYqDVyvdAy/9cZnqo+4lJOLENqtAeIP5yBPfe6jaxomgKq1hnf
X6seuwSG+ndjKqAZacbJqnirtMrE67qdrfgLeXGpTWoaduQVCzjAeqfwQM3DgbpkPbqOj0KV3ntQ
Yo+hUjW6ob72+751swgquLTxewF5XbDyVuCSg3yzoO3T3gqbvHn0Y+dYJCYkCPlZ4JvJqtViuxPs
xjcy6HRivalELi8s9B5c6l8l+GOWfxdkvjPvtTQBvw9oYTvBnu+Gr9VT+IvtxE6xR88UVjoX9cIo
qKGDv85/1S8GDSk3esSSeWS9L7yVZX6shSnCDMWJ2//s04S7nRINdzde1wUbuUpoc9R90KzpTq87
piN2HyBIKAwNMi7e+kHYaIOeGpWVM1peSraIkGB0bPO+niePOIYPc1fWeyvRxMHzrFSgzBVqkkoC
CFltFrN+90jI9cXKXLYlXF+lYG8FOvvY+Axvu53gUmlNlQgClwJcyk1DgTsqDagUvWyt9ezDzrYJ
HHUEXKFS07JsaNNNvJ/+dEImDDLypQgLfB/5W7AcCfFcjexYpNCkBRXxCPT5b4NY1veUmVOB8p2R
D23dxTZFLk/CoLpkMAxSsZYiVHoFQfHtOQiaA5jGXhe5NZD9Dvb+H3np3tjSIg26Bo2gkobRgp0G
XhOCvo84fOuZmnCC5Fp9usrJy2+lYTl4GoUNk+QHi8hxt+DAzzI9F9+6ubeoK1PpQWOh44P7xrxt
XY4P4MDo0tDqZUEDiSZ/EZ3kgOhLAFs1Q0Jp9nmxDXBbR85o0dpl079mEuUIUAGMQbpdSA5kk6Fw
ssvuhzv56pOD/Fiem1tIshKx+NFURUGW/DKtn989GtGXhxtk/z9S6d32OH4LbpnpvMB+zQEuiJLs
EwxRs1CvvSJBEvc31wtCdo3UneGpSZuE/qdmNnHY2On2jHsboJ4UeNWFHHiz24+NHzv+oID8X0Ih
w9a5cwADA85wwnym6H9K5ePIldYJwK37cRtr+SKZsEb5b7bBa8MZaKuw4uFwXnhfN6lgVhy2jWij
WmWu1KCj1Dp5XpqZZTdPiT26WvkcZWvCIe0bwvA0bpAjH4DWF0DMc7zZwWliJHdqllkIBfIrcdHV
J+/iKAhS7VlrMKyVf8f9L0Yv1v/N8dqom50xLfrsGBzSzPpJi5LOpAfKoQk4bXLY6nkch/poiEX9
duWrMJGEDSU3oikc/HhOnIdRyxTTYg6fNhG8WlKrrNqnpg4Gc39NoDMtEh9uOvIg1LBF3OhEIA++
0c72YukPLQFil4u2qRDL2kawdOLBVJAdIToFJ/hsp+kv6S5f0nRHAhv/ERr7GGJcWYUcb06Fe/1G
UUt5QGZKVdzodv/lekLvWAcu8LvjRHBWTUYBOKWhCulEkKU6QSZKK9l5oeLfLaVyiDGWCle04INV
zjsSHcV/1G2qPdIqKMjaWHTR5vXFDiJnf6UKPJOFJOt+AFSYlC25hpqXFO+MPccFkv4PyHcdXPOJ
swyooX2X/IxBZh51H/fXIVw6DD7+R5X3Rl7x4qJv9huLjgfeKExkLJDKIFH2xGTjePQD39x0P5PV
5+RGepB8tVqiOF3NW6UE+594DxAtztF0LFvx5DyB3NZ1qznNR2jdAxNsagR1g4ubJLo/B+m5F8KJ
9bP2R4yvQduvvYc2VgfNd/YCznfloyQMGZz6jGxaULNt6LeUpYBKfl09ztpVmzD8DtjllI1ptLK2
9WgpVJ/DFqww6oa6v8OD36eYhceKkWPBCPqvMjWi0tlYboYzbsh96wENe2mliGQTfT5LZayrCt0e
dDEkHpdkjUniH+qnh0SmHgCHT38Kc6zeG2rxG6ffeWjiDXm/dojOU83k/36epzuvB5SA9OaSmBNw
EVxBJrZTH2S7o30vqMPXin2QIAXpeKF8xhG1mgJQYkvcC8nKTFR9yIwi0fQdXffPWxUQcLetZvr/
bVhMwLkS96oVAs1hS80BJRZvzmheGGDItHm9qnAYmIqWtaTKl2QY/Md5IvgYc5o+Ko7gOX1wppX3
tZLWtlsNm9WBGSgA/EkTN1pGaAxHp/rnrq98J4fKNnIXIR6ZKiBILhp679B/s7aoFfsPDSDPgSSF
g9BWZ4Kdj1G+KQW6zbHkKZ2FZwKAOAkUin1kSzkLU+OrAfrcQSucTPgrEafD3TMQiskcEJsPHUMT
m25HamVknOLEWvuXqY7CW0DipTdug0z8UFFP8N3TvMKCu0XARRL65HwYXzJL0wfDHm6KipxS2QRQ
8D/a8w/mHXku1wNkdtpCclSlj2ozoiCRePIsb/Q5ttI02FDYi2hGT91kbmtbp8YIuxn3IUGqe352
c2Kt2ucfjUxnbM5rWIGGGV01WL5nBGl5AUghuTVTHJ/q6xLfQYuDkFVqprTtP4nqOscQkHc6GKS2
TtHGWspV5T35NGFRl2YbBwUUtkoKzK2swDkKOkrdRC/pRMRY+jKaBg+nuZJOC/rSKAOzTQAS4oFj
a0cehQM+yjv9qc7B5qkylRecrNxtrAjweI56rYdajv/PjHryBjAXlpLc/OUMvOQIjirvud7xF2cc
0ejO1FNnLcxzqN/oisPypYlqst79b+S7eXfCbzXWg2XJ1T74kal/vg6gBof6XDRewjHj/s0eFzPb
/J0tFpd3DZGNlmMNgsrmXS8UHSTeLoSg+VPPe1rgxu6hy5oTZ2IyKX5oAUR5M6HZoJ+dlBkyw/LK
wQSJf/sNBaIVG8XyG0HZoWdpHLTQUNzOasUzSpJrHb2/D2oV1/dt+owGBze77rXRVk9axkogQyc9
u6SXykb4hbU7/Tu9ixlGFtTbsznv1QeH56iKCWnjJdcZXONiNIaSuOVvH8dJdxBvEGs3a/PLVwEQ
W0DF3oHQ8Vx4QOusbe/9QRxXBwbvMsYBYozVtV6nwJK7obzTeg7YJQm5lXRo44NbteERWHGL4UKY
JM0EHX4yuMfRhhAiZkCaCgvax5VivHin3tlFGBdLBvrkqQZDcpl8J89rxGLlmN8wboaM04BBygEs
h6inCrbHHuCWH9L7/JwJZFlcVEKN6oKA4mDzba8sapRVqz+daDRZNOa4MoT5ZxNOtlwpr8qbq9GL
ZiMZRtoJF7yMgd24Ve01VVnpUgLTvkjiRDWm3Yh0TDI7t6sixxfthce8YHpF4O31jBfSx7WgJ3fh
ou5OKuLaXPHS2yppNiNI+B9CSdS4gxepMIhOj3tJFrYfWCjh5zK1rMWbrsQX9unoq2j6sZrp7/vQ
6q9pggnzMzbdgkMSD21r+v3W3Y17iVgrmE/T/OHTnbiNpiidAQO1wtk9bymyNeMSV2/y3yrlS0u4
CYs1RVxGFS4Ok8pOjMRvTonESl5MDPC+hd6caUj5+ICw3W6JvXdOzPFEfBuJuzTEhA2nGpfordAb
EPdzmsUE3DsX/sTomwaPWrtpuwUsHWQNDmQnpmbBk8Y1QMwsCPhk9FqrvvDUuK9n2OB6z3tBkQm8
AR2hdcE5ERPeJbrc1Gn3dwJNauNcU+XKHkIp6UOiKT5FHliQNZ/Abi1vuJAXtWaqf5bMieEp55Dz
WsUqp1ltJFfis69+AG62/7HR2PkQTA18eNgDXtS2dwQREulsv6O4QCFaG5Ii28VBZ1ixpFEgCUdy
KedL5dHpNJO8gAJDcouwy0hLrjfoChiIBa1ZHsswUaDdnaBs4YR60AErENx6FVH+rktg5IIenMNa
ivaE23LFuhzTsAuddWB55lL16G/uXL9/wDcL3vvGLuS0iAfek7HOVLC5632sRIZuEXXY+SZ0ixxh
zWWJUU5D3d9J9N5SAMYTHCDqHGrebFl5F7u4fmqo3DOcR1oqN14OG8EUfW6XMyKQpoRyJrq51MvN
Tej9mvp4ti2wOhekQFHeDziCSiQDoPZL2quyOgw8btXWVAVKKPqwIW2oWKj5t0OApzfCAtGff+0q
fO2JZh/zkh/pYYAdgyh1yVhJHgM/AxkjnRNlKpe9hXrezVEF//RM19t6ERmU4iUOQkX61mq+Vno4
lTNna53zVqA/mLw9bMdEXrja+Xg6hovKWLcRyJAI0YegpOFR8EJtDJI6/bcimL2NaHdjxEKKGMq8
Wdh9bHbJWQBUJrMp/zvwYVIRoEEpDG/MemR6W4jhxk3AVRPbK2fD4T2UHKnr8IERib9SK0IDqOIT
qspkWz+2bcV7T5MJJDGvD1MZiOBQFt4SWV+k3ofqKVASPxT9618olLDDQPAb+6t9GaL5QFMiS+XA
GKKQqB/rTgaRx0vgdIBVyEbtCPaepODKdeB0EzAI7tr1pePXx3BzrtodmvP8YmWtaxmGH7kYye3d
gj/3HSyr9y5gQddaTfgzFCilKZGx2GlYarDfBjfT2zeWsIPdBSsq1vSuc1FmtX+HOJ14l9W2PGZ6
eXlaMgttnCZfqEXr01o56HUkQO05G42e5LpzLmdw6D1uAvA/DP4dwnsAK6ReoEVZkqxEjylavGC6
/9riuHxf2stteDEIPLfDi7DLY1ODt00uNqiEd5Nysz0lTM37RCfGsWcqpGadGdI8xtWBr+f61PJb
DpuQbanwmdFit/dWyplzaO28MSVepwp8oP0cftWkjGRSlAEr+YJcv8Q6Aeqp617cK7hPrgodA8og
tU+JBtz80uVr3j0wpj5DGhHnnJVoknUcnUcR+iMn7w0P7F8f1XiY35GgNolGBn/VcxVN9BsOIh9Q
+Aa85HArCKTbAQ0O8hbB7BUCtC5pNyPAAbpSjSsqSXLshmTZ41UFEtUQi+RQHBOEn6XgC69YtMJe
lPEgsUrpIFTel3AHSpiJMNusl03Rrnp4plvUlNEIwTy0Ktvmt5/3AW1wzK3FIL2ou8PzqqbhFqqS
T6WE8mP++1I9TvWGEavqQouhrYHEcAU0t4CAoypQkibkow54zk0hmcpSXzSGR129j7mdP8U9liJ3
giTSR+7Bp9rgNq773gDHn7rQPIrsvgxX4i+fMVFSihZzcDrZlRZ1rINM8v8RDseUmX5bGiPB3BDv
EH8xiH5eVYNu6Ckuvt0WKFvpq8FJpNhJLjl0PSyN3zWdspU4CDOENVPqVtHsLP40BusT08ByWSaw
LoaowGhHHunW5l4MraYTkcb+rPo1Po4J/vz5fQZiLdrKYylkZipROrR+kXyEJScyfwZG0uIVoORG
BCKWx0/2IGQ5NfAhJ/4B0Pxfo/jeIPsmLKJL4a1Re7nAq6bEzQR4czhp/BtMc+33gzNxSvlV4s4k
eE3yA2Wgpyj4boS3aaq03QiuLYvXD1A4TM32HzKwkongTOWQq/v6tTXnloSLTQ8fY4BXLW56H+Bo
QV+fTzSLjQE+xTwoQdrs3/nkYkK+cej/qtUFFmljBchHfsT1t9y/XA9CV8/SfYU91LR0VpWjVVxK
5hYyk1Vj3DTWqoDjhWQ9nBvXB43QgVsP0G4orrR0x6wHgUQBCUWmGWLyafoVAkh6nheOHTpQ+6JR
3hyC72ilCcipSo5bDHT4wOx9BAm1nBLgdSD+UL7OSwm5qx4fGRfgaEaRkE8ONRV+N7cpuSLIOL3J
BLBEvAxGOXp9WT2+o2PlLR2tgkysQa4C+gSwo8xzVs5sBqW21xcLnmjIhwBa59CnQ8A+Ye+qgIcC
tQ/X/sqiUW1gRG4GyzXXqKmB4rx8n2XBJjE0QOCWAPD+phwASqPJ1hUc9K7qAoKQiymNkLUWFZHv
PFQDIfQGh7R5G/dpKG4GfA7ioS39X+GOMwydjRl9bgxM3kFGAo7nAVzqrsU+yl9RRg70PqN0PqLa
T06sA5tgpOVg6AuoX6proYuiUPbiE+ikDmmHqauL1fl+USnCCiDU22rxj9ruN/WCU85f2j05aTR8
6FJf1JdEaJ4EJEOSG1CaJHjWnGfat8GmX4212cK4QNZHPIqXKssizSy+VGpddNOnLWGhLcPsgjyA
JNJfGqe0gZXVUYTyy3jlEIIf2dLiXv8dGCr9IVGqOL2Bx+t9S7OhsCAATl+HD09z3/atPZvWaLi0
3sVZd7WPgcr3jVtrilwYbkY7CkSb9mVBvy68bX07cMVGqgmvyDj5eNcNiDyqOkQ4bI5Dt0LNOJoT
kIEYtny+bgg+Cio9prP15cKpca/DCU9PB3HT0GmboiKsACO7V8ZtW5E2b0AC3G6Op7huV7NSWeNp
Gg3GFNLJPDey/+VDiIXQg/NQXwxAxk5YGkcb49SqNoLto9bEGGnl77a7H26NQ+9dUxd/TY7F/nQQ
8i9TlnQzrO3yRehHaO7lR124VCDGWono88um+OXnx3K8lqN63TUt78tXz9l49Mb2F93z4O5XqR6D
jiG/cNcKPBxHFTCBLonJfbKCNAHVgksUpFlD9wxYn7sQZb1z5f3AYuts5QTlSEBw/kcIlJuk0Nk+
ZELEa7RJOF0CZJRte80o6L0NVYKs6QxrvNyHTJ2UuEpwa3zfED5/LmT5io3iVthFNHKWE/D+IzNn
d+w/B/kZEgEu2klUVEaJQ2/YR2Z8FQkZEHhk9bycfqT6ZeWnwx0Rt2xTV07nsnds5zby58FXtx8h
aZdgBdanoAvm6dAb1au3Izz+JMGuMg0+ZbzCHftlKg9FS6h7gq/uRa8K9/okdSvJb9fy0/6N5ukc
t4gpZ12E7BjO3gLOgOt2O3WOOm9xmQlTPubnhppE1Q77zK6GrJ6Q4PZV87fnaMw613uWPpVN9qKM
o0ekRd28W/TzIV1gnGaYBkxT6KiVPCWsOqCjCBITGBc96DauFKh15EoRUNYMtf1XQh6bAUCwUqka
IA6gayVzpk8qzv3PzjdUYQ+UoHmYBVYNawi4nMVG4mi1lrervJqOK/2HhOAZNRCYBVMB3I/fwi+J
L5DAuo6fPzwIM8YyAA2deBlAI9RouQ4TDD8bLOa4XBF///21B1MFStftQT7eSRy6KZtpkSqTk4k4
f7Eotdw3gaWPym05zSXCo8MaFR7ef5GblqVkvhKPhHG+8dQaSukFNOPmmvj9NefawngxaVEptzK4
RRo66sVeMAwxackcOSwOUTI5A5AqqF2gOzd3o7QxsjBRzRT+DuMYvIxfpWy1GPMehTpdwl37tRs4
U/LwFz1T2oEDPymxJ8zyC2JJKGEFcilic1QXPyOELlYjtKy7XtRAUF1WIRFMJpF77V6OV8j7S42N
59rWb18lTRGvzWgi51P0CJ/YYrREPZOBXkixwfK4y0Wtp5iLQFfqk5DECVwIkj24VzoF/MN1I/DW
eN9xM1x4Gb5vXAjDPtXJxHD/jP0ty6DNSbVsSn0umh/c6/ZyNqffLrtgis2SJaYP6F6/AT0Cj9dR
CiWIl9ZdEOjrNNSPEoEFbIFH46kR5Ju4nUp6cJoXkUkcFftqcACQOm/QFyL1Tj9b/ojf2lESmnAz
w/DxqKYehvBvQzMGQABsiwnlNJecErkOa1BzJhMLmin9PrHpXFcW8Se+8IVVUoznBt3ayMjtFHbc
x4O0FVwlMBZ8zhdhmHkV3Af9Oo+SGMFeaKPKPuZGDa3VWsMV88eI+Lc2WXtpp+TmmP1w+nurlAsK
+ckt37Ic7n2AKG6Vy75ivtJvB3hDadjtZqwi3chG/CUqDXKCX2ZPtEv4BPcafp1h99jRItnBo8C5
b+agIf61trugNTHp7Dk4rBRJXZPcugh/mb9JMuJmlXlAW9C0uDrFeslGHwZE8vdnpDJS05ZyX18e
a/OyUVdJw/DSOAAhpuvj9LUP8gGSYTgX3bH1v7OYmCc8EHfKMxh1+cz1Tn3h2hL8WZ2cpdyC5jQu
aMrhY++TLmMP91G8gY87OKir/deLXGz1+7RTP3Iai2p9UJGdXZq2oIxpZUYwsZG/hAWwZRv7C/oe
dp+d2nXvQwByMCCPj9jKbe7qQguqLTa3L4UFOo79btn7X/QInPYuuvNHvsd+WUnxMDmjoxzSwxJH
rscRIBe//yG73CwX8asfaugohcdaV+692Jv8ah1Y24qGIUjyZRuIqMT5GudJn8ac0XSyc3t9kNYV
4eWmSgsKNcIab4MH7DroW19tBIGnkopKKrhjzFYKHEXQ4KO4zGmA8aclZP6ye7VvlwExxDnfg7Tn
u9OvvwKXmb40uXYWX9lmLnmrk1OXizzWV9Ex4KNsS9vvwO53qlpPDvplh8mdunnWwOSHCwukWnzv
JFsvdMJeoRR86ccDaVBBkTkN9Rsfze4hjRZXiCww3CHUzz9+v7N9bAx74RK1TPkKoCiXgcbPKGGe
LpNO1/VHBmk1Q/B9UXW0Hefs6aprxO/7qYjf8bpAG3f5rzkbqzcnFuLw3FBzosVrVJa/VfRQOU1+
mIiQBjhXVb5dcNZehA9qg7xIMbsv/udMOCCGo1+Nzbsd8nP0yPj39QmqHKuFgq4s1A9j1o0FdS9u
CY5wmMyGU0QyJ9xIujber9deUjmDOGtQMLOpnXK8SDSAYc7ZiLFbBDedU0iEK+Xkog8vysw+cjXs
4X4QFTycWnX46VaNbYwoJXcLmEDHpzzi0CA1+HBtY7qb24fDZ4dmFVDFdB+fERUWLnFcs/glfg0a
vmwSVrqBX9/UGcBZYJHkbc22qomUd34WELMXH39aTDG/O7NChP+HnwRhAZkle4bvVliIKLN8JmwH
5IZvEBhUwoQoX+NNOBm7gBnjY/sxgB1xegzI8ZBnGW6k/OAfWXtul8i90d8NDAKk6rFgzqciWHhq
SEoQx0SGF2gDlFu3SnhHUOWYA06t1SyjYb2hqob8vBv36EBeVPTEs19H+KjHIz5oxNfsyrXdzLdD
zwQSb9DhyYTqq8FRduewzQNJv3dVeDsj0h4jE1nZwojbgtdwRCcA5FQMme0LY8T5qWLoyFkDLcU+
7KHyYAFx8l776ZcDIxe0Bu+SHOlny+dSS1mOCowgb3P60SiLzSn+Or4i4ixD1satYPX3Lbe9OIec
zMiLJOnzbRyvXj9La15NSGH0wMCXtn744QlUtsMd8VyoZy1413WJnmsooHnwyJuEciMlg+es4Qsa
AxzBGaYb+jo/8EKyIKTSRgQCPaU/4Oqgy5MQDz7GlJCuu1bOzYz1XsCb69sxoR7U5Lyfdhr2CYk1
6FDaRPbD4ncaIrk2Cmp6e2lCvV3Sa063GuWj3qYfYsaPGN7UX6dROSqQ2ivKJKkX5uHCo1p9WaKY
FKVVlQbalC0AtjmhOPv6boEX9Uua91yVVVHFBravryzh9djgKqIkO5RVTf4GR9tT+N7ioxtFfPnS
uFOL0Q+i3vLDdS2AmllWobnbh5eLsB20ia9/IwyRtC7JF/mi3ctVQ/McCTSI8RyD6FQqXJVfE0zO
jrzdO5yhecAotJ68Xup5U2PKbClhgkZkC4tRB3iUBEuPuewfB0VcVpcFNPqrAz375aTKVS/UEXbT
qz7PjZEWT1XWCvJ/cEvQfC9jRR7Q7qRTXVR1KqUu79sPhu0zhhFFP1AeMOV4rtA10bT05G5XyzIm
x39tUvYVbHn+XQ2ntE9UemFCbAA9If8xRq8rmXCVgzEe+K0S6MqrjD1nHqQjqPsBnTFuQ1yguoeE
gkCUm/xh3iXNMFBGCuu3++Tj7EXGPaTHwnd6/tme3XqXwLgCf/8iuHwtjZuWx26uV6/0GMx/PxpZ
Hi+WOb5HP6E9ih4MhVAPEUCS9Fg0mi0nhv6EYJ1wDSD0EyvScb7ODHWI2mYH1G9rq4UmvhIJvDbs
q9BHTNMHiGoFkXh8yiezIwDj8OOviU/j2T6YfHO0DWqcSO6qN21cr3euviaJatDbFTSg07ug2EiJ
d3nJ++8cAb9pPHx1+Xfle/ST/KBgSbjFTEMGZ2ftPe+U31auhzJlwG7hpxFW+01MjHRUCvxwP47F
C/osCWgXUjmpackq7HzQB+eZsyL1KhWekJYErXMu7T9Al9yqsmKs73R6uky7Gm2bVDf7iWA3WEDY
I6dIslBrT2y2WVV1wT1RQB7rRNVttn/iUHtS+lSFAkzGoKhEmoUAqUMG68eCJwpnfc9zHGnZWdgy
J/kUbSez/IkQSzGQwtJFyCRCcKSi7i9DVBoFnpTlIneU6C7xhQ7mCDJrSIsiXpZS10gTWwfwYNWL
VR56AuYLkPnASql4Q14tNZi0wKaq5smAS2p6nkFjM81V9KTrEDdGJC5QG7tnfo+3UIPl4R8Jys3d
TsRA0+arJtF2S+QqF8L/ru0kL8TpDN4MyCPjvOZOuQnGNCIfYQtgv9jrknauJvvuqpX8yFtUZCNn
7Rg1fYf3ryLd8PzsGdM/mIkGWocTMvMwvW2x/KkR/WFpZzEGzCDhWd2XNrwj3uwf/7z9d4BOWwuJ
BTUnPE/0wPZWPRXj760S1dwgnXRI/3UAS9CyKQqiyfL7NaJjMX8bDPUvfj9Dhfyxtwr3kL+j6CcM
oioFxxgl5JFLX6+gdXYvasdMlTzW7dUcp1Zdo4hWbXeGrgt1ZzNF58uB8ZQ9yO3qYw5NChSTIMYo
u8zx5lNxjALCxIHzI5QDHv+vF849d+MKXXMwe4RMuy+/hQ9fmByrKTdniN7ztvNTNIc//ffdACA1
EmjLi4N3xWMSIsgWQllJTzPV96OcJVYopVIo59stCvpVdpNbXTotsFfI5dKXZSTZq1bPs9pyH3yf
YCLQQBQqmT9iJVryr2dVK2t+OnlaSJ75tT2QZmOeNIJDHEl59J95PFOuiPcMyiOnjjNpvSDrzizN
1fDvHPH+Hf0Dc/ahHVEAoDiL7uH6UfhZlwOTrrqx7Zw5cN37JVPLvir/A7pbpR4oDflkgtIprN6i
aZkYDWC9ddsJHVjHpc0CvWYIy38/1m+2ZJ1/dLqXcATwcN+MCL2OH0355THPyWT7tzl5AQoGIR2q
pWkYPnRxATfs/YVq1ysI9vo3plmCHlqoOUXa6V38RntKRO/Z8BAwwuQq5yZeM0aV76nQo9ii3lMU
3igjhoC/fhROXFvo6rkiIN1Xn0LpuVHAjDuwVDMFp1bba5XIIanCjgeBXYWmwv1htFiwoh4bFlSE
R94OFc0rS9fcnwytvK9dO1IaEJRNM8mXpqObyRjhaFY/0a27Liujlxzc6qSxGXmCh+wEMxMB1Lxj
otWQSFY8/f4wJECydx8k/WuYoeGuYbIq/RscankdrMbK3X99i6N3LpHed7HKP6L5eb2jFWEo3gtP
Tik/A/UOzzP/f5xdZFwq6bJNHv5OexZqfR0mQy0HKRvvqamJnzoNclmEcZ+yZDR7B4KMC2oJUg9w
v7hXHRW3BMoDRl9yjbgJMMZQu1PoO3ohhylCzSkcGfP+iP2SrLo0Bk3g/HAE9Dods+bYPIS4ld7d
sLUqRKt6tnnvRZwJzjG/asqUbxQbFFqpYuJm1OEfXBCgit16MhcCgqmt9u7vv/EQuYi+Rg0Jlx/P
JAI6i2/0Q/w0PUY5HVQK95BMys6YfO50j0XKpuCrEbAc9J2Pg4IhB11DR1LO1W23lsjRlTEdOAvk
SjJrInUMqq1lEH5GxuHN/lwqIdQvUSKPDiYKcH+W+vmlGS7Vt3MT1/gD48LN9f5y1qrmYj3izj3e
NYPehpaNz5O87L7rEJy7t5IY087UzIN0w3ljaypIzltBRi3qAAtVe9TXXHF84MyXo0079GQfYwKN
60CDIF7gDXc1z/suOJru0J5eKW2YEZ8pkemYaifTr/eLufDHsZe/45uxprk/GeWepchOD+Zz9zSC
kbcOw+e+AE63ueGsdmtcyE7wwX2vm+4VGwJF+5Xj61JNGeOoAhJdHDrLORwK/Q720A57I7UyytUS
mVmWMucZMUyOzOqN4Zdkn4OS4+GJUbXiP3a+C2opjreEFhcNAvwLbSTETh8nSZmUyg9YWREQLs4O
TOXylGCo3uxkEMq+lJ0+TX6JYKP6rOLDea7htZHwEGHMQvK5z1161JAtPBH7PD3Dxb+7QCEgqXt/
OL5gCZ67mvFsQ344Pr+HOTWA+Z682HeLd167Iw7t/MUH2BTAdpXPXFg7HDzszYyT065KIx9A2GrS
Gp7Ok1nIWC4Z3LvlcxnKYV1NDWnoHLRgeYTzMJsJLf8e6X6Wx22RBvsbbkBuqymaABY4V0YuHsze
NfnMturMoTu5cjnzJ1o0cUPqGqxsx5JpIB0RzTinGFayT5hn7LlLToKyuiX4ojlLZQgTnaAzXW44
nZELZuO20L0pOwwwKZHRa+Y56zoOmipzr4rZybyKWYFrhjAtJx3E8dLfsZ4V047AY4LVF5CO1vsQ
g8SaWWFd0Kwstn2kErVOmLKRmaxyWNY+PyjNlGUyBIk5G3LkuWWVzT5VflyTyhx+lMFP4HO9n2U3
vFVE/zoMTXfNgIAwUlX87DlZweU9V4Z964F77m3jbNFQzBaIQQnMOF6VVIcSwKVg9J0GIo+cF6cm
+xHrk6b+clzwkiFy6RFyfvuAZIusa26PjYim2nJ5lhtG2QFuLXhF8StcSSRU6JhweiuYvtqVWTkH
XIaSRCvVeJLA7RGKjskbW8xNluS5quj0HN4VjXchzMZJkyp8qjRWJhLWjvACt7vK7rYo/ATvrXNT
ILCKf5s0rPwDdzHbH3IFWILZTqpjgwNaeQTijp0XBY4N5aiZjm5MmkIKDI3R8Yu2RFv+8BKl0w//
XWbXeCP0HY9bzX8n16useUbxyvjFZgtsTR1yXdvbPOs89UFnecm2C8POsVPW9gAzK8fLMISsAOgT
xj4HhUzPugCCFRb/cTA25HwMxrhP8Hv2Koxe+8DGbdtZrLbJGaaHVadN+xFsPBf1w2fEGlHcUs8J
IQ2sjgmc5yKYFoYn4/fRAWuoe6js4NSdM8pPKaViA4iDI6q+BoEW8Y95kwrUEZuxRFJP40g9HyA0
BIabVatGVkV3MUvgDccoJ6dqizlN/rGNIe7fPPGhvi1xjaHRH0KN3c/FyMXLaLvqcQjetIVoO4SR
lh6QojlsfXEQkpUj+q19Tnuy3TZ9w6CRJ9HEMyl/ne/sEVDBPCWg/rsem9YbT6zbjFYiH0D54yeT
ZffiGziikmheUZOx6C42gI0WsC6peWokB+HH63pjTHfWL+zUFaKZowgw+Hs2uCTCJ47uzu27QsBZ
jT1zmpcex2923+FZrsdyIw7XdR7LAYGbJAe56EFkiZZm7XNDiLPllocfX5IUk30XZduP9amEz9by
OlFtMXulNGdjJA11HKAP1HCzAY/dQStoTYJYUT6EIR18ubN+U8LITaWLPgsNSDSwHUZ1/VK5Xpme
SWSuBathIMtRJ8bo2If1/mVsJBubhziIZYC2resTpBWKWcItF+ZnJ0msoIpw54Np7pIvF9p3S/JB
2O0X/IndUHq1QfCvNOqJRZs0kFdwFsxQE3aGXiFqNIlL+JsCSYEROLsYV0Cjnr2hpNsJLZsSOzQC
EG9o5xPgr3lRs/kxxFLsukGXwQr0Z9RNMvLo+va3Thoa16lbOi0HqccebkHaA4yPoqoYELVoWj6g
6GnSBUagLILmQ2HDBEztE2W/1Yla0uvt6euCBvJEuVma8HJyfeoWcVpZ0XI98ovAx6WC8foWNSgv
ZsT/vHCe+JlmJUPMxTZWehA9H6cNzP7iCndJ6oiwEmNg+2dkNWJ1OoS3vIyzK9jdAh0tgOMWcL/o
vf2LKQIPRJ0i2jQVqNdlPWTpsoccB7AZkpIt7q0qw6hK71gV+oBZnmmSyhcjUtqOaOKPEetAB7rn
cZtH4Pr8PFf7tBKeVig6bc5xd+AwkcqXnS4cuGw5l8gpZNFyutUpMv2BmvK7R5XsuwnEWd1lervu
GM0dVnP6xwAq4lfp77yCg+lrtwl578gXF0lBBCKMMXMqSEqYl478qquRWQJjxkTkww4TMGILSyxG
6KKRGPoZg9HY+gVwzg+uUOsGFaPNhFVDrvDnsKKywdFcezHoLghe2JvQP9dDGA3/pEH+wwzHtrEY
SG6dAMnX/6L6ADHQr5FcSEmKcf1a3aKS3I/fnPmtENTtbB1OKd4K7iAmpPtXmDdsAdj7v9FfIqJK
LpYSAhT1zk4O2rdy4nh/jL8Om7X16YXHm+EFZJq7WZebWE0BZ0EGdoOtHr9Ki69EQKIV4nKGrae1
G/SE3lwqy+QxuasQMhu8KZsK0va0CEBzWH3XYSUavDj/UFRBRDMlDmlZWfELVZvYSBaKSQltD6t9
1oRHGiyyNrv5iCi+Xj4w+cS+lFWLEIyxRCfrRTAe77iZkum2PaaWs13sOk4Pd34yHzXqBecU+zJT
wOkp2yaCN9psJM97AevlEirf7N2SfuiUqd/zvAlNj2s/aFPU/D7JoEuCaa40wHgvAdRMdkxqdbWL
MXIb2EHjDl+xbaYfge49g8Wj02CyAIpDNPngwxzuuHPuUZ7SPTLirdAgcnt1dDn33MfpAuiYjw4Z
Wr19QVFcjEk+N2D1+k2FfE5XJUXMuGRpcB5DOrRgAlJGgDxyua3ev6pC6ZfGsS79vhRim3wlp599
CshWPhu6YoRaxippr1Ab6fz0BQOQTMargDB0m+50dTDidF9xabWN+rkJHWHTV5MTEaqOzpBsKj8i
mUF4oHe2vhJi0jfV3gdH38EnkWf42d/nsz5PMRhzLkeDRw9f2QIjez9p5u+dW+muWBCNrhFK8EGk
CStlZ1sycDfuIu2OYnSnUVwzDKr9k2zfLwtABx65OAf/Z5aU9AzpVJIj19b5hgtsqV9n0r9j2H4j
krHAO9FIsbB8aNQmsYwdWpSIIvgQ3A2CTEEhJn/hLqFCyZmEKityc9RO1DrlqqIVVGifbenCb+WN
gKG0L7zgjvY80uNNFU8+hEvmTEbj58w+pdmKcBQOvSxTK9AC1oJEoApOgqNDXVL4aPXcrGETHdOa
Fi/dTDpfv61SgWZthgQmZvJ45/xbl7qaEwcVZzX0ZvMzzzJMF7ZBzO32jCjN8Ut23RRcGr/Zkrmw
o4by203tPA76Bv+NOAjtzsbDtrAkPny6hWEc8UgeqSQHF9CwJe3/U8+pVO9cQKq3rHHt43j7aHJt
2zQE+x5kKlvmx1q0JFTTYj8fZBL4wvlYapvNaW4l9+OivPZZWcVIGrB3lSiuEKetnW6O7AR1UTw0
QlT3Wj924eCEm8elFRjPDqYJAkILvdc1rNaCrZMcldhMV0zwwcudoo3PujgE8bKW/Ad2ZDZtl2ye
iXxOJMpnDWiUnyrpkcJP8j5X6tmWHoltcKUSWvTSd7ySfSQIKYViwlP8CjIZWOQGUEisu7767iM+
G6QEyhGdL53sXOv3UnC66C1xSPOlds9qNYKbMbP1TJN1HjPDk+8z+swtvNrd4ljUgZIEhiM1373V
iUp3SWUZRO7UprRAlq9oU0oGKyPWS33Znvu30VNhJMvJVwucgdXlD9lzArjWDnET+BcYWhl6IYBh
0eWpruj/3xgGwGQMCcL9CIpIGN5/evTPvbR0c2TIE8d9QFbernGveKshaGK0tL+Zg6BxDkvPy5XD
EL1q64ER5Pizh0gO456ikk8V4SdZ+ckTvadEIGm9lPr9DmIRQDg4FZP5Skpeha+SrPX3hXZB/3vP
nKXR6HYPDF4144yMFtTACpCvfiZoKmUIbptPCf/up48h7yk4JH02Z21MeOC6D1d38HlwA93Dq5mr
BFrl6B96KeAa65ic/5+ShYqcoxCbno7I6iDSqYFaM2ju98VEwCeA+Uwro7Q4yPfgESfCYy08ma7D
exaidWOyMxYkFWIGNeqOqV9IIhNPH35a5HQalS+zIBjvisdYePStSxSI/CXqDRVhWnBQr7E+qIbm
NTvvC1H0i+Lwf2Yyg0o4tOwQ+DVlroHoSS6KGnXAB4gfFeQDnWrgn0qn3rAtBWqoZjRpss6uhiDL
va2CTL+zqina3WH+ComLEFf6J19o0IfXPqS4zPhHm6cHth/kcF9OtyBYtjxs+58l4PGU4WOjKzZN
Vq0Cy/NGbG0sLtNI+Nq9YaV3aAALOYInt1U+2t6QNw69+OXpT/JwpgBtXRIANY+O+SHWrYoY9vyZ
oMzf9kB1IHf130seHj4FG0elFAz+2ODTEpJZJW+2k7O6ffqUQSocnh5Q7bkgXWElqiL5cxOFYFqM
CtzM7cpLp9id46XaqsnV57v9V5aphzBrDnMUzLm2wIFREJHywpgEuVuoJdnI+//6lwrYD1n51REE
vF53sX8RFy3I3uFkv2Uk7q2kEJleKgkWOOsq0fuQMIHWTqCIL43rOPDOvkSM/0U8lm/NeMSQDKDJ
s8Bb1crFHcvEj/W+LwPykNyJ5V4eUWvXYXKcKUB0qtgijneCxQNX76M9RGM0M+zDv8ybQi4lFMSM
zwcUZzP55HuonJdpQyFWXIspTlEgvp2d9DqKGnaObMdSkBkYUtHIZ2mZE5so3wlinSRvu8vkTv9t
oCimjpioBT9dsJmo4OMUyJtKUo4CcU89U/ACwWZATBHx3jhbojtzNdwi7vkJfNxgFn+Ufk68Yk9V
IqdKLYzxkB2p7RzAZdNnMOtRJ6GPuPoTHwf5JA54fYDLVZ3J69gPvQsqNHC+oHtHG1dCiDhLRC+I
P/rZMrXGajlGkDe/ceANblqE2yGYvJKNFLIUBKWpjDyD62UuUIIwSxQ0JMa8LIEJ1J+XINaDF/27
Degsdx07HrMiyMOSCF4rAjG4Q3L95oWPjHxQMlADIz1V8V5tJ8XMRCWfOngW7fDn/UPa6lNbs2ve
Fp8CcT7dC2wi/79mo5c5itHnIA1/IP4c8IDFWVkCx0CHuUiNdJqR9GrjRSMobPLaMKylrVgIFNnq
6wcEDRc/CJF47zF2NfXE9atxmFsvoilwFMLZTGk3rAkk5+FrHfifQR9iOsc6io55OyBMCaZfa8xM
M0/pVew/KwzfPqO71D/VParFZmJXnKGSWAFhZASOxuEO8PtRyL4N0Vk3sx2zvfsICTYhu+NHtg89
OsXH/N1nQbpBgaiMEBOom25iC0igTZyB/BVm6QNYFa8dCNtCb3j/b18QFaVmX0VHX5To927hXARV
1XafquBqIKWF3my9glZSC4F0qqE8o8HxQL9twwMVbqguSNNeJRlF3SwTE0eSbgj5c6g7DPBS6cVp
alImc4P/ThDzd8vgOtjpNHRQGbP0IyFcuj7KQUPi/milWP0QFC7VhPyqL64oCj2zue47wA6CJ+RW
ts1WsHJ1gmM2vufSS0l/WwHnesK0uu8QujkWiSPYMX+snAWu4OS+ETgjutfEK11BArgKV2LT6CrF
3udcMOIaSs1wwOkL2pjPWfM7pkMOM/IzyMXFmxbnk/VzE3XklP0hy+Sd/ibPnpYNQx08XEl9LLG8
SISGEVzCVDr+bEAmH0pBDKuAH1fFY2QAtRiEq9760MTdsm/knX7OOoqBqz//MHQeTPP8XC/WJwvf
hOVRfudpSj0eG2tuZPtdlB7mLw/2W3fg0bkrhzO4SVAJ6EjWjj6n6lLYIpzLeq0YOOCNL1wBCJRI
SeUqwG9SOiABgJ1KZwalDN2zqMySORrgPCgl0qeHUcpCeALoy+026KMCQzE56I+s7Tf9H57nGlgX
3vhEcRi0HohNaLxiQNBrJHx3IGCjSkZF8jr3HxQKBuGv5YNjTGhYoharw346NIk0vWUZPF3ZKe3A
fYfAaljwYD6efWtR+4VRxicLSV1H6G/xxvBzucXBBX8ziUHRJNVWqAkRbSus6DxO/12fAa9Le1zq
r8H71VYRHBD9IJ61XltDgTX0Sz6su/8aX+yDvYUtXWeVlkknYCmhizKQJi0xMrHQ0vcUTKHWqggI
CsdSxgvXRuG2jc4iuQWdLXrUJIPgg3DT9k7wZjf4Xa8N2EtPg0Rb1iwomOI2vnAQAghp0Lq+JmlV
XxXP9SqpPqMrbZB6RdJL8Tlp0l+3OchCdlkT1qZ7TRjZWBSdcvZwVJw6wbnUldmCO4abwUmzvnpL
TWp1aXnd2jBKL3aaBUnBjWOBi8gbrdb+Izh8onnLXiLXbAePQzX8aVQYLjhL1rvJYe0gbzY5pXUK
UJ1rhmgWPrWzU913NQU/Hr8XA/dHeqTiTScVyfU6rmd36cBJ+vgc31seHzgzBVSPhG3g8SUyR1xU
OxYrEF6YysrxHxlkwGi7yQ4+9q2oYRmxs1Nvwx6esiiNmbQ3e9zikjvcJ3yRfeECG5O1rQHYx+Uj
fXDHbv9O2WdxNDMnY+IKdDIKRoSE8H0E7jtkT+YYXb96Snrjs0bXpS+1by2Ga7qOnSxtlQ1NCaoF
Ky9ygFKdNJXawdah44z/e/+70Ey4qMlnX6dnkDgh49773roLMHVA/RhKr3AxqUWGd3j1614XjO2U
1E+V9IR0SA9ke5eN225JK5TFriN/v/w5+Qr+wjLQDpkGZzYI55JzPKUFw1qHvvNgwrxTn8bQvXQh
B60RfyWcgDW+a4gLHOIexyM894J0A+45UR/81oiUEOWxxhNt5W/t2rBBoCAaNPqw76ozdXPprOXb
oMQWj0fKmixxackrsVXSxd87PUZA5YTBgrvPNb15sMtnE6t5b6KH0vct049NwAeukLBojKp5wWDS
sfjeKDZwRnZErlGs58x4+3Yq9D5yaWGjv8dt22VcCH6PlHX6Sx3A4tOixJQROjmymXkKHGaKAJYA
R55j9bOrgcIxaGhmRpr4Do3vV5iHvKWj8gwfzEXtMF2RXXLvJj2sWV3YdrAu8f6BZCr8gyNmMuO3
KeBnkqpmlv81mQIIFejNbHL9PMr+ne5Bw1IwwWHXPugNe3hBZZeS5zkKTQNjj+GFqaruZSXKcWrJ
nXg4CypDMruKyuRciNDoElJ14i49OoFqCW0coVvxg5e8rxUo5CueMx2ortPTsAClhfgqekFp5TQX
8HSML1NUkpT7wxuvlo0xVQcoXv7talBWKjy7QvCDxtv/1u9GscgeK6pFQ3yVxq4RHXJwZPpl5pqz
HVqbKr18Tf9rb/6+OHKZoTFf0VT3zYObwFtSokK+ietHzhRsDte1YikCQPh7byKQebtfxKIk/DVj
cJspS87ipRKlbGgARIjjRt30XsWky0Qi8PUppcyRW2K78Q2G2xX63cW7srQlInpz6fweKs+BDM13
qPIx0RI1Pkx+sSTz3efnzvMUIZVg0TAlS/3LkZZdrwgPj16b6+m1dJ8MZB0IK9F4spNWL94Qf5WB
YaxOLZu4NEOjD7sXPytUmFIVg1TSbdKueSNykJeeexdSG2l7u1HLAMJl3d78nEcQ6YirwfjUBQM3
EYgmpPZoPXoRjMt6VyrpaA63wCzkabQd/F9Yt41K2vqBwFrr2o8ezi5qIniDib6V6RmMKUD62rwu
2Z4RYLBhxT+JiB9cwe+bhrVFAxKDV1VoaoevwxfHG+ly1cyRjyc4v0rUHEdOw0lfyxb+YImGrI2J
SJe207+4QwHBQpNnxjFrRavpEBTdN1o+tzxM2gm+7z9USINLGCt24fGTZo7p8gdqnUyVYDVnwjv4
iql+1w54XAOH+xOqyMgs8l/Vz8HKK97UX8HOpW+11TtyCoC3GypunQBp3K43BEQhmLj7+xqDcH91
ZFTmu8SkWag4QJVaBWwcB5fnNrLe0p8vHeTEc2rm+Ur8AbH3X4X/g9NNp2EdXQC6HATMKIaK7u26
vSXtuJg6i0a+mII2s26zXf0O+I194ar+wsgYtZYbCyqPOQsYuRfbGcNfACHz+ouEteTGWO4d2DHb
3yeiqKAaWl1mIgb16j/nEIks2fec4aqFlm8VvM9HagwNN0+E8ZnpCnb6Zki5Inq/yt+nZR8OyGTi
uCiPZvT/42RLeV1cq/4KyWzLnkX7jidJ0QU8TbGDCHmPT5JbYhQXP9UbHKVh84y1RVKbYcS5QD5r
MkedDU3NZ0OSc/rcW1hK+s7bLFEZObWSEohiDrHg3WiCwRgP0O95xywl7ciB7yGFFr1kfTNfLfZ/
StUWj1wFWZalh7rat3UXIJkoGKTcGKdFc1lf4Q9AK6qtgkS7QbPK7V4tI3ELJgOkjn8+/qbfdXfq
oCCP7VVFLMMWrtoZ88nX56SyxNnu3fOkvd3JcNqL5Rt9PTK05uW//ingViJR5Sqp2yGICG8Mm4/y
wU0mdTOXzU2cflrUb6bf+14L7PFS5yJiVNK1gkBnmxQdGB1ZMuistWlNIDhhLotGw5Qc97twspzl
3R5Kj3NpycSnY+dvsIZ5t3+6YqOPEdnTaluyuPeWBcg9N99Ja1VWitkBHwcKK4fbjGbHZlVNab1B
YnGFbSXtGhm5kiSznbIZGPgsnMPblCszEYCiSrGBiw7mFmIw0zNlLCEuLSiGMkF0RNvEGMfZL52G
goQKe/zcLez2b6XOiJnBktnSBUDI9/2Rnbf4tSHCBfmoVYwnXQQzVynx5P7z0LCRWJS5IhXOddbD
pAMZhrfKUsXu+TR0PT0amUcscS8dOTKWGgcH3XLTsPOMWMj2Lc3U2UiEqBRwwi1RUuVJxIGOAkht
FIwAPrSu+G3dobsZlfg39+IwIuqbPYaA8q547IzqfKiLjWi1G3muQS/qwlu72Yfvv4+SjzGFgxSL
K1HhgB2yQbnu68v4aiIfnrL41ZPIoPr+FNjJC8MPYteaxwXbWjEwiziKhItMsQpurlwg9eaIgET9
v5PyUTX7MfThCSle7gmFhdO4pO51LRYhaJpwAm33LA3NCAcJyqC4m8TKlwQBYfXFXkR0ecyv481f
D1f4JxlwHp/Jmsb7ectrN13enxuCJmONHaUqcE1jroGxK8ZN/EKOVzhDq2lid0fgsjnuIwzpWfGj
dM2ZJxpcY17nZ8YD+emEKX9uQ8YpzMQIkvHFay4E5iY4PXe7UMW8cYsaLFmvMWpE/hN1McoiQ44l
wx1UdmqaYaSle3+iJkuTQPjzBKupFVh8pRuUG/62tP8hLlpbGUGEg+EUURdWHu3yxMN6gSwnbfy/
4xssb0IGpkY5HLLQ12Z5IA1spDT6EZg8wVhs1V1wq+lD1tz9iLuJAUU1bzfd58cFrZ2Iw1plAWn5
96FRc8z2vyP975rVGVDNqTm1IDOFeauMrugtyX2N1TX7vLDVNUxS+wZKFKNrJiGsCaVzGbM8CtCo
GFKrzPcsW1I4onrlJTItsDDwIHhFiUvFRABAVQs62GkUUXiFuJVDLdd0nbmO4LRqshqetwGZZoAn
J8dCP0kX6SAE9DkGytGXlzfMc5CvlMhRzzRjVkx4SpoA2TnRrLW6UGMMnf3YR7n4kKKqa1Vr7aZa
QzhwqJchicxggWZEgSTA+bwqEJ78UBaQvzaZsagmhHINGaHEDo6+TsCl31WHW/LyWURWvsQMkEYr
UMJnLaB1cFdbcShAR2+fwiN/g8j1COkDJOkExKzom0Y1V4SRiEWBcjMpY3VmoAcETg/TKHZ/XNCT
9g429nFfGbESaIxewNaz7YlyzKHgHGnJxNH4meH1LXJbsvJcjDBcUemky7OxPBK24BunobTsqCYH
mYhpLT5U6K6TBrmxIJp2ZfTfwcFWELt3jhIsUUE2zVpM6sx3JNZYJ/impOCDTYfNVcKm/gwo5v8b
f79+HdcEaeyFM/nb+t01fkFw1RZKHQ3nQ8CVbNGnefE7r3O/SV2fK/awTgp2P3voN7dbahk4Uspm
sAPjh3KW/gj28p9P+8lhNpghYGgvj92f8+/KQoEEoOn0TEP97AagTiI8Me2uYCPFMJGnrKibK5vW
/JHGVIRazZ+ADxF9+en8FtQOIfbENF+X3Jz5939XZlGPbrVdJ65c8xCG7kCv1kWNBm3VDjRcXLqJ
vjsued3VWXMuGUEzNGbgV8tH9uC0qCDdLG8B
`protect end_protected
