`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2448)
`protect data_block
zBECWPPVy+r54SMxygms3+l5Dk56ztXe7vq3lN0yPkge5pX5Tw8VVi6jSrWE47J7fpXmH6veKaN9
K2UdjIRVk3nkBOhD5aI5MYozK7GUCgE46f1ti0HvQqUGL0SAmW8HWfwT8PdiE+BYqWSg/u2u72uD
HZmgu44VMpfmD5Fj7iu6Bn1jk/PDfkcXGOewLfAHjvqGQ+LuiI1BlGZ6Kn/spKYHR9P5oxB4O1E3
v58nNhvefKhQ8x9sf6BMbgyW+tF0Yraly0YF2JPY6znx/8GgTBVyjU71h5eyA+LXeknqV4qG+EXz
eN/3Ds78re0ZmCVGVQCwccAdf+41X4v5tBy6xCl5WeLZG85BzE4fA19MBKKBBMRmuS7YCRVjbcSo
lFYtxGMN9xpV8Ov6jCLGbV6lAsiW3z2xhVQfTcuw1XtESQol9V/evtBFGxIcZ7TUvVMlqoUoO6rD
dnsgjMMOHLEbl7xbeHR4Vts4/32eP2zVycSbxcAgX48KxxVoXy0L+JC9nk5Ry8EGQjYZCL5aompD
MJmlhjqbbyGjL7UJCiPA6wMNAclSF9sNsy6AbNEXh2QMPNdPMKDEAky1KlEbuq5sasw1sqvWIlpY
e2yrFjOo5k6waHicKXpNhADU0raFKXDEYTAHIaq3zEvOZPUVPZ9EdHVbHumFEYACgpwbp7whOFmw
zSrr8Ak/35qAdVFgsgUifbetBOG3Bd39eHJWHixZSUvY9yTN8rtASAN3dgX92JQg2owXa4+rxUin
4ZqxLfdqzaqJqBb6vcEnCogxCyZY2oDKtNcA+J4u4g09EavOuP781qFPZQ3FeT1qOaoorgOkm9XS
Uci6pjyHuJNlTTTy+JlMAeVSNhkRMss/TyGeY9zmeopyjYiIwtWa/zuwn2ZZQrYgx/djZBsm264M
TyFc3fOZH9ShAUQiWWH4wgaEAhmAcW1Rknc4Y7DBVFwjJc+z+M5FfwCeXPQ4P9szevtr0fbXMeAl
SNjRM8QCXq9n9++ZltWnZKZo/0CS72T4xdKLjabaZ1dwz2tFtkiCHguBvATRc+dD6gRa0yiZcsiX
LBwiusBYWZbpAid/aMdJGhkHxIqt3GLgYGAExk//hKPCKA+2pMiPk00LVJcPqyhgu93NnzSj7D/D
oovHI5kapg/ULZbJ/xn549PHuFAtC355WD3AGdRJRPEmz2o24PkI2Cn8hh0VyIbTla6VcEBpdfDA
+gI0J+mXTJc4gZk7911ngSPf5vrXqCDP3xcJJpVx/1ZmcHh6yTq79iQI3RKqfPny697sstXfoL9O
Vm2dp4yoCkXy8pthOK6WsKm6uQVKVygIMcemzr1M/RdBWFf3cIKcuiv4f2Ys514cV6nl8pmvWcIA
dwAxnyiIIxmutXEAbdfJyJJ1cxnUBNUzH19kTJX4devrrJEre0vbkl3yIyK4mJVoCcHt5E5YeoKL
WbPJvQsDnDQ1ubOSM+VVOe015tO4BpoIGTMwovJwqkGLOysVsj/MvegRpEv23/cwEGlwfUUDoD7V
iHy0Grr/Vmd5bGa2+HBsftbKG8LRg380hkLqo6tEoSYuIdMkvVVk/g2Rd0QV392vZ5qIKsRuamMI
+c5K+NCCez7ah9kfHb8BzT42Jx9k37xS//Ez5bMOiPHesIN+8kwAyF10N+wZcBzwK1ClwktBWXCg
JnxeBSd9QPNrpxeABuxB353qiCx1mlrti77SZUsdbc3GJ81eUngwfqeZ0MwNcudZHW1g3KnTLeHr
X1AvTD23GGHfbVsp2dgkuCMuO2wM4doLysDL237xszPLsA2JdKYH1SkWrDvd+kTks0c4kaAoQ+fN
U/Tby+sgxbGe/GbInekw0Kz8R3eezVBHAXkM7T+YhtEtNy4UXMKAR1b3qC7qGHWkhsfiqY1f1R4f
jpgYNBSpZtneWF7W8FNb2rsZfmIOOnjkg4cOqH2b0QLwunFIV46zyzNNgm9d4cdjF/lOVErfIqSj
Hz+fLieEc7vukfHGEQP55MtkD6wspuSLXY3MLxawGHUIx+PQ2hoPEUPwhiiMTvvNodXEhB28La2G
eX5FiZZigd8SDGg98NUKua2DQbq2VUa8woDmYoE0vs6YKGoye+3IojErJT2ih0UnIAAHbVX3w7oT
eHyYTNxq1GqjYrlhizIaCLnQId4+JMYtF8zT8rK5Dsvbi7dCfRBSEKeQYPX5rpRhD//BF9MP0M5E
QVBrke3233SydCDopgEhxmGJuWfOULk1MwdyYaAJ6aBDNOG1nk8+eaLyM1QW0amcbxvlcUYyKFgA
JATnXURXW3NwIdh6lWG7USTHn2r7Aa1WHICCI+u+aVYfyUfA3zlqKxSJwq82zn2PvBKPwtMeM6o6
JOoifQJon9RNl9n4jwg5LC97OEosD5o3VYkuHmGRpuBdkeDP+4kfwCWxDBX3y50+bY7G/ux5QvCJ
/U7oWuaCyQU58VYS+B3gHjj+7XzEt5Z39mGJu06TcB8+KrhoIpHAlXkaTmyPa3hstGCBnc63PEyS
v47jL/m4pQ44LZgeqFGcJ7u7F5jim9Lo9uxSXxHlZaE3qD7oGU94fo01Qqr1TO5mgqlgLp/EAxXC
Gu83ZbsQ8+4M4ueK61m92dlwLTVi32kxCdQbmeXRnpAKA/UCkkS5+lzXV3CrQKMPree1m3WKJH7J
uQKTjltwl5bNRTnumQqtUfxZC6ViPRfeL2T4V2MpHZliHFhJTroQuoH1ZEaipBl50dk7T4blGolI
HoZmh30o0Gy08E7KDOHaWRSgN0gK7WE04GHajqTAEwtFlXV2s+Uh2wOJlWqb2NGy3b5XQgH+IaMz
Zdul1V3dSQbpV4m3D/rTzJGLVxaSD0uBVJ6WCMchQ4Pjk5w8qlOD0BiXjX5D5G8e6UnPzexoshVA
NArdE48Mat83aPyGA1OEQH6kD3wlIFPk37MA4WT9e84SHHA5COZGEyj4Lh7eacCW/+yZDXtaJR9w
hZPfbDHUGDrQpU9ZKcxtY+FKNyEAPX+3rnZXaAaMtodfvJ4nJw1v2BJsyDhPA/gql9nu/jxba6XB
ljsKg6XxZSjfP+irGQX6pj8H5UZmbTOP58la1+IzDhDur1hnLyLxnLLCm1AtwVpjnLRmDX6amNdG
7s44BBtOjETCaAPd1D9X42WsrNz0CUa5fVuhsDj0nm2Xu5gvAVjXJ3NaBI3xQYk6osPd2jHtyww4
CG+GYKG6JXRATgd78r29MQACUOn7ileL7UPhh2AJ2+BXONj81nEAPOGx3cAEYUjdR1XVlvjH
`protect end_protected
