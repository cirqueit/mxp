`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`protect data_block
qDbE2xGt77jvr7x1+n8peuSUKcPKa4Geu7pgvzmX80AqUaYgbFYrYAw7/bis8vcJ/OvZJlOdEMr4
roaaK2rWf8UJ+yqZvrQCxjLDMIw+g3GPm/5aKNmJrPMKAIVZHjlsCMcjKQCNOLKad8NA8tMdrqlG
RP1sAIFYityvNzfnQbuew4IHR1VDZmfthEVN21dKTjHfZjmybArY2teOVTeJ1/dg6ksr7n5kfAWf
ykKOUGDxi1Z/eouEr48F884iOuJ2qMTDUS0/7clO8nO7Su6tpwgowbjU16YBWIeD/Fg0HMrd3Kk4
wBBAEsUppv9qytXGvRHxAMqf4fqbD1jf8jKvUdfK/2R5w2n8J9yHvTRRiBA5LDfWGYV52hT5jD+6
BYz6qMSGHet/080w8Hi8whcL6hNIzqyVuW7Vw3rsSUbNPduNCRcrsRM62tDEl2bLLBAZ0OII2sKb
Au2QEms0ge88uDTcc/BRBjsMSfrKDyvudgsQUI+SIezf2eO/dDIkt9ZN68BZUkG6amfjDtciSY0a
bIySe+Jkfb7YNuFxwH/02bkgLhSefRk/FVzyAXra6RUuXEndir9wWN0luZbV8prBgdRxqF390R4/
swQv6hS/g59oeYuKt9o+xFJU8Y0GVLCAB26HfnLu5wlUvF889vaWTfG373C63+dS9GAAk+3C4Ztp
5TI9f902bIhIsFHX3auwuXq9yvbnWgxAKywwk7BdGLEWNADO7WStsFB7Vc4luDazeqa2PfUwecHu
A0e9S6AWqNwtjBkQ+eBJOdrBD+na7arZvt4gxwFlByxDY1EMnPD1lcdD/6yZjI4e9m+wEHaKQC4J
9+zCh9pwh9XWt8LM8rEMy2JOgR9cZTNRB5JR+hbtcUWa++kMUR+1AO/hKZl4BUHx5qwWtbU/+uNS
67zWC3A2u/uHERSW6ElqcYW2wCG9bmvJSk4bBT0eeRqbDpSTVxOwMy9CFZK0ONP4jac0bMc5cL1C
VcUBrj5C6Kjy9qFlgvTAX69/6oaBGrkDN7rEwyc7bHSFJJcJPybOllGy/V+wzIMDr85j8ekohovi
jlJdzCYyKynvjRWdCAV1aff7DvCzMvDefXycHsiI6cRqcCiJziQGGplokttAxVMsV0Z5xS/F1r3L
/jY9vrpO1fSOS72ZxQiWLkNV6Dbl+jsEnhsC0eQcFJRAFFheZki3mVLRzHyfT7uzyYBM2j/Eau73
Fb+5ngQMxmIbo028062wUJzmbWCS1CD86WXHyJHHz2m5xiLypdEcg6Bsvg+GyU4VaT23yhrqsoOt
zVX4eqSkHgpRy8E3R8OsS0lFM8PkYFhIc1d6+QLV+Lfw6DAM4e+9QEzkzvy83y31NffJNVHwX40u
wZldGKI9ro4QiXWyWT1CpHdOxZldr/Ql8vAVEG3bGUKIjOQ+0qkihEijaNEAHZigEtlUStb1RJHt
hxIvJLNuWbwKEDvgeh2gC0BBvZg8bvZCrLi6lkwAiboiAo503Ki/fFidP3sdcAS2ocMmpt486DAF
//m/BKpcer2nj1YVvmtQtCQk847CNvf3N1GFSNGVocol5UIntWqIxXhghrWvlU00T3vOSAcJaFnV
8xAjDYhrVds1BI2hzinbb7jeI1VLJPg4g3w3E5U6OydVRh+u6BlbB/OftgjHti0TtIiAqt0+uZsk
yMLYcVMJkTp6i8ZctWN9B9WNq6riYiR1guSFRKA+qUC+/LLfGtvr7k/WBq/uZ8Sd0gsbjefJhk3W
/x2Ozk0B6bbTgScGqsFu/jcyprZ0yEfTnruLFK+OTh3L18dxtWTcEKTcFaH00fNHhIXApK1/J3Um
eMoVWMNKInmzyYx47qCsdfIizn6qZnwefj3RzhmZWDy5gLsaRPD/QCFJykHVS0xwlmM9RRb9CeAz
jnoO9nqgj5u8urQm1yfh0hdunDeQRXiRZjgv36rWloK7UtMVEEwga6n/+1rzjQaL+Ld4mXnJ6+zc
1nXvEpb4N/rvZMs6COnOWhC9cZ2Ld9b20npa1iv6uD7jGnv3SZeDj9rH/gk+LbBgYjz0Itx+eHew
+jW+Gi5zKTxqt7FM9rPfG6VKpWZ3gXyVRnzjhlEl8rT6I8yoqQ+VLi/prXoDYh81AesI4/081pLP
KbvHUZvXu0cK09y0CPNckZxzJMgF8mOi2EJNe/N0RPgrBnyYhRgGVecVmz/+KT39fS4Wv5nbayP7
zkS8RJbhmAt8jGBv1WeEgg3kMV1VRgNl5rUHmSgoJEDZCyny8bZqmsSGKq/uNwsioSC67jaeNewz
tI302EkR7XzMrb9Bhl3W41m2ZITxVKjVCaRzD+rDQLVcblijA7LVjpng+xJR5hpL371lubraFzEr
9svxwOk1GYh4SJXR9yZnI+mOMj26qw0V8ZrQV9jNgVs4fVCQlCdBXW1ezEzjnQwvXgKNK2Km1mw1
UlFHxHjS98WrFwylBE4+OTecrQzZLusm8xFBj9uQwZq6QHK3JgWH0umG+I7UApzhBURThsIlhqdw
skZcPfHnXeo8pE8k4fQGFKiJhXMBVo+5Rkyq9LZfaeVppDQsA/+a910w78hkf6KM2dyhuxzu7Nrq
uZi9BfJzRhXVuB7/aKVRJ4awyzqql6sTaHXKquo6aefeCfN8WGz4Cc9p/pfj/V6WA38X7zy2SzvN
SFM/29enoM0YJFi17SQXDlyP8LWTRMRvJXx3ukqhrSGWmeJZ8kxIGkcSQoSC7NVk4KMv3omLN+FZ
Tw4vatu3Qkyqw/+dlshcVgYki4l1+aMGrwgLMYkzW6VzP2mYd8sNtCZ5Il928hAdBdo3Kg7S92Kq
zae/InnUWPhq4xKgkayJi3I4sdKo5Lp6mAysWmh6DLYnFwxypY89sxxLlBD3evmM+Rv+zzDWgf+L
RFTvKKKzmpesnAOtVC1CIKwqoc9OjzHe9zT3GPhcXMJdmWCQ3kwMyPT+b0rF8d6aBMWkiArtE5C+
AcJ2DshjfJiFUHgVZNFChQtjEhWPF4M2la4fYUwwe5VY8KWY/KEnO2pnhrXMe8DoxEzafk5ojufI
ez2T9B7+X+y4VfFBKW57/q4nwXtLxkeXyamwj1fP9AYrdHjOLUWZr+JDPQtbwdMVc/HQZgghjhjC
mnaSNyC13MVtyTHXSlYxSo26Du3MmwFqpSL7dnoHWDNjftYGYaq4hp8J4ETqg8n7857TgMvz+TFa
JDEYqqdvkZ1m3GbB1c2/pp9t5L4XYrYcF4x7IsE7LJ1BNrDL8n2ddwsxZBQly5/HC8T6G/Wi68Zk
EbYIJtvKqwuErXTEtq5ew+MXcg0o5NbJlfOEDbteUaBywXls3CEmF8hLqpzKpL7jpW8S+muiWYfp
OPK1hFbdQ2v3rCSrtuzlqMkMPU3pxZOhSoke7n7B/j9U8Kq8pwYQxiIpIYVJgk3Qc4fwOqsoJBLr
b0JKrykCY5ljzbToMDC6R1wqMEHk9nCZueFDlIzdEeIO/1m3YAveoIWsUKCT9pyNUBmZJZgILHi2
DmHnj55Gw3uOdwpzodZ4fr5ywolcO0HqF+tRtoLJkHqnXrsTKFa1q2arrsGhLWfV7/BBBReBD9Uy
XQfoLV699GITjNkmQ+BRpPbbzrqS/8u81+2KbKWEveJLlVR/fTTgGOwqbpWOQ8VGcQVq5wYX0eud
yLL2svN1YgdWIvHPz0ZV2x4BR6YLCjKr4hlGzGjpxrTLtBVKB7CaYzZ5LjWqC6IO8ZGN6OJkyWjw
7FkY2f0v9ICizHfoPHOrmINO9VRVgkQLBR2dSWoa9DTCKWXDFySknn/6ZxB3QUIPg8a1s/kAWoqm
NM7C9LgicDcrhkI6FVOE6dG8PkgyxW4fKQsDX1GHP1Q122ZV2ino1DlIzoZ9p8S7NlIWcpHAGrFl
A9ap2FgDlvOVKq6GtBes0DHbH8uIfSKB+lyxrcYEQ8IhjPSWNXDrOs/oTYm6B92watnqD2mfrodw
py/44VfTIqG0kMFeXZ3QPopBJnyBL7wUCJm8l2xvhQYNAZG88uGvDIT78DIpLiISd2KaJ3iidBqe
rI4vY3KI8PhOIro5bqsDh2B3+gQDHpxWqP7ubSz4dGhCSy9ykChnigdToGW8bGo/ddl4hhWybX02
5nyeiUcPFGgN6XSDtoeqAshRA7r1dqFUJWWQwlplf0Lts22QZQN9gpQk7GSvfWM8IWAXy4K9VwCm
R2NxImQVROPNEDmnK3nmFFo6hbSktEeB6vpJiVC1s2z6cd7rlAZNUDiy56I6r+COUkQ1i1r/RtTx
Y7os1RArp7vZA7BFhDKCwoRhFuwfTYEfAUajOFPN5zc6WW1B3lJwdT8ABXgZebG1JeGX92qz1znX
KPHzDs4Od0FhjqXoXerFSJ96EukHlrD/P2tk0Oda9Zu2Rc2uSjx5P47EIfyuTS9/KuDbO1omm85n
35N2JJdDPzCJ6M4JNZfXWjY4xXy7kqzmsqqdg5OaUo/HqULlwVemDvn83UWMLBEJaWjpc0AqecLq
tHeylEar9l2FM3edT7xDSoHLiEeEwfY//CQ8u1ZA6rclWrk5vN6bnqnuwfwP3T9Mi1eD0foLOf22
I/ufrs7s2lJBj0TyPuXIOkkUZ2/jx3+ms/tjTAXK0HRuxIrcB9hAXgO2FnjmM4X5LQf7AIoWsil1
bPMmDpQ0cp0e+Yg=
`protect end_protected
