��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���(�(��BM�D:�����7���q$m�5�׎��P������x���a��ZL�2��0���e�վ���^�GU��g���,��#-[�d��F\�~����������1� �5d�=�����Q�5��~B�>���b�^���	����T�\x��~�{e����A�s
�˫�����ƙ������Č�wޕ�[��\[ Ҵ6/�w�u�~hA��u3D,2�(n~���6��2�����4�V6Z�$h��2�>��逞�dUT��l�q�ts)�����u���/�^��g�?����4/g�0�$Ń�F��o_aey˰��w�_-� ��^�ݏH������T�Coߡ<�;k�3PR�+��X�1[� �~
Ѳ�I���f
�7�ݶA<��Q&��L*�!~1�r��f;�gp.N�p�b_ӣ��85돝�N��xz�[}yz&�+�p'�?E�?�����q.I�yb�E���]�4o}���bҳ�AֈS1���h��0�Q���o�0l��I�!_�.�80�7 ��^D]f�P�ǿ]Ri7��O�տO<s��p��ώh'd�π{����W��w��<<x��E�Q@+�!��#:p�q����0�������{��O_T�1�%��3�XR I�/3p�Ql�+P�l(��=���q�r¹������I�V�߀0��\b��-�b�`�o/|y?�<HT ���O!�y��^E�1�u���P����ǋյux��*K����(8&^M=x�[S�Mkxc�
`��ii�:�ģ�1���e�v�b�hVP�R�Z�j�שVX/WO\��dS
_�F!4�O�],��/����Z��Y4x^�,��j�̍�Y˕(Hp��Q�~�"e=x��`14���)`ݫB�q�s������> ��Ոp���q�	]D]
n,��tt`0�F/I��_"2c2��b)�%j�ۙ����;vge����&(8��\͜{E,��!e�z_� ���K+�� Cʔ�_��⚞����q��6�否}�R��>б�m���Yj�d������ ��wߝ�XRc@P�v��R�?��qJ@��M�kʃ���Ǜ��8�0H1�4p7&���Εv��#�u�>��g��g62j �L\N>�q���k����>�ɮ�Z��'��M0���8�9�֓`-7�1ɦ��JpL ���>@z�b��,���-�2�|��qk�l{E����J�w!mz���%]����)���ř$��jZ�C�� V �K�_�C���M[�Wb�;6�s�`��s5I�����~������:����*vnԥ��>	[] *��6�7q�ǖ�W `K���i��f�u�d��Z+sYqj�-9�g��]���a%�v�r�����4���=F���@w�*�^����d	�S��J�Np��ec�o�5�T���%|p�g珲P8���CFB�ځ�*�4���tI�=�˚�FL�{�D����3Tu�5�O��?1)���[R���d�!"'_�dR�� N	b�MZ]���"��ʼA��6�b��a,���`�Kb`�~�@��=5��X��W��i��J��<���I�7֩,�;�TL�H�p(5�GYwi3�n���V�=ƻ�d<�W�L՝I�[��5��킀FLl߫�c\�>�.�i��,�B,f�DP�e��DT|���ʻ�a��d�pcCGv�w�m�ې�oo�ɚH��G��ώs��wG�]��W���	�ɽGV4�2����8��tq��)�ò�!mݦd�����M�y-Y�r�9�Y�D�v�Q�c�=|M?�g�_b'��"��:
'���ik6��3f6��*�x��QL���s��d��]9�^Ee���%}�{�5���`_�ޝ4dxt��ሳJ@Yp,�І
0��bv�
��I��h���!�h�Ԇ8�Q�:'�,i�da�q`�3r�Gc�=jKV��W;}P���{�� u=� �Iybv䃼N�^XN��9�$mM�^xX��/�:�A,<d,��b?�o>[V3�g��v������#_��ǜ=�a?�.���UZV�^�V\��8+aQd/�+%��Èz��