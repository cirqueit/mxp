`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2448)
`protect data_block
b2tUSTRzMdkhuSOta3Pj4f3gb56J1g5bbzZZTTH2fu2Zh94RLimFR78m69kOoOg6iIQgpu/t4o6h
F5+TYVk30eYzrtBSgLFQqlypZAxQTJp+TYc9NJhzSm+3AvktSYjeyzNj8xQFaPVplr/a+jvE79qC
VlNwW8TvWn0MPNeQkOCuQ8DdDXtpMJbSBciYyzLzAyT6XeJVBygFwqq2BJ9kDZhuCyO3aMzcDUws
alrmddXBacxFdoLTyG/ljqvFSRD5Hih4N0G+1+XOFj40lX9Is78VYYM56yOkgcyVL90/xHfoCaJm
zrcnHRBWKYdAJFFsaHTMIKmNC89oL01vT+bxRa9A+HJHClsB8ST75wB09bi+ccBAd7TxCyvUexMi
DGR8Yn9oe7wc3c/OwfZ6SDf2nzjmx/1kg6JMAPmaHjrauJovoDeQD4xiVxogUDXU7ri51MnquSOY
gY+dfutHrxUVxC5I6k+RjcKsZcJ4OXVZEwth58zrKgFcNELiEbwL+9lzYJcCHRv+/4j8na3z4nZC
tfMGOgdx9GFrQ7MyZLz18ggxxak+YDsS9f00fKnwRLyUD5Iut73kS4SUXvmp9GHORrWludN0kZKg
8BR37q6b8D/zeXfHCQhZs/MuhQJS8sufNjO626iOO3XUJR1QIevYizmwVq9qa486ez+a/TlWrVLL
ht4uCLmewkzLaRy1NndZeKubCh6/sZiL5eCewnoSeW7MPiYrhLxuP75ZhmWBTZRMzKm2X2RsOGgt
RIrOPKo+kBl4zDJuaG5ewCkOZ/0G1oG3DzDXl1FOcVfZPHyJj95xi1cSIndceAik8lyA8Nt8UWQ4
AIUu2LZ7KCirZLXrCFO8rIq9gMixnzX5CXfReAngcZRbqjaORgYa+0bSFJrHyrku0ubTzz99jTAN
zsqDyGr7S+lG+N5yO0RDmit7XaYY2n6bc44Pnwfp8Dmc3w/97Lacz3PWzRMb8ET4aSZZ55NSW3Lb
TvkEo8zLpZMfdb0gfRjGXsquJLUP5Rqagi0A4pN0hie04NS2J/DsFiBiKg2vd+59QL9FOekyTYCn
RRvZW+6GGZJZ8hGSDgf8RjzFK7ZN/gjtbCyfbpuhK8lSl6LX31+0Rn5CMVJZ/wlRlXwXwlxib3ZF
FhzVRZWUi833zR7u9FX48nje1JkytSkNv/KiFwf9sh8aX0fKO2aq7BLWvQ/d+TZx+ChQose8ZSN8
695d+u70tKL7z3w6B4q9T+MCSpNSI8hO+BeRsXhI6KK9+extG0BzO8Cej0JemHQt7vVOI6s1PBSP
J111rloHqryJsyYP2cD3PdvaCF1ZjZ3w9VA0xLVB/JaGX3qcjy4x5XbRUA0w/5mBNoJPd3wrJ8h+
QHdkHMmOmRi+56iohhtNClIMUDmvrdjs8CIMdEzMPLswidBA8IdPckH8o9vq98I+gd2cOh72IB40
4fVOLsQC4id2ODadWM8EMN6oWIxP+IuXXkW93ChvagQEgcZjB0q9otUy+VM67e8wV9N2XkwmrLKS
7BXjBJdHoOpjE6aMeFet9qCEXOqRaeyqARo1XunPjns8i+vAgfuVbwc/DoaOPHP2UNndBsXLJL51
XnQiLX45Kl+1p0XEX/ENUDmx0ojdi2MsS8ZpT9cvRkPMTfRhFrEsAVUjppogMNWEYLemtvVEMqKI
hpFJXAtTLDB/YhqqRrG0RZaWarY1xDDv4hrfSwla69RdwlB/LB+6xElzWgU02mxr2aVma9eZYZ+V
zxUF57TbkVw0XQtfIvZWuIDZW48ZvBpd6iAHJDtzvGydd2fh28rV6oq40DmOD0L88hDT8B4wRYPd
586t+fgt4X8wqT+c4c0EuWU6CdHo83wwH2F/AzMOtO23OFqN4O1Lxc6QETGNS1yt/+toMUPH05Bx
dXw4VOsXSA+NyWy4EdzsHKpmMGSfbgiKCkQs5+U4x4f/mfPDmH0uTtiTA4PqQhOyRE/TtY2IReP5
BYup/rQpW7dAMiv0bFQiE4xEI+19zuZkC1KNbNoOeiuXuByp93KBjgcZxyoAi1wuuQffz+kcZ+ns
psSeOI9DByw6Uww49Z9jQpWNx0qKigzygmgzUcgfoJU9XAionWuAwzd49MkXlaulAk/KYww7PI/E
i/DWo30fB2GcpM8R+0bHIQs0RXzTeGQVlvB/bRJtmnFpxXhNGDGr60njbS9Ma91wtVQUeD5cUZ0S
nHSyp1w7CXEYXvHOnWG6S8CT5OgvZTm1vM1CiKQq48dUPWjMF0CUZ5JKazJgnWok0xLaXydnSwtd
UFQSdkiZX4xExJhHFnKFD/O8fXIJK76gOXkHi4i1otUC5DNL8cPGfGTCXwCKwGVi9sOgt0eTDwE2
p64ItUYpQgrWR48n7NU40XPx6qk7LwaNLfjdnRPWwQJUjgDwcjDlbu7gP6jdz7SfgGBQXJWb2+OO
lTC7i0Duv/HKHj89SvUNDdsxWWZUCZQtxVw977HPpAt82TRZw1e7PY6fL1cvONQ2vM/jfsT2azaE
4nOaGyW1wRmB+pThlxbc3msMtZ2nYN3/wc4bLZbTGWrDZ/UitmhZxw0phrhMlLreTmrzPwvab14t
/sFUB4BYgNSqaN3TYAbK3HLdV+ElJzGJnhOX/QOz7HyPbfgijf3/ei8KWu+kYosrHGZU9KXbJa5R
qIo2CKfyxOHGJtI+ZHZT8S53Gh7CB2TCsFS/SyCbnIaoaoeiAPRA5XDnipRuSSaSBxYE/JGZHnfk
7S2L0V37S/IeRi67Si+h2F9LgSEI2TNykUya3OXNKvw3f2/FhswD6awrfywGIKhUXfexeco4i1Pk
tC5OUFPCS5wXHnIMFc1/cuMH06pYc26YHSxEkdeui830hkIpiNXN77OP0Npf2vfyWhPqi8KXeezM
ku7O4slsNjv7gdobgrcG6ADNNiNpKFPsxMCepjMv9NKtbv4Xvh3M1O1CJU61+VAflR0dECl4cUxK
CyxhzRm9eN4aUuYbIu1TSqxY1hd3HhQ1HGIPj2u98wsc8xCpH/Y7NQX5ewk+nIz96OhFaa5h8I1z
mbXNv9tT9EOrV9GJ/ozcChh7Ro3ODD0S+qMl4sS/ZIJmoGVO4WsNFZuQAcTYfnw18l8bwgR25KI/
3xEmuMSA6ZmaDnXDeTiHWaLeDyklgLg9/BLXC9NCNcpgff/Xw5KLB/jG4Pw7w853oVZByZS1OXV2
kineIkgYZb9FEUnVqUe6AsXrvJGLML2n/YYGEBDMtr5wXM00lY079MhZVgJQg63yMpo4HO+W
`protect end_protected
