`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
ums6m+PqWoP0BqstkXdy7dXXlZDDqcSKooP4ZH49CbOp6j+jIbJXf0L7Tnq7Wa18CDN3Q31IqndN
1C222ld4Q1pj/XrFD18zt54dsm9e1oy0b2N+8krqnejanV5D9kd7bFli5AuqCDmlq/KP03pXiAFM
keL+dI40UXtIx+hcZUaW79Yrg3pO05ut9nbmct3xcU03ZWRKisrYEyTXRHAdF13zS9ED2v8B8l5r
BnKeXQ3iDomAPDSmCWBVBHhaDJe52JEzQ+/UB8shNoNEFgbLlyXOzvvGqyWYMPRHuMfhPR1x8Ho+
vGHVfCis1jvN9I0jj2uFRL0QQ/tuiLwCDtE6RbGmkIl3R9o0DmH2LzYeYbMPMoo+psgOG0pBDnWT
3qVGQ5NkV0kavoa+7YOMCl0DqWJV9j+xbULew8cnbjaZKhEsMVpc5os/3TYnfLDwhDqsKNweVEvR
WTdk0aX8C/2gAOEwIN+8UU/t5J120fI/TQnTRzWG3IRYK0IHEPK6X0/oKeBUvY19YtcSkIUjejct
beg4kJXqYCk3dsxhHnQRDQkLD30i1gPhwHSSAFya4kEyzdGagfMEld8DqJ3c5/6I8aLsnyQC7GF8
5377wtA385JT4TDqCzUjcM07C7x+1j0vtu47hG5SksgEEZTBOoaktJaNvf8UvJSI1KBXbbgldWdr
cko19Qvd/FDqvsicanjYJsdTwKX1/ld7J3gP8OkJImiz4u01KUjz4dKQKmWG/lOMKlHTsp2skkea
V3SAtOoK5BZ3UXrEHuwXCZ5/s40Xstge30/6PKQ1FveXdXg38csK+LEDEBq5DHYhWsb5kY363ULi
O0DiYhMD4ki1ZkxoEx1FfKkNAGXZumJe0v6YxYeSjiePTy8uLwo6U2fzcr+5gi7otn6xXJmjzM//
WMIMaAdj0LqdPpAvtigP4ilnYvf+sKL33lf4yEPvD3PbGiRy80FxR9N0pP2AzBJeJSPZGOp3C9fi
NcNoDEXTgwP/2MWRx5Xkz+wtnrq8oF39A11isWS8tkcw8WAe4bVqbBIM7ycvPY5O/OjaI4NHe1mY
PNfojK9lp6KfKHE/le4+W32eNz9jXJXrMJB2lVP2fcH1c0fmajM5zWn28kL3e8Qh6zDC9M/d3xQr
NTWJr/Vf07iL7Vl9utfaOtasYl0qBmWBKhITOJi7j3WndVnMGHE19kZv+sN8y+h57yehVbqYa0No
pM3IXUPhaBNHmAQfUNQ+VOD7uIZAfdgm4btsIdCcZZFxVtMehiFCjjBX5SdEaIR8p0EpdsAC2wTR
1FCxeDpIQGTUFkbjpxtcik1SBlYPL15BxkRGIgmFGXH9bL8YZKsc+0VmHP1YtSqdpR8xV5LpDNNK
59V9+Bay0h8ImRNuPk0X5JYtT/x9L2kHlg8T43UXiKVRpkp8BcQOKCxCBHATDTT65GtKzXkV5+L8
JAF0yMMusSMIvJ2015rewEtCQsONb/+tCTM2oqLIDwGAKEKn1p2rpu4ObEcNjLSh9PY0dLjiXZV/
jI7iAC+mkpcICUE9nAuTfAjTHDngPD76JgWB1TG6woJqUVVW6i4oTkbCBR5ghBtbi8fdXy4yzejl
KK/vgJtOp/rgWUa1HcJMJYPf0PoSF0XFSbfMDLN8QmempZL1oyqHjwA7IUmOrivxhGd9oFn6QNMu
ZfV9Cgi92fpanV+gDZsvS21g8T1LEAYUvW7OOGXHS0U+GC3I2FHTAy8PN+zeYuvf430D4jidkFwH
z5uGIGUrnf0gBAxE+OsL82Np3+q7oUvkADb3lYShLInwnREbTrtPGRUkX6gp+iDtrzyiTPcfeyZS
N2Z6twZm7cj7se+DVFnSO/woFnW0VMVgVscrLV2caKk28o7gCvb4l9gqtAT789MouNdJGTiQnTFY
9BMU80izHgVlqXD6Wr7LJPmeaZTPaa7yS7J0BdWUF+i7yAjhm19m7e6GxdKJbwAvhlzhWmYciq8U
nsl/y7NTew7FQpN8dBZgIGV8vZ2fZCVjgmNPg5WTfplwmIvijKWHB9lDFkmt/dMHhCHj0TNYYRb8
9Tj/SjR4uwol2vNmbkQFB3C+hPHiZCfTZ5T40YIru0wh/a+l+U7MtLR+k1I/Xc7PzCBoiO0/KClv
xaNRTbufnQ0o2FYAgac7lMdmP3fWDrszJDWkhaq2ha1Ekz6bEx7er9zNY7HoVTOaf6ZvcYeisSji
jB74nBFPm95HBtz06HZir93enV0F03ArjWgZXKBqaVt76gQv75ldRkRHL35nsEzgu1+bc5rWPXuA
wqLGjOzDs7bBTaO9cOuM0XZLkd8XvR6Ji3h8B07ODGXELle1AP500TIm8utP9O5+eJjxkE78yPIQ
GWz9Pw3+f6hyBbFvpviM7Rt5TVw8jTBQE/ZCJ8VFgxxNEb6E7Tv0X2yupWdl6D4XnaQsZrzk0qUM
hrQcsyngwqq61llsO0ZI6TqOD8LBVBcD+tn0OjYcosVbSL+RXbKB0gXN4ogOTSgrsVhIggMz9zG9
DiOBxUbdSIbwfdLGLngRnmFz/jH5HSUxR18Eg5hWqwY344TKTcgDKDYApMAjhLXjDeuWMEhkQAIu
cgqqK0uhZJLdWtV+e3B1aw1K1vqzNZcyxVccpi/4jjsZqu6d4wazQSwNoXfD4Yvb6IqAp55aFJfn
agV9nftD969pYSvOOPv/6bTUfdccj0Ow9ZmpXHGXxyazK8QT5kAWMiG9Sdak5ZFokikimfR0h4iI
4tTc4BPazjRq5QO10J00RGW6lzaPshQ534B0jm0qJ4NdVnsSST4d9gkNeYcGrl9lYuzdGLFSZQkG
bzW3A66DarZ3Pb0PATTcvahwKfqRe6cEky5zWoXopJN+it/wcl2nHna6AdNu0mReWPOu
`protect end_protected
