XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����}����z��U���0/�l�R��M���;)=��^&D������=jD��aɣ�Q���y-FLHA�c
k!Q�Ӥ���+4Ϛ��"Z�4��f�p�e%D��cB�|z��[���F�
���4�Idu�m"JM�嚗럹��,b/�@�U��ɠ�3�����9�"C���.�[��4q�*�h!Y�Rw;R�d:�MC�t#�W�?����4l~��(�� ����#�}���BK�nT�׈�!tL�̚�1���b����݂棤�?X��������J��^�$*6�^�^G�Z�kq��Ț�[��&ҙ�3�Tl��	�l'.�����Mgx��+L`oN��n������<�Ww"���w��yS
w.!����J��U䎰M2�T}թ8�qo>�+��{Ty�0Y�|Zb��E��xc �ӫ������i���Vs��q�SA~mbWX�w���[�Ay�@Z�nQ�V��~D��4�7]`�g�� �/h��7xp,�o����f���m
sjU�B��5`1i�3b`�����X�b4³Y�b�p�,�DN
"����)�c+��#(��;�P�[�@��S����ĕ� d��_y/I�!Y�s��H���ԺjL?���� }>���U[['����A)Pa�3S��FW}v��F�\ �����B�O ��M�~d�(��T	�o�ku;�=U☐w�Ԗ�J`�� �n0��a�-���,� X ?Лs�[7=I���XlxVHYEB     400     1c0��5�)y��6�'2a������t�́�{W�o50��C��m$�Go�	��8�JTg�_n�d��zDD���W�q���5��?=�	����x�nC9�c�d���pK'��G⿣1[g�b��b{E5��������U�{9����c
����tk�~wws;����#����m+�\�!�-�L�%��2�HS@gum;�4��,���
`<�k��%����%�O*�ʨc������<$)�Ţ�8(*� 3��a�F�(Ӕ�,�	v&���v�W��~X�z����e"����#����r#��C���eq(M#9��0�qBf������j���Ҁ�T�2�{��Qa��K�U�=�~�;�&:6�L��]PO�/�ѐP�>r��/�H��t���Fs��ݒ���5w��Q�kĢ�,jYQq���_GkN\��clU�=�{��XlxVHYEB     400     160l�,ϋ<�"�V#O��V��9����[o;�W��:�0n��es���"1FvG����g������?i���? g��\�]�U�딖���$�w��������Ɖ���I�IBU����8���7D~���8���t�B�o�L��Td�i���Z@d��	��P�B�Րʽ���g�k��t�nδ��<")���1�k���߷�{�#�b.�ep��]ȩ��ޑ~$�;v�^�������e�[��Zu��1���/r�6�ia�6�������?C���=����HX��d�ҽ��_a��u��f��I��1���=��le��[}�l�+'�\R�~�8[[�����:��fk�n	�XlxVHYEB     400     160����y���o4�:��Xь(�蟫���Y~s�����܌NE��-����.6>kFQ ͅ�t��+	\_������!Θ��Z�(=Ă)jj�V�X&��M��SB�(�o�Duf���Ɵ�y�O2�6=AG�>��n>�n'��o!`�܁��E+��3������v��Nq9h@[ ����^)�	o[�Zz�1'ݝ�:�ō�^��q�]N $���~�Y��X�rb�M>�S�@$�I�{4	�@yUlb����\vV�:'�:k����-��}q`_�G��w���(_���tZ����u��8+��v�G1��ʥ�`��|"����$����S~��EA-��!XlxVHYEB     400     100T�/�)x��"$�z	'�&*���y�k��ں!¸u8�wg[��@�8�i����9l���[�"d_o:�AD)�v9����Ņ,�
]v�;��d?g*{��δ&�ݮ�8��D�e��r�I����R`��`#5��f��r~
4qA/*�M�[O�� C�t��<U;�j�X�� �mD�>
�W0 �\�͆��m���Y��yq.D/�:�JpE���qP��EgI����O"��3k���P[�5J�a�y�?�D��XlxVHYEB     400     1a0��_i���A�R<:aa�D�h�}{O��!u��1s(�q�9������y�$�p{{l�w��3���s����.���Bς{J�T>���z~�������ȕK۝�w���|}��[��F��ɽ~��A��*$�5�YZ�Lc Q#-݄*�䰏�!:���mؕ�-��TbD)�|�������������|�[dO�Օ�{�/i�9��<%��zL,Oy�w#D�m �p�Mʑ��1�yq��K'oY��hn(�3�S���ЖQB\�D�>^p1gl�8���S��C��6�;z�i�N�[+ �x1�L��~ѻ _&3	��j*k���;9���B��>捏�h/^���������t���Z��h�iޭcW�<��){�V��X���N������e7%cp0}W�
>�]XlxVHYEB     400     140�=Xk��Ƃ��e�m%_����Xg.�6�k�~���-7ˊ[�n��.�<#���,�|�����~~�-�߬P��p�;�R�U) ������Pܨ{������Du�l��/6��0�I��Z�D^�͍�W��0]��H����D�9���0���!��Bk��O�="to�j�{��h�z�d�1,�Cx��N��!�����o��Ok9T�l�A�|v1��c�^"v㧤�[ǡ�������C���^!]��	��-�CΩ���ﰭ)~j�ݝ<��	�����N0DF�f� ���w>�����z{V�xQY�	V��zXlxVHYEB     400     120�(��*KoA�����ӷ�G� �8Q��Ifx�s��GS��j!��R�lΖ�z�cG��R9�g{V�IB��5�w�Y����R#5o�I�&Qz�Ȓ���}�Dy��@�	�n?����+jz)TK��F_��#m�1�-k����$o=a��#I��As�`ԝ`����h�g`S�S>�8�\��,��'�诉�9�����+�cK��\|��^^"9�Y�O�w���uDn�wZvBٗe{��3�����3ס�j���m�Ч�/~�ѧ���uΖ���U(!XlxVHYEB     400     130"q�`�n�iU�!7���$�2�#ǵǮ�=W/N�w?��H�+�؃i�Ñ�Fۼ���(o�s�:1�b�P�
N���hͨ�3�;��4�w79-��U �>k˫?�?�q=Ėn�Z�Yr�S??��ʞ$=���*#X��2Q���E�ry�n=)ǝ[��z��1����`�y<�ԡ|�()�fζ<B2��������O]3C�K��!��@�z�J����T���}d��<����7O>0l���b; ]��c�#��/u�z�@���$���O����k���!�i��PV%h��{XlxVHYEB     400     1c0M2Mq��4\�.k�_��Þd��������bh�?_�}�9<�Ӕ���\�]8�[��y��wma��p���r3�����C��V����J,Ml9�� �+�;��Y��gT���:�� �8	u��s���Q�8V]����0�b�(� ���n�I9~�%d8,�x��S�\> ��>s�Ŷ�@���ŏI<�k0P�� �3�����a���$�<*����Ua8|�]VZ&�A�YE8�bz�b���&eL�P����P���S�!��k���7����@~��x���̓�E|կ�Y�kH�9���#�`�3�O~u
��7�F�[2�,*Ž`^ �2�ە����}S6�5@*�]2	[�����b�0�����JW|����7 [.\X��B{�����'�a9Z��0K��Nb(~Uܷ�d�)-��H��l|[���t��/��<XlxVHYEB     400     1a0��	N��2�^=�ȼ�ԕUR�W5g�p� �
��A���ChM�$tM�R;x?�a4(3�-�f��?��ZW���k_5��K"��x��N1�.ϟ�2Iv�� F�E�)�"���0���7(X2��/vx�@Pzl��e
��>N�~y*��t���lH�9c-	���" r����rt�S�M���Z;���T����ȧ��v�
_���q�VB)�:�@u��+���W��	v���L���I��v�2�����
J�qtv��[d���anT�)bW���
4O�BN~�q~D~G�=b-�N�r�:%i(��2ͥf�P*
@8%���)�V(��;Id�$T��&����7baGH:����m���N�uZ"4�J��cw�@0�7)��*Dz�¼�5���l��~eCXش�{Q�XlxVHYEB     400     1a0���y��@���k�2��-V����$��ִ>mQ���n�y������y�,��Nk.e� �"�2hS�~d|�C!G��GF��)�h����Hх��43A1"i���	���M���-`w�4i����k�Ь���C��p-�*���O/�cr!�g�҆.�h.D,1�K��ku���*b���}�k�V3�*�0��v)�M%��o�<���V���
ij�3{�I�A��C���HP�i���p�L��Ġ:}iS�h�S�^����-�ݰ��>xbC�����z:3TI~|�vz�SQ�7W�Rn�����[!���mD���疏A�.�r���|@@�j�K���7��(��P6�*8�Ŕu�J���2I��ʿS� <I��?�������>��Y3OA��"�猷Y���G�XlxVHYEB     2d9      e0ԃ_ˣ�x�ȊN��ؖ��ڷq�<�RAm*ĵ��s�*C��M��θ��� N�4h��ms�}�������N�ÎAm�X?.QԒj�8�,*O�Do��z`K��9��3���+�5�=>�[M�0U����}%P�M�ٗ���#fLƶ<t��P��ݐ��M�p�E�8��d�S�W�P�T���
k�3�|Q����,�0����ܳ���?~3�om{�q��W