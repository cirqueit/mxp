`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14912)
`protect data_block
+MwDRPnQQ9I818HrcOABY3304hiH73FN7HeZcSab307kgZVweF2rlwwgemK5gtZOYBfodU8yCvmD
Ydjk5VqF5opraEEL9yV74EquoRDh5ju0jldt7dGsY2kPesSmnLkWMm74OFyWC5T0pMoc/lJOj6f3
ZDk8xACMpRPo49IRww7Om0cIGGSnKvdXhjyR/hA8pYUkWqtzkxxi++jZqWuCMufGIgHBaFF0iUQJ
fttaOUVOYo0Z+NzMvm5NGi0bvTDIKTtBGDRakZi/8Afv/Ck5t0QoRVWZHxvJKkbvOhG5uYoW/1AH
b6czck6MDcwDJfWveW9EL6blcRAdm1rS/tmB7bTtI29mV8Uycf32Y10aPB+Gt9f63TqmVHP0rLNj
Tj0uT1tHRw+eZQ+FXhqtf8lBt9rsrT6xqYtKJh6UKPQ9tbrtztQXaVz3PAgBEIH1ADa6SMhSMECC
kupwTy+J8W+8W8hxCg3cd8baGvt6+jBK/ZkhD2yLYEwwMA+lGJl7UT2r22sKov6kXhGJ9zpkWn3q
jKw0iQw9itg1tl5J0s6BpPohbAocBMOJDruLePoRABywTop9fVuDO/S2IjJ9htBQdeEw00wbTKfm
IsDWdbvADCUBJPGN5J6WcDP+xGopWbEuktmlhtSsYJOO6RlUsquSwjm8ho+0qSvURHjGVDYofARE
AMfUOOsN94mW80m5d74HKuzaldioI5zFySrhSd/oCDD9iJ6h75iaSSv/tGwtoOGihddTH9Pclsfo
DCyzCrYqK/GZ7js3WWewSaawLpWiGi9B1A/U2rJukeZIkSPU5o3gCLUN3GA8zYi3pAWssBpFJXnV
hw1V9FCpzgcjqn3OurNP61E7vJuov2c+9NkXX0W1ikMB6dBm0bT+ZzruBq9MQSkR8JrUwBbyUlaj
THyMsS7y31DDczigNjFyR5A68vSNbox7btt69Fx6hRc6XtgyA6A0dmqGr3VXn1V5C38Kfphc1AEo
vEIDDtwJwpW0llvxVrfQvZyIjV/xumCDP/0mcEMCVol/mMTWBhe4lDfUW9nqeS1pQJRqEM6Mndmp
5o931ngR6XxGjLm7q3m+Xf+uzsjT7EAplUX2ZqUpo0OB9Zxx8zbkucqOTyzU8tlDcUr7rZmWJ26h
Ox0w4PsXGRNeKjOqh6A+G3XUqrGtPbA4LCHvksPet6JadZJaOBi9EK45ycm/5NSnIrbEdlXKFL1U
nCXew58u03hx/+Y9hYgWHXsibDrjLDxVCNQUYVnb7Km/Z0/6Ozs01IwJS2o61x5h5tPtE9rPVXet
Drr5R/hcrkzYZE9Ai8dE8hst4yQkBwGgNqZ7hqTqnVWrJSriG0q0XSB+ej6OjQPbQT/hikpd6r7p
KB7s+ocDReKm/d7XPWhTuSTLbzu85+Y6aCGFQliOwu6wiY4hnN48bONqrbsbOOxuN28VjXR8JVtw
FJSaAMvvRKq2vzBa1M4xWluAVcPMzbZbDUkoPKTPr+B+7WKBT5kag5HaKaqYOJgRDBU81lf78G8O
yN2Jag1MDqSvtyj5VuGl/VFnOZYgL9RGreDgJ9UtsTXTjOXLPWRHmLmNuhnF/R2r0ABi2j3sWCEU
Uu3hzZh+zVBeTeg947yOfvBL5FDL00lrKa/qGJtdhbl3Xm1FcGdNKVX/f8g38CQ0dlFD4MxajOjg
aUSVKZq9bcTDEOM5ZBolEasqlqeC6Eji2NAM9JCk0WEj8EdnO5WN4SLOHEMTobiVp7tB+KpGqdbd
Jnq9P9nvMMgNlwb+fzYub+FVpKNAO7Uz0EX3hjcJEW8+uN8zRZrD5yITDJwyH2pwzr45vDBxwIR7
s6w/WcpzL7Vs/jAd3zqDyPm+8vl8/Ij1nCrvRUgl+w8c5BqTrIclJWhDBORAWI0a/bU50hTwrHEI
nmnHO2TqnsrJ+YaweYBSO85lxr9aQj5fByoVJPInvShzbItV64L5HRzygF8EhLf3r1Yei77kBkgn
l6D2d58OERS+4SlbbuO3eRt/uXvf14NOJvvowvInTkQowsZ/r0JUzor5t73T+fx4XUKA3C4sTo/J
zS6mBeg4J5/5jz8FUZIeF4IyewJ6GUotwd27HOI8ZEHKygQdX+HMsLTIBn86iAxwKM2C7zBRG+GB
8b5oc2tzo/VjZJJRZoyDKMLVXqH7SNGBHSLlGp7kcPTGD5MMQx60goV9zWmjKrji3MiT8fQVGq4F
qqon6nXdt15JBNqs88f1ZgjPaAgOxVtu2c3AGkHNeoZVMaZTaFDz+DxxszQmG6IB28Vh/E/fCTFs
5UUoyw+jUa2w+DbBls3dIqghU/On6g5Ej2RGEyWdChWcMhxy94czeVmyqaII33XBMiNX5NjlLBTs
I52ro2rrIBApaY0cQLhKePX0Aycxgj8zG4pDyqu7OlpNzlyeKUK1eX8T6HKkvtcUct8uYdJCaH1w
nVCyv0EIQbj6KZGlhwGRH3LcxWiP90TpwzibphlsznAZA55Mqim6P4tdszUKVHGv5IYi4dfu+zU6
gkJEXCVYHANlPOE/Zz+CclWhM9IsSw1LrzuIeeUYObowD1iZ4G8KQO30vQg8zag0nUk9ndkwxi16
YHFfGUvucfGejetamkjabIGIGhSAJi9aBY65r9aD2H4Nz0dcAAIwEWJT8wsy4R369R9FZZ8Rn8gM
Dr157pxeapPx/ArU+QwSVg7Cyt2UoNMxGPNg9J2FxcgJz9ezQu7qWj9+pnjhYPHGQuTk2yOofN42
XR/8Gmy9baeZgRxnS4ODQqxPWlibIVMSaYqdBa4Bdm3jP3p9mgXFu6gt1mtEyL0pL6jcHN0EhgBc
9rcgcBJqwKWjuAZWjLor/qDbt5l/N/UtBsfMhlvFxisn7uWFhLf4XJVSRfh1wR0qT9ApPS5AQ98o
XElbB3T7nQbfGjht90LceVuysdrVB3vPOnB0CFdOC69UJ6WYJnOsQ9nvSRjb7EUxd85wZEs/yhn5
eO05AsrZpP34wf9oLcdI73kKd1uxo7Oh2NtjzetDLTutEpzHNtXt1VTb8SEasuXEJHjXb5/IlABO
b8MZDKuvS7D/xDw3pXJQ8Us85kGbuGu8SZ5VRGX2rnj4ecG00B33Dr+FfcXx+QYVt866JcxbZMAl
an8AHSCfmS/dB9Zk2dc1C4WlEG9z+qIb7E9F/UNeJnFrJKQ3jIfdWLQHKLeNwsNIhbqBxECq7Jee
ERB4eAc4YF3mLnatKuYtcPKplRCOBgQLLMC6lg0XyivWbYWGF4M3VOnxVL0+WeIjTcQgLQwGkj6g
WjkzoFNpRa40FqGu9bsWdwoG2/UERBWAIUv2y60zpkSVnh+CHwqKnGFCeyRGVxCVYSdypG5ItSsN
UbTsklAbq0Y7DgItmDk1OZZ1pwvcX0O9+5wQ5IDnlq+mhU78m5qvt31POrQaCOPoL/u4mn0iL4rI
yRCBhSFRQKiYtxemENtEv1ZdmiIkUkObSStyddjK0lsixkt6ghoHF8miJNAyZaFp/esKhZwAvVYA
mj4Gu4p0vB48rIzyiOfAfLuMO6F/YsqbUsk+GkTWJUqqvc2VEJJQtFh9b0guLTYVHxt+K5eyWYgF
U4pxZlFkSVgdMVWyFYrZ5uNYSVOp+E+fHl4snnngNfPq6ZoYnHLR3fEWX8xOqZb4zL82RW084mm8
dE2A2UVEO79XabYCfr+1HTgqmIJRnH5W1r24qzb4IUj0BTvWxibZYHqaZF7wyM7Bm78XuOoExbKE
MUCdQt66KjDRJb3L/6izxmDnm7XgIe50EcZpYuD7qgtSekWZvpwJHaC5iFf4ROfWkj+EwCTTPn7e
m3hCM5tQzVJERXzGH/iHxiQ0c8TJUNpLQCFRk/KD+BZBV2f82NczkOSEgEgnoDv/zQ+cI/nF1cII
nRxI1/RB1RYc7q3Qy6wXHtGIxVP/KSBiCctRExWY+ahoYVCES4Fjpq+jZmnlZDwI0NLW2XszqmXD
DhkD81iU4fdE4hC8OMZXLFFIPMMI8HA3csknhpYUWXv9sTCDFXSvoJwZWrdrfcpSLA2PIQCyRHS1
Q+OP/RSWv5JphNAsfcZZBQqDA6hATnOX0/92hdxavVWw/II2qHD6OUWkipeb+l7xWNlEPDbshjfm
SlVh+41mAD4JQw3rj1UStdPg8synifyp/KK7HOmOKVizIy8qMC1jdDucwLDMjrly4WG/pTKgfIgm
MNkFDoM4Mp16t34YDle1Ruk0mRWlRk0vKu9xcr6KdN2PGi+7nRpgeIGDpB3Y5mdrDCz/6lNbSOBO
u4Up3bt2XjEbohXNfawF8NzqGwiEzgS+fLc3MoOa81Flfx0WuAwiCXPhhQ1fX5Php6SQ4++L0eSk
b7f7aIOHUstMrnJ/JLuKWA21ZLiEkC33zlZcBEWoq0gAX8qjJParYvVTBKpLq8OPyO/UfZWssjqq
BabiulhcKw0L72K5nlO1wuNSYnkNWSQq+s+q1vhOy1DF8ttdLJv1aIuA4RZskZEPnBtBXjWFg50B
Mv4W7pVGQj5QHfsjLapDQE9w2PBCRc5Je/x/G+96PMDKLizely0YoAvhrj4BcfJsKzIzprC4kgu3
npMpGyAjahF5+yM/N5icEdt0NiIx+XPOh2clhfgJYcoIZPc/D5uB9rxkW7mfec4grLHTOb61CdeG
mt+JlZr4/z5Fgi5ANudHjV0l7SSJrm+4NWvzhCiiY/2Usc26t2VKyJqIAaJTuJcCJcMxT8U1A435
AWTFL+n/OeOoFWoYV/lZwVrOGeH+e8sdYSe8qzef1EY+OifAcIvf6E2JVpGXkbVZNQPmIQP+GX/b
sSOW2TvyzpkGFjEHaG1eHOEgWY6/spDdVWmcb6EaXYk4zop/3yp/5eZQ/GwDpFsBeBhzBukIa5EL
6jc1+7A9WcuxJvEuOv5xE3D8MNJreN0uAgiJykBxHcsTfdi4nwvFSGsbT12scWJOWmcYD7kk4SGW
BjZ/K6RGarZZJKhbbZyl5EhToQox+PH4rq3oVQoaxwD3HSh4zz5I3khCg5BNyLqaYjWGALI0j6OC
A60bFwTrwGwq8gmIqjsOSzrwXfRFrx5DQ5eA4fYcKAP8nCIiFyap+16Y6Tp31JLXPqq70NLoPzP7
tdlYdgPb8+1fmaR5ZumS7XmFVq51YZ9sgw7LzTHmDF9Erdi6pBOlXr3AEL2ITI8Gt+kmsGqbvJXP
P6X1/cmokI62GcAjHSGfuRFSYCsYvTvygw5b7BbMMwroIC3qNVTnGLIPPuLzsAHvdifMBhLXZKXV
UC+y5yMYolnQ8KM+HxQe/EA6I11U8qiH4muPbtL6OnoUoz6oXXrxfo4o10OzlH7AXCb1R35NdPu8
eb036jGInaH6NchzMsvI4IHPOJOFqLPgEvWpQOoklM92OwruQlr3+jaNbeiXeKRj5QDOQEDE7tmI
aYzrojWUKCzgn9/KKaI7MgQ78K4/kCIBP8og5SJxWyFMyKcrj7Uk1U9eiLaC3INtHYuiZS9d3YCm
yGtCG2JV6tPI2KZefczN+Z1i6XxumAnKggskOVekRF6xzGM9iBAKFWllztUq5lU98GRg5xBNDegm
o4pLGimeznVFdnbrt/cH5dubixwZA/mWqFwmEflAI7vw16p/YM2KOyTTCLdjvhvq/lkFgD3UOkTG
Jc2AjAMG7/hUAGyZ7ePRiC2i1WRFW3K+hkkaJI1XAJporaDAzUJcvAXdRf9pNq34M6V13F9ELobr
JYxk41LCFAluuL1ZPvFgoforOy0IPYHdeXxCPBLph0QECAv1yI2OLwQvQk4b6afhs4+H8bO6klVD
iiQ1DviAOgcde04VqpBdij/ksu8gMdB2xHKKHMIoAJGMM32fOPPlsufeIJoak9XGvuPit+T7fmpV
32mUde03SQs8U9Rp6tQ3WM3wttC5F7s1s1HiflOpC/mlF4HARcRbeVGbrYvqsAhzEr9o4cTkeG9F
qA97/COY2xNOc/miNcG6hydmswzGlqIlHrDR7z5AtF+2kzwfo3+T7AnWHbDdczMDcs5bUgxNm9XA
GKStr/V3on8XKmeghVjwktEG3rG5BQJra2fr5kBssbPSl7G5yTcJU8Ze9o50Zz1+wcL9m7wd64Pd
Ol8acRVjM8UjXcBAQ/FUbMuOZIRjH/nJQqvPUM6FwxgdZakoOg7LeVHSS3oyabliHu8kHML+IKXA
A5L5wObNe5xlmMYofHfhT2ZjZm8RULOUldDVy65SYSeFR4owa/s83IEK/+i30tuB54NJA4CJZyNO
1JyARycoQl65/AmCeN/yJtv8N/u2By5sBAS5QQ+O8RAk5Uy2rPtX8mVsSqiQkyv6++dE5BuRpLQl
xMcUrBV94WEObgcv+m6OXol1j9Wel1NzeXwF5MpioxOtWwhHuKT9Sh4sb2Ay/FppqErwA5GMs1VW
eurPaZ+jkQPt90twQShWbgR5vLU8YyvqOncQpHF7MabSPykbT2pbGV/uNnAKzyf5eJi4TnpT+3En
iUOL/Izh9AySRiyWQTl6xo44elpFLlT4NjtM0oVoI6cAMrfKvlCFvloT24zTL0UvZzmhP0QQECRH
rCXP7c984vCFCOqcLVb3MHG1wEczD+KxL/dcyvGHyToN9qWwCQBdv3HxcpwqmUvkwJ5Cl2nu2qPv
0A5riKHBqoPt7syEAhwzVltOKORcBSkmctqnrEokyv/4A9mYK4Uq7QAdv6NAHG/uKlRnr3XoJVe8
v5hkL6E7jnLPMkDw+LvwW0GcvEs1wZNlFXAqG0NF+6GuK4WPPCzY4ncufV64HoKd3JH/pMLlkNpp
WOt4qYcjIeWn/flF04inLbn97gttBirH03H1lQcLlwe57pn2pIm+zhlzaq8U1Itk3+aQGZpcPxBm
zvmK8alw76/HB2kL0NKawG6cAYgp9IL6gzTpvYw/9QzBgQrxuUzTsJ0KRm+7aSRMEHI3W03JNOBp
HGClRY9GxXnF8AbaDQL2Kz4xy0HG/nUMn5Fr/HFBEc6tMC3vjFUaT7KZyHchmBSCym0vqKndrn5P
O9gAgOpWb7q8LpQTJzWhoVfqCXy+dKJlx8ABxzTRIKz+I+GFBcYdS02Y+6pGbLgFwxyL8M2aRSpT
KpHoSeMvkskVtkS57D5rCbHQ2qzdiKzkSDiLkxfV4kXf67WtRdH42HctVUq+eZOcBz3SVLbInGB6
8fxMfkRplTRbd1xezY69ie8PXLcZGTMp4PbImPfrUOH7PwYutrl8nt27ZrSyenK9CP6xV030a8NV
b9YBNAXywrJCALwkeODi7dma6GMVvl47N13oCFupesrWl0kuf4A6SKiXf1SyAS+4jzJq9ykxSn/V
kiGeUmtG0bkqbQht0vkCVsp01iRmXxoI2WpAoNrK8ZmbvTkpp4cgBrE4Y5UzJFF/5OU0lvnoa1aH
Zu7xi3PuDh2lWHHB3hHZrMMo4q6gv5n355l1YNtzXxqWS4BQPANnntyvcuAIRoX3GOVjVJLfq3P6
ST3BYov5+CWE0jpFswMdRpfWkbf/HCyn1Xk8+mAHWUpr89QvJk7H+/z3WRqOFEe5fGhWYPzTHh6Z
989axy2PeMJZW2yYFAOUZz68NgirZTejWk1ZqN3uJx7k1ckqynWnGMN5NRYngvPf6V1W828rZt6Z
XHqTELCO3iu5R+OOpHxzxD9qOjSwlEC9VglIKKWvkE+rY3Ye/LHNHy8ucZDIFySZnIGL30K8dMhl
1ehERYr8QYYqyGEu3RM7mVpJHnExFz/mf/IoL1Coj/3f1Ju8sb9MpVKfMZ3OGaDpnHJeY6fpB8wZ
pNPQaK+G3dYMKpmm/qAQt+ev5gDkg/rgfJ0LxMjayaGI+Aq1MDgSeyRiiCver0loWDGuH3rMVOZp
2nZHXLv35lz8PzgHkAi1PCv4wztM6br1Z1DdaHg4mAxwJJMGh9FCWxB7Wd3cjP5n1s5icIGY2LUp
2ZX+MhmG1N5oLdTCuyYLIO8mEnLLhKIiY04b818FRmUG7h43V431Uwqk+Nyy52Dc+GN8KcP4Z8Pw
nbNNRHUnbQXJmx0sH4IeCAE4HHKaAYXWI5BHFFCkE4M/cvHXXBCGgxM1exG/fft/+iTOWW6ccEle
kziNlLcC8Zj08T4l4nysQkfexAvcQwlpBUMYBPGLwn80EsbZ5hTjy2EfB02dD2Ea3kjf9sU9EB5c
tztV7mPWlcfRdUmeNQVzPY1fMUSg4/F+LzVY3ESlIFTpS43gsrAaPi7Bonvf8SWCN9/+UGctHjsJ
HRcijUYd5nXK20BinMllrmpVdJL5GsPuxhfsMe11Ify/I56VZnXfhf/qO6rMs1PyLJSx2melInE/
A8FAahBML2EgnZdd45Ksef/s9lEbLf/Dr8wt0gzAPy/CJYFvmRCwg2Skzh/25EVOcVpgX3Q11tV4
ds6wcoj00nxa73tQ/ne9LDTm8ukQ4cqR1QyIs3x9n6DYv6tGBUULYgrele2q967q0Yp5emNiXmEu
+uuxW2aejImxcBUjhq+ZQ01Iy+xLQiQJdIuV5Oq/y/dZSKYvVy5cIfh0QFdd/dWOdy7N2OcvWfnd
ad28UaZLWycOVlqoC76yUfGquGo2ayE3494iUeBMPN3pyP2L7nCA6jUycDkefxJn4PPjN6hf/4p2
pJDO5QAeS4SnGIYSeTB5ezI2C53ayblJ3UPv4vHUnojnTvg2rzT1LjVrcq2BcBBuG1YRUT3gf5id
VMFI4BwEAbm7YzHPRjjtq8sUxAsxvtl1BIDLD8IWB1PS0Cmjsp2yoAl3OJXi/hRrzTvKNYSuxfOM
bb/CYEvJFEE+tlA7RWtkDNSeoUDex8ha8SK/BGzoi2/OwjsoyoLS2KltkkeQQ602bojwWjLJC9vT
6Nei7y/2AqFxznVDenkXCRPN5qpwNiLqTr23vR0gyLT28Hpl3MBt2Mqe1R2gc8WT55fN9lq530f4
iI2LhKdhHP6BD30K3hw4DWPpI9f+4kGt/bdeA2iT7EAjAlRbpXd8qutE3TSE1a9teiApptBuOuPM
T7zXr6M+TFifK9dIfKEPYJ3JVbaGrdCvFsZvsqRT+Po/oRKNFb8afZP3SaO5ZW8QnClOv9MR6OUL
1MGT8DbRa4ISZaBX/HDyVNtJtpG5wnAVZTbHmvabCrL62qlRwuAityls89+y87AKw2iU3ki6N9WT
znbIdrZgZ2Jen8eGOwv2gx19tq2mTNuj8U1bcKuWs20ogN/cRrluZNT7tnc2zhAzjW6mmXy81t4b
0igQdp1J3eP23j7i+qw4uTzFnw1riSklDlOAWPBoduGkbdPhAOwLdl5q9mM60BIYt/Axh6mRqzwV
Zal8LT86QSBiLoqfM54XHfzpmosGXkbAZfwnxZSh0zuX/Zftg4qNaqJEH+outLDe4ulMilChE9XO
yAPMBxVLP5j5cMUlPLpkP2Wv8g0jp+bYHCtxgvhmlhPab+C2C3RnuqNFRjEJARX9xDuAT0vtkduy
gabeSF/5V0P2LyoXJuTVCXn1QHpHNBK8/nCNWUiu/C93ROSmwUDSQoV/oZZCjHTdVup2GV9WzaOv
F0BX6M/HpAaNgPvm3d8gtEaEurU1DzmER74OZTNoOt3+UDx+tqSoHIKzYA2Qs9eXQlgdOzB9m1kv
YHah+6ZGk9+qic08kMOZiJX6v/zTqI6YScWhpFw6HcmocBkr00HX3zOiBnPMEB4PzVBMEC6mdIH/
YjAxYS+grypQRgm1/WV9tLa63VtLEf6Qv3X9ubJ+YXixS7v5RUINgfiAHE90zKceDoTR/V/NglrG
ykXC5BW9lfn/5esD75gjjcVdnQGWgkhEaUVslN8Z7LJfgcAfdPRtbPCIBFAiqhxPequDBQMTmWIK
QjGANlZuM3g3ZJItBUSHGmKFMLLZEnecnOPfE7oBd+XjU7mJAOd1uo8w+biUlbjIt9+2fkYpo3gI
X8uTTchX17AJ55FHJwRcjjvHh0b5GUdJa/AcaEnzLUHelaP9IAzVdt+Y2wE99+4VUTN4urxIx/Rl
DgUJ1g5R5M+LvjfW4XrDD6peJbQbp7VT9yoM8P5EirBtMKZdxYgCEi11mQahDEssUk37xy22BSaW
rVG9rXBJzF3oxx2B2xVEKZAr47wCBVNlyncaG3odJvz9xJMXhJb+CSdupyyvItc0dg3LA9faU6Vw
PbHz2YdRhCnuDLkpFhyFvtwmmuuyUDFxYKRm9CYwUTlK7FCXuLNOpaCN+CfIVHNlFj6UBPOFBPX9
iowPpMqip0GRr9HCb6nfy8UylREsYX0AnniIQTz4SsYUhZUlTfrNXYfPKTYIuLRxuBJe6f/trIik
CCwWeF/GgcB5sVnqvyJx4oI9trEwC22N+ziP/uOm2PWxZQD58jXzWZX/ZpmH+a3xah2p1Bo6/lHL
1ARv3LFQxyy0Iep4eslHl/uC30sAP77a0BEb8cMgRIrnfbt8/lKcYnZ16jrZ75Erxh6z3EEH1pDC
ofeXX9v568lAemY/5OA15rGio4a+w35j3F77uCnnTORrDx2lXQv62QofgAFOx2j/5KG1/k4lzPvJ
gVy2uff/boFiluLPwoXzA7A0x3G4kN/kEG4cDjsXUQUvKNjgrcQ3mWDIGULrioWBLUPiLHCibXIM
0dPni663KTIN1oR6ezwFE2TbepnnyyrKVY0wmT90FhMQxySrBO/l0aFJKUhl7HO79TEP3gZDyHaJ
TkPo3AHIEzUfWyqyPFe1TPyyqPvgk1GsiV/b2l+kIizkoGG+C6VsuYXyiw9VrSV0fi6Yad784VB0
cKCCFBXI7QLP0NuAF/qWVdmm/NnFFd2I0xWFjSr/kQT+voKb3NIiNnKF1St5i2WKz5Hl3Iof1qlk
J84IoEQQXrf5xBM08fXDNHMghdF+Qt1l3YDNq5CeI1EOUguk83kJAIJ9qi/pZLRBqokRTrsWRjjw
qFY5erZn6D+Vt5/vGh3dHB3XZ4+DiAza/Xcy+NxR/9zL0soDmhVcl8sEy8pXbq3psfmZNU0dMZce
n0tQays/SnxeWEXqlQ4DZh4li2bGJ1BspirTSQW384zkro2JAIRW8sbnrgdew1FpK/z0H3lYrvFc
UDQG0Bf9Wx/kiIwpKlxgS7ko6gR2I9b2lBs+BCuHeXGcA/QRDWmknW9ZLKfoqC5T0f3Q2bY+weT2
rUaNM8YnKbbZKXdqBL7NKiADAjtwp1gNzBR4zzXXHiNI+mbC8D2p8sos5Yd1pdcQhGkVyPZ/WSOW
W00qeJ9L+yi/xGAxIBDz+WzgRFbKxk+BJzwiOUwfqnGHQPtlHrXbXQrGTUKJZkPvNNVTzXcSY5TZ
7+d+36oE3yh2dgqerCiYWUd1bM6aJJVjyTqhRYyVW6Vo41n3WNKOLP2m2R5Q+Vm6PWUXRvsIcBMR
tFOnHcZ1qfro0qHCDiPc1WmMdrORlerfP+dFQxeRuhxM6/VCZqxrc2WkL93/dsuOjnZMiffpk6gs
1dODaJ8SKm+1ANVeQzqAhmGJ6O8bOWBNsdlFFUhSR4ZMh+AFfAkHxYRP8VSE8U0rcJwpHhlHNZQa
rrGwJVLZyFmpzH6DFDJY+SsY6VGhWejUCNeJPAXSugajb+R6ADZeVN6NDpQojdYdQRzkvKJD53gs
rnMaqAu4qm4ddq2r/qtQNP3Yu/W7JoiyTfR0TUsjh89HrKjFvQzjxw9u/9bPqwkWW+UMBh7XH7Q0
iqNezXvRmfJ5IzORN5xXtvqdPJ+POxnK93FmAJe+gJ6oUoRRp51ZE1oif+LoI64zQaNt2RbbCr2R
JScAwLUtlaWBCaKjI9vdHDGc1CWVW/f1mXcahxysQXgcguIXJMUw6FXXJmN2VLYrpHtG77jkPYRX
3+U+jxFKXo/D5pZw5gBL1mC3vMtVHEjb6u2eTRqjMKQJMgl0w3g2O9In+JeQM+/pVrKt9lxG+9M6
ftOqeGn11bA0P9Pk3AbNBIilsoH0DWVIaWcjoDMtPj7E30eUMivXxHkB5XwOMtDkMm0dn0D65yIp
E9iUX1ZyXH61UOPKMGihuiUZWnKuBcbwH9vZ/O8B4KbXZJecCh5SW7B7oa3Vhb7LvCJbbti7PTTV
kofhXi0niDNxdRfCvY9IsmO7I0LAWEg4ML13suLlISI+yzC7SPE4oikzwFCghiBzPA2aB2N/rABE
Axbca9QK3O22rFO6P1QyYUu1ykNMeS0QDuRu7sTdS91YYoia5R1jUUzGR60ZZbW0EDQ/hSvs9nZl
JxpuwHs8GXI3UwMIMAtRPOHCVntN7FVBqkDVlRb9XIaRWauQRtPBPNF4JsZ78hsKuf6UcwB3cM4u
PltEDo+pgOh8/hIo007wmnbZH9lUV6xEW/TanWBUYZF3HBwWw5M2YFT8GGMWKeeKTS9avj8dqCb8
Yd//vOwB2AKdpH2dNurn/wiZOsXvAvg6P9w7zWk2LPsRK04NRS4IPr80FNgBAv+ORqDI9YvOuUqq
yUccU5jA1rlllDp4u/oXEiuouokTHfL6xW7TYSFpade3Kgnjp0X69xoguWoYM8cMLA4cLkqznPwX
hsXKXKEJdzwAIAH23QGAU8NRS15nRCkdALdgf5ceKMWDUOSN8I7K1jnS+OgJrQPjNF17NqctxCbv
xrn5DakkUuyjFSPXuwbv4bWCRjgC0aGevtdOKpNrBPBiRMT29ekAOmJ0774+g1upSOG/ChWrvCPr
JyjLo78nK2JuWAwyHnYXN31xTLsItzQ7O/eMm2hOm+lWDBsobuAfi07Je1394UGPYMmiow7MsyTv
gyjWKc/ivwHxdEwoZ2BdAc14C1otLhyvYhalKNFB8vSI4JWGGqtr73Cu/zC2IRg/0flHbqp9QB/v
T2b/lAW4mfDDcj3TNpBzrUNdEuG3h+3+8J3BoepCJuiR8/kI1d8bRu7uZDutFm+tBXEY/l80UkHc
xlh17WI4JzBOz2nvRkjjD4Ekbhwu045kUjqmg8xRqOjqNZS/Yv6T63kF6RoHQNgzZhG+6aQxj2PZ
fNPeNVj7LLDgkKR0WmahT6ZgMwZKm4sdSlyzVKyUO9WuBnmh02oT3qTlGyzAZn1mnx6M9Ax7BauU
qh2hOZX6ISrvwQkxZEfdISBw8K+1/W6SB0cb1ZlxV7vjMmHC8wXFLPybFEtPVjccP2qPIWjajjKW
1ko1qT1DPUdfj3Y1QmFIrvdydhZ02fDepnNADEqtLFeWX5aWQVJXOudhVyPMhwD5PRosiIncQeQ4
CLlZY/pXluV3/6uBnlJRULPk1Y9tC12IJffqEaaPavLEn0k/tfe0mCwD8kAvEt8nP8rlBgKICe/D
0n7JoLvBtS74Vt20KkzDAFaeJDEfKXxbbD0tFq66KjrYv0MtdUARsrIy4Knowh49pUaS5heVdQit
bxDzg9zx9LwOcDvhwM2VLo+TznuGrpuWMLZ3eN+BR7LIVck60JTWXNchZ5jpjc0Vs/Ac3WNdj+UX
NjO8uu2SNzAcMeO5wlznJYbszm3xJLF+V1PrkySiYfbfJncPBG3roQ0wkez4XO6AjqFEuDZ2Mxsp
RPG7Bhp9AUFBXoCfNg3a7/G/LRgcqwI5Qj0JN0+yLsECYWyPwznkkrwG/3O6a40vPq+SmVZxhE3d
eDgXVlQJbeAHqVT6L2ln6hXfxB1I66u0df0T5PzNNcBaslWM/ux2d5WUXYvCeMchCYdTR52hbrFo
NW32P/ieSzGrzQ9MPoQswALVFKxuP/7FmmAY70l4A1B1BTsgbqHVbq46RuEfPXJQXcwPVoWC607N
Djz1PkJ4K1yu4+tpWYIV6gG0xbwCPkR/JPc5BfDSU7rfcBQsg669Gkl+xwgGC0Ry7iXNDKSPuiJ+
zoakQggA89YO+lpDr/9XDaZ7uZGCSWOU4+hr1FEGU9+5Pbb891RTI70OtTk0VOzOQ87jJpRLpNuv
zh3nGdxPdJ8ie4JHzqf/kuP03u97qegfj2FDPYWAh/yHARDOIc0eAMQyzaOq7PUKUY99djXMJj7O
5N2tFNVvT0QvY8l3Pw+IyBnB70IWpgp+V46Ch80qtT3awMPN76adoR6tbnUB6VhBSKjRA5cmXU21
/JdcCY9ozKke+clFuOKBPkhz4rhF7+EY3qWS/7Ogt5jlAi9/GDo0EulUv8dkaNI4d+UE/bVFhhJB
LLF/gHMOwJXy0hw6ilkPsn0Xcw45wSKGw288nWQHIJS6P+1wcwi5VN/hdCMh70i7/XOxqB+PkFBs
6oGgo7uT40qmzUEUZhTyr43/sOtyaa2v9AbOEk2+EZtDTe0vb1ka5bZ3PsnNGCG9tF4SgGgTkRmc
f7B/7cipUMtxb/1jy+VDND4/po/RrtKGnX6zaBUsQKOBEo7BWCaGJ6WW/5FhR2xgVBq/BikTisgi
pfsCj/ZA5tK8Crq6fQClwPU4pCh6FMvCMv3vT/XYUi7cYWPfx6VrTKXlptoMaxLzAaGT3gR4oHNe
XljKQ8iFWHcCalYHc/YXXmBMIMfszU6vE6jbOQRg0OZPyOZD+furyW6/+t+IJ5GWz+DBMSeKpgdE
qqEwJv3wSBnrftLEHV0YCKGsDUIFM/rg2Ad1YAHazBII1hKAupyur0SeH4S0v8tJqUFRunJsVFcW
4LQWzsy5lHwW+w7ZGPtjwsb9orJGa3JIXIjFUpd6cpjTBG3rW0Ndmwp/nFgvlTnadyPpOYmb+unj
pBakdJXojOmqqCt2mjhzllQJFyft528u3BJlmdOUMzA8iXREoYXPilu6/IcgrWcC1smofsrJP4B3
65SiemHmwKPJZXSmi+F/7jyG0S0TVajTuyLNMX5bqsi7vncfc9V+NRX1wmlg38TzeqrazIex2HP3
wWfo0EaL5URRKYURxLPMl5g41vWabNiGKE+ntX5KobOqxmoSAfXotiKtqRCGdl5odI/J26E9zV2b
WenKncxYqDnX5sjfzYc/jT2XmeCQB8S88c7hb37GGKxOatEVjMLL31mcpp+qd/daVyz20NXWmoIr
JX1YQDY7l4XsVa96QYEIp8GO2PpPgLxIzeXePGbol7VWQkaiM3LAm2n7yDHizawVW7nJgmE3dDsx
jdA7jrbpD095aOVMWt/eF2QWlCOeCUXrSLTdqcw50OA9qLfkmiUoxmoelNTg/wlm7vxZ9Z7Mf/Mi
C11n1mJnzNO35xOiwx8gGqQTIa+Loytkaj8bEro8+rRJbAcq0V+nKEwlkvRufknhNGcUCyU31eaJ
cBpYVGoIf8E4msBObbX18bK6fDu9XAZerMxsZhHdMOpSpTOU3gTlYJLxYO+/gr5JSjVE92UStDOg
TDcJpvpPyxzwoUtroXyB0M7/ObJu1wbdoW8yTq8fcVRkfRbiTKcvzwJnCeKKPS2GhiX7KXP412dW
pJqRzHQtjZPGWafng6UswsD3hRiqKgdRe+i2nvgjRKXLVYBCHPywGp707QgPNZ54Thb5Tz4Kyu/N
ElXgTDrH46C3C4cqWwemEnuiYYSesCUXyoMLFCvi9U0gkFDrqtlXvwyPlsQSCNvqKcutfgSdnRXn
WaKziRHuSOkYn1o5y6POQ1UkdxfpwGNZx4axRdmAiiFppeEJqdPmzC3m4t06HyNCpMlZDTx1n39s
3RsfsMRmqu/tsrP+04nj1H+1y+hhaLLpQA+Y/4xAxsVhPZU0FJvfFUONqn1WkXrf+gMyZZ0Ik+HZ
araWjzqANlMU7SxpiefO6XbVV6iW7OY2Ajr81GIIVs1l7p2xxC7UcH9A7+x2J1trQYdpB1wR93U4
vTWTYpU/eB/5E/08795NAg2A50MtYiau0JPY5/yzmnYNi1JoDWow6j6Rl1+alP9Nw2Ms7C73RFZS
knH4eUAPlyjKxiLHymFyxH4HiPRusPmju5DHbz4gabg1wZ8UWw/F8HBkJzdwoP8FO71ejA8o1ARB
L7lh5cS34j6+mADOa7G8bS3r2fjOtp+9ZLpdcfRzB+G+dPcDppS8ZacwxbEiKvMsW7yodLH9DXDA
xc3T9MqOQbO6zWK2HS1CCEYhmiZVLImOO4JvWfuWbcEYGO347bkolXVoM9ArGdWQrCr08m5PvPYe
Hj/JP4wjVO9fsutbOn2ZNBCylcLN7qLd6GHLAVQ+iE4I+hf5q/y+VI6XeEVK8pcoowWvxBMoQlsO
HN2saRheObeBTtelSmFtuMZwrPA7QNkHTQ7PW01kLTYwGugPLo0UmrHJ/yawUNO9XjRiG+e8M5qv
hVlRFa4zcDX96420mXEAQFhVd3OgrtJAoqWwR5VOtTWqmYtaCeau4p8vrPt7nb1BwR0poPbQcsKj
D4PcL2igMmNhY7zm5V7RRymCA/rayDFIz3rAB6mLGNZ+wf2dQVp/w1d186zTuFYXvMoKfXxqRrJs
da4vhMRfP5lWJDuZoKe5sGDnwNc1YWnnR7pGO5cyGpfG7Xz9DIB00VmZ4Schlw82G2PntXsK5+Ax
SPfXz0OGymXCcbndRYHsKR7qjZfZaCtp8AhNieVJqBbh9ymkaF7O6HWyhSZ4AdcVFj+H2cajQTyJ
fldP1ZqtNTUhHHSjkrm/d9MBlvUzLReA9h6I72swRjKkvYk0iYaSV1ZvgyaArLwEXL9bxL3aqfdO
BooSkuN0/20W0KCjJrvTMvxpKK8/q4KR+qGPXTfNITlr2fhLt8V73KRjIlsFS6poGfhzg80iMgo+
/qzFXlRCJWqLPMSzvzFHEXdtnKYwG2h591O073jy4eT7q8tG62gMxjUJPkvMXLe5wkSQiQ1Hw1Fv
JkbZ0YiEEZuG036LQJzry63lCJKk8Z5Dw+uRjyTC61rqLi/b0UC5ZtH1Mskijn2iOAre0IuLs9gX
By9/9tifqRXtL+zzFFPDsqvLtTLcgeRJWtTvjjwT5EiDW15eg5lviaY2Lim3I/wYa1l+ATqkb9YK
fNd8cK+F+TbaW3rCMBW5/Xz+vxoSeuGLRGs7xTejavJbIuuIhYVXjpbzeWTmsv93MzS8h7j8IbP1
hzLTwjg/eV1hhImDdcIekoNuJqeLzBbgmUJogmINmU8o2eVNvbQkL1kF/Aj1h5Fe6LtyYf4WQAfs
ME68BQbMoPoWWQ0PqIsXj+cWplxgS6WyPUkpytaiFI0Ebb0/fKwzzIQSjC73hwaza3QMXIpLLaEY
goxEHRUnmsHd2e7STVQjPNOoR94saJ50FYia6Mfyagem5DTUnQPO2eV+FvK/JBMb8D0VhLAGPA4m
dXjBw1RSZOVMbT/sRUJpx3yJ91TfMbG9cf4VTxzDEfYXpoyWeDVn3vgebmOs7ppsQ1ykcAML3w6e
nXbAZ134o2JWpz9dCbUXA4rhWKnComSEatf1/2uCYms+Ihb5Iyevwu7lOoj+yBn56am9TwSCJhzo
6gTKmXykEpGeGVJycLejzpHnzE24PeSJeteJMgTI2rvl5zyrUjoe2bjgUf/4b2TnjagOH0aNoBNz
VQcVnbQJF6HujOccYiXYdl1jaEI9XYj/xyS32zDqGgACW0WLe+3dJ7FTlYsnqy6Xa5c4mu2vYBkS
1gclPUL3LsaOpk6cTqLWXbPSdQCGmXO1qYRyI5MMfDIOh5RHlLNDj9b64+dt2R/jYsQv9V23LdVZ
CtKPLJwLIF2lPYLq1wt2lJLY8sl02fF90Ds9V0O3Aslq28eEqJI3HvjE8fw0oHS+aehHMgkVtvTu
YQtptfCRwrykibaeuX6n9xXqLSV3/3sdMU0n9s3EYqKwZ15SWqaS6O9FsvocdqGTyNCm061n0H2B
dlZciAAkLD/ROYARLL3kFMPP2RtPsCPmcGvlEllVT6J2NllaqRQfeAynymmTrDXHt2roEcl6BIjV
IgeGgo2moJRW5cNXnsuBef14oVphlclsqWqiwwpCf78io9Sz500du3bVYCoZFIrlO60rl7m6smc1
HidroZKAoCARkePM/6o7nkzYAxJba/hMY7UQZ/5vJ0zeYlQj/fx+vNqak6ovcVmrYZqB79+ywbY4
v2BLx86do6csZY5GWQgXloCbhtMh1A6kkreNXEcG4Y9Loi6FvAYhwMac5LcOzkmsV+r0f587wAkA
qfpWozycgd+JeTtzo8pWxfe63QFqLnzvo9+OeT8xaLiGd5KaLiMBpECHgQE7Q/oa/KuTBpibAHgG
yK0mKlkWjrfcnrdkCktK4szs4be5x4TQ6TxJFsiilkV0K/ExAOYYkOe2gwh4TPROzVKsmlgH5Czd
6uoxm2yQWMkrSnxDdy8pAyssUOkFffinhf5SHbwKNaYQXs69JGO3LtIbR1v47wFagdni0cpdvN7y
SOUvgk7rcL7XDivVwUtnu5iyeGc2xwxdXXQ5EPsQJZglUKC2WUtCQv/7aZVqaI7uNIs0Z6jbSXuY
WjNOp8PnfM15ViIPIURFwgxxQ2/NOhlsYIOvwVWC3OGpTD2x08PcodmJ0JikfNRgPBq+98GNITuC
Aun2YYQpOr+EMiYJ0fnYd5G3kW6rqn0heSoH8QYvwDVEGVjpEiUfFxzC8ngySdkG+ejJXLxUxSzm
52fYniYXx/xIlpTVNIal6TFKPir1asEujYlv01euwrl/09pOoUanM5tQ5ph584m+7CJLKOjUKjul
W+fqyWGf6aA123GACqaioXq/SgxdJyc6qs5xoWwwdYAkpraXFnONpgxxz+oIlApz+fRkjSeQ/r9U
eoWaad6LF4A5JVah9yegc/S5Xu40Vq4htntp0qQtQmSHvQBqdPb8TtHoj/CJVr5oVOHmtwwaAx5v
49cB8nhDNAHT/sikg2FM3zeWyL1Rn4S6JGvNj9v3LVGXAw+8Qo5x+Nd88V+w1m3UZBlDf9vz/Ql/
ric3nZmU25uiBp38WbtyEwafYd4XYBdykkIh6g1xIVpsomotHil9T23EgWbrAvRtnlOOx565ZItS
cUmyQGeztUuDNV3/5Jf4C/ik/m2HrCQZPL2ZI+6ewLviB+lGp2oDBOCZyxA29iyizZF9g4XuxlIt
Ex6PQ5y9PqB9L1Vh8oz8JSQ9Po+LOPr8gIpwH50nlJjMQL/lXdeM7DkvfKgHuzLemTetpOhYNW32
HzNPNzBBmhNSxTZsEWT+dljnECfMowaRhEnBRjfqLsI2Tc5iGEbQ9nPWYK1AywAPc413S1dVqAnx
EVVkgJtUvHRpjd04zo8pJ4GT4XvExEby4vk6I3+yJYCiRyxcCggWZlcZ6O1QxgsUBgE2mMhl+Imd
eFbFbw1ZB94c9pglV4gmatLAgCCskBnakm2WfHtTPgLXISek5VlSFSlzMunYZUksh73YwZNi0E3Y
+w+wqQlX/wfjlg+RzCfdaXXj5wqGJLmPpevT1Yk9smHTzDKf+cXTcnymoiV5hVWvZdFDWdX2FcW3
4gcATPdgMVXi9I7r/QQAI6WikBQhUK8DYi0A1asN7xRCgHciHxrafFeUonn3RSi/F+kL0McEHklA
dwd913RKI5dPzTx8yQHLSKlnLYCKzb6aI+hoNfdxAfzJVfv01nU68I/avvul3TINoT3BIpqznCnK
QfNzB5xMF3glVG4/2Rq7LFtI4HlIuK+u0NQxs8GAJe7H4Pkrqahr9MTOgsWM/RP7UBnVPxPefuXX
KjYRI7S40iSt/jIAaD6mtKDdpZUWyd64bkdQSqQ2r8jjbd353dYabIqDY8P+ZKw9mcU8AuDb5sDh
b8q3smcIqv0NUAK5g8zYV984pyyqTOIWscndtS58nXvbo7E3RibsNepexyAsbxFYoKCRZwuTjDd1
6GMtMoDFpn6qy81Zh1AFw5b3F1PZe5gxt0DGeojFfjJ3vezAWCG8y30BurAtlqDOhA4Jmc6xyK1j
BWy+9RYp8R3HCZ6i7MN+5zMr8oCMUSaaeov+dBPYUIvtAqmBO2SEnfqhX+DXN4+9ym8h1JzEp56h
32XjK0jjNBrlKhiXNyXEEa6x4fveHZhy9ISonypDy1vvcAryoJDgogM0SQUo5L2CzZbUS9qL1+b5
2YYle35ym/ger6Wdlavha8KqQx1GDYC2y9tYy3W+Dq2lOH8=
`protect end_protected
