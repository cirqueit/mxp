XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����� �.���׶`����[ghZΦxVMZ�CfAgkej=6��2��X�e�_�U����F�����*P��8	�X>Yd�5+Yr&���n �2_���c|���Y@���[���z �60J�YoZL�J�hk͖�Ht�f���%,B�F���m*�Qآ8��Qt#}5a�ʴE�~t�>vK6�8]��F3�^ ��X^��.��ֽ'�/1��(��H�5H᢯lkI\v^$'�O��
�ZT'l��/I���o�Fn�1Y����=	���;�T=h	]�i�r���^� ���g*Piv�䗪\�x�19�tBM�g7L5���בּ��r����׶:3��G6�Z>ӆ�u�Da�@T�1�<rDua���b�fo�8��666��sپ;���[�2X�>N���?��Vb��� 3,�hd&a��.*a&e��l�)�\v�;�����	lV����}��;Z�����뽓P��[��Xʦ5�_�'��w;�$�{��XL�&Iq���p)�ׅ�3��t'Ө8J����j�R�ۚ��G�bY7	#ϋJMsh���i���`5�7Y�떕[�ק֞�5.���1$B��#�����|J�_��/ӐH��
~\UW-��w6�KhH����|S�ax�{d� ,W�K[KL�R�t�R�OA���,u���~X�*�׀�[xG~����ű/���j.��m���K$>Z�J���"�O �*J�0���LR�e��E�7��Sӄ2�����6�� ,XlxVHYEB     400     220>	���?QV<QϮq��tX"����q0!��,��"N2x��؛Qޫ��i7nt�����|��W��Ő�/���P7|6@�8�ǉ������#�F��,��� ��*U#�㤨7>����`B~V�	�&Fm|GV���f��k�<��=�ز+���9F���܆�[E�������/�5�!�D�9уJ�/k�����v|����"���/0@�p��RÀ� ��4D\bVA{��%���z�P.!��=cS�gBX�d�Z�/>3u��k�,x[�<��C��ypj��N\�wN�ѿ������L��@FZ�4��>r�:/��;��3�t�K��� ��U����sQ�.7���xY�GB�SfڭV��He��f�W0�<��_G�g����6
]�b�ꄴ(S��h��`����ղ�3W�8�|׏3�8�w�)�أ��9��%�+��UzF�S��γ�ڂ��G�#i=#�t5Iiqρx�V�]�E#����6��(9�W�J����& 2�G�bG�	���U�����-��Q,�i�(XlxVHYEB     400     220������I8�<�nw�@;�3S�����S 񍗟�j��I�x��O )"�<� ��ӽ*��9�m3��ƙ��킊�bў��9���q���#6�>5 ���{2
!�%2�/~�Ml��l��W��{����ÛI7��+��fl�9b�n�t�mh�k��A����P׈KQy�&~[�1��k1�)=}I�z� *�/��^��l`V٬�j"挹fS�b�LD��弅�N�3�GH����k
�vT� +�=��e�Z�h�*�ME>��z���2������W�T�Z��f�!r�������6� �_G�Y����s �:E�f���]��X����f���m�#K-�A�A�b2|yy�G�(N�?ߵ�7��o�<�ܵ\ʬ�]���/�xyWS�_�#��y�Լm
�<-A���x��o���L6�0qј��x��g Bi�4 ������j§4�pZ���J���ݼYe��Ɖ�dw��#}=B6�J_N����(t|��)�{��}qѫ �*����w��0�R�y���l��k�XlxVHYEB     400     1a0>���Y�40��@�zy���߼����|$3L9`�4��{�s�_��_��o�hQb�f�6.i1������ӆAkE��M�S�gd#����uf�䒡w�għ�F|_���z�\��Ӝ����⹑ ��Z�^��hT\���(�{�q��Ď�O�p> ��؎c���h���� ��+��X^�>�(I���B���r��;� �1��6��ej����
_�;�� t��f/d��oh+_M"S�n(9����%'D�;�s��.Cm�#���C���
+n2�t�rK�A��;��~�-����jޚ-_����o�G6��a������}@7�6\�7�k�R# e��=ϰi~[F$��a�Q��>��X�jA�ggew�:,~��S��`�ǐ|��XlxVHYEB     400     130���$o�c:G��=�>�q�xͩ0C����̌C;�HHR��iP���٪i��4w��遣\)r�1����&&��`1��N�0�@c��yS ����[�!�;�nׅ��M�Q�u��}ߍ�[�^u�o��{x[��*:�8/��-;ܩ��ulY��J��q���Ѓ�;I��R�����R�����'W���P���+�9������_A��b�	�a��^y��tn"B6�y[qfmi���=�d�*%0r��wn�'W�`C\��y~�z��aC���P�l#*�/�b�Y2�XlxVHYEB     400     140�ďL�2B��Mp��lO���	,|�A
M�a!�f?��4OY�(X�5�۱��r�9�[�7K�� �>6�w����q�G}�d�<��Lbw��]�2O�Yqپ/�f�.�{�連���J��Ff�f��On��C,b��F�Ռ�3N����;�-���l!?����� Bܾ�N�z�p@;���.�,�5��&�}���5 {���]�͏�P���9P��Y�[�_o˜D��Y����[|�Ģ{�WyxA	���]��-��> �ԝg8k��ڶ��|m�'d�+�J�E�*|��5��
Ma�_:�r���,boSOC7(����H�fr��XlxVHYEB     400     1c0�St�Zf�K5>�*$�^��tĸ�d]k�`�Y��Y�gY81�䛙��̫!т��b+����7�Vz���fT7��J��x^<C�ˉ�\i��Y�m�%%O��kT�'�p�Ӂ�)"9#��.&ަ�		���"��pk�"������t+�,��]��XiMTb��'��_ll�`���������
�;�`{責]�A����]f�D�^�96�(/���6n�?�\��G�A-h�V�d�[���%�T�椴E՞z}j�M�pB�3�ǸsH�G�`�	��eTg`�7ܥe��l���v֍�#� ������H+7VԬ}$9�l҄���Z�~��ϔ��u_s�@�=���6�,r �O�<���!;SW>��� ���`bb���2�FO*��5+�-��MR�4�g �-��j������[ g'�1Q��8�L�f�'X%XlxVHYEB     400     200/Aogb;yg���6���Sb�sc�`��o���L�"N$��㤼kd��K�����K��('͍W�%(䤮a��L��*�f)d�T%+Ψ	�Vl�	$-J-����?r�nȏg���U�֒F��zC)��G$t�뒖���{����ɡGF���l9�ulusZ{�m��8Ԇ�nPl���{��:� �|�p�S��I�%�m�R{��V�w�ɗ�<n.y���evJ8k0wa��g�S�c�4�(�V��6�e�%f�Xs�r
?�F�D�)�'�d��4�ݿ���x��̓6��O�:�b���ukɷ��iz+.ꋡ
 Ñ�1[V'���x�C�
�E�і���^��>�c��}��P�@_��΅q -�������b��:+l	E�#��05���S�Y���F��#��O�O������EL��dl���!w�m�)�'��m��-ݕ�[^QЧO�w�QȪQ�uγ�/���F2�8h�ܰ�/�#���X��.�w�=�j/bXlxVHYEB     400     1f0	� Oa!�Qr��Jg=P���s��&8J��v�' ����N[Ƙ/���q�QRw�o�!�[�L�o��]�f�P�I�>)n�̮�����v�Dt�b�{0D^��׭Xq3xM]U�\6$����̵�؏��ta4Q��|�4hK6lㅯCY�&B��_a���MҶA����?��4A� �Wh`B�&9�;Ķ�r���
���&�<��#�5�p>���u�*%3�2�p��{���dە������]9��E+�v`s�aLq�ⷉ㓋1OEy�Wس�{�E������V�Q����ڷؑ^_w%ߙZ)�lxo�ɲ�t|4Ǒ��V�*[��Gse|B8�F��bs���Qױ�P�N��Sw����î�ٰ)j�*�aaz�<���4�8��2L����Υ�R�Т9�z�S�-���|�f���+��_?�p�h�ci?	��%������Hb���+Qk���@��{s�#R��T�Vk]��M[\XlxVHYEB     400     1e0��2���4l��#k�>� ��p���¤r�"�h3Unܓ]�a��}A��uA���P3�	�c� ���7��&�5�V�i�����V��Q�l��߯�t�b�@�2]��rt��:�%���>�?��-oy�ٹ,�=� �NC/��W�C5��X�`R`�$$�<��� ��Y�%@;1�0��a�$k`�ĵ���t�z�<��5=�ηB��ec�Z�@�؅��e���I�V��Et,��*tNF�P*�``+�x���?��j����t����
�@�Ο��*�݁ _�·�7g�x�ޯo�m� X��F�X������wѴT�I�����_%��6҉t𔕻nk9p{R1D�j�-\�@�Ȱ,�L�k��-��ܞ��:zP<Zl����8��o�[jF�-�����At��=C�-��?�b�>l^O��;3�9�����A�矖�{:��@��k�XlxVHYEB     400     1c0|S��"�IxMCd=\Zj�!G&E�q(s��0�e���!	�ik�& �f�T*�حG���3iݩ?S�ݢb Z�F���hp"X�6Z���*�#�[�ji��9�?��f����u=3vI�s��񢷍H��6xp����b~Z$��d��3I^��ہ��$
>*�zo�U%�Jٜgc�;d}��*@���ܧ��%�Mp~�TH�,^�,e��zB�����(��aX��"� ��i���E*�m�,�A�̉��a�?��w�k��r]q���j�ۗ���Ԁ`��3+2��U��Ҿј@����<s�i8�B�3��:�m`��e��&v�y�z�j���Wy�A/V���@6���@R�v�G|@��Xb��A!z�L��4���CZ`'�\(�6�ڠ�����c�
��%4}�ؾf@a=ߜ"��/lO��HD7���d|������2�MS�N�la��&I�XlxVHYEB     400     130����7�k���JX��v��-��@�9�=@�(���cE��t3����D��hh���ns�x���.���;�dj2�c�*�U�WHN3k�_74�C��˳d�Y���n�:�԰� #aˬ��������v�iҲ.Y�0 ^�K9�\���$���F4�U�����b�#��s���PB���tC���iۻ�����+JKf$���dN��|��ҋwPÖB�(i-������T'�@�`�"���keTv��X5��	��[�*lA�N�`��z�^��C39��eA/���X<2_XlxVHYEB     400     170C1�Zԝ���%����db���'ڜze�d�U(c���O�X���Э���96Z��\�dIC��V�>�y�NAb��vN��$#�k�}���A����8���̔�y���@�sG)`l�?��\*T��(��Q<U�V��C���@F2�����BJ�)˸�������c-�B�G{% �d�%�i�?��[�L��0���)eװ	�sKdN�%d@_�^3��(�,�,O^~wQ����v�d��T�)�nD�C�<�&��~�t?To��_�;��*�H�f�y~�7%�������#�I��si.�C�&U��v+)t�=�"HD�c��B���3?;���Q ¾�`�s��:��h]�<Kj��;"XlxVHYEB     400     110H�;p?�t�\E�'Č��V;�S�"_!`:����բ"��:�W4R�qv�7Ҟ��YL���Q3��f?�#FqN~(,g��i�ռ��^ۻq k�AWIbP��5&�Wd���o4����W��{�;?��v�����K���tSA�R������a1{A8-K؊z:�wF��ΏM����V��+o�z�rGAr����V��^M�	�$�����4��`�S+(��p�'�=0�c?��GWl���8	�Ҍ�^/���`4XlxVHYEB     400     140L*��^՛jQG�Y��d�B
8��Ҟ�y�gޠ*��a0Δ,�Q��./�p�T�\-��[�v%rB�VA��f�x�(��MbZ��(`<��9�U�K�<?{G�(�3f
gǈ'�����7��������q/@�E!8�Z!�m���o�Z����$�ܖ �������h�L O�t�X]�K�����=)�yH�/&�UBY0$1C3U���q��{m
�2} �[����lk������`�U���4wz�������I}}S7�RqZ��)c=���?3�ÿ�u$-¬�C�[�rI��[�ݬ�*�Vh��XlxVHYEB     400     130QΖ�3c��i9ݻ^�0��Q��t*�����ّ��e����1_����i�T�o�v-�����Ӻ�{k ���\T�5H�8��R�{(v*�hQ��<�Z�N���%���H�K�L<�S�L.�bN���F��5i��'������AF�|WlH�rf2��i�e���Ιp?�s"RfqQ��/�[����X�������[�3ʬ,^]�*�Ot���1�^�;`kߵ�rQ���U���iȷ뤷5rT�ͥ���BIy��ɢ��l��_u�k_�����ż�w0qXXlxVHYEB     400     130\fy5��M
��Zo,Y�Qx̪1�����ꄱ�_,Ms�w�.�o�z
����}H�v�d��/Lexf��J���BBL��{Rql����i��)֥҂O�&qL���" ����"=`K�I7������GW*�)(��(���~������{zk����"�ޛ�l�� �>i�kG�R�M<@7wi
ł0L�f���2�qH=�7ܷ싵�K����br�t�έ?��*�髸x:�a�a\��6�L�z 8/��� 7�J���`��Ea;2�KD�W����7:)�<�}����[N� XlxVHYEB     400     150Mr�o�XS�ꗁ���ʄa\ｭ�@��@�nٖa�}��rfV'=PaI����RKd�w3:z!5��θ�'E�d9�IE*v���E��oYw���*����_�c4 oK���ӿ�p�{n1���Q�?�H5r�O���#4K�fYp�9=1�h�"�lG���ͺaAm��]g�ה$f���܃+����pӱIK	:z"0SQ����<gS��K������.}I��3oAWvS]f�W�qب�V!��@Cm����p�A��)'n�����'14�n�FKM��!K�:��6�����c%i��=B�e����5z��R}8cɯ�.�`q�v�E���XlxVHYEB     400     180iB��?�%�IYg�9|�=r`&L� ����қ�0']��������ș^+�uI�S�<ڡ�k��a����R��@��w\��)���|��(l�z��S�81=g����{���n�/B�X)� N*m�#�mp/�c���#J߼��֖׳QV(��L? 7Bv���L� y=J�d�$�m��C���tj�N��ܹ$�w\|/��(�����Y��?Ph6=��8�I~=����ơSY��%��\Wc�2���%#�~X�c<�!�E�T _٘6��(��bH/�}���4����5T���cR�C��c��S'�)	����V�F9,��y�R*��CT9{�r��cH
CC�Q��I<)Jp�>��v�E�-��Ό
-#�j
��,��KXlxVHYEB     400     1d04= }6��~��V�G~!G7%[[�I�a2<��Tj2:z��A�^3��Q�~�6�/F$��9�E�GV��ʹ�ky�Vcҟ���,�P�+�?�E���?�
Mb���1�}@S$AU�Փr��θӫI�e�yT-T�*X;��{�%Y|�Nĉ�,�'���S΋h�Y�ޯ��6nCPu��u���z����I<�r����'j� s#��顝�B�)�L{��c�k���>q��T���5�g�Bᔲ�	]s���ذx�DрA�Z���*�&�uQ)���= �l*���q���֫2��
�7v�5����m(~��'�j�fcfw�h��i^õ�!��{^����Lx�ݏ^[�鉊U�:;9	�:�,IQ�v�ҿrW ��>�l.��t��{���ԯr�G���6����'���xTWk�u�O�XDS�.*��Ĺ���hݤ��C�dv92��'XlxVHYEB     400     180�j%��ւ��il�O�����XK[�L>����U�	�W��_��ނ��OKP��j9�$��ת�S�rM�iw�O��})��A5�Q̩̿���.Zk}�A��|�~��������~5B�BSSc?����8R"u���ϙ/6��=��N���m�ba�YT��;��� �чTN(
�gH��8?���2N�BZ���m�O�[������Z'��ج�\�@v�g�xA�;U":<�sQ�PVϵit!H�;�DX��+�5���*#>�BR�m��E�-���bqTl���ԄW�"��9E����ۢ��8�o0�'�,q6�5?]�J_�f��k�4�y�>��Bw�>���4]+-�ó�Y͵�Q��hݣHC;w�;/]~���XlxVHYEB     400     150�Oշ�gȃ>՞�f�`P��]w���zM�yY� �!X�Z�b���~w�Kn01��rc�+˴��y/X����r/�n��$ƅ���`�����#%wr�?`���}NQ�~ԃ{�c~���\ ��b�К�:��mS����idL4�!�c��kӛ���C	x`� h&����D��zU�x<i����Yz��Z���|�	�Oʰ���O�ʏ&��	�Ë;�Yz�sS��ѕ�8���`h
F��T�*v������sV}ո�%'�?�2p<��XK:l�-�3�@��M�\�������͠�o��g��㼔FD+�U8H������XlxVHYEB     400     1f0�ɗ�>a�ueF����c��ǚ�L������VR�cK�zw2fA��P<}���g3�.�u�� ���F�� �(G�-��Nz�P@��w��ǟS1;[]Swe:�*��?ҚW�*%��c��jT���4�.��
<X�x�����=�~�-_�O��4��R�"����l�淆j�Մ��W���(x?� sb��'I��X��ؘ2.�.�l@֙.p�e�84zw�x�$�F�mc��������閄�>C/ԍ�fS������;FT�}]��uq�ʛ���:L����L����n����%q�EǓ��˷a��/���hv��,s�|�r���h�����Q�|�%R��X󎖾n�\"�{�~/i��[���.��3r�!k�5��(!���
� Β� Z� y�[HD��-<P�p F��#���}e;�y0�X�����4�FkJv)d`5����Ü���v=��(:.����<${�W�"��I1t�ʬ�XlxVHYEB     400     190J_7	�BM�l3K"vC+�?^����1�G�S!�ש�����3��)��!�I�@��(Sȕ�������+�»(�X^�+�� �6'��ɽ3�ŻC�ѐQ8���=7�]�pV�-�ľVﱐ�����4	��w��Q����í��޺C6@+#>����ص����CDzD���P �
W0�dNg�� ��m�;��Y�q�]�$�w�3A�ή�wQ�S�,����5<|m�Z\州+Q�ph!+�Z�&YW��V5؉?�⯃K�	�x�y�ٜʧ$� �;"�=.��,��hYF(�E�cɾih:?&��`0�T�����M�T%���bC��D�D���J���7aI��"���f�_e��b���_EI��[�-����lVN�]psd��kۗ�*�g�4eXlxVHYEB     400     170�3������7�D�{�=��8�n�ͮ^���m�;�+�
t�q!����jhR�:~�GT+úk��Ht��������#3���F�+�qƷ��[g*S�S~��;OCĈQ��!WR�"N=�>��,/;Q�(��d�m��z���2RzaH����^�Jw���z�E����V�����ncJ�fy�e^��\����a��pX�0(C�Ux����屸�Do�����9�8t���O�M�<�Ƙ��ʓ�9��ȷ��p�����$���G�G4_��:��UmN�p�M��oAJ�u
Ⅽx2�_v�:{ݩ���j�|�^�EnJ����}�fo���v�z��fL�T���{�u�����Z8�;��!YXlxVHYEB     400     170z�b��ٺ�~�T��	鶬X#R�j$��6p�*�������7�h5"�|���i��BHn�Tɰ����eU6(Fc��Jv6�2��F�:��#��&�s�-��<�1����f_=�@����l�=�lG8v�����r�|�M��V�g.�T�]� �Tʙ�y4���OAo�6���`Qx c��Cv��n���48R���dn��忌�K=7ʽ�����G�ұ&�%��&���(sT�K��U�f&�WU%��w�:�o�ѽ�M>L��[��5t� )#�C��D��N���_hr�Р��76\
,���^�k��!�6s�L��߄zׯOR�"�����So��VA���~��Y}��J�ע>l���t�����V�XlxVHYEB     400     110_n���K>�hB&���Ϲ�lmC�0�F�6�DR�T����m�����J<�:�I��%�D��M�q=bJ����<�;���Ox�}+���\���zR�����������C�G�E�y��f���5;�
�],�=�S����!3���WL��%�d�S��A��t�!�ť9�s��E�P�)���F��Ȣ�0�����k,�s��9�).ں�����A�`-�!0�
�k�vՁ�극��v��lo�Z�J:g���wO�7�_�uP�A{:���,�XlxVHYEB     400     120��b_J�M�qd;��ʲ(��NzZ2>pݦ.��!c/5��r�_K���Z��emQ1�oj��m 1�}���.�,/���r�
�>��Q޳���(�^b�l�����.����B2Y��\J�9���o����z�3=�U�kQ�x�����m����� d��,��`8��u�Wk�R�y�w�3uԛ��t�/T�h��_���`]ԸiI�:���R�i�qW�70��?�`�V�XE�ul����p4��!���\��0�Kh�F�¯��=�^�O�'���8+�L���'XlxVHYEB     400      d0*���/��3��j��z�Zm�N�Q_��R�U��'��|�H�i�@���2%6&d�6ր!_}���+�T�[0�}m��6� ����j5d"�<�_��>!��ebݒ�ٲӌ:5�<�����>Ab���ճ�C�����z���N`���|=�]\���M�Kl�j�mI�w�ѕ�� $��YU�骐�y���XlxVHYEB     400     1404�uc`�@����J�\���Ȉ����R�����qTnm���jM�`�uPhi��J%���0!�S%2$�5:W;�?� ����vf��T��N>W¸��5\���E褯ٮT�jQ��J��Qݭ���_,?�v>����H"�j�O�ҋ���4X�6�2�na�����0)� )�W��o����?K���6���nA-T��n�<�<�������^X[��ϛ�+��F_�HM壦:�JuMi2C�RDL�ˣ''�?x8�"[0�0�>	�G��V���Ä�����(U�Z}���ʦ>�A�*~��͓�XlxVHYEB     400     140=�;����?57:j��#�"񳻟j4Y����D�/)_�?�`8 �Iۚ�F�sqH6�Y�e
9Z��6*O
�gn��3��]�A��#}�iC�ޯV:��Hm����w�����]8�:���s�ko?���K��Ф��Kr�S�1�LD��F�sY"t��h������
��M5)��?L�����0I���9L����L3�Td�*����OŮ5}��U*���P�~�{#��z�Ġ,�m���S!��{\Yr�k����,��S*4���#��Y��kd��Wlk"�1=[�D �p��|M��|F^3c'���XlxVHYEB     400     120�;�%�薟�0��T�ě�5����d�oF�H���dm�+q�� =�ؒ����JM�9�G��>#/���b|�!��
É�i4���<�FTL���ܨl��W�k�	ȃڽ�>��i`�>�����1'�$��	��[���Q-��N̰b�h�@�^Z�+�. �	r;ة@�{!� EIp�G��+W�ݦ�c[�V�=c�3.�;�Ll!��X�+�N���htd�g��J����o.�ѾP��}C<4k���,���b���8!��bg����y�|6��?XlxVHYEB     400     1a0 &�)�u��w��7��w��g�, ��}M�N�c\�������qk�w�@���hE���2J������$'@S��b17�����k7�q�v�2N&� Hts���
):���x�my�f�ܲT{���:Ob��c	E4�h#�j�&pv���s�7W"�:	*��v;�6�ɳ���)yw����Qlȏ�S��u��-�.*�mKc9ѕ4��Ѽ|��w�gB\>��hM����E-�J�I��=p]�+~yp�i��B��Tv��!�
YE�[�&��U�}��}��\��k��)t;H�V K^P2�<zW�.H�zsz��mQ�=`J��PuH����t���/w��\W��a���r��G�Ao��<���h��9d6�|�l���5�¡���B1�l��QXlxVHYEB     400     120t3>����㜩#� 3Dn��������p�S2��t�2ii�ki���us	��ן;�[��(�ʾ�q�o��1n�;�w4���1>d����i�������1$biW�B/Z(Kfj�����f7��H�Qet}��{�ץ~	�
��ߞV�$�+/�=���'�wK�����o�V��M�-"�C\D_�e�Z�1�l�>����qxLZF��S�\�g��+���6�ȇ/��`����M!�d����('w�3%26�-���,T�J�Ҟ�s����W�XlxVHYEB     400     180V$���2�m�ܱ���M��
)����i�g�>'-04�a����Y�q�ܳJb�d��Q�6�p�^�
<|ǟ���MK��k�x��ML�Ek
Ȼ2������_N$�}� ���y.��������r�Rt]�I�s��P(� ���S�\���{�ڪE)Q'���2/��r���v�fO/�QW��qj�_'~^F?���s����^�&���ѴZ!G�T��rs<Q��a-����<S�{�C<k䏖� ��=�Tu�tש�	��Q+\;��.�h_X7���\���+Pr��C�Լ=
.��2�)_���4�L-#+��a��B/5`!�[|<��i���i\�@Ī~. ]��jӁ��K.�iNXlxVHYEB     400     170x�a�@�m�w�o�%)ܒ�*Ip�Zuo�-�G\n��Y�R�����y�{~�2X��6�_
NS����QU�V�uVZ>x�'���*�
�ߙ[J��0kgK	������N!//,�v�'U�½�ڝЁ��m���ֻ�~cx�����	��{���ɏ[����}}��͊"�ɀ.�"�Ҭ�����U#.�� D�J{j�_W^zC�l���4ycI�ע���r���)��A�������f7��p�8�g���v�s[�B���a���D�DדPܓ��9�"/�)M����k�۲�K������8�`��!��O6����v�d&�*���9�>瑳/[Q���I�B�+���l�&l�R*f3��~XlxVHYEB     400     1c0H�ߗh�K�[D�b���4��l�a�c�'���kc���
��̊e!tǛ�ZUxЈ�y�1r�V�b�x���>�:Z7y6�{�����H8͝�tGkZH\�"��斧|S�4v��~��P�] ���z��|y���e�.I�H�� �1�8�ւ���!�����;�U�q"�/j+�{he{�C�`�!�2����1�|�_�{R���8ߵ�V��Q�,:�;0պʫ�'��
��%�� F�����\�{2�Ǔ�}�׊����,ݍ�� E��\＿�#��I�փ ��Vb�r	�����(���{K���d�E�z�-p�::���㞌�=?V���*����v���
�o��b\3<F,�9ӟ�����yLn�����ߊC�B�����j,n�P{:���=y�Jj_[��Ґy_���I'��O���0�xquXlxVHYEB     400     110c�n:c�h4��y!S8 ZY����(�}υ������a�k���w��ֿ��<�Q �2�>�D�*ZOC8im?�QY��,_2�@:B	�b�b�(��\��m��6� ��69hM|�M�q`���QKɄݤqNw���^i������Ő�)XT"��	����tR{�xoN�G�Sț����4;!?�G(��;îp%/���U�lΝ{b���-�$�,G���xj9l}A��yz�:B����pg��l�V�*1�
�I�h�hE7n��XlxVHYEB     400     170���GjIHϭ�{�m�r��"��ƚ���m��èwH(V4xRrl]��5������̉M���{�
cE�7���捳i�&Q��x�~.RHۇ�b�s��Z`��+����W[Rd]�m��֥�;���(�k[����J9o����+�#��#�������Q?��3S���T�s[>rw��-�����-�u
#;'+b5���� /������]��n���o�=���$'��	`��%)�� �a҃�xP�*k#��NT�(W�� ӧ�b(���r�?����?�c��a�=/I��
���u�������@'{G,�lm6�Q������� z��P�J3���_�x�l�^�3��%XlxVHYEB     400     170#,!V=��U�����$uj֠��?���c�U��DM�+����Ru��z�$vL�Q�`j�G~*p߫=���Y�EkT{�>sgs%\]{?���?Y���uH����k4��U"�Bsސ����73� 2z���ɪqR{)�pE@�gtd��d���͉�� ���؋d
����vBXXF�s:�>�Oy�!b�X8����[�T�,�>k�[��&8��TY��Z�K�0C�{1.G�d.<@p/ �6�7w�&o���P^r�tI�#�	]i�ߗ�<D_��'y��N��N��J�:�|�;epA9��Ba���t�^젙q�����+�!�Mc���D�`�{�5�Z74ҪL1�=��/��
;j��/2XlxVHYEB     400     1904��<z� �v˲�ȁ��F�͑�\1Ԝ=��ά�.L;�`	cw�a�9�2��>5�(o�%�]��Ѡ��E`�,O{�(�$N��n�<�)|+��g)��m�O�h �pv�%6�m{��
4��iL\!�� ���Vkq�m��"|��o����v��҃꾗SW^�Oe�����7�~�仛�����c>�_�4'���R�Ü�9j��aE=Gωc�����E�1��6�߾OWu�����H�`�T��Q�Z��IЙޗ㑐ص�����Ô���� �0� �~�zjmR3oB=)`>�f���r-H,���T��V��JJ��%'��<��w$������k!����]\M�X1��J�Ǉl�+����GBGU�a\����A]ԯ��
XlxVHYEB     400     1b0P��{��ns���]?]%T�Q���Bol��j+	���O�2��O-Ӳ=��#�$�Cg&�p@ �oaO]��)���v�>�(��5�|�E��(������[h@�U���K)�]7W��Pw����.�7��㗶���k�2�Jb���3�Qo��[�h����m>��)'�$SɅ�v�H��p����I������y��)J�.��@�Yդ��j2�?V�VF���ږ�R�_\&aӠ� \gnN�bx�lO ����uar�Fʊ�;��p\�!�/��ЌV�m���c@�K[a����;��G�k�7�[�=�K\e;��x~;�BG��o4�NA�±2��D[|f
ډ��w��:)F�8��U۸=�BI��$��"I�j�����Y�f=�NPb�:������)�N^+j`��$WpP{���x�'N��XlxVHYEB     400     1b0��o
,�ӿ��7��|�v��T����()g}Ў�ӆ�z�@'
��������Z.�!K��߻mo�Rt���Z��4�X�:���Nd߃z���r���8sډ*��.�ð��Emá��D���Kr��	�~���ǻ���a���쫜��&M��j�"��m{�p�1�\}NF2_6����WL-��6"ǃ�W<��B����<�DH��'ӵ���Vv18L[��Uk�Q&���O�T�	��DUnJ!��}�3�d�����iM$rr�	�GEv��(^V�f$6)��2W�j'8s�}�o����s�fO*PzK�L�t�.ƶ�BP~�`�k��pswؚ��ϱ5+����cVT�&=T�=5����Mw\XJ�|�
Z��y����S�=�Ѩ�F����7�|6!��B�E�⧸&�zV}�����^��=���XlxVHYEB     400     1c0�]�e,�����xU�uS�u���s!��[Oc�1z�@�H!]?��f`��\�x�<d��/Ow�g�j� ������,�G*�d\����ط�3�n�E�Ws%��� �Y����W'�����4�.*�"w�\x߼3�[�ġ֖��0T���6���Y���m^���xx�6�Ğ������ʳ�n�������4�g���Ь~{Zȍ�{�z��qBFC��$��)��p2�G�dy_op��^�8w��ȟ8���w��Y5*�~|�o�o,�Q� ��pz ��!�V�B�l�]C����y	���[n��XLHR*���F��{1�>��{/�<��?�C1}��ۄ���3�˙ԭ6�V�g���sA �mMS�^.�A�yRx�D��8�\���+��W2�H�n�*�TyN�/<)9Y�:cgXlxVHYEB     400     140�3���]U��F���U�h���Z��v��5��(�T��׿m�H�������W;8/#?�-����m���?�oyzB�j�}�oў�?�K'-���7��=�1�x�&����'Gb�?_��l�w�����Y��$�`��L�i��;��Z��,D�|���E8�a^i��Itѐ@HD]���E��r�ߏͨY���5���Ƣz�pa,n|��	⣾�f�m�������X)G&-�Y.u���;iB����$?��z<�7g5��xl��Q�y���X�KtT�-QeB���ƫ���:�X��ѐʤ��XlxVHYEB     400     190~ZF������e�0.6����5�k��\���f�����5uV�,��UF�0<]�4��guMO��8c "����ҭn���Kk�$�D���M���yɤ��F�����x�:Gc��UV�&ܴ��/)�إ�R�����K��ߡ���J�Ɛ<(.`��e�#Ԩ�s��#���@��v@o�$��H��)�KWɂ%��������Dʦ��B�H��`D~Z����P��C��)�W��!�<f��MLX|
́���� �Ҍ;��c}�9��i*�k�"e�7ߐA�i��^9
�s�,-ēn���T'�цd�D�茨ӌ�Я5�/.H��}��
v�ޛn���&V}X��rIm$��)|��$%�,���µv�Dtqն�j-�2y&��8%XlxVHYEB     400     130�7����=�2�Sޅ�'W0;N.�����M}�=n#�y�(3��t?!���W*ORA5vBB��C�"*��� Gv�?E��DKG�7nFE�g&Gl��e��W�����z�9lY���l9��(�X�	�J8��#�@!��x8D}�GiY���搌
���Vb�<��J�k0������/2�q7���Ά7*��4ϟo16�*����L��Nn�D�$������W�`D�sPn�;V�:�A�~$�/�+�h��'�Η�᤽����<h"Y�[	X���N��������hL���
��s$4	XlxVHYEB     400     150�<Sِ-чN~��\�_�	��)���,Ly��s���H��θyʣ�k���׊�m�S��k�t�5����n���oK������=	��K#�'w��׸}:����M�-�sL��
L=��p��#\-�����v�8����U��A� ����kz�h�.��w�����wC���N�C4���G~��B�;d��<5�m��*�pX�ck_������lR�꽬�<ב}��?Xm=
�
:{�x�����E&���oFj'��k�Ε��ȃ�sX�8Il�<�e:m]����h�Q���l�J5�g t�٦y����6�B��XlxVHYEB     400     19048�]f�A�[�bֵÉ�^o�\6���2�}�lgԶ`(����/[L�"�ϲE⸗��`徤��N����� ����,���_?���i��z�(����#,�e����d�c9u�z�K}j3�s*�7P� -�-�����i{*��3P��۷��t7~�ιU�M`NJL��E��8c�~�@���$��� �e���q�[� $�J���e�����Qm�#�8���D5A�7&W�����yxj��i����	h��lW:I�Jȴ�Q��Ch�|�1�k��p�?��&�4�6/��5BӸO�O:-�("kff��7(`@�]����������e���8�,�Y���3��������Ծ�P�	��=�L��~��#�>N-<�h��[�1����l�EdXlxVHYEB     400     130c[^ᠸ
�sP��6�Y<����¨��v44u�䧽��L#.��śa�)��cr�`��8�N�дxf.�~-Х��=+�V�md�Be��'
��f�j�&=���2N.����k���*���&J�A�(����dx�bJ��+�Ex:@��Ǝ
-!	�J�I��bB{�2?[W'q��Kj���ft(�7)�<0��h���Mrcp�ޕ|�`=Qp��:���ʪ�8��+.� ��sHUְe��:cS� �aõ*�(S��-(e"���.�?U;Pj�;^�P<6�I�~�?��X��RJ�lXlxVHYEB     400     150�;�G԰�l��3��b=��-e!LdL�E��k�JQU�!���;��W�O�p�����
�O�T��z�:��m
M�pp\ �Hƿ2�� C��1��^a��o�R��>o�]��*K�_@��ם$Gi�I���S�w?�=F��,�����-��N�.��Gn?�pC훭�כ��5����v���CN�KmUI������*a,`0HjK�qdRo�LM����K�I���3q,���6P߯�}�F�d/�b�q�Õ��/� �>-k��'E��1����@v�{�u�� �t>�f:p��;%�i�^o:Qr��7}q����<��7�Ǘ#�qXlxVHYEB     400     1b0�W�!�\����!��ko���R�4Kq�'����X�w�
��7Q�
�Mgɗ:�N�U����_Ѯ��+�n�gV[�,�!���ʄ���ж����㭻:���L}��3s��+݊�����P�?�1�4IT�+?���+6�mXP����H��/��I��) %L/kD_
,V��L�V�}����;0�5�h�p�0/|p��<=��T[�QNS�'�%�$���1�{��_��᥿�i�*{�;��0���
�[�PG'�b�*t�ݔ<�83�����tFz��b|Ot�c(g�Z�!J��a���9���=@�`n6cS)]��v�"��E5�9|zAۉ�E�J���|�|Q4H�Ѭ��d�س	�w��S��<��by��T�l:�{_�6:�c]���?Hy��|��'��XlxVHYEB     400     1b0�+ h�\��s,�
df�tjhF���o�ρV@0s� ���
�o�%�Zl8�}�eC6�#�-*�ND�����|�1I%�����; >0�z��K��P}�?�t�{mA��`�ڎ��ґ�ƴ���G���J|����(�vf$�7���"����˞�4�V��Q�}���(�#�1u
��(���d�s��5�xb�;(��=�l����Tyt��h���gm�ڐ�]��]ڥ��N��ȝ�1	b��B��%�W��)�5�u%w�O�P��:(�]�-;�KJ׺"�Mz�?�-M�\�J�4'/��]�Bt�ϱ�����Z�O�ǋ�xG������6QI��,Th�]�n���������O��B]O�f{8��n����fk���6n��*��^�𴐭[��@�>{��H޲����2���*"U�2�:DXlxVHYEB     400     170�rK	j�Z�'V���3�
�f��6�/P.�n3#
n�W%���B�
Ľn�?+])����jv���띳F�Hi45�_;�*�VD��q ���;G�_M�y��fG�f:�\A&�~a�	6A@�u}6���r]�o,�g��2����Y��W}Uu8ΆB0N� ��ѿ�V-�g���&C�<���ٻ�۴��+n��̳a3�w+!K�Wx�vYv�Y��HS���k���99��gMp�*^���,�N��7���L�%�n�o�p�1mH�EX;����G[<�X���7T����HG�kM��ȅO�z�Z��q����Z���r���2H]�"r!s`�~,�DEr2��)"�5����)�mS�|�nX*XlxVHYEB     400     1f0cNh)�&`�P�+�\�Z:E�2��d vu�Yr'�&��N<��#�F\�񠽷q��]}��Ph9R7\�����T�D�	�uP�{#�2*�v֟�R�F5�<��Qx�����|�;�.��	���)�?���S�>�O���҅�����R����
���<�3[@!i)����u�y�ڲ����u_7U�����`7'е�Z��`f� nZ���gƕb�]'.������{�"@�����%��@��xS��-&m�%��.e�>�}pi +��K��\���m\W=�H�d�خ��ڡ�"[S�S�Rm��|��ۛl�\ՂZ��H>O4�4ɞ�r���TX����Q6qE�q�P��-��l�V���,H��8�&W���b,��E�Yh�>�5�oD��
�q簃��O�#њ�9a/�`��F�L�O���a?U��PE��NH���-}`��
y����ga#"����7D@/=m����2l��M�XlxVHYEB     400     130���u�t��4QE<V{d�ߑd�����X2�+�G߃u��Q���?��E*m���L��T�L�7� �ɍ�x�.�[�=ۀ��2���Z��M�"�"'ߩi�f�^�@N�p;�Vo�oL2�ȓ3�K��U`�km=����u�/��(kB��=�����e'�\����7ه4X=Ħ�P�����KՋ~�IKx4v��J��=g��՚�(��Y
�7��O�~%$�t�+��E��Y�����)-��k���c,q�\��f��zSX��8M!cWDK���^"۽
�zu������ߜ1��XlxVHYEB     400     190m���9�*�� |XF�V&�,ba�~Ԑ�@�u<P$�9�X�k*��
���J�]����;�*����!��om��<l	D�a,�D�����O����?,�������榆7Zr9���82b�_r�vJ.\�I���~�ga)~)2RQA��"����[��llyq٫hP���=�i>�^|u�+:�H^`p�0�t��_��V�9��T��<Nd�H�q(U�~\5���Sh��L��7*�	Ik)g�3���7���fꮎd�闇D�fe���w��h�[.�ՠW�6�#���}���r�E�E��*G�����d�.,菗��Y���-�ܔ�JK�ZLg��c'�����|����T�Ŕ�S�nA-mGS{���?;q����<XlxVHYEB     400     190���<m�sɽɦ� �T�V�C����dL@��8z��;����I
D~��
�b.�aj���r�Z�����c�kfb��͐�*�A��H.B������k����%>������y�.�2m�CZ�z�,	����2AD �7#:�}���Ժ4��a۴!4a*�pCq�8+~�^�r�Լ�R0ۉ}�m*/Ƽ�"�qF���W`9�*[Q�40��B�Lc����"鮵r�<牀��٥m��4p[��%���̌�GIo���+{*ǵ��M�f�W7�����&m!	��ԕ�5����c#�!aִѠ���NV࿒;�_G�ZR\����-�3-�D�'������{�-Ū��  Њ�S�*��;LGR�_N9p���r�Q�maX���!���"��XlxVHYEB     400     120���b
#m�g:", W�ԍ�23�����)�NnR./�����f}�܌�0}9� �|.��!;ۨ�w�xv	+�f<jXB�)Ӯ��W���T���z..��J]�!�h��3�e{t�_ȵܼ�]8]8'ݺwK�Q/=�+�Mʳp^�Z�cY#��b崘 Nj�Ct��l"�v�9�aH�X�T��=,���<s(��:�B�K�P�Ž�� ��?�����m%�(s�ڻ3W~��p���1���F�[�t�X��PF��gV2i-u;��xmĭ�gA���XlxVHYEB     400     170��n�=-��Y��
F|�'�5��k�h�j��W.�\|*aw��)5S�0���Q��-�Ѿc6�t��v��#��h�{n(_R?D��k+Q'�
h�����?�Я���&��J孺+7���69�.�R�v��[��=}Kt�W�n� ���&8�y�$߲U��5j
��jUR���ΊUQ-sQf������8���/��i&�p-oK��E����xH�+K$�Y5Sj�Ol֞ſK4j���8�ʳ;���m�Rx����{��l�beH��c�.m?�j`��S�/��,���N~�\?�(�+߼ײ��d&b�=��ӷp��Q~xAp��ܫϑS����]�C���A8W�VW����uXlxVHYEB     400     170�Ͽ�S/4���i�̞ ��|�Q���0~[�m�ڱdɥ�l��=q����t�td���]�+"W ��W\��s�'��ynJK݈���J�������e�i�y��Z���S���d9�y����]#Qb����z���o���A���t���\/g5��a��u,�h]�襞�y`kQ_�f�#�	��V����#c'���P�}�n�aɠꅄ�,Z����K����#6h�=�½�$�%9vK�Ed	��ډ����H�&�q���x��N�	>ɱ�u������#@㥏&5�6��t�fl�c�F=�J���Ȥ��7t��	gZ8�z��ˊ\wֵ�6�L3=��l��,�AXlxVHYEB     400     180�FO�ߦ:豧�U#���!���ߘ��EC��Cȴ���48�g��7��c���G�"��i3���2 rL�i]q��$���J��_P�@�Gv�Q�/kR��ǟ�D�(:�5���>4愖+��X7cF�M�K� @#!;FEwn��L�b�^��n���)-)��ɑXM����F"H�E�/���}��ݦ<��?�U� ���NQ���dnc�]�hj�ޡSc"�j�������$��ld��y<��b]{��>�h!����ND�ė�Ϲ¿���B^1�Ж��@�&�%C܅�6G{�߭t�1r��ZgV�������?/c��x�c�<����'8�T�ތOѤ������/!����^�I��uXlxVHYEB     400     100
Q�\�B��}�A��q&\U��U�'ч�d��oؗD��#�*���y�5<�М�����ug���%;����m��`2-�hN��?�j�ı����Y�9���^��XO�TY�<BOs�V����8�D�I�jY��(a�Ѭq�8�phG&W�d��؅郼�����r°s�#��sV��-g�d娭{��y��QJy�tO4�ML��d+�.P�ܜ_`W���wQ�ʜ�wx�. �5z�ch�%
#���JXlxVHYEB     400     150ն?�~�{����V����d?�M0�YX:��Ɖ�1^Vq�=~��d���+��ē�:T�|--R����f�Ј�����W�閕��ҫ��{@��_���r��kM��Z�hKh0�1�%3��e�}�@�G�^{��6j M�\�dl@�A�tA���jW�%�2��D&)Msp���&˪{N���2$T����P	T��I�I��(����n6�s>��B]��NP������`��g�D�:FZDY|�d��)�4V��k��\Z&�ސH� �%%�3���w�FR�� �LTx����!�LH��.'%xMDB�!o����X:v��(�XlxVHYEB     400     150i�Τ�ȳ������)�Z���j�Z���ϛ�:�R����>�7��(l
�ĕ�z�o���	NV�.�9fe)z�AG��Ys���}>+��ݩ�������`�s��#�@���5�RDN�tN	'�o�g�rL��E�7D�&	�N3Û$��RH��JT�Q�y})7GN����_��K������y� `7�W��5+c�����A�)Z��� �^:BBI/�V2�)-����"C&k�W.��Y���(ౣ8�v�X��� gT���-���3�,ᐟ"vtw&�|o���j�Ż�uK&��U|\0t2��ae�����s��$�;XlxVHYEB     400     150/+m��Z��E����fb�����CH��i��F�l
NZ�ⷠ�Qɗ��ù;K�g�l�ʙldȰ�a_2	�YKA�8k3�:[w�a��337�zrէ�5�	@����%ހy:=l�Qz"�$�ꆫ�G骐�c]$��qYUtbQ�#B�ݡ�۟w[C�L��s�7�!�ҪH�VE�Ixd�L�&,��f�� \ot�@bw9�J�36A�����	���.�zX���|�^��2��;搵���^����OWn��P�K;¡����A�DHC�V�����dV���,�/5B�q��A�_��\�n���wSօ�G�otvR�XlxVHYEB     400     180�P*,�Js���8�δ�!f�����Q2�jP/�5��u�{�T��"�,��Ӳz=aUd��`���j0q@@��΍Q�4�r�~�̽��C%5���H/=o)\�֌�~d��U.6���6K�����a�Z���u��,��\~5>�W?L��s˙�r�X$�-��pP�t�*�q��RՄn3N�+n�%�x�Td��cLsO��x���۠�:�y�X��"M��܏�҅j���f���>�?�/�$�B�Hr�Lh�e��0ke0 ���_�yǏ��Y3M�X��V�" ��m�o�}��\#zN�;�˵\�D��[�y�p�y�����v�$St��wQSzZT!=ϐ��@�J	����,tb�!��Wz�j<<�d�YXlxVHYEB     400     160*@��鿀"�{�,����H�J6���t|ۏ��g�`3��U��:�<��COʓr����H+#�90
�v�/|��ظ-c��(+YU��:aj����;����gr����u�B�K�Z�-����^lLKLؤ�(<���A�M�(�+��Ο!o�pE)�ѤǈF���Đ�%h0����X�Ξ����ry5�yϏ�'�)u������}�+ɢca��u~"ѻv��M�J ��+mRIm��ߟ`]�,O�?s�F��yZ�[�1����	���/�CTƚu��|-���o�SF(L��'�љ`�X��pŏ~�4yR�$��S�4��-Yv���o��ġz�W��JXlxVHYEB     400     1a0�.˱��Ü��_��IH�I��yWWR�k/���`=���0��dwO�4�� BAB��`$��xP�ޯ�:�H&j�'}}�b���Z�^����v9qT��l7z��DU�����[���A�u��_C�Mx��Q�A&q�����n?���fn	/׼��y?�[�^��7����ۉ�&x��qL�P�gT�
t{���G�c	�j�DG��릾��p-�?�1Ev��DNX����^%�ݾD"{�D��0�:�m����9_���>&�;�À;��L�.фuΦ�k7���j���<��������m�9�`�3"�Bԣ��
����7�G��H���e��>R� ��Y?��|1!WL��8@�ٙ�!�2Ӗ| U�ٛ�2��wE�k�%E��68߇��,��ƃ���k���KG!OXlxVHYEB     400     1f0��яV�!U��i����%���p1�5�-�-�xd���jL�0�������㳌ʣh��Ⱥ'%�c����(�!�����_�(� �_i�ѓ<���o� �)RS��k�i+�cR�{I����Tr�K}�t��L6b6E1a�/$0"�ݤ�$�$�kF>��dB:{�"� ,��<k�L���$����K�m�+%Z��GCyA�џ����P��?Y�pAhx�Qi�]D��(��̖��.�1Z��A��UJw'��BO�r���d��������W��0��f�q�L"̏��U�$1�K�oɫ����b�Zn��0�BϹ�C�K�(Q0 5�܉�MN��l��i2�4ԑ��?�Y���~!�:�!�.w��U�+��/;����9;�c�f�"7a����2�fް�����W���)�� �ωXl��dP�{���sF�����QB�@��h��y�1�����E�0�"<;�m����M[�!
����j�XlxVHYEB     400     140k��R��bVu�}�w|e��ypD�ny$`�;���w&C/�c��Lo����L42��N�Dn�4���֮�Pu}6x]�w}f��y�ۢ�Wd�@�����:�~4�N�ReW�c�д�J��}�t�Z��y��;%�^&�V�@�V��W��U�kt�M2og�G�%��r�x�3�����۶���E�����y�+}��)-/�\5A���\�>�qrS�k�G(X�d��~�)�cu�/�38���g�x)��m�wD�הN�r����+�������p����=8��
�EҴ�UM<1��)�n�Эӑ�k�񑞣'yx|����XlxVHYEB     400     140���~���J��]�ߔ�nB^�'h���=���*���������?�T��c�if��q-��s�s-��&�ږ[�X�"N>oTW�kV܌��Z=۰!���B.��*꘧SR�
_pM\AQ%�.�0	4�!�+��ړ���M��0/ ��X\ώ�)�5������p,M����;�(�n�X��kZcQA�F+����.QT?�-0�Ui���:�l
�#�:8>��4+u���[�����N��)�j�ԍu�����0�u�F�T�y��i�B9�c��U�{LDx[��*�_,�
��*�~�s�f}Q����XlxVHYEB     400     1e09�B��I�O�Oq2����5�8MP�G���Q$$Ĭ�|��
��,pH9:IS�Ke����R�!�`�Lxv$���~��l3دh��3�j_�G���D=O�B`@Xf8�`���W�Ei����Gӵ�}H'�#��/��Ip	fT��1VCEl��)���)ԘZT�'����Js���36���
�R�*�
�t+�[�4�Z��a�B���ͷ�)<�S�*Z8A�,-�\Py���M�8u�e��߸��F#���X��AR]���F^�6T��؁��3�(3'����$�������0B��H�?y�����$�z��P�+uF�3�Ы`��)�{L5��w���	`'P�,�(�����h�6�a��6��C�"�:V�ƞ����>���8,,-W1�H��C�Ѡ�%6iഃ�=�c>�) ���&'8�t��5�v�kV�,�y�&8���1c�3���\d�H☸;௶zy��XlxVHYEB      90      90�u�Рf4o{��g�J�|�62�P�Ɣ,��$�fqE���3S~�B U��Kt��=߾���&V|����Z��w�0�`��z��S����f�c#�֓9�ϫ,�a�8/?bs�p%k���IѪF� ~��tx�bĨ$¿