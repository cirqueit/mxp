��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���+���٦dD <��YD6�!��&�J����Z�'�9 B#?r���qt�r�򙀥�O�b���jISI #8�q3��ʖ(\;�WPi�k�����H������t�F� sG�2q�2Pĕ\D.{��2<ա��]�#��,��o�N�D�p�U��q�����ӎ�N�H+��ੑAW#	�Я���W5��RM4b�8(��O���gb��7NY;��l����bR�:^R�,+w`ZN�H�4�I��1��Z��!��7���y4�M�t
)���&05>�`���x`c�w����l(�&L� 4l=to����6� �֔��C�[ށ_3t���?��mE��j��Rm4O���he�J3hDܟ�v��	O����KN�ݯ��ڤN�Q��JCf�]?z�Jf���b)�e���s�Wo=C������ϟ�V!-fbX,mX�i�'�p��Ӣ��v?�fC#{�~��/�6��Nk�����Ix �9��Y�$7ٖE�'�j�i+��Z#PE��'P�ua����au���Ku�[	�E>H�P5z0>��#��H*��DԄ,��[2If�2QBׇ�
��z�'�	���`+V��@��ߒx
R���&���VC�5,� ��]ȫ	�!�/�"ag���V�[��SV����639�7�&*�E�hV�`2)9<o�
�n�S�6��&tR�<�SAApڅʊ}��j�H"#@ꩊ��Q:�s�
]��mKr�y�-k%�)}CYab^�n�̖L��� ���AZ�	L��n��Gu��yi&�U�Ձ�IJ�3��K$hd��~W��>����&U\�	˲'�ǳ]��ToLy���p�M0S�+-�i7����o�{ �P�����]�<6͸��ka-�Խ��������1���字���^�� ݚ��
��(��f���"�-|&^=�eKG�pU'6����T��epN=xc�}�G�߀�!�v�:6����rxi�&�U�6n�����>}��6�����?�I��Zw��ԕ���?��_,�L�yftN��dyko��Q�V��?���F��~6����Y.�o�lᅋlӭ��o'�1��B��Ü$�m^}��\�jr��ӂI;��m6�ⷉA������S��I�^��T����,��h�3��u�d�>y�x�SiA����=Is�^�Ȫ*:��vܡ�%��a���f��W+{wR�^q�?�V����Ǵ52gr�L5�0�1�Р�3��Y]�CBT���R����]/p����{���J��:7=���J���c����0�d�KP[���u��MǓ�s�8G���D���@����P���mt�]i�T��;L�>��k��y��L��f�U��5�Q_��������C�����'�i{��9�Z6L�D=kv���V�����������Sb��ٕ�M�������W���k��?<����3fjL၃ ���̢~�4-F�0C�$d�S0�5K�[��74��w��.8��>M]���TK&��X�Wb�[Jk��bi�{$+�_�UK�zL6�L�� ?�ŀ�Ь�*�$�5���&��r�M�-�KL��@�~+���R���e���g;�yϿO���� ����:F-Y�G,W8�t]� �N�8)��e2�����)Y�|��w|w�eg	�����4NF�:Q(+׉�WFk�~%?��2ύ��[9|�JI*��8��!&�n�[�-��eUjϗF-
9�����\9\yiճrU��v�!^�1�YH�<ں���Z� !~g =��~�!�z�U
���d�sdvR@��%|@Qr)4L�p��QjA��C.�����U� ~67�*hn�d�A�j�sb���S�!��G}���-+�O����-�|��g�|T팞w�j����#�c�-����n?�g���ܳ?3�3�D�&�@Aka��(�����e'��n���˨-n������h��0� ������v�F_��'�4��D)�WB� �<�x�38[tL)��3������+�x3!�p�	J�7x%�7��JЊ�fct�d�n\�g��x}��}P�
�`��S��-8��/˳���|Kr�io����N[��!QN�:ͨЏ���7J�>V�C�ĉ�[0[��1tI�Db�߯�KL'߷�4�S8�5B����
b�8(r D<���	0m{{s�(�f���&A����
f����C$rg SrS(�i=����؞�;�"�c�H�`72�HK�rؤ�{ ��B��KWg��^:hR��teɢWNi H��$�o��>r���!�
��H�o#���6P�`h��ΛdCf�' ���~�y�u��,��瑼p����7|�V�\
�,Z�J��P��%����R�.Q��݌�p�������2={���5q�F��Y�)q�z��`�~�3ikKy4�w��H,�e�E�J�2})�o����y6��,Q��i`{�aT�"��Ҥj�[h��eT���fo"���/I�\l\�o��D��+�-+VhG�ZqQ��	�B���(K%մ��P���=&Ia+��/���V4v���ǀ<8~�K<���8��RE3�W��2Ah�̌���s4&J۹��057���CH���`	���V�$e���t�Gc�5 3z���2��5�Ǌ�-�|�ң�A1
$�)<��P"�9����x��M��s~�N�^Gp�Z])�q�aR>��
�$˧��k[q*�-J\9/P�|���d�&�Q�Y]dB4��KS���}��9��e5v=��3;i&Xv�*)���bNf�}c���<��ի,q�~z���L��ʱ8G�[�ج	�UtX<2"\�p�j�ugv�w�Z�s��̂�l�a���'XjG���_�$�g�u�c���M�I�K) ˛(r���Ʌ�8J�+٫��u��q4L<��ώ���;��d��a�_A��gF6�|���I��j��'�հ=	VzO�c�R� �K�6���>`�d�S(oC�t*G��	"8@#T`����ƥQ�ѐl����6C����-���v���i�A!�� �f��&Q3䍀?����i�g���{tY#��!�QچC�5�%`�g�+��/1����tU��յţB� �����ڌ���j���ї������v�)��*�X�G��ϡ����B%�����تy�V�#�e��7{rE&P9����W�Z)S����8�d��
%v��P����mq�lٱձ76gh�]~�E8��ܴ�w��2�q%}��?�쁳YΚz�>)�sG�
����sZ<���,����5��HHN^����Ij�q�e�B�����0�g�~�}�9y��o��g==���dB'��ꮝl��I.8��"�����~)�4U�ڮ��m�	iOh�n����ZA	f]��-��6ZEkTK��+�Hc���{��`TMX�us��6��zԯ�r��S��&���_�?�Ѿ����Z_��*�^���@<HL�EUĴ�������Fh5�=�K��5ľu�b졃dY���<]$���9�pUtX&�$�d��P�I4���u>_P�0����\Sx&\̀w�I����-g�:5����,R����=�c[�g~d˃�S��i]��8�6i��ߩ�I�o�t��a�dH�Ys�<n�sb-'��"_)J�&��s�\�W��[
b�)z[t�.?+�J��Y>�`[�;��_}}U�h
� /���%�0]�޹#�R4�u���a�aB�����B@6}�#����l:���xŮ��wF3�B5�R��\J�{L�Y����ՒI����^EN�3��źS]$p'��C�,���g�	3?�Mm�+�ϴsI�G�87O�rW��G���j;I;��C��xc�gzJ���i{�c�c��v5|�0�rP�?²UY3����v��vC�H_l���'7�El���D�n���堨���L���a�A�)�¸S������� >�$ٷ:�ӾԾ��]7�e{�ڴ�R[e��b�ަ(���ؘ��KK?.k�1>4�1��&���.n.�oZ�$6�Ǫӓ�^�K��9��^Ս�75�Y}�tӼh��)��C�7��iTz����y7m�СH�$�|y(p���*�IW)5i�<��E78_|��z\�#*ɯ��f�-̶�8^�'�o����C�_s���B��̐��Ɣ��O�m6�ϵ\,��O�G�s����k�/;��4�@���Dh�}Z��/*dy	_�ǌ$�T.��?�A28�t�A�G!���PB�`��	��xV-+��_q!�D��H�/F����U߭��5H��18�e��cA4�fO=hA���z��l��^?fA�cԻ�J�T�=��:^��8�w8�Շ�"8�w"��G�ʆ_�1	h�*UvM���/�U�4��,�\	��L�@*Na���i/0�S�&��
���Wq�_�%�%����;���"_O:�4$���]�³9����+�e{�|zvg�xqT��~��o�w������J���>�����8��l���(H�D�+���(k��
]��� q����'a%��*���d���~/�KD�q#��	����k��ª҉Nl9` Qi���D�4�� �ج��`�;��M�9g��9)l�K�v� �.�U�.Z+:X��Qe��	��_O�-�& ዛ<H���������}�1��*r`�-e04��1�ݕVu#sD�_t:�N��=d�l�;l1i��Ǽ�Ǹ�#�B�����Z��������ڦ �U&pȺW�8�uj�� sZL�yi&��T=	4���Ma���R�����v��9W�v��&F�mF@��q���X�L�������ڬe�%|�Jp��9��=V�'�Ez��m�'X�4�)��н_�z_4����9���!�ţ����%�C���쓿b�D(�2��Y����u�u�'�}T����s]���a>��}6����KogHց�� �%Qiz:v2�Ǐ�/_�����=�E����;ꊤ����N�S��(v�R�[t�aeЛ���PI��hL������� $A��L���w�O3����B8o�SΛ������o���)��zzPH��~�~�D��f|F��T��Z��/?���^��屡2�d�2?G(�팯0�^c��_�l��q��]؀{,I�X��~
�pN���e�F�9h��
��k����|X���s��f8|�D�M���{��2�#x���i���#Pe|?O�s�P�3,7^�Y��B��+H��䘆��G�)֓h"�LP�
�!q���Y���~5ļ�t^ht�y}-B��2��r'
�l��cZ��.1'��.�+v��Z�c�7~�������Ζ� c0P�W5o�^��ޢ��;�|1�<�Sd;�\�bH/��8�!�*콻�
6�s�K<�4x�YQ�6�/�Z����0$�߭v��/ �Z(޻_��\�x&�J4��1��p�ic'�D��-�ҤU��ɬH��J��5�.�A�����l�H�)y�-�'$/�i+hzS���׾�Ӱ��)�J��dA"�{Ogn�q#�-i����{�>O;ԇ"�ښ����7�OE&�(��'���X	��Fƪ-�.��Ġ�+s��E�� �����	n�X�K���e�4n�pb,�T�v��޴;E�I5��/G�Hl:׶P��S��IW�݉���|��3r\��?!������ՙ����k��v��a���2K0s�Pt�?�(�D�����.��%u|0<g˗I:�]c�%��y��6�BN�����^����gr�,XDP�V�_���B�����1}@�+}�'��N"_��n�LԽ7d�YUn�Cؓ���vH
���te�7QO)���a��\D��oz$_�A5`�����4��7���q�\�Y�<�-��j�Yu؂2�%�#�����[�&	���H�D��j�I.V�g�u6�?΀�w����2F}<�{�	n}���lQ�H�7� \�y��z뷓Ԫ������T�����f�c��[��4њ�۸�@������7��%��ݒ��ٓ/�w���$菅.�@�h���<u�݋nt���F-ux�߃D��ƴ�aCF�D�����hX����/3M���U�wMg�C��o;��sR�]��m
WHA�8�|�4 2�*����/��A�q2DZ��/� �s-��[{�V����~���
�Ż�̠E�ћ��_�'8���wY������Դ����j�E!�o*9��c������bX#���'��Xs	�P?x��_
yH\ d\��pAfp����G��Bkǹ��� Saغx�vUE��=KR?-$PQ������k�=nzR_k�q��AՀ�� �|@7}���aŬ�к�&�K��qm)Rl8��ľ���͡��k�{�����W�Ѵ|��D�f:�H�-�kq��9�P��5e�����9E��� 8��A�_i)���x��j51j�>D�RW��X��!̋��X��Fp|�ȳ��-��L5Z�W�f�����;�ݏu�0��i�ղs���!I�R��,i�ݣ7r��j�����!���͑�(g�B�(��n��V�>���p����2��-bC�(���mr���o4$�;
��+��0e���ֽ�R-w��#��*h�晗-
3��B5�J����M�fk���5[�����B�	ܦL)%=��4���z�)��$]R����덶�,��k���N�F���1���9��p����Ц���|�V&|��\�aDb(��7�0����)��.��eg��`�ρ��>_"����A�jv�㫧ȕ}��0��$�������"�m����uz>X�z�V�PO�ԍ�g��p�#��|��-�.6^AkL��N��
V.����L7Z/��MP�wƢVɧ�#Tۼy�}}"|�A�ֿ��.�.��KY��\�֑������`����#�9�{m�w7Z6ֲ�4��]`��⟜�3+ǀ5r���M������DޖƠ��d�%�&2��3gU��	R{ ��,��_fj����8��.a�Or�RqV}#�%	�u�3�k%���˲×*���6��Ju�FP��C���K;(O��}тٹ���u""B���m�>�&\.H�C���-O�U�Fp.����XfN�'�H�$�z��Z߯�=�єQ��8V;h|��i�"϶��ށ�x����=.�fҳ!FC+z3|%��ܦez����;�����ɣt�c0߂q�/O�_e�lR�?v'�M]���K�؜���m��ھ-6��#O� P0M�����䙽0�JTXg���L^e������D��"����K����e�=wr.l<E�Ԃ�r�B���a��~"v{'�1�aC]��2�#vq'F�5��,�o7��p6�9@�r���nn���%<q���o�J:	��rΉ��(w�Y�ԥ2�H��H�����h���$l�"����jj�ǭ�c�#���?�X�,٤}��=vc)�6���LƱBNl�uR@A�=�p�|MT���	��fٽ�c��d��(D��1�pJH�o�i~p�>����w��/���(W8��4C��|�j��-�mc�]�y1G���it���cÇ�<�l
)}G�i��T���=�x@q�(nN�\�=�C�om0�[z�bJ��9�����\�iάZ��l��E�l@0o��o�o#/�#�0��;
��$`�;�X5����Ѥ�']��+AvBK���s݈���ƅ_lϦ�`�	�Ҏ�����S��JTgN�#�I���J���Q�v��h���(9rc�����?�o��Jfs���U"(�מ�i�i����ݷ	-���R�Lp�oI�$T�#�q��y��H�#i��������ra%�*���L8S����1}�-H
?�������2��&��v��J������!qf���sP�t���؟�Ђ["����U�ǁ��l�S@[��|�*7hy�����X��*7|�?�C/�>J�J�������[��PG>SpjVi�ی�iM��z��*�ۼ}�dJ��Ò�=\o�f�C'���r��(�ru�BQ[�(�Z�= �%�hΥ�h�Dt��=~�5�m2�A���'�{��}��
�/���Z�8.�r���v�_�e�!4�@ȥD��ֈ�l���J�}am��[o>���g��MA��n�	>cՓ.Z��ÃŎx<��(bbC��"�a4
ÞnM�Ҝ���8���LA>"�)_� )�ߦL��X\��,-��P<�.���h�Y�RbM(?�iNC��4��(mN�<�����Et�)f�9��~���,f��p5IJ\�s9���@���>E�W��9X驖C���omBk� ������_��Jo�ʾ[e��{���	�h7Vm ��iCQ�� ��'~��>R�7umC*D9�}-D!!��;�[z�c(�%����2����Ѡ�.s��j��%�`������'x»�0;�{r��v��n�����*U!dV�7�b�?bR�Em��U+�*�3-�;��V2d�[��aS.>ͽM�qZ�\VhP�1���sesh=b]
.&�5B�#�����Z9�@t��c��ǭ`��c�*Y�{���){w�+6Z��	���V��5F��g������4$�(ty[,=������Y!�U�pv�4�J�9�cg�䧬%�hQD���Ç�[��Ŵ}k׆��X�o�H��-	6�=��%�� 	�h'��=+�{�"g
�0?�Ӕ��f%�e3��iO�`���@sm;�8Q�~��m1�����@Ȝl������g�>��V�3Lq�������9��S�f����b��0�\� �=yq�izt�AKO���m��zm�Rg��ϧ���}�o�A��z�2no��
2��G� :Go��4$c��h��(jVa[�?��W�8&PB�TC�K'��d�g)��ƺ�>5��In�?����=%�U�������U�OD��"/C��N����ͤ�&M/����p+��H�4�D��@�C�I����H;�'w�Lpjy��E
��\�&��s��k��ʓ����L?-�i���wb�L�0[끦@�Q~�@�)�x��)�G�$������H������([�G[��x2×8�
����9����J�R�af�1|��\�=�#�Ip��_�����b�V3��O����>E)ߖ@�����
zǕF� �� K��7�I��ikTʉ�����6Y������fE9�1(?<Z��+T\u����Kz�8o"˺@{e�E۰ǁ������ڈ�QѢ>YW�I$	]n�|��T�V��kS����z\]V����������Rե~Q�ջ��5�MO�DC�Q��%[��*3�(�Rl��CTc���*�#���������m�C��zty�d;As/�����e3��V�芽ΙpoE8Q�DF����d��/@mm/���,�0����/G����y�\��bݺ21L������u
��N�U[�	}ﮠ;7�+�������둒�
_�Ͼu�\��Y*r>;$j�����]Z�bAザ4�&���UE>���.���W����i6A�����vu��;�;j�/�cS�Y��Gk <�	k��M�����YH���Õ�0�x-Ʈbȡm�|��h���j���b���^��E��G1m�w����͔�NR�Ou�kݧ�;ޙ��t	�J��\y��-���w��wee�^��FFH����K������˼�}��t�!�.U��^n:q�-\V��FՏ����lmS����#H��󟻮I۝��$ڛ���9o{O�I�i%�����,	e�x��̃e�
]�+��	�ni����+f)�m�����S����(aIR����{gMY�U^3_�*tR��/�}����i��I��Г��n���
+а���V�(RX�w����4��>%�Ѧt'��k kB��rw�ޘ�]��L� &<��Z�[�7;����V���x��O���I�`����K�ts^���?�O=���Ţ�Z"%w�T�UѼ{���,�j`�_02=�S�*��Qߗe���Ѓ.*���+����y�ؾ�c�w��^i�g�iCHo8���{�&��{�(���E��[�����������VL���(+��(�b��NY}�!\H8�#�8}5�i��e)%���&��>硜	r�rIZ�O���zƖ:������^�dȔ_�]L�O��I�mr�(O������p�c�`g*Q	��`&r�YB��oA8�+o1X-�P�Oh����?LLJ�z���;8c�<sb`0i?k��uU���f�^�4ez�4�X��Hː_l��.FW�ڟ�������2�,}h_��23���1�7�S�͂ұ����#�R�~ o�������r���Ё
�á�ɰa�� �c��
b�z�[�|,�<ѕ��VƵ5A{�3I��&�Z�����&p��B@G�>�_Sr���yշ}�,oЇ��/�fπ�c�[�h��8i7k	��k�f�dȐ�N��|w�`T����?��J���_���~A���Jo���[a�q
�4W_��z�N*�~�?O�K���(^2�ON[�5��U���_nf�+��jx1��'�Z~j�!�
D��0���\�K�C�3��\��OP�-��NXl�=Qם�)Za1N2�}�o;G���X��<�(س�P/J����lQR{�)3�'
,�iS����F{m�9�_8Ete�W� 4�~�D.�sYT�y�¿��gߙ��ި���LՓl�m��	Y6y#�N�˲�7�]�����iD$9@��i�xZ炶ڰ֑��'��źd����7�����f��d*2���Hh��i�$�����(�l���s`���V�@�vlU�S�Kd��ď'o�0�ǩ��ܨ8^H�3V��ѾDH�����՛*�A�6�Y���Ӡ���� �l�Us�1^��	Ac��ZX�i�T�>M��:U �;X�S�ًV�il�i�ʀ����u�����ݣ���,��m�QǦ�R!����:�
��y�qj!���w��
q�I����۬�sZ(�r�2��/=��4�FN^J'	�Z��z��$f[��FL��[�h�ń�G\��:WGT��i>i�EK�@����9Y7�3�'EK�'�S��6����b'�0�Xq����LJ���z<=q��}�6������zmmO.��ʎ��cj]�I��V۶�,�IO0�`@��m�e��ޗ���=�v:�t�^ֈ�_�\�UqӼ�+G"�W�>ՙ����TT��5�2�*����y"�L��\�E�uY��d��#�k����g�����A�o�
�y�M�~*�z�yY��	Vʲ>�?���Q�W1�p�nQ�[�O��o��J��4(b��x����O�9��^DH�� ����]��v�}b:�6nf＞w��6�U�-�Ͳz-sI�ϤX���zZ ,�KY�ڄ%t4p�(��#�ޕq!���R�Z䭒���@�[p�yķ,8;L��"-��x,�^8+�G���j������Dr��*>�;�
Vo:�7���>s圥��� �X���O��;	X�mM��0#>Dǅ��6�����VC_�(�K�hzx}%��N�hL�$)ի�	��ۓ�{5���U�?N����,�"�)\�OMMi�fc�#|u�\g�QiՏ�c��.�����(U�l��R��a@6������],�x�P��`�����$?�yW�����.DP2Fi�O]�δڙ���$�#36� "��ǎ���?.,O� ��H ���q�vI�ZJ&�H��D?ԞV�*_�/�d
��,�wb*
f�� ���27�{�e�h�����;���y?B�D
�<S{��u\�����M��~c�������L���.Pl%�>�n��bPU�o5n����ɛz�x�J!)#���!P���]�D$CgZL��8pK<+
+��O���o�k �S����\R�H!��e �|J�8�oK�@q��}�?6�-���vv���_R��ʩHp���%��P��H���jA(Y�1Z��쇵"[ӎS<,EЙ"]O�]J�"���E��H�?,�LI�a��P-������5���vb����}G�2,��U���˼�//6M}J��|�vL�L
�8��/Vod5'lpBv^H.�@��P��X0��-����c������J����3m�����(���l��R��0��-����tJ������1a�����R�7kzV/�1��\�d�*^�u��z���~�!8�����p0s������h�'���,̉�#i��
�C<���cA˟0+~S�`(���8��'\��Cs16`ɴ�aW����S<��.F�IU���\|�&��5�*�~��^��(��� 2q�f2�@
���ޅ��×ؿ��e�"�U*��߻ʉr��\�>�'�H�Ń��������6��� ��P_�3-�+D�Og�sߩ���q
7�8ы6�����bu �oZ��S�(_P�є:m��{��Fh%?yc%���9X}o�🣍S���a'��PS^tH��ԱoL���@ج����j��w.IۋD_j�A��T	5��!�N3�͖�����.��mO�:q�,23�C��Q�ĔE����������d�eu�n��@Mu�_*�c���cM۲���\(�T�Z�ξ��J$bS�,��� /q�:��Q�ާ>*���FFZ��@k������J�7���S`�+�5��qW!;�+��/wb���E���q�v��tXX�ӱA>t7l|�oGF���b �P�B�1:��nFe��ӥ��dZ����N1�с�8�_�@���v�.�HT�ш`��e�E���A�d�,WI.TUͰ����Tⷡ4F|#���)2g��Kw/�Jk��t@��f�}���"�u���@�^Czª_����8e��z<0�l�x�D�w[5��(�e$�A�4��8�%��ꏪ�mC_��Y���q�R�D ���i;E���.��.���b��V�v���ՋTϯ/��]�HR��m�C��z*�g�-]���&���Bd�X��c?�B�}$I��Rt��(6�����{�8]���^ٝ�G:�ݹ��	��i�Y� D��G',bw0Q��(׈���R:�׳���CǙ��D�>-�$�*���BU���9��1���+��q�#-q2�ʺ>_��������L�,kY� 2��&d�D����^~�CC��/�O��2��T�4�Fl���9}��Y�3���(�˱$�6�+�j��?�-�P��O����0�p��/�mY�B��s�A�+4���,�����ǻ5���]����<b@�~O\C��a�ߜ� ��qh�R5���J�T��4����1"���3�m��B㯁�"\��֚�
?� U��i�t-�%�Z�>�^6��Z0i�SP��d���f�����g����V�N� KV|��31!�6��o,�:��~������P!�w8�Ah��3[���n�=LeU}ꭖ�9&'���j����ǘ�̈́�0�Ɯz��`r��|��J�ޮ!+�ad���f�@A[�^�Ic>i�����g
6[�I]��Ѡ��`�6��z?Ǡ����b�jI�3��^*�|�]i�^xI�*������b�e��ke�V�y�nq�K"�L��,���U�< -�%׆�Y��#�"cFԃ*!Dz�PnN����q�g�;l,Ʒ-���N2C5Ú2���o��;�ڍ��G�����mW��i)i�^�S�>=<�&�0�ܪFr58rɲ�H�!��\�>n��m�p�i�D���5V���2|M?d�W`����_#f3;�}Ty��>g��Ԟ�)�� 9��w�g�V<F��6�P���O�w�!?�<��t����M��I����t��7��s�պ�A�녶��jq�Rn�B9��-��.��@'Σ���2C��{�%�벎}�kP���1��q��̤2-��w�i�y�D�.��Q:�-4%7�0,�ȆoZL�4�S+�Z��P7�.y.O9Fei0y�o#���5�����*��v�J�]9�R�<�i:�	�I
��R�$�){^�GK������ɪ��yi�TζR�*�:���%�H�u�wrGf)*��\�?��m?�N}U�z��\��k��T��'>ʻb�+�^/�����e���:��y�
З�������v"�LOx���4�������J�~������/��R	v1c����؉�Ѹ/%�[��r��*�3H��xԨ�͏c�G%I�K����s'=�iv��y/��,��g4*	~��A�"I�=`Z�`&e��?�����i��=s�b,���=j���\>TUUC�p��+��՛\���`"��Z�	.���tZ�� G�))�`8�M)��t�����y|קQ���3z�I�"�V�����_���ȳ#�-ļ����ˈ�pB,�=�g�"A4��/&IIl�lq#� ��@`��	�s���S]rF�5H�Y�XoIG@�w���_�h��MXi���;[�q��κ���XkE�o4×�E?,��;Z(y{��̍m���ts�N����z'�B�ڨ������vҏ>�%%nSbws�p�~}�`L�w!6}��'��z�X�i�Z�(���)�����0d�| �\fF��&�(Ct2�3[��5�Ux7�<y�,����|M�}��	[?cހ����i�T�;��-:΢�ۧ�h<|\�ߐ�ioP��^ӄ�S����KZ1D0tdZL��ڕ�ru�:K�b�3%�-�Z�����8o�}��3��y�����6eN*� ���b�l��Y�����b^9���~S��Q$� P��t�CA�u� 'a1g�A�{���LK�b��>������a�ml�~�ؤ� j%lK��ں�]�?��(.�9���_�Gf&%�|��#D�L>	ߏ����[�a�AW�6�G3E�52�:��Ȩ�z�88m�^��"Η�n�H]M.4���"�6_�N n 9���U���O�sQx`��d�xQ7��+)�ƕv���.)����ٕ�I��%E,�m����`!�7�SU�4�hS��BL��g�p�P^kX�ާ}-3�Ǹ��Ҟ��y��`��4�	��)�Q�焸渡�%�]竑�s@�(%��F+�;,Ty�c-�ǚz�h��z�U��W�A��N���!��v��%�4`)�+� V�:�A�/�E�+��v�����l-�uj���Z��g��nh��H�j�MU�T�|������)a()�XA{�d�P
(���u� ^,@ (|RІBՌ՜*�h�I0��ٻ��	(�7�$( �^F���\�X��m��n�+��7K��ɇ	����6�͒q8�;M5�������Գ*}o&�AA��t�Q�eRLV;н����BT]�'�-�I��kI,�״�1�����!;̟���|�o��%�\���j�$�G�D]�r4�KM��`��I���$G��Sx��f�mښ�?6�ݔԐn~�Q�.̑�E�#��r��	���S��Á����J�N_��*��u����_�)~2|wW�֩�'�kd1;4"u�-�^ߵ�A�]�yFj�5���Qu�GԆ�0ġ�?��pG��C�D��em�{r��6��kXM5E�,��w�R�r�Z�ì��1�1l*�ںV�k̡͢�zba"@���h-kS�w�+=G \8�#�B<aZ}�͓ձb6$r��Kx��?�q�A�c�0�9�޶;_���<�2�}m��MҾ*d�8�����^:����L��f%;����ɢI�v_|�'��(�dl5�%�?�n��W(zN�,:�e>�L�	!؏����m�]�B+y�j�\���ϒ&D�s�Lo� �
�>d}g�FX8�6D�����F����z�٢h�K��'9"���WV�3�Z��lEOm]�u�̀���B=�i��Q�~�qO� ��R���Emx}0�m�p�f����q�6���C4;q�Pbv����ޥ�u�\i&n$��'8�h7��2;vbM[��!Vbb~4�C�=\������Qeo1p`m�]��%?b�J�z�J�[����`�ks;��r
�q��w��&��8��^Sf蜻L�@C���G�t�qL �
��]�y��k�7K�ğIK��z�,��ܽ�e篑do�[�_RJ�Ϻ0��A=.�-�����7ϕW��bi���,Jkr�!�v2f�FV"��X2+�y�ĉ�@�'��"�K���S��AV�4d�m����b'���_�)�u�8��ۓ!� ��W����M i�Ǣ�X�Q��5���=�gW���0{�\U!<���x�5��2E�G�_H������w�b˨�I�8~��ڂ�S��U���M_��Y�L��0`�C�9��^cY+�s:7Ի{sw8b0�'E��8"�9]���m��Z{\泩�O����3�(��������~��}%�L$�ܸ�\�֭����N6k�Z���'��#��9��N*�xI(�Ij�7�b�8I#%��b�����8�ؓ���%?
�l�(�L��(�	���t+��]9�mT{��U_5����O���1徴�b����^P�W�N��Paջ	'�9ɐY|a/��@K�ʎ��\�38�B�S nE�x�!-��BBe�L6��m��F,W;Z׶¬�h��1� ]˃�������}
��L1fE�$�i�u��z��2*���0�>|��������:��K4���"������9M�mM&@���HN�W�+���S�J�i��
z��H4�?Ŏj�6���Mz<t�A�3���V���9�d��1$W�4H�	�1�~,���V�L	��{��&rGE�9/0�%J����X��.���^�W����5�9�"P�5�}>rE�I�z�w7�Z�ŕ����]tSˁ�f�9ǖ�48�����{��'&W�{�I��_o[O�׸w�yj���z~c�˲`���&���P�y��Y\2��, ��C��䭾~��}\G���ȱ�(`���t�6�lȠu�|���@&3g�D�z"5��7��<�\dCI�<�*3�n��on�Z�)�\V
��`��Pb���,?|^v��4���$_���+l�{:�����	� ���
b�[���wP��|m��ۈɟ��1q�NnS>6;�)�Վ4(a�(����6ȣ�3����S.n
gF�!_�+�K|6db-�,s�H&����/3OL�s��E�P8�|��UBg��P9,+����i�q
hG����g�/�n�AU�LAB"��Ǐ�:DX����%���qjcU#���>u �̾|��	D��@'���+��w�h�i��Ax���X�����,�h�m*��t�ٿ]�<V����u�����񋲛��t��R�ˮ7tѦإ��L�N���	�X�2)?�b�ā�|�A%r�?�`ʞ��r"'�#a��dk��GB����_�\N_?]n�(ٕ0|��D�{$���(=(=�G��c�1�Seխ� ����9,\gR��d����)�/1����ҽ�(��2a�I[�M����͞(|�Y���Z^���\�&j�4��F�Ŋ~@@�n���\��M�D�泒���Թ��4LJ�$���o�����<O&W7���K�X+3xdТw6p1=z��Y����p���������;B�\�i}3�).��7�F��:r���Eі��K�5��bE�Q� ���ΪG!aK4<"6��bq ����c���zϡޑ��#���[�<�Գ��Tp.׵�&[��/9o��h�MLC��J��'�2��������h]��v��񣳊�c�(7x\���#�4n�ըV�l�FA��w����a˥z�aWA��	��{D�KJ�-S�`p�5�;)Y�[,d� i�W(�sa'��۷E�_�ӆ��`-�E7�_�$�78�z�wY[zZ�����l{�O��8z�{�'�a�QM���eD�S���<Azmb��| g;�r���Mb��7	���Y���YS@pk��j�%9Pe���s��d
�܌��Lq�q(�����Y�ʮ��zb�d�3O^���6 3M�"4�<�jJ�#B�nѐ�t��;Z�|v��-!\�|_�X�T�!���`���w6'����s����%P�M@�5�6��,V��:��uS�K��T��������*?ꤱ�B�d�Bf�,x�-�
� 
��]<��dl�Uל�������`�p���xk�݇�*{HNug*���-�HG�R����"+��:��h�����u.��4&�+W���.�t�gI�H�s��!m*6�a�)|�?`�ѕ̈́9QWv�_>@H˧��m*�)�^]�zֺ�����Wg�1�W�G�*���&Ϝ��]i��5Tm+{,	��8���1,�0��t����wm����\X� ��$��Mȏ-v'0t���w�t��)�!<9��������,��R�G�Ά=�²�DP�E�wV0��,�:�7��_�J}���Ǧ�(jhB?�&��=dR.�	�{8zC��5B�j�&�)��w�F���}���~�z
W6�H��U�R8O��Ɩ&�_:8�0F�,�[~��>-ڍ�E��G�)�-ܳeP,��s���+3�'��0�]���y�C��]��wV8���|n(Nwf[$�5�X��Ibq�3m�����L�(8�k�#a����ޞt�؛⌡�C�Kҵ4Q(�#��cR�d6s�L/&����,~��^Z�<�1t�d�2�;+G2�8[K�0Î�i�z[��o��h
�&m&�'fq �9��cN�����e��d��ݰ�OF����g��lt�a8�@+�n��Q�(	�)x�N2�lU���87D�t���7��n.<�bG�/6��"ҕF'�s�>�ls����IU�z�=$�v���6Z���XȰ|rA�L<�,�\ڱ,�$�xْ��~�i�ϡ�~�P�bh�ݑ�� c����%��eI�����lg5�?C����}��m�����,
QǊ߻W�R��'�@����\��Ox;�i�0]#�hx�'PQ�I(dXs�����8�b=���19d$��6�f �fv�������G�Z6Y]A���躦4!KrW%DyM	:���6%��n�0|��|�:�pu���Ǝh���Ȫg���3v�%�tA{b	ԓ�c�{��\0/�ų�>�)7�q�
�Z���.)N׺�e>(�<�k�`͂��q��-~�Ƹ�N-�K:�l��p0��֢͙NQy���j��Ց�Q�0�x�o��i-cy\��tqzݜ d��YO�3EZAlc�e:���g�}��Z:�\�R��&*xR�b��S�o4��n��l!��A�l�"�ת��%Lթ6�eD�&s�0a��>W�$Mc?=�p�Z�=��U��.Ia;�	�Y-����3����pM�Mژ�c� �L�6o�cVD3s���ZшAFPB�X`�-H�zy�$�\~Ԏyh�������1�7Wa?a��-���~�^:�����	pOd�g��*q,2�d���x�D�H�Z����y-.��(�P�O��Y^�!�jA���ww|[F�ê�
�,�`�sꆢ4�}�n����I�Ud��O���-��.����E�)�ޞ�O�h�/o���vN�D�8� U��D5��p�.&#��M�`^����Fk�DF��2n2��SX�ld� PVG��6�o9���`��+� ����X��MħJ$�Z�M�[EI�%�����gC�{���,�y��~��H�;�����9���=�v�6�a
k�LhO
��O�:�~y������gʗ9.ip���.�R��x��G�J�G[j}���<��L���*�eY����
{ܱw��x�e�e�][��'d�T�ި��>�c-�T���d�W�04 \�N=�#��R~ȳ�y����a�����&n��Ml��;I;����F.�����X�R��r�(!]ksy�Y]��k\�p��iRaU}���ÕEw��G�)n*6���wHÑ��O�Wݫeu[��zC�b����:���5���V�A�^R�Cɩ"�O�fْǰG�l��_�@6���S�r��v4��.�s^ΐE���o��]�1.fwQO(#
�Rx$ �ڭ�s ^�*%a7ȇ�	)-3O-�dr�9�T�J�"�,�2���`k����������W�\���ߍt?���(��k�KB�f�Ը�'�HbV�{=.ځ�=�sᰪ {ɯ7�[y��7���5L�S�m	�@����N��R�R{��{-����g�$�S�^����
^�%�m;��SS�^���a�������Sa���<je��osp�! �CٴB�ч��N�˺����J$���Ab��FsL���&Z�D����E̤;+�e#�ح�����k���F�^*<#�2U��_���c`/�^���O�G����lp��W_��`�r�vӖ�j�'W�0�eI&6][^%%ܕ�Ru�?��Q8<-0>䦸�Ҿ��+	 �;'�.��oJH���8��ΐٚ<����=rDn�a��S�Ql˙ ��!�=�$S FZ�T�����֩]�q��n*4��V�o������3����,�#�������h��i|�c���y"�6pO��R��4��l�>l���� Gj���-=�9w!7�S�gK�>�b�u�d�p������V����k��?6�.�I��#�䶗� 6����z�Һ/["�Z�i7%Cz<^��D_�Tנ���P+fm���X�b�ɬ��\����4~"�<yV�Ӂ�{��� M��8������ԊO?E�� %ؘA4˲T��R��$]}�w�̆�H���{%yO��|~F҇�k��CS1���Z�Bi�)Mk�D��Ő��� Cq���b���YO�ǿ~������w⶷[�B�\'h�0Q���gR�ηsnl���P?��t�+]���ی���%�=����*f�����䗂��KB����:��[�~���S��������r�60F$��B+h�	PkIl�V�2"�f/&�:�z5'��Л��;�
�*��L�V������	�����1��,�K��es茧�܅�o6PC�'�6zQ&�F�@̏pϽ�%�L	���(ڞ���I�ꎎJ@ʕk_�M7��0�U�23�>�ڤ#}�{-��g�d��j��_]
�!bG���K���3��� pkx(�s2�u�qirT$��;S(���a����Ux�q
��l�������ĵ~�,���O�o��u�/�9 2��T���1�!&��+<����$���.���j�>���S\wm�8@9RW���V���̱{��9���>A�.Ց�BC0=!�H����U��ŠX�-�ƀF�q޳|�~9�[����Do�֭�}m����ҥ,)������͕�3��ې�r
�7��d�2Ir\@��)��'�]9��.��!��5�p�,��o�r���{;��s(���o�OQ��� 7,�"���	��y������6t����N�.t��@�A�+�9�3�l�Ƈ���v7t,/+D���(����87x.cc��ʣa�.��J�Ь��=4_�D:wk�[��e�a���t: J��j�;�/+�9e���W�Zz�;/���Q�kH�wr7 F%I�7L��j��_������ 貴��-8�g���}`��'�uۍ.y���a7�M�>�AC�u����lZ
�P�$�	Ĝw��6?8�!j�5N�9��6}'�󓚩;u`��4T�37�y�����l-�ͷ���\��d%��8�3�|������D��E<�T�M����1`��}k�`p��E�_[�H�,H@q��y���	�!�1<�%��Z�{ηb��R��Xv�A���$�]�h>
���q�_7�rt���3���h���2�涌W�(�TѮU���=��myjk�ǚ�6�Jq�U�x׊
��� :��1�bؙ=�6�#�}:�r�9��	��=�k*��W��*��j�EG�	���S8y)Dt���Qm����n��sxD#�=߷X=�s!�@2��뱽C���r�K��p`�̱h��w��D����v��f=�
���J`˙`܅�)�"7�ЃK�c������K��,âWx�'B�x��{�T����O%�
I	Hg��g��	��6� �1�p�W0q��4�����M����]�h��Q�"FDZ~�@���ȹ,�H4|S�A[��'5`�\���'��< ��d�5�'�G����홏�ӌ,0��$ފ��h_p���<Z��N*�ޜp3{@gz)0i����'�*�J��QՉ�S��T�^�k��ù(���>����''عLש{E�<�
IX,VNS�r=�p:����^o>�G��
�(�k�Xv*��#�~[�/H�����ݍ�Q^t�C}]�P;�K�#=�4W��sr�#�6�ƨ
�SǮ�
Q�[!��?�2"��!	l%OGr��
a%}i��6�񀝟){0ik�,�	��PѽSk�\1�3�Q�d�T�HU-�+���0�����u�ER�"�G��Kcى (�"��[ƂN!�6���[�(�'L����J,��~Վ�+ã�H��_�#���22���xg�x����jp.6��Í-L��O��Y
����bE����&L� L�F�r���H!�Q�{�=ܽ�x���k{;�T8�Y���m�����E�n�G&�:��U��-���<�uR[2r���  6>��1v������#5�nwo��9&�%Qݑ�9���g�����l��УqC۫�����WA�p��܀�{��I��(��z0��3�Z;��������7�6{������ԅb���ATeϓ3�sX1�!&ɻ=M�DK37���%�i�������8ڟ�I����)�ڇ��/|[�HI(zP��Mu�"j6rs�@Ғ{�[�F��q��d؆�dR�'槿06N71 �E�x/7ݺ� �8L�/��(��W��V�%��ܚ����M I�#3��w���`<�L�r�ŭ�	�!	��9N�^O�Ӎ������o�X��>���)b���ˁOD���U̬��P|S�����]�	��D>�]F�Z�$G ��c5p�nt��!�qܤ���"���������a�0�����c�PDP�[m�Q>�Z��8R�ҕ˘�9��m�����:����#t�]�gUp��7�{�#Ƕ�N���M��� �Dw�^��o����@�uߪ�����1GR!�8���i/������(�ʓ�ŝg���ڸ�^��i,F=�"����j����-�
�33H��Y��s碕��o���xw�f2���hr1�(�0GUn���b$w�NM�͌V�xȚ����/��>$*���� c8�[��a"	�#6��ϲH���	��
!�ypM,��(fْ���5����~��� ���5�
���I��V!�	��za�����!�-48TF W"��.����t<r��}U�����(u�n���'Aݙ�3k�%��?��������U�f�ȉ�Wt�dvd��BO�-��by<�!94:Z����n�f�^&�-�!�.G��T����]��v� v������PP�̦��T�j��s��S�g���9�"�8X�⌟,'�W��I:�	="@G��o�P~�
:�F��!�p6��ՙ-��` N�!��%H6p��G��˘v�\��S��b��W�s��ADz��Do�#�lrI�(ZnP.Йlڃz����!�#�bW+��3��T���.8�BT�d�'��Mqa��;�����QG_���˙h@^$�$�����o�Z��^�"]�LO��Z���&ɋX3�8��#��{��,+���̒�<��s��f ^�k
I\��X�l���K�ɰ�k�$G�6�o
��de�LL��4&,0	�l�P�`��~�S�khh{� �M�BE÷Db��D�?<�%��ez�/]nNݙT���9ʅ�]w_p���b,k*��(�8�}���nkM��� __���R�2a&��GN�Ù`��N��|��)���7�F�Ivg��g��Qe%���� �Ϻ����3�S�؞0Q����+w<�Efk�ϗ��.6�뽪����E8:��:�����P{v���k��7��GS�{�#�eՊk��R����T�:�7�U�9����V�~�/�����zS z�gR.�s�=`X��G�X�����փ���4*{����h �䦄Y)��馄Y���R���OA����By��(c����]"�1Y"��\:3W�ԔE��綮�[[X �G>]�s�LI�_?/�q`��]쉠�:�xi��\��,�d�>�p��D��ja�G�F�ϼ�w�����I������]d0C\[ǡ�-ش�e2�����Y�d��r����H%���˲-$�c����Q[�^�1ե�D�q�ф5xD~ӠZI����	�q
�Tn���f�zk�����Ze��x�g�%Y���$��
�p�md�ZO'+���"���YK����?��I�f�:��
<�ה@&��wK�#�i��j����ݣ�%�"�I���r2���S�.*�Ճ��[}/��	��ў��>L��x������j� �8G�p,!�1c��kH.�[skW�e�O9�R#���9���Ra�$<��.� �b����MS�Xv>i>ۢo5&q�9��� n���jx�*�o�%����>��w���J^�b����%���25�_�R@�KC�i%1�Qj��lA����1*1�����)�z{��!��O���=��'�Ӈ�1!Y�o�wYo3�\|K�Ƨjb_.��\�!�T�T�W"u�/�>�`��v��<��
ey�����*�7���7����E��!RN�y*S��fj9��Yf�b����,�؂ )�7q������*^�h(qGq�]HŻ���Px��?l2����މ�r�r���h���O��o�F��W�ӱs$�-����8x�d� �/��t<1���]D\^1�0&�ʐŷiI�à��p]���8�H��L����C�9V~�S���l��ۄ�
�?��`Jx%Kl��_q!��pU�#��u�*L���ץ�L	����0eJO����Ɔh� �oY��ñ����	�Yɞ��FpH�;��)�Ft�[]94�*�/=FpO���7	������>g}�c�-W�g|�nä��q�Ug�o�o��E�3<ʻ�-����N$t�ߓv(��=���橬1y^�����[�������O�� ��=EG����!�lKs�2-���i����jtKrڠgnŶ��Sxڜ��zzB��'�ę$�[u_��A����2�d�[�hG����Y��rΝ��T�-�b���Ȣ4�6==V��;�1��Y?ֳQ���Ez�`̍�R�W�O��7��Wߣ�L����X�[��Bl��|��)�K�[���#��j��}^�С�-	'����m�k�����w��ND�=<o0Z�B���m9���B��Й��x��Y��$��֧�):-���(���UE|�q\�D.�]PC�\�&��@��A���5�����æc����	}�d���k�z�,�F����h"F���w���~]%��1;��p$���(�Р4�D���QdA��{G�k4[�&%אcs���T�/\�$����&��yg�8����g��\����)%�U�T�����N-���Ȑ`��OJ�lC�n�Xjp�^���$O��rD6���FuA�Y��੥����T�'".�yl�>��	{5]M�K�5�B�[���߂�k�?݊��]x�]��TEL�s�w���M	�L��)ڮ�9#Y�V�vB1��9�q]�6"����Һ�5�OG������)x�����4YM��%	[(��/{`�BzJ���������G.N�+QK#�'���D�
,��A+[�]QN����W7jJ�\B�����d�󠤡\�i$!���g�q�P�k���Y�{�ZFch��X�K�J�E%6$�����,��-��g����ߙ����o�d�Cu�Iw��v�$��ۃ�5s"�j����[��l9��j��rS|��j�?V8�MC� �Q�\]rDVRC�BN��q���苑sb��}�+�}���;g����Z�����-W8j���V�_0
;�aZ>���w^�t}D��"-ӑ�9����DV�Q�M�"!ԨLi�����{z�y ��7�Pu`Q��6W��ސ�D_���!�lKnlI�~���Nޕd��n����Yʪ�N� j�%�2�x���jW�%�U��x�k;^�t��0��,jknp|�NdߌZ��+�֗'�&#IuJ��~ǅ�"�é������4�Z�'��i9-�ag��uX'�k�9��#��i �ซ�	H��u���T,��]����7�*�fT�z�t]�F��p҉���=zjQǱ�����FD]T�M�a.�C�3:?a9�����{�Gt3�+���(��ɡxLYu�ƺ���O�`�	��,q��`H���h�?s�s�`����S�0��n�W踹�}8v+ߧ��h,�m@t������,�M��;�4����v��K�S�=ԉ�TC��v!-[�����D�˿�`wI�V@�b>#�i� ���=!��q"O�I�3��;�ԅ .�KCc��xU/qGp�\VG1T[��b"�6�a��ݡ�.Ymj�����ڡc|ҊQ��(�n�=4z�B?��sktt�9h%�i�Ħ���9���5Y ŏs˛5��MA}���F�� �%�kC����0�����COC��vm S� �L�"�U�����.y�St7�H�T�7*<G�Կ�~��9��Q��8.˳�8y�>���p�psz6n]u����Z{q�X?B!el-�'w'�n�,=��bT�������$�y6��j%�}ɇ�r���z�cR���Z�.ԑx���廯"��5������7$����
x$7����A�
�����1+CT]�W>p�{��Q������s]+}����mM�U�ov�>݇����&5(OYˌ���%���rI��-OX��m�Xr�1�G2X ��+m R��J_�
���(�Uw������Cʾ���h��K�.p5]��YV�+�l Izkݬ�6���/����T��__><����vK䊊�ڔI`�	X��LUw�rb��4fQu8F�I�%���|�(o�'� ��=�uh�dF�HKr��� ӿ����_�(ФӉE�Ewj���O�9G���"�'y����$�#B�^&x�9U>�����D�f����-������ZF~;Z��9�!~n�.�6q�GR��ҡ&��]�ϑ��9\Fq��	���H5���6�7�}�q�3,E<�u#��~�{�`����"Y����ۨ��D���N7ǉ�#���~G���SN-�g4�P���D��Qy�~D+�R4L��ad?FaJ"H[��b҈����]�b���B���ݎ�p�@l>�Vc}2��\���6[����+�Ge��K(����7),�|aR�kJ��."����ZD�9��Z�ln�W1R�0f�P� �W��<`:MF-�Ҵ5�(��ܻ�r��*$J��xQ㖾(�t�-m�P%�2!����1_TH�prUM��(^>��)
���§�V�Nmb�?@PO�.�CV�s�x�����(�k���%��D#8�	���F�*�X�QЪ�@q=��4��ьz+�k�'I����*f�Aۃ�"8��h��,�y�/t:T��;�X̢B���\}�Mj#�-�cb�MԤ@��t�!,  �>�]B�s��(u������r��Ygcʶ�@>2�&� QԮ�󮋀q1p��\1��9P���N���O1�l���՜xo��Ϝ�S����5x{��4q� X׬.����6�1i���Ja��Nd#�2�aM�X�������}������t3I��Jo�wGE�yQ����1[�ᵵ̈V+�G%�!��T�y���~�ji?�����|�!e��@z�] ~�'I��n�����6Xx)ʼלjqo�ůJ��b�j,W����ۦ�)}�����2z;n`�哧Y>`R�*�<W�j��6�z!���y���[\g�oD-}@��s���
��5bH+��Y0^��5��X����Tȍ������L�'d�Z�����tΚ_�O�]��&�m�S���+G4�U��K۟3���6H���9eX���k,8�}(����M$&d����*,X�.ðҔ��nT3����=A�#�������t�Cc��N�;�9�N�Ǆ�ٯ�W��� /��j}��*��F�h�5%|/��25l�QO6f8�9p� ����d��=�s��6��>=�§>[$���e)����nC��ؓ����lsI��/�s�v�7���7�����S뻅F�V�D��f����hp ��=�2XK(u�m8ڭ��hSVH���_�(�m�&�*�a"��a[ژ����&�C�{\fϦL�>�o�ۉ�w�Lr��+嫧J���r���慒{zR_c�3Q�p�>����Xv�b���O�C�������t�m����)�[I��cb
����wtN����hJ<�<hA<�u)���3�;�<�U(�V��+���H	�o.��)����w\�G�#ӵc�5�*�`цґ���N�{���Y|�U�,D�\� �?�H�ՐC&AX��k�.{,W��X�T`����_�hH/��2�DE/��3�jB7�`�%�;����V�=�i��.o�̜�W�f�@��	�ʀ�'ƜB%���8R�r>���x�}�'���%��p�B����?w��S�x����[j�T����9�IېJ��#��kL�0(����9�<�c�Uv���%��j����3��7<���jb{3EtBR`�z&O�������B}�NH��]�v5uB�Y�T[K��R�q6�5�)��"�Zk����7��h�"h	)�b���0��yg��/��r��	݋�}W�� D�	U��I����Y�,����XR\(w�l�2�!Jt�o5K(u��̷�����{2p��`��c�d�Ԩ���q2SŊϋ�4�"p�RVU��,�i+8��Aw���"_=��.mxT��Y���@��5�`���7b��Fu��k<�� Q��+/R*�̽:�`:V���W�z�%qPѭ�%O�L,���񝳯C&��`\tS��
������q[�,�=, �M ����f=:4w�Xq�K���es`y{���Q���P B{� rġ��BBG�8��^5��/e?������+KmνW�����E�o3������鳦n4�J����Ż�D��+�tv��U�ՙ���(�	�0'h:{~�}�oCQ\�Mu��8����c�S����%�T7k�|�[�Xīy?�"�ȑ2N�F�`�����[�J��N%~�����y9����lR@a�#���8��c���
1*��`�$�^X��w��o�K����5���zATεe��q�`9QL�7�)څ�JW��?0dn},|�h]y��8m��X
��)T���O�"�6&�����ٳvm��xd-Ǘ�*B�L�e�>u�=�>�!?D*�{B<�n�8%rZj��	���X?�~�B�]|�����\U:���n
����.|;B�f�/��=��@��n���X����ph��g0�QI��<�ax^g�|C��Ap��T�o�܍�?w�iSI钚e�E���BoFo;�D^9��
0�DD$�+i���6��q�3�o�C��7��׫9 �۽�C��4�Ȑ�51"��q7dL�\�$�Ad��y������NNA�`al[KV<�t�)��n�D��G+���w�k��5�;�<�%O�Tpɯ���(��VF�	���b�4ӗ[�ۣzp���/Ë!At�O��y"K�/�.:��Q�	9�����|�3�9��$p�*Z�F����8L��/���X�#?����Sm��tE�*������HJܷR���~8Hq�[����l#,#����)Py5B
����-����|�?J���g�qu<4�e�0Ժb��[2ڼ�R�!kӏ�����ϝL'��ݱz�6;[��D7�A<5��yj�0bяT�a$��>�o�Җ��0eC��l1��}�{
�<J2b��5��
e��/L���
�S�T"̰@�N��5�V�U�C���[ �D��u����$	���(M�K��|���9���>�^�5���1�nHp�r��;wi���C0"�uD�yѐ�i�/�PE\���wD�b6I��o�;�{��i�#��������B�T�P9x���!�s3��fZ��M�ۃ\����!�"m���L�<ĕ5E��03�쓯�q|j��l�9�c=9����5/�g�5�����g7�����}02�Z��q�=��-;�z;;=�&wm9��u���}����.M�1?�ݪ�9���U�L7K�A��}���SdHX�2������bZ��Tng����:��rG˾�^���X
{j�1��������c$0�� v1���(v��ǩā�v�^�|=��h���.�Q�z��,&	T@�l� ��=��yj���ӉY��,��'���N������bl=��
VD�7�Z�ܭ�q\�CgAL�G��%�.���N_ ����;�v������x��!o�^PZ{5">֯�`�z�PWF:������SL_9������O����6Z�Ԁ�o�R ��0�έ7��2�2�L��]��G0dj�!���� ��bit��KOX��?Ǔ�c��/����IZ�yh�,`'w�<�B��n����E�P\ko��[d��n�Bam�����u��)�{'�k�$��@a���Fw������c|�������u=v�4N�^�4�&�8��KL��-�,�e�s2Mb�~�:�ś��@��XH���C� |�f(8_ ���
g�����a�R	�jhPL�9%[0�	/8�y̅d.���Y��Y��m��B4�~٨l2����u^�'	A�5c��,�.��7:��PP�;vچ�;"�>]K<M�.<]�:�Ӗ�l��6���
r:D�gc�-�f/�[�h�,��Y@l:B�w��v��<z#����j��f��8 ���NV�����CR��:�}JɃ�;�l�/EH�Y����р|�y![�C$<��k}M'_�<>R�ѫ�2���/�T���X|���gM^��%}GT����=<'�'��I�T�g�5ΤE [Rpɞ�0�{����H�\�\�˞ЋDh���40�n�4��w*A}��м�E�n^H
Wg�?\g�`��p��h׷���4�K�v��t���S?�{��a�y�m�}�h�xX���a�9~�
�7�n�q�љ�]fQ�.>uw�<���gWJ��2��j�_'c���C��'���r#p��Nʆ��̰�I H��^L~W���JrHqΤ�>��8o��%�tњ���q�1�H��⡨N�*8�	�\��]�ܣ�#�&��1�#�1��* ��Ւ���Y�v&�yM@X�M�%s�>p촕m^7���x��vʣ��]ܰ �(&�l9y:�ͳ��*0��0I45S��:��ЎD�B\�A?�����ۮ�r4��<�r��+7!t�ص���ʊò/-��R~�?��lg�_)�z�A�Rs�~!d �,��T��@��	��=64(C5i����WIh���U�%t*w�"e<�}��Bur�b�jݪ�.L�X� ����4���Fc��8Sc8�u̩��0vY�d���5B���ӟ^�k��$DMҲ��*4M~�K�S���=��p}���ˁ�`�L�����V����9xqOv x�b����U����^[>u񂮉�Ц���N>��&6��R�z�tHCU��@���2r霙ҫ�5��l���@,ϭ�<��I��uz#2�N�����G&��_&�/?9�J�$��@.�G'*yc�ńC�L�֧�b�мw������$-��;�ȵ
V&������{
�����!�֪�]�Ss�Bi���Ï�����(c�~�d����)�.]�#��5�1�/�����`�.(����Rw�H7�t;�j ����dh��tL b	0D���̐�wRr̪�,��V�'�fd,���G���gB��ɤ�����8���T��U��t��3����Eb�q�Zp�2��l�#��}W�����s	i�m�}�K#��������;�w�Üe��$����+F�7o�3��!��ت��!#z��C�����y&	�v,��c�.�����]�X��k!���#�?ZK�A�*��g�w"%Yݼ�wE裡^���A�y�v�1u��!����q������(:�=�;HpI��{���i
XXz$�rE?:�����kXv���4A��<�_�o���;�>k��ƚ������sj���V\�RuH����x_s�]2V�e�)c����jWL�g�1è���P�ֱ�fݿ�<�� b 	/&�n�xkM�x2=F����OF��e�r ���Q����zh�#1��H����EK�X�P�k{�70�^�ꢛ�����z��:�}81}~.��ݹ�k��5�JM��A�l����y�[�y������&j�n��f��>����h�d�{���;i5�)��U�r4#�si�ź�w��Јvy�E�B�8�1��jB�'��ϰ�{J`�UE%��.}����� ag��>~��/�:0���8�h�)�����oC� wc�>���VѼ�t0m�R}ï�p�'Eʢ��FG�P��%�%��6� ��¾�ٺ��\�Ԯ؍�p=RM�T4&���p�d����(�!���	�ƕ�q���;�.�o��h�/s������5�����B�*��bLQP#�F��%| `/Ԟ���u�3��X�i,��������]�h�KP}&����w?(�Ӌ��vs��D0�s�8 ��9jΨ�Qހ { �	����O�ȁX������R���d�V���L�i��лV�<ąW�/�nF�T��WD`��FL�]+!]���x(w�!	\��7�Y��}��v�2��W5��^O*����.Ȗǝ;�)��ҏ\�TV��G<�p�U�Y�M�>l`b���/x<��|[�Wڭ����u������s���O�H�䃰�8C[���w ���O�^�N�'���F�8E�`�N8�����i���O�4�� Ǿũ�������?ff�L�C��^�[�9�(j�����c��/�v�Φ ̉��_�b����]>�F�'�� ���_p�2�s5Ui�l@x���w"�甕G��xE_�3yD��6��<$QJԩ�H9���S�-M��t���������n2ls� ��5.K����'zۥGm���7G����	j��G�}w�3In G�O�P����G�Q���jR�.��-�R��b���
�eC*U�,b��(� a�_��u��>;���w�JkϞ̬TU���6GD��C@�EV��iT�#Z����\̖�����9����c�	/�c�e&jT5d*�=!�'w-��'�~�i_�E;/�v�D��s:s�+��m6����޵Me��0Ԋ� ��[0's䠇߱Lt��P�;�%9/����7���J�4n"�6��Dg�u�N�E�ޓJ�1���� |�"�Z����Jea�Y�>�T�dٗ��$�����J#1�bRBN�F�紣�h�m�C p��b�JLכL�m���o��#���Xƹ�N��!"qD�Q�1a�<�����x�)�6/�(��|[�o�Ȼ���[��G�v��$(���4m���n�ƒG�}���}�J��R�T���1�dn�9���:�7 ����`��>&U�������)�U�Z-K�Ep"��Q�q&�[�5��~�q���$S��K:�JuT^ y�� /Ŵ]��C}�q�&G��l����[�S�J�,��f���š�N��4t�kl�;3f�wH��}�B��i�����AR����=�`�"y� 09+�f"��-}P�M�b��+��mӧ`�b~�"{47�F�n��1��@�Cu�H�W��������9�����|N���kJ�mvb���`1hHYf��r�O}���C"��v-����H������vŞ_��0���~u�A�*ٟ&��|;NW��B�i	��j�|�8n��)�*t�!����NmD�2[�}
��k笑{�m��,"�c#�!_U�AF��x�_f���^�(ެq�%o���L�:�"�1;p�o��O�X_]�i/D'�u�/],yY����a�r��31��}8L���(�n�,$����i��z�{�L�+� �����0�l��=U���F�����#��4/bM�4�=�$��*�PL�8��rk3�K�r��<y@d��wp�S��ȼ9ȯ�a _�kO�.�%��$fOY��`���Vj�[%`��v��#���p�E������~s�ES ��/m҆߼�~g}O�<�v��p8J���@�7S�|n�Ƒx$:'�}�Y1-�vѹ���\�j�m!�w���s�(N���5�x�0;�g��� ƥ.���$�-�N�\~{gp�GV�x[C�19�n���$ M�%�\�����6*��s�:�`������~.���{��O���Y	X!S���WB�H m��F�<�BeP���ô�BKn)L ��?���y8������r7CoJ�=�򁉎������}�I�!�_k�f�:��״܃���X����� _Nk�v������vb<�p�[�!K.ȃ� Q:)�vcVF=,G9�;�3����\h�#��)7��T�C Zuى��h*���;vf���r�{��QM:(���R��=��&�ꋋY�R�R�/�4*"��hR�J&�)~���}�!d���
6����O,�Ǧ$���0G����n�^C@��IO�=��+ﴽ ���kcΜ?�� 쳀���* /����Nu<\����&� �X�_f-V�Q]y�����ϱ���[�[)nZ]m~f�[XkOC����<�������G��:k٪�M ���Ơ끥���7�l��L����4�����u�>�2YL./}3��J'z�!��z'ǯ�^}��#�t�9,W�N��S0;�����h)��.Q�8ݜ'�;?��w�Jꔳ��x!� =��\9Z�4Vn'�_�"�fC���thv���82�s�I�	�)&[�Xlm����8�/߁M��Tշq�1d�d+�Q�q�[6?��O���� $�ɫ(�O5m*��Hg�k���~���D�R-Z-�l��]����z{ۑ�Z�۵�9�^�eS�&z����v܍��(�hFG*ϱ�(ku���� '��<ӌE-9T(��wk&JWu=M�����~M�)��Zl<[��nF�����8
�c�;�A��l��#sI��5Bo�jK��%:�W��I%T�F%��+[�- �b.<h	����؏���ri=&8z�O�E{:b�n��ղX�����;�Ek�ѻ����2�&��)0��ޗ�8�e�4�I�9�<F,��n�?и�=q磢��ۣ��֤+>�9�� e�K���4�����s��?�R�PPSq}�7��~�W&�g��<�aMU����8t�S��ھ������0�T`\=��Ʒ����y	����I[9LU���P�.5�p�Ef���_�M0(�b�>�V�B��c>dv�J�����r�eEj����"kդ�������n���䓣�F��Z�J�z�����Y�._�R�e�c�H����l�A�.^F�X���,�O�JZK@��Yj����{X; q�P�b�2���Kj��g���-��k.�wYCr��0��}���H%i�Y/�֌���)T���D�cJ��(.����"`����dN�����CF4V�q�z���zЊ>n�GT�GdƜ��rAz��X,z�c[C6���ss�nH�Y�P3� 5�>�w$.�%����P��gG<���>O��ֹ����,�RQMV0��/�B��B?g���y�/�*&�5>��Q�Co���Ƽ)��C:�)PY4"V�[�8��z��l���^�=}t��/^[��X�E�z�CCL
��W]���z���D�	G��$iG�t�.�-P#�X�N�:r����n��JA ��`�A���e��a�M�eƴ��G��e�K��Qv���F���z��eK{s��{�m|�TD|:��m�*)R>3�o����`��T���
E�gd�qV0��0��:"��Kk��{:*'�f�-��Eg<���侤`����>4D�t4K���+��-,�Y�
)By�?^�M|Ei�7�!�UP&_��6T~�q�s@��t������*ƚCE^��Z[��n�9X0Q��1Å�c5�����,A�ZBaD�+%�l����	ZJ@�� é���j[sq�I3��؜�[)n���D� ��b�;���&�<&ʸ�d	��^�/M�� 
?���]�¾���6�!M�e�^�N ����ZRߒ�z�5W���
S���Y]�pXU��O��F�װ���3�_��6ڃ�
9ų(
|���;R�y�z�뒥?�I��|�=x{O�Wk{M�췃_
�Hu�7��1�;Uq+�|gn.�}��h����E���c-��Qein�q��(E���|NΡ{^��t�i�o0��b�Xv&~J��ԮmR�oQ��O�c#�y]��Ȯ�:�C*� ኌ_3"A~�(�����/ڀ�MvYa�.�.�;s8	~�遈�HT�P��?���_n��)�1 �q��I
ӳ�HY��fe���bds���ɇ5
� �	�\4*#�Z�����3U�{փ�\�`�J��D5�WV�������a���l�̨p�5R�LK�@���È	�u���������F{�� ��nMd��n)��� BO�JSR5�cy��N_����UD8N)����a�J��<B�o"N]FD�g��%�i�%Ū�������n�|x9�a9��3�~�� ��/q�����U�W5S���	a���0�ۼΐ��_��O�c���h33�ـ/ӗ�l��	���!��x��r8k"^�G�E�:vƬ_��6}L^���*�\8��J�bz�6i+�yr�5Rnu��R�7¡^u�fiC�t_�&|���L�'#�_�����_@�������95cy��P�;�܈�C"��"�U�C����m�vC�9��E�,U��?8��x=��$9�	�a�����R��l�%��|{���Vڐ+܃�7�(8�W;��0	���.�_b�	[���G���j�vir�탓Y����/�+��d��O��վ��?]�M�m�����V �z��;=�)�F"q��8�c�dz�L�.e_Ʃ�f]`�k�ԧn���į��2�������!�L�:�!��Cc���$1�H���s�id��$�5�\C��NP��A�f<3���y�{�s�gR�U}���5��&&/��l�W��������z\�����b2�sOd�(�/m9Wu�d��3�K�[׽��)�������p��]�1��ds��ArD��A���̈{`���ځ}~��4v��VD�[%�I���L������.M����g%2�A��K�NѢ6�9Cp���;��.&;�Q�<$kh.)�lM�"tk�5��sU����S�<�7x�9j�+��AӜ<�y���<h��F����_��:oA�I��gBns�"�io]L��>��F��_J8T���>�-5 O�2_h�&���'��nCI𨳟����{[���]'x;(r��kRt�C�`�[P2��3��W2����"�2��sKE1�k���y&����_�H(���7�E38U� ���'f᪌/���\��6Ƀp"�u�88�1����Ί��5��e%dg������Q� ��t�Y��T��e�V�4�{2������������U��4䦣�^Bד�����,�L�[IF��+k1�j@��m�Z�D�2�v$����l�.�<�f��?�=Q�L��|����#�<����dz���0j�XR��Տ�?�s�G?=�F%��ү�O���~��S�2��\@���R R�)U.πV�x�\>��Y��PU5��	���G���I��\o����׀��5����'��oJO
�˧�G���`}��{�E��-~ �>D�dV����7���m�E�鼝�JQ��\=ÃŶ(�H�ӧI�?T�$Y�[ď�}u��B1a|Hd��N
���bx��o&�4��?֞=K?qE��lYw�2�5*	Zؑe�J'U73�y<92}�式:���4�n���o��;�.b�_�����&��Vt�F�SR���0�O���-���8�6?��
B�9�\ݖn���4���t��-z�tR��N,<���aQ8��<�D~D���$�Z�ja��.#����GD�����W���氞o�����K��R�v�,v�s�E�E7	2�t�ё��Rb� ��6E��b$��#5V	����?��I2�3���$L��2����u)�+��N��E��[!
���� �YlN���w��`F�в�:ןq+=�d���A[p<�����`b�d�Q�b\\����A��σya���Q$*�6����Ys}.�z�T��_dK��JպN� �F�*?�וY�Z�u#�8:,�7tc)���L^�::���c��R?w�K�΅"����� ���NΞ���o!F16�$պ��O����y�e�\9��x��9��=w~O��@4O�����!��@ ��d�m��W;'=���t�Ђ�q�a�IAQiv�Ԑ�Dp#��oλ��M�=�-�����gU���~�U1�}7��u���|;���נt4x���m�uIj�qt�?Pk��o�����ļ����;�Κ�@��YB��e[;����#��ܯ©�1��-�qJ��Aҋ�9�m�jq�<��E�y@o^:�gi�5���	L{��B��`��[e6Pp�o�H���7�<p�����Z�m�ﴭ�s���0�px0Ŝ����p���k�w�����	1Oͯ��G+nmq��pX��钽8
��+(x 0�@�9�@aV3K��J�ӎ������-⠄�o"3��`�ws/�<�{����|����1@w.�s<K�G�v8K T���8��Id	�wc9�<����8�Y|��S�};T|ϒxv������ᅨv9���q]�����`�]ǫ�ѧp�:ʊ�ʃ�N,�r ��L-�d[B�k�����9�]h��j�8��D��`P����_���~ɞl|�G��_]�L��-������tN���ZP�T�M+�^�OMe��h��Uq`G�6�����oe�+��ua�r��G5�!6�,�'!�>0�X7?R	��zs~���m�%�=G�B7������~��TЌƙ��~�!���i���eiD��{�Y���O�,�o�!��Z��\�rG�]s3$A�Yc�����$ЄU@ħH��5Ӎ�3�vP��D���Q!�oOF��2���yu�_W�E݃/KgH���A��w���#�p�'/�Y���g�Jdr��i}���F1��Os?�� J&D ���O�q�V�!֊��("+���H� L�2���bJ*n '+��D��buz;I�.�
���������u�������9�y�!��j��)�n�Qy�AG/I�M&C]5;�Ȕ}��Z�7$�Q�q<�/6�qC����m��km�y&�s����5{�5��<K��+ʙ[�C����tU�ǎ䤜g\��B�˄''$~� �o!� �3>)
�+A*.'Û�s��Kk�/Tg� �,�OتX����'�YW:���X�d��_�%H��O��Xe��E)jC�<���?���@� �R��I��U	��������0Z�y�v{jw��`H��F�)u�D�#_ѐ�.H��3�eW�l8������?�@f�[�:k�zez����8.q�}��޽�&��@YR�NU�� h��=�؈
���	�ޮ�Հ^Rmu��|z@��ѱnk����;��MB�-Ի���$~W�d���n��Ю���E���l�LV�CeM`���\{ЍW�l���ڶ\շ��tO�!�(�߇s�3�z����2vu�@��;D����΁��v˨���ZI;(�"�(�oY�Jښ���~x�,��������8M���YE��{N��{&$i�>�4J��*�5������4��UOG1�񓖅��4j��5�8E�w��&��&Ji��&"[k�������[x�Q�5]��u^����])L/{�2)zQ������m�S��<�����i�rjA�"�V������=P�;Y�|Lh6���#�$��D���0�-�.cK1�����NcQ~�g��)0:��?�LV��p�3ȫ���i��+M���35��ií��\�b%����b�(�u�1� h�F��ʧyk)	�	/�!�G+u��b�5a��O�Q�a������-���p��t;�ܠ�HG�*y��E
��
$�!���g��UhF�<?@��v�PK�Lo?,Ot:��`������'-m�;
3��O�4?�?�����_:�LF��)e�C��(|��w�v-8j�͇v^�w��T���˝����	U���c�y9\�I}�
�ܸ���-؀�@�,��,� Md�@�QX�g͟`57�sMR7��A�8�$^^%T6v:e=�������I��<m���ݸ�E��!(
6w�!�In���I���w{1�=��aߠ]�I�46e���+�w�n��μ��ܧ�!�)4vR�iޅ�({��5;�q#�\�0ٸ�t�dN���q�M��~���)l�(�%D|*`��z�9�f/��KT���	�|��c:I.�sm�d�^Ҵ^�u0�m �}8R�=J���.�\��Uf�uF?�f�?��� e��Y�_��M"g��n�(���<�X�����:�̈́V 1���e���9�~>����bj}��"�"��df�5¯V�Z��3 ^QÙ��x�����Q�a���X#�5*�7,�!8�R���_���Zm��j��ʰ�0�:~��M#�����~P�s�����^I�e�^��l�߹*h��!�u��-Wj$�EJ)�d��}pS�6�$��;	Z�$�.�� �Jɏ46�S�t������'����b@I\u�A	��3��)��Hu�l��5!OJV��sw�i��b�[Y{f�zo����g,�(a��u!ͥ���s�����e��z��Qrܳ�4�𘶧�+(�$w��1�Y"��|���}~�y����t��h5��š���!�;���a~��$+��]�ba�T���o�9D44>�[��Ӊ�W�Q[�%���2\� ���^PP��;��}�M�!���o���r��K<jI#d�a´�5��C�=�-S��� ���Y��NXk��3?M���AʜLo�4����q���;�wJ���E?XM�<s���;�+�P��Ǆt-��m=�J�9k�u�a�:�VB;�gQ�졪��I�g�}ս��ь�7�$es�p�~4^5ܟҞ$qQ���v�ht�B�z����2��׍(��ҙ�����ȿ8�S"Pq7K��ɖ�ld��e�E�ya�v���bq�-��!��ZUIC�L��C���U�y���q^�5�&��eD��>u;�B���Ö|��u�U���}�I�Ňe,�ba\���� ֝�B���K�����S�k^]��C�����1��_���}�H2��{E�7-*:Pq䪺��ؘJa�B�������+fh���ڀ�)�ы<g;?�V�zѠ�"1��X�&�Abz��	����� �����ri��2
���ǀ3�|\�i<�Ԃ[�A��z���@�k�6�wT��W���Q��j�����b>�D8*\eC�R7yq������5)]<��3.�ls���lԵ9������t���هR�*�w� HS~��Σ��u�y*D	��T lY�����߼q�	�'fP���;0p����˥�Ix��T�����v�;W��n2��}�Sc5���/`[�w��k��N�^[�ǁW�s�J���R�z��l@\�b�,ޘ@��RC�,��^�����5u`ILU8U|ۥ8�h����Q��tL7��4M+A'�+W� �Q�dO�_w��Z!���%�v":7�a�z�W�WрR��	� b�gw�$�I�U?���o�T��	�b��  �������k��{PVB1@:�k�m/�fL׍��"G8���O�Ui�+�V�On2�b�6f�,&.7	C鍾Xh����hg���4s���/K��L�K�lț�6602��dI���X�!��su�$J�I���S�|�$�Х�ߩ?���7��u���-�����qdepD�?���evٟ����ooM��^E?��z�F�(��(��ʰ���N�*jb��N4��W�fQ��z$�m��P%�U��+;��ǖ�^��S������^+��buEF�#�j�z�/��]�?��H0����4��'Q�ƒ�
o3�/wj�t�䛫����;u[65,��p�K �X@f�;�|�(L��\�0�aW�OC$�v�,����m�9���x��C��øn4Je�����aCG�H�>c���}��:�~D�H
c2P��H^�_�#W�~G��SD<2��p}(���t�[st`2���(AU��Yy����Og{$�Z�?�:�J�Z.�$K_\;~�Y��,U���P���C�Tůc>J~�[�O![O����"���#�shL���r��SE0��2%L��vRdz�Lf�R$m2ȉ���j�#X��HO�`�.%�'O�	��R��ǢV�%'�������=���o����=��d����N
�zE�����6cU�T\xPg��lM�NFm���8�����vEM?��E>���_� �X;�������X�A�H7��ZR�j%!%��T���y��!H!Y��2�U�������́쟝�f*�^Ѫ�)��|�\pg�'�c��_(�35�Lٞ���zz�%\2���ex>�G�	��'(�Am2�D,f
��ӄ�s�"�5U0�x��1 �q�.�^ݬю�fm	��Ƌ>�n��:�*@�`7���Cz���9?_�Sx���N�.a��eg�u���\F��D�8�ʞ�\#�Ff�"2H�J�M�0:u%ߚ���[ߩ�D��h*�j��72�Aw�~�N�b���V��.�}�^���̐G�H/�IBR�{���į�ա�;��z���6�IhԔ�+=��\�i���4��ߓ����ѡ-
��7ǚr����w��JX���r|��LQ���D�j��X�"Nʶ���}�D�a�� ���jF�J�w{P�X�z�e��X�d�����X�G�[�R�	�;;uK����cyF�����,(�SL{j���2�Y�^5�/D�G�7۔��5�Z��׻�;��Okh(�n�Ԣ�h/ÿ�c�+�u�A��J2�q��Ch�K�!h��ܙ��`Fbn\�Iu�,��zC�	�v����꣕9^��\���F4��(hq�.�e�X.�J!�G�[q��Ed%��a �OSA6�c��S)"�ɗ-����8�OE��8]Mru41�Ѷe�������#������@)"��M�6�	�fKr"�B"�>�}����x��{��/:�"(5_zi�J��o����0+��	���8S�x�\���Q�
�����_��!�%(c;���!:�J&��..�$������R�b5y�el�\aI�U�l��$�*�\P������$0c���=�#��A�������?i!əp��4����1�5�S�N�.Ag��ݣ�S�?�Ѫ7,s��i0�e�Iu[�B7��^A�k����)���2�Z|��9N���u��t�w3d�!TW�_�aN����4ag�[���Ȋ���9,��ā�gʯW)�o����3���\�`���,U.YC�2�+B��z������WYz���ft�L�f���C"��'�U���ȣ�}��xf5u�^�#��	,tS�q
�;�����9��41����u.9w?����8X�8�]�9�.�G�lUZ����Q.�?
MZ�=�IJ]ģ�5N_d�4�<�\��ֳW��*t2a	<��ܩ*3�'d>����ڣK����������=!� �<:�8>��Xb�b�w	�=,+�+����
�!�&�I�$��rug����e߷�����껵��	P�~�����y�V����}�����@q{:�G~(D8�.�����#�G��N�@��4��	D������!���x�7"�i]�߮Ќ1��P_/�%00��T�n�̃�Ẽ�b.WXB/�u�(h'�ZʅY��e��:���Ebyf���C��y��
-�i���ӉX������GT�ث>�d�ј�VPC��Y��|{�A��jOy �̑�ta������O����2Ӎ�a1�[��ʘN�B�f�s[��P�� �-`F-a^'�܎��"l� m�K�<�!����%	�*fj;�X��e�~�#g0��Le�n���_5�qnd��Y\�7]���p���|]�\ڥO�[2{T��P$[d�TICN(���&|ho�)�5H�7,`PO�Ad���w�<P�!!���&~wE��1<uw��-
�5�(�T֧$q�4����N@뾑P9JQΎ�L�1�7m����u\��:*_l�3^҈�x��`��9I/߷���ܦ��ɮm��7l�����Zq<�p4�� �Æ�Dx��tQW�j[*��ĳ�����YV!�2&׬�e�
����	&/+E�=��\C�����rz]�{wfn.���W�H�Q/rr�l��~|�p1	n��<1-IAXo��mq��3vaG���W�mW�G&�I:yfL��;n/l U�m��r�\R���(���Y-l�^5�; �8����qjR���k�2t�o���.� ��k��`��.B�3ҙA��ecF�uT�1^#
1,���o�L.!�h���^���^��m�/^*>�F΍>ܥ���tInW���π�D#�W6�}�ܪ�_?�;p|�z:̔���k7�m{�Z���=/��v�w���tQ��R��>�Q����׳ޑ�����6jK��	��>K�<��5� DpE�BUج������@ɭq8�$���J� �Gv��������\�n���3���{0�t8Ԁ�����J4~�	�7��׭P#�n��h��?����jF1�!����q4�3���A���S�#��15j)+C9��{䎐Q�|�p��̧����Q�\Rc��f)�'3���ˆe���(��>��|� �s��У΀w��`�U�<��cp������
g�%DX�-J�4�z��q�����n�a��z��C�{	ִ�T�>��I�$}�Ƶ�7_H��߈��G7�O�wL�%���?���C��I���)�g_*��������JB�y���匶�^��*&)"���cq#'2U2�So�+heE�pm���2�91�����z�t�	�Db�����SMpݮ��}�_�^��dk�����$n
1=)*�+�(� �-u����>���L��険�6w�k�#���c�����ڭ���h�%�����]1}$���}V�J`��sJ�4{�U�a�I��b��c�/D�XnNy��LU�1�DD�Z�$(���K�8/�7{�.C��HQ\��'A^&b�bWPV�;t�W���_�h��
��}6u~��ۼ��(=)]g��M��d7$�lml����u{+-'c�́_q`��Ǵyy�O�6���G�e~��|��P�97��cs2mOI����d �Qx6�Qy�����.���Up�s���s"�����R����}�C�H��H3�%����/�HN�o�}�樦�t�c����Á����n<8�#�U��b/�ć���w�
A/P�v�K�:�U�ZXېÏyP�6�ܛ��%YM��d�F2�vV�>A��@,����]'�ˇ/(b���b�b
9t|j̈�=�d���F������J�f��0��l�&�O��߶�2���-��Yq��l�^���,�ܲ8� X��vb��:��`P�ٹ,Z9�U��)f��3��̏���s��3'�d̄�gG��d�K�	�y�4�UR�`2�&yAa���e]���6q�X� ����<E����v��ʟ���c�F����H�	R���h-{�GIDֱ����4ǯ7�-	ߐЎ��f��=�z椲��}.��r�q�E�;�����<׹�:����'�Bҥ��L+C�q��5��v5c�:GC#<n\Z�W{��w�����w�P@���e?SK<���^l�����7��<��P�ዓ��v �׻��tёS/��C,�m:Y/���˃Q�t�A��a�o%�l������?�l�kf����<B�I~t�
WYS��?7p�5@����[�)��YW�}��H����'����l���w����d WN�в\gI�҂��zx7 ��Ø��Ԕ �y��	��WW��,�#�Z �\VpY:x���.ruP�ѧH�0��V��@J���^�-��\9u����P&�wC,��ٕ�ڂ�d�U�y������+���h³xS�'���W�1��-˯d
���`��A�c�[V�xNCӬ��Fo^��/�Lp�{?�R-$�0Ʈ�7�AU�] �uqĲ_��0C��|;����J_�F:�j1��g�e��'i<3��Uk�}���+D��z�9�g�pߐ���U��9o���8&O��|>���(qC?|�)��x`eI��.�?��(֎��X%h��ځ�=<�H{�Gs��N��@��q}s����D�H�L���ת}(�����G��'53�HZ��V>b{O�Y���(Hx޽S�V�ٲ=�c��u�W�R�u7���W��O��=?��Oﱧ�W�^�.Z��Nw=-��-�/��!��j��/E�d-k�I`^'�jgr���|�i�s��'�w�i�6k���-�Uh��1�$��{*{�kdcd
��Y誰3hn��Q|�\I�!<�}'�E/��eo��ؾ�E[&0����,(���}�.^��+�_T1���ʹrCI�"�5#,��k*D�l��ذ�~8Ĝ)\DϮ�i�}rH�+!z���!}O��BH�P���E�L�\�N}P�%�[��~㕱�V8�O�5�b"t�q�I��t�<.�rP��Ļ���	ter�7į2����ƨM�ʓ�uN�/�#��qS�zT܉@?�����9@lS}G+�gX�Cy��o�/��2�BZ�X���2_t[_o���T�1W5�:�x�����}��e�M�5����L�����9�M��U8��i�H���
%��B*�"��J9�%:�m��USe��z� �^x����~�;a��C�ʤ�z��6ӕ�mS�=l2.F�g�j��R��ل��ԗ�6q���3��%����l6��_m�!~v]()���i�JH#�)� ���Ap�����n��㗗�u�=�d	~ӈza@E������Lp���i�/�l���b��W�V����m�cif����S;������x�r[?j*c|D�7W�|!
��-]�JF�B$�ӨQ�v_�+Ȱ��bs�Z$w\��R�7�b~��2����^/���E�[�"�Z>aN��*+ɐ~1B>��ODxW���[f�ϒ
���k��D�\z��y�yT�:\(���6\W���z��n���[�)Hy�ߔ�X:sÌh��5�E ��DOd��}��(WՅH�D��(���*$ί�"��:�˜6~X�Ib��x)V��yDv�3���jh�>v���T�W杺�V���4~����w�:ܻ�k*B��-��e�JJQ �,��X�YD�7��b?H�c�d�f^%̧�L������&��'�ղ��5�c�?i�KeH��Z=�gɛ$uo�p�m,����Պ�L�I�>f��q��cE����R�$�H^�C�bar#a�YǢ��Q8[�o��՟乩ca���w�������*�٩�Z�9��u.k!�N��_O���%�Jc�!A׫��S�f��lmq�L�����b�*����h(Y�U8��.T
}����r+g�v(�ڡ��1�����H�I��+P]˛��6���8�P�v�b��З�f�6����!_�����f���Nu�g��k�Ib<h�)^��s/�	����?	����p?���玀�ʢ���Y�E���.LL�K>R��Vi֔P��P�P,��i�����Oe�����6��N�����s�9��J�S�=����>���#�
���>��]C���a�kuqh;�qJ��oYȮ%g����W�D�e�;�s	ԼҞ�.�f7oO����:�4�H���x1�l�����QlQ��T@t8��AXT��1r�k���$6�zJw�1;����7� ���Knѯ�P�GM�;Bxr��3�E�����WK���1�o2�L	�c�e��&�]�W��Q�h�i%|j�d,[z���KǇ�6��I��a6z ~��xΜ�Oq�Z�@%{O?hZ���S�i����-:�i�u� �Wr����{���5����u8d�J�i]b��A�f}ٙ�H�:RߙE�3T/9Z��뛵�n%��:F������Ģm{��2�O�:s\��5㳹>ϟ��K�E�mY(�>n\�~��]@?k�5�Y�Mㆲ8׃7��:�3[�Y�)�6|��E-2I��3 
�����+к8���CB�Y��䐭���l�zN���b��ǬS1���M��X���hn�5���|�A����x���C/��5s��Ln`G���hF�t8#?|x6��[�i���ZƝ�`t���P2�НV�-;����U\
���U����>h«���ֻo��������ht��g��Ӵ�d��Q����Ȓ���gJ��p��V1�U���"�.�� ��#R�?;��|����Fm�r)��S?���닎)E����w9r�r[i�����;���4� �����⑹b�3��I��R���X���R��5~x��rƢ��$ߩ�.�KN2��b=��
ޡ�ӵ1�/��]ծ.�!�C��dv�ҘJ4��&�s5�[���9u1:u�뿥.�n��M����W����8���:�!l�J���4x�zZ�v�au�0[օPqBq�v8o� �ni�(���U�h(�P��.��͡�K:Vۃ���A�S(m'�7���h�97�^9��zuv�)Ƹ#:L�\�?�d͟ �dj5kY�O�r�ޑ#Ж0�
�H\����A��9��]F��]�q��˸Z��7���� �X�.�����"d]\#�Nis��P����"h�iMc�ǫ� 6��r�`����2����6] ����J�{��yp�I��m:i;�PK*T����\��r(觴x�d�l�T��R^({��ۙI�ZZ�v2�?����Ю��c�����6���.�8H��T�\��V��R�m¤E��gR~���k&�d�t0Z��BY�ZA)��){�CUЏw[��`�G��<*�+��kBy�\�P�js\�0��D���,�m�ڛ�E�nm��}^������YJwx1�|��Y��0?��������)s�w�R���@L�i)	���>ٛ��kPsL�`��h����87z��G	�oM�G�����8�D7��R���]�C6���БhP��R�S㰂B:�@w`�JT7p�|��y��/�����/��U�e�X���5@�_u�1�Q#c�b.%~Q�Ȱ���郙M��i9l�l����Cl��0�V����fǓ$� G
�Z�S��꬙M�@���d����x>�q�u��~$(q��=(��;CY/��T��V�-��^�ܛ:������{���.թ0��.��F������t4��y���Qd6N7{�oك�&� ����[]MO��c���� �����L)K��Z��?����Ҷɰ�W)a�#� Y+6�X�5QW�cgt�=���Y?��f
��B���������ۯ����9���,-5�A쀧�R O���l�I�����M�:�MH��r����Z}�I��_�?:$�1�I�f�k���.}.>P:Ŷb���DqsJ�4q+�X����P��u,�Bv�t�l�ߖ$�������'�ʉ/ƪ;�I��n�W�Q��pJ}�E� l	�A��=Nz�~еg��e�g����<����z�Tv�]­5�p�HM~��5��ٽ�)ȏx>E�k'�j~����Mڪ��]oBL�L�Ր��pe6�3a�2�â�棖U��e����.�є�t����m;��w3s�J���S� ���2��[~�߽(Qp`�A6LJ�8�j�nȶA�3�|�Ë́��/��+w���8�2{2����V��>�����m�J�H�T���^�PY�o��7�E҂��y2�G��"F�Y��0���\9 ��6��,-3��-ܰRCh��ì�f|��� �g��(��r���Gr<�݅�1/�L�{~���Lt�9Z	c�mbT������	��í�`�팖z��c|�X�R�V���Ǌ���&E�׎}�����v�8f�S��V�Wڦh��Z��/q��'�=b�$"[I�?�p�4SJ,l�I�{#"iYs���!=�o����s�,HQ�}�@ƠάQ0����mC���{P�1�a��W<�Jy0�h�0i��E���UPT�_z���B�A�y�F�*��9�"�V�(�B��{k��`#��X�out:�~P̖~��٭�����\3ܰgx�1[#E'-��Q��}�I�8��]��DqǕ(���Ž�o�ק8*S�<��N��A� �c1�����z($27�.�=¸�Q�ߩ��fA����8\��������g�2��rn"Ȱ4В��E[���gد׵�������^?�h{��@�2����/Ծ��(�(��3>{���L�|J;4m�/Wi�۾{en����7��0�"G�%����1�Z#aH�n���O�r�6y�͒a��{�]Q�D_{���� jV��|ȝ�	\�Y�dq�8!5��a��X
���x�ϴ�{�[|����!�A)%���[]h/Έ��c�"A�l6a�w��CVfRГ��r�$�7�?c��y$%c�p��6�^i�=�����=)pip-��T��4S�i[�ɠ��i���̏"�ޑ�C&FQ�܀3]�g�Vm
�ؒ�϶��N4��1T5!����	�zgA^`Li���ƋXL��ޜ2���PQ��4eZ��6��hlv*��O3Z�.�0��Y�j���;���?{z��)�ц3h&��H���cq����c�?�E/վ�e�ٛ60��<P5�A���A�zU>r%�L�s]x��&�u��$J��1�0S7�3����s:@��2�;Y/A�(��,��9�o|򆄲�]���U�J���M�v�K�3z����M��N��{!=�/X�XWX�����44�����<߾�;%��xa�§6\���������5�[��v��B>/��i���ѩ�|å�@����3u�ʸI���Kko"ڋ �h>f��TCjw��Gk��I����d�#�o��i���9/
�����lyY41�*�On����X�Wչ)u�c�[c���b�ºտX�|_H\�K�z{G0_��(�&��ȥ�uPAdm`9z��X����m�=�����ڧ?�z
�qhz��	�PUŹ�t��1J��!��c���ٯ��rM�T�D��(zڐS���z�P��j��Ư~��>wJ�
$z��%�����d#(6q�-� �1�����a;'̓x�&����N�Y|}� ��R6��{Lr��z��������ƿKE�:��B #=Q"u4I�3	�ꫜ���͂fm�,)��E��{BȰf�*�a����7ܡG�Q�3��Z�[�g��ڗ5#��X-#�:̢3�cb!����D�"Ed�!�%�P���3J�]��}u�a}� �,����hV_G)��s&r� '�6-�Wޘ�(+���#y樁�&�l�KZ�5*$,��SnB���4Ǳ�����%x��w�$# O&��tp��"�����Jq�,�S� \f���L�[�Wj
���v`�@	��V'��B�m>�ޚ���*���ڑ���r��/홺�;l1��A9�,e�О���*�B�ڛ�Pn�t>/>?D`g��@yӈ��|��Eo'%���1�IP͸p�52���EjS � �YiI������~�������.{+c|��DI��"��,����D���B�Q�As�k%��H��J�p�`5GϤל������?ܽ�I�1����	1�}+-&�r�ܤ�0�]T2T�V�����%=�El�|�	�k�K�7FV&�F7Z|{#��f�l����@/��B:w�3��jW���3n=��u�����)���J+.��<�1㡚�u��+��	ƚ��j�!H�w�'�@l�;���U�WRq���h^G�&�7��������[ ǻE:���ٻ9D� �+:s��f���G9B�OG+l
���*Br�$������ר;#�,�rl�r�=o���&�n�N��1r
�_���Ӫd��H�N"N�ځ袴�l�Yy4��DWC���3+�Ҙ�l����{ B^_�?K�Է��#�wxtV�2g*��M�BLv�|Mz�AZ�$T�_Ѿ�NquX�4\KIRߺ���.�Ԅ��p�f.�d^�fXT�n�@$�YV��M3����_��87����������E�N��J�_��6X���wQx����z]ٴ���~#�=a��u����H�\M�������n�@όQ���5�AfuX��Q-��u�B���ʴhX�卮�Y������F;Y	��;D�
�š$�.�O3vp_�f�"m,6=�^/BZphğ�q��}<�<B�3�H^��G
�uF�(�IQ v�L	�'��%ɱ���}D�[Z]�׺�z}��[�V��9G�¡s���M{Mʂ��1��Z%ad�˶��[�9�eS�Ʈ�JSG0�
�֖��.������.«�^�)P����j/���4���g����N�ᖩ'�ɉ��E5*'� �<_�4{�]BvQ���&��	S���c�=f��k�31�gi�-�P
���Y���q��w����p;K�հiD2m�Y!|���jU��"뼂�|�-��G9�XڪI�i15���`#�l����֊,�7j����w�f�1x��ġ!��S�uo!�?'8d9Ч]���r�4�dT�9:0�F�[��� 9�����~Yq�s�!v+�Q���<R�����*�ߴ��H��6�%sCѿz:A�V��]I��EN��x�!�uы14fA�ɳ���v"��3�H2Ҭ�Rm#� #�b�7δ���k7�<z��-�a�c)�a�K� 6��@����i��b���u��Z�@W�_B��J
�%מ	�%�l�^0?�4���G�ؾCIP��.bn.U��J�=`k22��Y'm�Z*�<
��09*���K��;a��V��*K������ǟ��V��g�_`��7�7���"���`� $��}��HM`�;�k�;�t��8�9�F�B��s�]�0�6xw
a��bׯ� �S��Э����.�	�Q�װ�.@�ܘQ]�h&�Ҵ �XIk`����yPs���mŔjD`VMF�񩶶���8G0R�>ȶ�oy�J�JPWjQSk��-%�1���c�y9_�����a}�I�)=}�jog<�K�M����Kc��¦o��yҞG5�4F.��}�����'{���2A\����f� �R2N�hw�+^�	�{�U�G�3�U��G~����Ų� ���d<:�#2�5�q��Op9��n��^�.j����Kl-�5�rS�m�;��"~<+ad�C��~M��٩��>�qCC�\ȯD����CcK#X#����:�zB�|������5��b��'�,�^����~��4c��9P���S��+jo7ѽ�g��������w��f}f�S;��4:���pԁ�O(��$aM��`�!�����(���L�!�.���f^�<�9JH��o���`ELd�)]��,� x��h�&0
X��t�������l�DsK���*��K�	���#����.����d�1�衆�3��MS��G��pU���� �"�籝�Z�Vrb�В\��>ʚT~�W���>�����x-�ߚ�4�bvL� �������y��L�E;����N�v�$+!���)2�`em�G=�mr,KU@~��᳇{���#X�ɽP��,c�׾M1 ��I�p�5n�^���_�-�i]�~���b�ƴ��_D�� L���Ï���ݻ����4ДM���XZ-�t�X� �޲������W��l_t�c��IU6���)5#��	������̷S��R����&L *�F�:�t�ۃ��<��}dt����.q	�ij&�b��5Y�(;��/ץ�<���;.��ٜ�������	5>'���zc��:!�8�=��`*�f�R7G5��k���t��=Z^�0cy!^��Z�0�bz	�쇘��N_3G����`�Y@��=#���w�n�
�C���2hzL�h�7���z�| �z��������~��*���0Xˠ��?��oj�M��T���`�M���v��#����z%VmL���@���sC=��T)��$�͔�Y:gx�T~!���[�������5�ak9�^bh��=s�;�"$��|����.;�'����~�����J:|9D��7ȗ�9���
I4"C��	�$o;CJ]��5gã�JL��yiC%t��K�//l?x�_2ݜ��ݔA5�n�v�a�`K�v�Q�0�����Fa@Rk�z/+�&& V���D�qޘ4��ԓYu�8._�n]���j����AZUE���d&?�ggӆS{����ݒ盢Sؐ:�������j�hp�!�fj�G�f�a�d����P���I�Uw)�l�(�y  �J'�<�J��&U�a�����l���"�Mf2�mk|c�:D�7~ٝ� <��c�D�$!�A��h:���/���yh�i�;>�/��ޗp���P�U�3��P��3�u���`�ku��ѿH��c$�هK�@U�$�#X�5������͘ע��pX��O,p(�l;����Z$rbo5��NwY��߯�P�������B^
0�}	M\�r)`u1�"ʺ�e�-:<).�ߟ��=�Ԋ�[��pT}F�X���&���^�@�
�<��˩��fVʢA*�L4���?\m�Z3_q�EA���R�p�&���h��#]I���z���g�K�8�CǦ��|&@�"�Z�#�c��~�٠� ��3ȯ����� �"ӵG���+�ې��s~��l�Bk-��]�ػ��r�[�=ϴϟ��Q��%q5UDv	�
�����P��G��eb���}�  M��^�@�`�$��>X9�E�Kh0�p���&��FȬ8v�d+�\|�Fj �s�d�������5+���.��K��^V�o�sƭ��"\�X�:[fS��g��Q����<Ɯ�P�N�!,4�a%�湲8%QJJ���;}����V#[8[�~�=�����El���Z:��ҳS��\��bz]+�������ʲd�z��ܶ��h��G�=��3(J�i`��O�0�g_]����	'˪d��g�U!�g�?�C�*B������t� �;F7nj ���VH��tr�D8�g��Oi���,��m�����#:so���I�Y��yu��ٚIc"����uǊ$�r	��풜�kl=�<�����:���l��3�$b�H����� ��hfe�=�=X�J�Gݛ0}4{��n��n�}�vD��B�BȤ�}$s�s��P/�e}���̣[�k���c�쏃�\|��=���j|����\~�`ȏ�/];.�cv�fK��z�ʠ�l��*.�[2|.V��Yc/e������A�¿آ��L�sY�KiW��6>c�;�Ep>��;�a�iT��I��~��5�c6�+F��ƚV��Q�: ࿂�Ιy})�OO_�[ �9\O�M�l�� ���fG��apSڀ��m���le
ňv���A"nZ�,7�����Ȣ�#����E�l)���Q�k�?C@���l.�F)���!�NmhJ�6m�(���{('"���c��ũ��j�ڔ�d#͡B~��َ��\�JS�4�FqR��i���iA��w��\h�MګPjd*���C�:<H�x�V���=c�$i�{�����2U�a��#�	����ANh��Zj�pc_��F�VوO���iVV�H��B��w;��7�����;6ewtr0%�����d� �?��/��?�I<��Ei入X�nL�^�9�^�ïy4U/xn����/`����Gݳ�0T��h[�m��hP��*Ԑ�#[r� ��Pb�te��D�Z&lL��j��QxX���[�R���M���j���ʘ}c0�s:��G%�P	9��%f̑U:�	J�N���P�X�G9�p�؅2��?�lM��m��n�?e ���K	�F�b�:⑓�:%p���,�>��+�c}ȏ-��x��@6���k#N/��Dn��+���v����4��j��m���tb����[�ک�m�z�GT�1�H�4��Axd��}��دZ�f=���e#ǽv�`�8_�&�������ҭjw���Gɂ3aQr��'������_�������aS�|0)F��hJ��Ɇ���g�;��
8k3��g3�`l����|�}i�*�����Vhx��z�sDuR�گ46ő���4(�1�Q}�ڡ�QJ$֩�������fG�� cT�aǭCK�����\20�Y4qҍJ���W�J�ҳ���&�[�����^~
��Ay��e�5B��Ŭ̟�D*��L8�p�����2iQ��7����`��w{�>s���Ro\��q'aHv�t3�qq�W�VJ=�&�<5�������aU�-�!׳��=����Bl6M�h=Y��tx�������*�3�#;dN��*6�3q9����Ԋ����uN"nV0_�&�<j��5��:}{�{.�ev�)���O� ��^�PEBԥ�
Q�_S�;pI9:k�N��%�$��TZw!����p	�w�FN&O���ɐ����X�.�!\"��:4پ�"�M����S4`���$<�'{6�Ӧ��7~N�{�Y��f��M���~?�4�fk�b���].tX��������>����CJ�V��������?�]�&��a��\�H�僳���g������t����!ہYJ��S%�s�]�*f���p%?9�g�e��֧!󅷂ku�BmO����8rbp梉��KS�t�{���� �C/�3V�#�]j_�cy>�z�t��w<�b��Mk����~\�R����I���u������@�CL*o��/ê?�E�E�׼��!��)쐎�I�K��s�I?Oƿ��s��D֌�f7���|4:ɡɤ���4�KX;t����&Ke��.ƨ�F2?)=�j��c:�W3%��5�O�z2A�`D��I���%�w/�8{*��C��@�����+�C�+�{`.;��RF��p;��I�nl�;��ؓ�c����M����L`�S!�7*��-���#-��$��=�5�"��y�-�]B�&Jϸ����^X@%�ϭ:�L����~�sCqղ��*�e:"�@��k��6��W.9*�>0�M��n����금��Bg�[����нu6�6Y��1��@Kr���T�a�AݢR�fv���;F=���*�gW*�e���%��D�Q�K�=*��;�y;��Or#�\yN���Z�ڿ��b����z|�4���D�ES�7���rw��3&`iY�q��9�V���������A�j'�'�꺳c����Xvr���.�)m9-"T�ŗ��N�D�<�4y�]i�����Dj�x��dfJ�b�]�Ӥ��En64iB���5�ž��U 6��!���G�Z�P�=uf��9*Z�̇�b�o&�N�����CЦ/=�3����������8I9dh�qm�C#e�K�9�=�x���%�V�
�Όsn�f���G՗U�M߇�	0��R��R��5���@�*�(I��t75j�
��_F�B	���w�$����dYN/;�d�Ay��4�̵.�_�{j���⤬��^�j[�S��>*����B�:W�����"(#EW�Y�;�kh��NJϗ�cp��}v5;�mf$�9s���`��E�w��,�D:5G�ff*��UJ'`2 &q��nP����Wl�uEƲ���r��܄�P�v��7Z���\U�?��ٟ��u�-^�*z��\��wW}j*?)�l�	.�pw���\f��"��L:ވ�"��ɑ�-錈Q+�$h�n��i�x���B�i��|�'�����L�A�P�������PZ-������%�6Jg��msD���RS^A����x��H���܀PG�\�<f�WY���ܬ�f�MA��n`tM��FZπ�ˊ��� {�E<ntk�JoZ(����/�_7��=�������6k}?��CO�U2�sl��{wtpq�}���5��ƘRLV�j\�z�',�a�#J#�A�����L�S�WF��]��_��q[t�f��B��8�IT8�cV_~�����5�\n�E(@(���9�2���Í@,���{�u����	���(���.��V}������,�^��[��ڇ����W���6ޝ�e5�,`+�r2Ԅ��?sO��Y�|��ۓc!��QY��?R�9M��0�q��s4�ō��l�C�7B��!P>ɫRG��1I_-]M^�TlKd(9Y��"�y�����A晖d�Lz���]^{��B1Q'��|�]w�r
��)�W�|R���ʜj9���_�1�{��B�o����m�5ٻ�X?��P쵣�kg~Q�����L��$1� %Xh	�;|Y�u���^Pq\�ӫ�����͆�vI�Mo�]!���Nf�\��h���3�5��QPE$E
���\R�#z"����o$��>p}tk�,�(�v��̃��xf#��ܼ&��T����|ԏ���{q,�%����fE,����X7=��x�u�K���Q�S|���n��o��NcS0突� �w[�
�K����(��d.��cH�R����c�A�ny�=����j�����G ʢ_�˔RF�/���^�<k��<�1�g�`n�P��#�/���*ٕG�.�D�n�i��q��t|3���n�.�ݦ��lX�`�7r��x5�� ?n��s4�.K]҂�O/�k������Mz^`�w����Q���In��l��k�FžkR-�Ysԅs���]�jdߘ&r�*�s��E�w� ޣ���8V�<C���)��,S�I�NE���{���ᚉ������-��g��=���yE�m��ʂ�w�_�{�FC^E�!u�}޽�N^��.>s��a�n�Y�\ؠ���2�ؗ¯�x�+҄M��g@q�o\�uxgςLR[9��GmZ�E嬻���l7��e��+�v����{��]�

��3u��kڮk� �6���pʹ|�ά�`�������f,Jj?�Ro͂G�4HB�����dԉC�`�F�*a��)�̹�f��\� XN'r� �T��9�[��x��,W�y]u�޾n��Y%���A�i�	Q�hr�j�:�Ͽ��I6�](�?��%�rI�*âWaC�@���?�4���O4� ӈ����U&�+7U n*1�����u��̄�%kX�[D����#.^���̞�������ʛB-5VVi�@2��M8�����A-�P+n�O��7��=�U��kf0QeV�&%2[���\�M��#MC)��$�.�t�[�=d������q'vN���o`�r}'o��R�Tj��g�jA$�mo����ݾuѽiT���0�W�6i�'Z'�Y�FA]�7����租��"~�A�[�C=���8�`���z���|�l)~�>LZP��)��I"yg�^z9,Y}B�)�~o�U�[V\o(hF���E��]^��Y�tT�L*h�c��rwL-��=`ꢦ���5�W]xL��:��/#���@�B�vl�<��Y�c��6��G[�(M��ʊ�茷�l6��]���rP@!�CO�9��8 ���E�>�Dot�� ���Ɓ=O��]��?�hX:��0@�)f�z�bb:�D�d�~.\���0X��UBM�ʃ��`Nś�9��$����ܒ����ޥ���|1Ⱦ�=�#9��@��N���6����x�h�RL��Z�!4O��A���NA
<OH<�Hze������s�E�_���D=�i�b+�V� \�M�󅎫ݿ4�|��uQh�S+9ו^����ED?�8�;���j 0��2�&��f���� �lz6�Z����X���,3�j�3�:�O"d��I�v8��ӾboF_�xݽ���_K�Vҫ���l����\��z(UD��[��@б�1��}v>w��*è[�0Hx�7�}�c[��Z��;[��:���q�0�)�-��_��b�H�錀�ߠkӌwK��.�L�#i�G�Q���3L�+H�n���p��ۨb<#/���3�I�?��ߎ�����������ޝ�࣐�rq~iEȴ�R��K>��q�#LĖݢ~ȡ�(=�����5�+2P���{n��ً� �:������M(�K`��mۢs�PtC+��1�SKJ	Ȍe�
Q���Vͬ����Ց5�"5=&,"(��5ĵ����މ�c�RK�j��g��O!�B����}D�ߞq��s����&�Oy�����	��a�"�T�y� �jB鵠���W[�,���X�
CI�F�[^4d�Z�ҿF�l�#�Y�>��-�����d�����+"���j�7xt��`k05�ֶ��kp�'�#sy]n�\T@�>�,B��S�<��Qt�d6t[ qD���r}���I��ٯ�� -h�V��R&�z ��U�+����:�Tу/�5},ˌ}�� ��+c&ա޽�c�s}�j���YU�)�ǎս�M��O����el�C󼏜��K/���۹c!kA�����(�{'���dW/Wgf5>�s���A^�����������ՠ|�����j�����?HU�];�q���Q�^(>�F��5�04n(O�2�`b����#���x�E�������e�c���ӻ�����Á�����q�����f��H��ךG;�[��%W�t�F�8�hς���I��65�&_U a�1�B�X�r�Y�_��t&�#�)�M�pqNR��#�ć�Lt
������zJС^��d_�k����c���W-n�e, �N��@i�/f��p��$ˁ[�%���B#殮����?�}d.��F��w� �;]��,���A�j츦��L�.>���Q�Q��ǣ���z3EJ���O�a��*��R��
ui�X�NV��I�6<��!��m1rX�ݶ5C�o"ʠ�h��y��Kܦ�?Ɠ��H+_�-N.�%W�[�y5���a9h6��/���hIf	���㪉{��3v�ʉ@�҄����\�6�r2����@)������:�������%���x�uW�.�)9/�^v���>{\��L!V�+Jo�lp�^�v֝��=n�	�al�πOq$ҍ�AN �\��)i5���f�w`��ԱBA&�~�-��4ܵ�$o���u �h�c��{x��>�p�Fl�ر�V��>i$0�6X�����Ijȹ�0�Ua{EuǉŘ�V����_�E��0�9�[W%3II�B���<�=�5��fW�����8��c0���1�'9��Ϳ�N�}�@u�}���ı��?>��Y�z"Y����P����Ѿ��������	��+�� 6�jT:ru|$Z��N����yGk�Jd�t��#^l-K��	�=d'�?�
����>_�)��2o��]���y�j  S��P�_���O������谪���TƆ�{Rc��uـ%����?������Ӛ(���t5����}^��(:�����.�~>(a��B0�зt�g|~�g��=���,�.�+E�=��
B�y�[�F�,�mT[/qi�Z�jD��l�M��5�'bS��T��:��D�D��Q8pc����������kg<ST�~��Ǿt�gi�P���yD�
)�bVУ�;#�� �1��ԃ�{�w�%ֶ�As�'�q8i,�6wVB*n�pΆ�V!R��V=���ȕ'(B@��d��1����]Լ��F�s#U[o�6�r,�U�/�����oP|�Sd�R��U��#�/���p�ݢ) ;F��/��pP<Y��NHCGi���v�(�'ֺ�qiӼ"*���.,4������i�D��V`@� |���Zk����Ə�I!4�)˕�c+�k\v��۱��q8��o�I�{>hM��Ċ�6Mj|>gL�y�6�G&����EՅ��UB�ڤ�{g<�$nf*��ϵ�<����Z�!�[:��՚Ǐ��"�!1�W(k^xk�Eş!���؉��ҏ�!E��=�%XCQ�ù#�:6͆]���a	�G2�ݐeg}��D��Q����)~��#�[�N�'O�#�9�

v���8���NkY�l�ފ3M�����1x�Ҹ�A�csT�F$ȶS����mŜ�d�,�!��@M�07��y�ƒ(��c#'��D�`֬�S�lB������:Pjv����hv��,q�ɂ�W�K�wJ��U�9��ė�g����i��=���&���z��}$��߯H�X�`U�뉖�,�]�!�]X��|��R�L��p�6	���k���{jw�"�.�`�?���Yœ<9��G
��c7��+�';���*�6khDS�@�7-8�vㅶ&c��V����;cM�a����C�zf3��Q2�T�:-����د�Qu���j���8�d����� �����dȇ�"0)?� @Vm߾cZp��(�K��]���+��E:��JY\��4t��xK.�ާ?�_�o-�d�h(���;-�~��Hês�����է�"�'�N���b�h[(/�Ƽu��	��#��}!<�+�EQ�R��0Ǧ��!E�x�f厞B5��:��Ι%�J��yN������`��6D��oI�K���.�E"�!�1���ƕ�L~#/�2� �l���+ǩ�׳�$f�I��xKKȗ�i��ʰ��a���� �n�Y�ތEz���Z^1Kj�
lÞ���k����ԆE��u�1���j����]�?��m�� ��r��Sү@�;�!b����Z�,�Y�~c�u��!A��(-@�����6���G$��9|�N�"gEO#��>>ԁ`w�ވ���,/�Y��}�4.7������<7��h��m4�U����e�%�&��8�4�	�m�����S���]����2ՏᡋWh(�:�)�'q���6,6�"����w���jGe:o1�'|��9�Ndn鷵�Rd�� ��=�;�RF׎�n��%�< Q��?'z��&r��#��2�ߣ\J��\\�z�%��>yÇ�_6��l�Nb��7������H�i�)z|�n���=}���6�<jI��zߡ?�7�R5�׶�S��V��-�����*x/�������N���:/�LY	Sty-P��5"�3=f�oek3K�6��YE9��F�)B�dЬby;���6��ò�����ȣt� ��o&�6xdm��8��8Σ�z�� z��ҝ����G��D���x4���\�kꂵ��r�d��Y뿕R��I��Nr�U8)@���e<^�a��wA��?�GH.���oHc�D%�UP'<Yo���@�93�C�2�s��x��,k�{���ؚ��d��i��uԹn�M�g��z��]��_#�]�}I�?c�B(��UJd��	�����s�R�1��i}�6��q�w��,l,�X[�>�S��M+\�絛&����k2Rw�j�O�L).V�H\�v_�%�-s~��<�5�Ӹ��؝��< a�����ߤqO�l��V��V�q�ynqO`T�P@+8�i���G���),�w,<,#8�p��\"v�?Gr�%ъNyh�|=����}&o�$�����q�ۨn�Kh� ��Bbx֓8o�ܕM]M��.5v�7/b�mw#��w��ާE����7@�!rϸ�z����S1�-�38����GV���|H˂���(�p�)\���'�@٬liGn��f�ച��=�����/Ǟ�{��#�a%4��s-A�>$�=�Yh�S��(�qQ�M��\�����a���[`�Z[��S�3H��:��ǚS$*f��XF�Er�yǛ߰v��HW"ۓ�����cA&���4e�m��qQkc�eBKTcO�Bf��Kf�������Hę�ۣyWVf�&�5_�VA) J<u�M�a@Մ���9yx0">l�>f�{0z����{�O/�?jU��X�~l���p;���FЬpʯ�0
��'��_B_�Ęe��@f�Lu���}Bd��,H�헍"muc� s]�j�2� \�5�>	7��P�t�y���U��wI5�xލ�0+RN����9�i����P[�T��`����;���v$<d�9˕{��nS��<�^�١I����,�˒��?��"�;U����$��]���Rba.QG�aX��P$��d���M�X�|�E��&B�%+���ֆ������ނ�!t�-�y�b���6M=��"{����$����$c�p&C�=@�*�0��I�V���E6�.� zoeJ��^���F��9���[#th�_(R��.8 �g�E�=p̏?��^ڄw�x�k�@�Lv�/	��O��u��2��YD�hG�-�<C�(d���=����C����S��mSZ������&4+�A��[8�.�#��N��jp��;�ð4:󵑶�|��"]A&2�������bej	{��R�cb���N$ŵ��M�0��텷>�	|G5f�;����%���^�K�Z�V��1?4?�B9�?�a<\����rd��	�f02���}~�a�Z<���$�h!��s���/1�<:�>��*��$I&%Hd]���%>|j$��Ǜ�&4��Ѳ]�OR+���bc�v���@ �X~¼(L�s3�>Re+ �iM*�[�=�Z�2�����ơ���Q����К�~��n�ӈs�I��Sپ� `�D����9���f<ubp�2a�5��B��X�����j-�*�5���X��J������I53���9�[����fT�r|�f0���	{��<\7f)lC1���*]Eũ���T�<o��Ϝg�R�Z�X��TD�s�G0�d��r,S��f���.��-=�\�#~�W�TҞL�fZ�cXL�mG�̄į��zA��g���-���B�W
�����}-6����[3�����W�a��<
�*�vS�����P;F%犐MFa�L�*E�󬙭�kWoj$����9Laf�^`��	sX�X�)?��\�a2���6�/��K�{�ޱX�(�/Q��C��%<%����c�:��o��o�c�hE6�����_v]2��x�ം���'�&ec�������FXM�+B;���,JGD^!Q�+�L� ��zd�U�Mt]���fLF6��5"�L#�yl�mbK�J�b����Kcr��N��;���Ζd�v;�@�����\}bT��$!yF��n�=%di�E�u9n���-�ՠ	V��]>�K�����fq�����&膸Tv��i�̤lG��R����fg��}�q����B�Bo 1�_?<�(�"��.��>+����۸���o{L�Y�H$jݱ�!��V@�%�b�"bF����y��� ���'�)�!���F�>
�z؅5�C�4u��LLs�8���x5�V��1
��\�oV�}B��C����z��1n��ٌQ��S���vs���%w���Q];�2!��E��dIU��ηV������7�m���`ȱY$R��cT$7����P���n;�^"[�bU�ݎ�K��s�iFa� ����u��� ��RR��u�.��M$���N*=��Ɉİ/�+����S�3a���L��R��^����Y�O�F��]�-[�0þ�[�cD�z=�d������R���SS����$	N~Ἆ�T��=wP�6tF�T�qUi[�CjdRߗdS���������֘@~�f������`L�o�ϧ��];�4��aU�2���|�E;mBE�n���\�`�B
>�I�6��z}��C�ja��ǅH�f�ۡ���J�*x��4�L������j����*�J��
�=��PO&�x{7�ޢ�#�R=�ƝM� ��X��C���q]>k"�R�c1�)TPg�=2s�;��`��+xF��������r���X=oJ8*g�v���ݣ4�B���Sj��F#���r���b=F���KH�eklv�~vy^�)�e����~�/�ߧ��=Q����o�Į~�'.�Fi�Ce��At뼋#J8_�:�kL?Vꍋ��������n}������z�@����Ⳬ��o�r��'T.��۹��j�F�����?�Ƙ���Mxt�`�O+�L;����4��������߆ᆓ�`@�H�H�DAL̽�"�y�nm�#�<*�>����d��" ����;ԅ6=`J�^p	ܔޣ��I�3}77�UJٱr=&P�����_78��!bpP;9��:�@�2�U�
�R�di�Q6��>���ی��^�6��Jp��R��z�]�3��O��a`Ԟ�h�q`eF�U :47��5�X̾�ƫ���y�IA�Y	�T�v�q,aP��M�0����Hܯ��@�#_SE�R�Ȉ\B�K�O���z���-dr�g��1�fb��Q��}7��b=�V�S�=���zD��RP|���k��7�a6�FL��0ܢ"8ݟݭ�Q�n�p��ov�e;�z����~:�X�A�O��"^+/uZ�[�{�.j@+ds���x�P�y����`�=��'��g �� t��N�ܤ���m�����m@���m�o��#��{sw&H�ş�����|�0ڒӄ�ڮ͊���}�h�.���HD��WN;��ʽ�J�'nvכ��ox|~?�׷!�R�D/ֲ@%�XS�Z��Pw�4 �
���HE���|�g�~�����Dg��S���]�Hܚ7������,���t��**l��$_���e�FI�9��I���{f�\�L6��y�R��>��E$0�r���5
0�2q�� I^u�i�2�c�{؟��<6��� �K <8�Y��$1�"��Ke��Ƿ��>Gİ�"���K�H��8�}��>F~B�k�,�-ļ�Jl�AO�����<r[���2B��-�[��湐J|�� �z.g�P�7���C���~�@!<����ƚR���K�&�