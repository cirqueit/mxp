`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17984)
`protect data_block
hokRqtyXri7z/ICrWp5deBZxyFKyvOs+JHXhpaU1p8vzqQvuUU7I3TDn26C5AW314zgRf/QBkemy
a3nA71p8ClWhmIrFiqjBOLZFev1Rwq8RB2+d1JMYGd87HRZx4w5bZrO8QZLvmv5OXE4vzs8lq9DW
oXLJRQ3MXcqunnFdXZAZOtE6Qe8UcJ3+bsA01BvxHs92HzbEwyiJM3HRIBcVPK9389Zq1/jUZWW6
oCl130SWsIaP1fzVeWJgq+G2xsaOsR/BVHr/wSYH+KJcTMvMc4bqU9Nf/OiTYnMJWbzv1B7bds1r
SThWZQ65B4Ope8oDAgsavyig2tDqSmBEpyJwyy1pp96SmqYFP5fD1JOxrDKqM3AQ87z8BJaR82ov
hLpGiXMNjIcWGZ/8lKl7pkS7SySk6D8yDS6r8EkMyCbn3faxe5EIzDaIpcTS0umcK45uHiyZLGuV
fswE/M9i8bZ+KC/pXxcmaIrD6dyggkboPBtECP5Ky9SOdnD70BtGaLUCCQsJkwMJ+kTdcCs478Ib
60aRFrgWBcGYU3Miy4DojC034SonQ6KuyP87tOsivu6RHjJ7/cUqs7oUcVqFNikLjec54qAtCdnv
+uEVfg3M4cdmt07VS0lKBt2ZsO9gNUn4mm5GHdFYF8YDPx1idlMw45ugZsCHKvftoHTK327tNYM5
nErRva2YiY5nMnizEP+9Yme4CHCAe7V1yNo3bDA5PgJQ5pku6KbBRZ6y1bLzLy5c3laiqYjD/9Ap
8mzJguYDMldfXhgfigVTpEBGhE9QSQD9C+WRMXMU+6erG1fa6eO8sbwHMk0KStojK4/fUfW8Owvl
q93pQNUASZAalppjH6vOm/mM2y+6rEVCdEBbnrpicpni982zG55BOQNbs3K28SWqq//8+TS9Ddwx
NCP0Dja2Rxs1J0gbqWVTGO0Mn2eZba43fUXFvFgapsYvrFYIgPiHSGYw2aEWIwyQbB/Qq5aS1vyF
a6AohpT/Few5mkkrq0KOFZTNnc/zgQooVwTCYLrAGzNhJQraBvp8UZUne+Xn4u/nhj0FxNBOMxq0
fJI7xi2eLQ7d5B5bpGs2w0xERU19X371Ycip5Z1bufZfa7qh2YMHeNHL11pzXecmfTAGTfruUQBb
CTq3ADIjVHXl5F+BIrvBKdJqTl/3m1xQnafq3DcbwFGMX1TxU6+cmT0cGljaWXPY1WwRlpK9/C6p
OBvsJxpPCB86F6hHaNAKzDGy/RZUzs7iKMLVwO7ZiR0opT1gCGeuec5hElMp+bgpZ3Xx+8yN8ps6
V6krGtYDs8dhURTD39NKajVsUWAeKXrj84FDsu2EeLAsDh4L+5ZNRNzil8vycUisoO+eWiTlr3xV
3i/dURD5agczgVkxBse7NVT4jF1o1m8V8Jr18VKAAo3ac4UVjc6SN3gC3xMu+ykW+T4Lpzte22kH
Z0iaCKCyKYoCCQMvyBExuGTHo4+lH0F6/p1TKGC53wpRC0kvqXJRIQS0iK6UnUWNSrxUNqxSkW10
n2E3e1n2XGY8LgRQGD1R+uDkwefiZO8pFm4qDbvLd/dCbOdO0sX9qKQH21gabVqWpF2lIvTl1VI7
khKOvATz5Px+yGXDJWIJmt1KKJU4DtF3D83B4PSZM8RP3GZDL32oB3XTtWWblxCpX5qH1JsSLKEa
dR6vcEfamz/Qf3uJ2dwyklUIaywj3IilGa2JdZIwwjOPjrSU6Sg2kI0ncqVhVBvZB3WNdHe8CbJO
SxPFBM8NQjYHkWfcJyfvdDz+F4hMgj23geq3Kc7PK7N0KDGXCjc2xYPUUIQTYbNTZsVZGn6jISA6
YIcUJ4PfN+hbDPkM6HMgUzxSHryD29ec2/LesRDD5BRZwpnnZZKm1UZbfdaK3PzoPvXj9CjJT3XN
SF8i/vBabIvEg5N9zWhbouphKEqYqeSRCpVOrWGQP7VwVvP9IvJDRS7uvstdqWSWKy3oPPGV+8l/
pbkXhpfbTfsOdDQY7uQ2ojSOCBxropfVh/ZWHA0+cIspUgsJP5t50m6W+shMU3ZWch/9vDB52RnC
0JLtXk87EHMcSZJSmeK0xi6OWhEzJGAhKyt1mepFY/FZ9CiDjwc202jQPFcsLS8nkW9/3qjoCQhE
OP2QgOUiF8Hm9jIRqNCRSaeozItiKD5JIJRLr0G5NvJTr+rDliuyhhC5WmMv7F+2A/LdQGT6FC8a
SO+08A3IVqqnZBlY9oTadpJJJgNkDj16em/tfITC2EOjiWgLTONljtKEqlSi3PcQzS+g9DcB4Un9
KnfbU5ucHtAHHkdMaEpD9PD2zjY+DU2raMima4VBpxyPYonIQn0QHugj4iFD1tcO5w3wfLg2+6yz
AdzV3XxhqHzX9SJrnvGFo37snT2GztJ/RLJDE5KgzXZN5r6gTQ/5ETEBqudIHaO3HkGCym91W6G2
prN6cEvPUjFvn+DGvW0ZiaGCVXNPsfVByouHBYK9rL6QTPSIZrCDYUd8Ps73Sddcyz9kQJew7j9X
sknP6dQFjPqbafJXKS/VRIPFO9EFifg8XTVw8PSTYk7zTLtRUWCITLEAl0mldY181DcIh+AxuDzc
Q2pjTsONrSRl/H81kqsWOEaE2ahRYWn3bYpAo8h/iUsvzfNFbv+ZLBq3IRsq3v3Sydk2EVdR46VD
KaVrFf+Stis4GooMrZCVx9K9j7+UHCDPtZerUaiEzocA+h7W2kty2cWfBBNJEuMiLivvnrc+XxAH
3+TwyVCyispBKSEKVkxLWMU4RkuaP15kLM8Re66gXE6+vqDXrVxeH464/dBUUKsyOOurIBWjibbH
7U8dAmhQC5AENtLbHwPYSsuXzWRcmF9E1XZYWppwftUqzgo02baKyYC7/j9kisbXLXUwoUwnVcDF
uT/hBjCTEfMp8hEB1ldk4Lnp0muV9AWCL9uLFabH8JE0EbhY8Ul4ZoxzZluO1pZRNDmFTjtZEvQP
+U+o+8Kw+Cl8vMmR8MNOf7sbfF9OqSgJC7eUs7kQunx+WHnIW9qI1nbhHyE3x994O9drecM3HQnw
zUuOSy/JLGUOQt6bs64eB9yWvs8Wo5cUZfNe/DJ9McbZk7ZhT8myjyu91unCfEPbHthtnUBNZ1cu
5APcEJJf573ESd0g8OwRLN+RYu3ljnuVQuxus6oBOag2O64CmgTG7yijH7YKRdLTO2/tGdOQVAFg
x45K6ik7HAwE75fsLC7lkVdppPcW0BQ0eP5c4cVz+j9SlMgdRohUTYQ+58C6kDbjAERn0r0NQB4x
1waZLtZOeIrruB/xHvZA1iORpHFOJH/7/F7TrszcdLJyJIKmXPwwcsdIDTydmGnj7++hhlg56cps
NPR/qcIJwGeXYVP266pvbA/x66DBw6eL6JoCbkXR+aZ+wXsDCQ+zwYhXCmAjgqORLvz4SVnT3O3p
U2ochCEa362sWJ2NL3TEMNs0b7f/XWSlgeXjBokhLM6byTBYlfhA8QeI6w8gN+C5Pqg2FNoU6RVE
jKFB9SHkiszA8iJQs33dXH0U4BPaif+PSaoXpryGm28gDe+WPvEM3ZJSP0aqURR2juSVgHNb6ViW
FhrkhqceRoPE1h5Vv6team5H4BnTv9ZQg+2QNwzaM/LdYeO3mxrxY/8LtFYMpDysu2sqWD7LBStI
IibKCN3Ql4zK4mysXH8Jre7Dp8WmIYvvm3IfSbnrjYNJKUUPa9oVYI+6bcZVRr6JNja+hPf9kUmT
b5GwJQoj7m80/uZFBmWFp863YQOAuWfRpQXhGxi+LNEMi9mBDMs/+td4SwRkpBUKyU2J8JrI6bXk
s99HYrupuAOZ4rCO0VcZpYHh45+gTjXBnC91iMde0qwbxchaAa7IDpxLn9M+iloLcfMcHR0fpvIX
AVVSOdPtdanbNSDFuUhnDwmxhn6ZRGYzsazbOxHT5dIm+JbMh+2Pky9dpPAcx61m1HHP7h9E43P+
B9uoC21p9x59JQ/f0FBaKCC5eE92+N6HjVZ4FW2UEMBVHYz9ORZPZQk0YZyE/L8tPD98AdiDbkaR
CYkotfbPXVYSYLCvNeh7ezCHThqglkWiiYEiMjch7fGrgm6K7/IpbUSEYe1lY7jRkwR0ummg4Vrw
Zwf0qoHaxdIeMRX15cu0AtNc7GuDkh/uQLPHTvrxLigUGFN7l7FU8bsG3WKYGLFzIha/Pc+AAHqq
CyIB2KquWxK6ZqRtf5JTh6M+XWUaz2R82Rz3kq4QRWGkptOfnLeI1JGAJq9XZLJLCMrmQlFSBJfm
iByTa7aG8DXf1lvjOADKmfldGSlUYQBceXvSXLvB1mIla3/qTD0E0IKwzl3dVMBSzu/6PnIiWQco
bLMP50oXYQEbUnfbMioagH6rKuC/B/ZcpoYvrhbIaG0IJ+jQUGL9cpsjKwKPX66Mlr4bq+s74qh7
2+Z8Rq7pkP2DiSRHGvufXlmSsAeEsKahePdvgPZVVbn7dt9XC1aWraVyMvSKdp6XO6xDrlj798kK
/iEdj+euoovEwZxwAD4Z2HuoXTCtrp0B9T3/quhaPlwALeUPD/Tu4hqVOioOHXlkggHBnoFPbLa+
8Tn5NYgHtdSPu81HP4WdvGfvXo6O13kiOJWwHtW/JNFeHUk83BBWNvi8BMDqqIq5F6u4lbxANSMQ
2bNqwTbF0Kq1vspE1i6uGipnu4cqvDt0OVffbnTeldYgKVt+Smhi0V3McB0rQKTEbd04kYT4nHV9
iEhmzNlUlbhLjAP+WdY6r7XLNAK8b+KXucY8F6cpWBFLFaH+zcbe25oRuln2nI3bJbqk7SntUH8u
m+UVqHCdIK8td4jXFzifWXEHZWunWn7PfNHbaQJ3N7G4M3YhMF4Is/g2JtdedV32PEjmR71X+avJ
qAoFXM82Sv4KTrK7niBLxy33QoFJdX9NubtSPzSwS4dP6mTUUkHp5xRztYSWKaNfkEM5qGCdltsg
4neuFgpm1UWKINagTzsbxhU69xSfr3+5wGjwAljiUxztid6Bph9OJc/rjVY7FdFAPpJqPKEYWc9g
k+UKAf7l3GGR4FRmQWvdf2TFGenbGOquerm9XnWfOarNPju83CGpPM4nwiRpBg6fDRi8acIeAjhb
PwbyJdNqteZjP5bMvwicbKOBZDIWQ78hr+dKiQaNWmRWftFtch9p/EbIvPQSGjxv6K3IOWm2l5xz
LmlNUDY+YJsHXyaJIs9f80qeO6U6yhISDFZ5KJe0OhVIl28C8+XHNa2Y5QSvBPdRx8JcCRxT4X27
Y/+rZzjdYh6c2IUMSDc0I1XC6fxlTj+89rKTacmfY67xfS1/Z3KTZhiTLLbPPpdzf7XDpqG2oi0D
SjXUrJ4GMVt6z204ansIT8Lw8QIf7qs/szrHBWFvJsmVqs68x9VjvyxW+jmcmIFkolwxZpVrmJjG
HnUVglfwt2FB+F9diWklUJDS0cSTkHVZv95DFTWNIFl0naH9ubMw96+9DRq/JEwgW1jn7pwsCQ0o
FPYp/uab2y8WPQkpkxCLJASMZ0uMLiG1LfGBcGA5ukGXyEPuAzoMwIpcXc+9fg1ysz3ePFiyfRwS
NmxIoa7A3h8vlmTvDkFpfMgM8KaJliFHJ1XKs9NzGmpWD1s23Motiti/ItbarSfZQYgLRwnVG+9/
HRWNmj0KluZW4yZQ1wx3OQ5fJD2osxmKS7ULrWwtyX729qFJf1O0aXBIY7VNXuTv8vNSimbVo9Rs
shGD4YFQQO2aQr3019IBR8NcYtPumGCw7U4TZUUoLF9quIMUWejhuR4XfXqFMVud+pRt3s1a6/eH
oPepWqV1d3jA4reWg21x3+klH+wlrhrvMDjQJUDotPggPRL5Mv86gCNVU8rDjCIrnqEPI6GCi120
xJNH6ICYIqxRF6cfK0wlCCSwytZeb37+o/VcR+kKJnByB4tnGohxDzwxy+a/zP1RgIAh3adcplDE
6kcISDKw6BPb8HnAUSqUbSMBRv9hF0zaN9eMeNxwCsHSkPU9w0/xNsjeBvmxRSJSCz/11LbnVe11
8yei7HlqUC7fkpLBF0o/6EZSDaXrk51kjQNQk4/RJ8zcb2JrYA5G8uRnLxBA6aCIgu1A4GauoykR
cRs7MgsiabGe9ozuXPpLcuUSjO4G8JHF5+Risihke10voeblcZM0LYPtpZnGV/zWlC0AqYEWE5C5
mHMb2K/nIenkKMD6xHfE/GJTqkpOLQ76VR+zcKPlL0Op8QSbHggnf+TO4fg4q+Xe1tn+QYpLrC8b
WILy1Yu+py+2ftmCeSUHV+UYnnaEXJ69o5a+CLVLLAJT+NDMN7/v0Bn/ULMo/6plH6jz5zlvT/hz
Wj6xjT1AiaXs8v1QexJ9T/mCKc2RJFjd7HqpFyf5FJ0iwrhC18DY+3mzU3uWg/j/gD65gUF/EAEp
8HYPFAsXOZ3wOWs44B4I4aqojNzP2MvMIfX7LYeLS8WEEtbqjd7TvC8N+JsLiOvJhbENHhUbwxns
0tqpQoTX+2amzu4bwM2W9aE05e1dm+BGqyGwgWt3j0cLuOZ75Agg90515w9Mb786xKMpvbK9KBQv
8MDoBjjJCZSCqyoMwF5H1+GhQ2KaI86iNI5BG19LTHFuseKFA0HyeywXcEikz9dJP4u+kXv8E1aN
V8hNfnH1lzVAyhwXciwa8DAAvgs3w/qKX/frOSdpi2+f8gfjcqTH7BhpG6npx9vAUMmSi/iyGR7B
wK59YXPY+nB5TKHLhilLj4FDEIiEFxO7bkZH7pVvQicX6MdYRyRLJJ96pvrYU2gxxQI81G8tTDWD
s5uVDvceEZ8njPtoG8VUF3i4N5AiR+yrNcM7JOimNea5kKF8aBqz/HLU9zLqN1PBWZL6B8SpnBTh
y15V0T2/0x0PdOdSZtkjEja6lSFDEYw3fx72HrKwfGwPU3MIKO2ifuY7Fqx+dBExUHvreYpmLMZ4
rua05eNAoMjMp9X50Y2+YzwQJwUa5FeyGhyqr9iLeBPkXlReiFngr3rhpwu5pK5mcrRga6kU7ZWU
kr0FK+6B1L/nqf0D09VmTH8/NzK35rtZELtrZwQr27GSBx3W+MowdQdEtUl/C5WJuG26Sh89vWLz
eyYAnj2vxpCkPivYPldH5+8937zqGFM5Yb8eI6XeCY1Mw8yYLzTOyfcSmTW3LbJgL7+PjDN1/TjP
/sDSUM7oVMBlE1Ph8vRAN/yNxW82MtFAVkzSTnB4ssgEqPVuF0v6E9m+ZduH4AlGIBTV8znPzFsq
avmaDsSZrHD0rAx1FY5fmobO9lgrIeqEoO/X/jCds1D1PyhwNLsDNh24OXPfUtUIOs0THdQpaFJ4
vI1A01LyTYKi5k6KH1UHHPozwYVLgU8VcKIij11fFHq8kfx0hW/sHzevo8JumCP/fdUxHc2bIpNY
jmoyIZwTjW+z1LZpGSoU1F6Euajtl08P6+JashaCPEDh9naxPV1111AgC4WgPMoLUkj0+AnOC7VV
e2uYa/J+HG+OKi93QKCu5NnRjc8v5+O/QQp46SNLSEug49vorNW/JV6H+WQVPIm0ZQldGZkM1E2D
UDgy+h2C1/rp8uNi4x0pGS+SlXJxaLsfcY0m+e81bA3d47OUF/XyEEh6h2d2rHUqLxRcNGUl2ebh
z1u0bEoeX3S21NKUo0pzW27gV9e4XzZDzx66veAORr6KxTsviBiCBQGy44vK/eYLTOAfQWmSlRbi
l4Te3zmnbAu0RfkTwpB+mBGc66kRs+xaJo7+5wf25dsFA/lokBnFE3mZ0JwLncXVzkD0IxJurZiQ
FsMCWU7F+hjzs96VZZ2XpLt+r3kuP9Q94ziq/nxmpMRSevKf0O6uUBIUPCBa/cQK3TGgmkial/ed
JRx4HcH8s5+EJ/abrkMbQPzJISV4Wj1wX/2uaiAZt847hQH0Fo7sPrRrBuNcgfL+Q6Ycb1KAzOlq
vjekVydsmH3HLIKhURgiM8j1zJEqECpcAcuETA/rkiH9TbhBZvFBXLCrSrWzWwAeQe8hGm5GR5Kw
9qDmgy98RNesI6E6ugGfkyf0stPR0c33rL3Rcm8QnhAeDC+ILxKHbc4HuGUx5ejmetMk0eYDTb6w
+KLJ/C1wzNstcmA5lPE80kwU0YJfiPfh2enaDSN/PFUfNrW2TplosCgqz9lsJ7RzqNNaliCP1vb1
krCHITpXIXdge7PcKrMFptq4e3gJ1QlNsNczeXB9Gm3ZycLEq2flcjv8DMQs1lCDdX1Ow+GkX1Q0
D3tZnY0AGqtjWjK1yWtG2D35lyCdbKkt/HFJwhaKINhP9Om3iPx6GYVZqJnc2PHkWXX579V0CkCg
QHKQq0SWeGPhQEQoGr08sXTcQ+sYZcKttjCPKNVHKl4drgKVywqrO+JdS+uLMqLO4QW4osULkGix
dIQ0QTBTnCWPUco88+3ukgaOn7bNDtgV4hgqKqY4qIsN/YQSJV/InlI7T+xEL1QTuTP7MkaKHcvW
CtyEFvyR75hXj9Bye+OOaiSe8jzQQt2KnPZQ0jr7CuXUyD+Od4kmiBEAMOSFhPAjZZ3W3MV2JnP4
6E6k6Fn11w2JdJpgu4eZQwhgX+KQAP0M2bWm+FLpEDJpOEZ7sG8LGgevrFosJ4SXMEX07Bjj6u/m
beBitAMb8UGFxkKJ4PWoBgYYFewMqV2UIxbf6Z3B5jJrJJrQs9iOphq7OK8s5xHppLEtyxqLxjnm
ou0Tbs9uAheSiyPbiBPwDEG/kCqxUG+RsRNlS5OMb+LWctamp1HF3EjdKmu6JtHox1oKd+r/hok5
YoirCeDUti3Y7/D6tCQdFtIkBZrsECxnsKRmJch65eC3gcjQX3VrFAGYarbp7Vx7HUf/uEVUTnoB
AgiYM27u2hjK26bJfQIfxE+luzIUuuUVTYj1BBlRSEQbOpYo5buLvtGfWSrlmVojVhnpSCFXyhYI
jTTJDSBZbaKovmkuNUPxqhRd7552d1rwMuNbtaSqxc0J37oQn7e+9cL6bFlOXTQ9QKdzbVO2TUcZ
3SG3fWEAUS4RKhjceioEdgQVLJzn6e9ma2liMEVdEY4YJfKRS90I6+BecJqXP1t0qTcqR8SR/IZV
n16QS1V6KPlAl0CWIw/0auT6NBNe+LAlelU1Y1/0y3nShrGZoPOaIRdbgnLhi1wi9eTDU5JN4kpa
8er2ZOtEWGVAPrMouJNALsLtk6TvRA0ynp2+srIlF0r2sCgL/IaPPmV4k9bTAo2sp0ljXuW04nT6
sKEpNhgvtS4gp1o2duoXFDv01zSI0bpX913liB8iPDAnQUa/486eBs/d31eI8k6/bPhKK42omce4
oObDulZsjtvGN3UDDY3iPiAvjWV8UzOGQIMYTfQeN1HX7pkUQBGhjKwr7PudOTVw3d1631pZ2aaG
iIjarb2NrzVlAq6FtUIx8AFs2o9sRuH+NFyNtZpAxqK1MC+ES1G95WJff9WN1uYh3izXbgwC93ws
tgBSDyB1QBcUlke51/De/aCCU+LRCSJmxzbJHsD9mHSK/0q4S/oH7nnKZuEY0E0C417GXOKt0txI
FytbfcN7hyPZl9aWG11qpUsUgDpLzw/hy9R9fVzkoK/o72q8ShmHIeVWRFkgwrWn9K2VlDGfKque
tWCQCvzWhjcZuAxTRqPWgpPmm3qdiQDZGr3QxTSS1Z0WehrV7yblgA9+x4mtdlGqNSFB4TPbFZDD
AldUpt+xT8bfzt/Jkobz+QNYS0YKDbmHulizOoQ7fhS9y0J6FwN+QHcNK9dVLn1VxRlBnEciOvlf
HzPLpeHIe2B1wJ+OcEet+RqvgpM11LYR5OvV17UGut6vmTXCDpLwTZgEsYJ/G4qGU4fohHWNNYeT
MpWBolFiEt6t38Je9plIHomJpUe7bH/85nxxx6gPO9t6B/IYdKMlhGgE1jk26cwFRIJBBNfjDeqV
LNJ/HoK2zPXef+F9qhK5uQRbGaXmqinEzQGNCIDtf9DlobHx3kHOTfwUZyLUDfqLY6LLpyg0dl2C
BkApFL/BGtd+mtE8WWifxINKFGzTyBnG1RJet/VU3HEGwIy5cbS33z2Yda/AWc+82ttiM3IMA60c
wIJETAapNnT0XjVjViIL4yBkb4T0w30mNf4UccUMWdMi6KB46lFGrF2V6aT10xoDtSmmCIr7kpPm
9IR0yvIKjCAKOcpwIPhwgZG5vGkdpwCWretzqIn6BuZHMl62DmKeStA3nfeMK8jTyts7bSmAw17A
3h8dzvjKwVJBiWX9UzmBb3X9MVPVGZw4COYPuzpyH5LMuyTPC8iANPYfU0ZWZRWjjCvUib0jN9O/
3JpNhDqVe4rRqJSyRLimdCU7KM73cQ80SPuudXa4QLDDTZBjMSuGgjsQSCPQlP/qOnj6+tsmg21x
soLvuWe67bUXvHoOzjCFxYkYxTlt/q5u3W+w42l9KYow0ygyuos/BkdeBBeY01BJRey6451VFDBa
09NoPIPVH+FarMHrUAsqxhdl13qme+4/oB3tf9nlOV/oEuRNKP5EvJ+QGekBG40et31jUeleBiNN
tnJxTB/EH8ltVeeNnFWOIa5PI4/C4o1WJ/4p1TUzxYsZ7IlIGKMlodumwWDdUzjJLBhpV940AOJe
hauwk72H0r7fXTR8sdnXPM/dM9fyliFy4PYiNNja5pODzpJlCi61/pP3eTNXSbMWPATAB8xkf9hU
ccd783XuKnl8/EvjVOiYRDUua18uDp0mkW5eOqfwFm+9qebFxMzrHQZSYaDcYwisINU1GupUvXdN
53diuJW/8a1ig0nY/Ekxz97wfL4aNXHYTrwLe2/0Opul+ubv2KE3wHO+y19mFDD+zc/YfJjuJih3
/4LfocN1e0WsDJn3lOWwMpSRTxueBkbz9JJNBS5an8YeLAj1oVizxd/F1tY624+Zapr65P7gUExV
g6wjF2AjHW0j54UHGRMDvp2p5QjvkGgAABnMp4MvJu9LjjrsoQrJLLTSzdhsU4g5Z7y/uLs2/gjK
cFNgC3+B2AJ62nH4wb3Q16oQgSf5S5B6xAuLVpjssqvs9FiWBMPpwqXL2X0o3bQaT2HTU55Alh7J
y0WEQqSJfXCRTxkFrLJyXHbxp1cnWXjhnne6nVJ/UWR0zrep+3ASpujgvZWqmhY4ysdImJhDkqLR
s8T968XigpL9l/jtkMJtO3kSVzp3XbiEINf8YG9h34KqkfnEkXdL0r4+f7QCCh9a7JROo4OqzFqF
87snYrKMwx1Qvp5h82+biJJ5v+hksG22jU2YREitc38m8XDrlkzKVx7wqHOqEUFyIQ8lwA+SPHzf
O+YwZxdTTg1RuNCzdpidC9x6v1HBMUz2ifjhi8G2ff5ERXJxKHtxc2ST/lwjikKv22EYh2Ok/w2C
nLfVRPSTOG/upfjoZ37H7gLsfC4LZsE//QN1Vqcsya9s6mqIsstt20o/QKBj1LjofOMEJiv4kNnO
Yj6gEHZ4z4YlJg4jmz4WyQ3ebkxqYpikEkBkeL3gC52qVHXGAHS0Sfsog7qtTh23OEj2rDbr8/qG
naYGPAKtt9alJdfjV1BbwB38A7mUl8uU7PLQDQjrqdKhguo3BNPrHUFXRUXVy280PYryxLuJDF5D
xK7ITPKzRcHlkmCBF6rgKaWUNYB5fl+s2jjPKTe507P//Mg+ipjEv3tvFc/Xmqy/SNtw2Dh26ARe
LxgMX+u6vDZgB5Qsk76tBzK3405OUiijoLFFkfjJhq+SYGwLtBwJtoC6dUiYoTt2uuEliAg1OC9j
IIvncgO5qZ8q9E8K117YhbQkrK6ZIivm5Lf9F/fW6NxrrIL0P8l/i8X1SN9WgaIK7yZDIcPM4zBx
TOW+QTA8ARrvfdjz+n4cavLvegMk9E46q4H2eHotyf+dXnIy1oGKXZpBHB9fNVWeeucXx9FGhw4l
kdF4+uAAjb3POvYtvKSIHRG5Ew3skieg7x7nR0+O3imAKqALAPEZHlwqDjWg52RlluPxGCbsBh/U
R/hd3VCh0ZsrB/hH83LIwWkUEKDtV3VCL1eInUMGTFRMGAeK75HFuOUHV7Axv2s9df8gwzhXmY+V
hxJNFU6Vb6TTcoV4WQ1m39NVG+4FtR/Ih5x/zF/R7LJeWeZUORp2LruwCE4xIZU1xMyYHV7kFlmU
a4bk4j6/oix2cTxzq6TVTMwYHaKHAZMvZ06YoQJS+nntoIDpZNsv6oBRskA+UNQUgZbNDTfKeptC
xgMPu67SqBf/y9ZWkZEw0UtRS1NxmUmEBJTI1d841aQXEA4c3vwL2PmbSzmHPo8RYnc6o8kzlf6U
6RhN+Qm62adJQg1fHmD6YAc23oz51WmT/5IFGx/u2g5jLhuib1IZ+7oi8VWfWBvt7se7/U7jHYot
MszcH8+m3Deihp3FLboCaeGzIyrNlKDMuRlfS4SajgVln5eLxhO2HxI9waVZTld8JQTku+U3JD46
TsryI31y/jUlm/N+Hhb9m5AEgnP+vvV4cZTo4vJf2AUGsCIzmXpTT9fcAhO6ux5n0Eo6Bz3oBld8
cAk/OePALWu1/42Qr7ConaZjDztCms29mcH0Ywi4+3J2MoVXbtYjUXTuVZcNuo/4cT0iKwKGCvhS
7Y+W9LP/sqZ/avnEAbT48GAeBi6oQflqSwPPgT21YoORvUtPdb6YF3vc5WDliL0CJv99HRRDPjF6
7Ln+NcA19Og35FLtIL5QuzqYSaeBXnosS6c2mx5uRoUopTce7OK/FMIgsBP0jftheQhAVSrhIuDO
FUP2mDPQj9y7+bXSrdgDRm4luR3O1A/XT8Ahof+QGEiJ14Evg9bZlBgf/0otVcLE0JyaJ4oNXhB7
LNjUwcaSPgko9zK7Wn5d8zm2gd3S4dz6o2pXAp7XUFtz4IiTtIcI3e/uBFde2k9+ePhT7kZNwxOD
j3jk6N18qZhK5w4BZeJVylJr/L+CakSpF7++3FtQWcvBN6X0AQeJhow2ZcZ2NajlIYAtBA17oIAI
u3G26y5tdHWPVfofzZL9KtExlTFYTsW636JTN8HkQds7sWAHk62iYaJpimn8xrqg+RplT46H3g2M
RJdzQDgrUn2C763ZZducqZVeV8l/TkYW82Deb1TSg6aMgcu4iWtTFiBqSXNIVQJIUM5cwaa5f6zh
xCfTI1wAvuSeA/Xl4AdYP1S7dj8nPfRPrr1J+IlBn4J+OJt2kegOuEYY1R8OJaE4+t+HG7gBNbGO
UUWdV7mCNtKyiv1+tkOLQ3RDiBOcAEXxrbHQSjxJsfPMqf2VTNVUQ6jJtiRERQTzZGoYMqQeNALs
WCVq3E4JP4IfcHjHQdPsHrApdU+oPFRAujQeP+cyJlC+nkf+sDsmfncIjL1Jzg8laDdBM2T+LfxU
kkMMcSaN2q8u/T+Ou9862cpI5LhFF0JdS5pcf0YyJsb3/5ndiebh7bWsFkMyY0G8rEoZN7QPLSu2
/I4oTcDZvLvC50WuanWvjdNEHyMOIBzjARcnqCCo8SertJP3nJPI0ccPzhYdgu48q7R3g1EQdrow
NScUrRpDSw2hmBr8jQFvhkWA1YN38Vee/H2MlyH6tMIwbwi/hMAm7cn4w81sXq6rQtsfSl4weguh
69R9ZJ/AZ+fbaIrwWYeNgeZY5V0U4FuccGdS0dYCKoBLDHkALJFx/NoDEQoyo685/sPjtDoAilPv
r74XSIIi0XF0SZPnrfM/Euq1TvNmwSsbsoo+36ODHX3i17C5SpsxS7gO9sojkpATsItjMoROM6+3
nLz0xBsa3ngqpyEnC35/c2Je//yvtxDNXaGw06hl5NaxZ+42rTE2l5qLXLQ8+Jk6AVNpw3RPFa7/
/pT0kuFypr6fg76YRN2x0c56TWeFhIZErLquo2ZmT+YUHzd+NjM+03wonKw6KZSkgWJ+U8q987fb
fX28lfcW4uXarQyj7m1JSoLcNkqFyhFmyG9aS4fUUf/NIuSVfo9GAFvzV1N/G8lzxkMfy80VFUn5
4MFysCiW4A9dcU7JdxgtBzzQnxngWilBfqa9PYghlO0D5fzD3LJ/q06586CNYx7LWwikqpHSyi0/
OS3WAJR4zumg9eAySMBk0lz7I7TeJWn5n65R783p27XM1NaZ8Wrk5ggyfUBmjkIEdEum6sCQlrAC
JcHn+QMNm6ZBSWay+FjxbasyH3vkpRcpbjPVcFyxM+A2JiwW3eBbC5EXKSKBCuQJbID5XTlHz4si
uqsz5OOSUks7yraYWdzgmaOgUfuWI/5ckZ4ryLvb0AbP1fwSYW8UlHdNU9qNmBvHxBG8P2mmN4sh
7aTginWw29z/p662P6DCtZN652c3hqKFSAnATUHe6BIgIJWRLYBdDcVAIl5q6g9COd/38ONdkAEo
pdwlSE+nfsc7dzG6s0jyY5eq1/rDbDawfhXBwIbzcujiS95XY8viSH8UUzsv49KMVIuBX4K+nqXf
Z+bL60ABAh43Bp1FbwcfJWETwxCwElaJdU0KEDSjLLwXSmrTneuaU76WLoXI22ETfeATEwAdV/kw
Uh2lXMJo+TrEk/QlgcxNaWfbCHAs0WzGUkUAhi7NVqe7yFzQCtNZirjZ8lywa4tWZrIGXBnUXQ4i
5ws27u1Oku0Zyb8ZRWml3P6xBkXA8UMwRLXTngtCu9Xgu63249IOeSVsU8t7cWoglnGmtvBGXMYr
BeOAvGe3UmpvYpdSZeRptP7KrI1fSOb/4Zq042+FuhFCpEuhii8E1WBpUuV7z0rrO4iwusCW4CyY
j9xDk7yUo+8wg7wXAH5IzNZ054klWHbZgVpus4Wtps7qyS7Lj2twCp9AbCS7dpjLioxo5eF/lNtl
qTLTwvklAl2y9PMmMLEZnJI2IW2odOyHUYqBRuQM1h82r1v74psOq9ZOOoIKVyLuBLos5DYvEMRB
vO50qvHsjlBHXpysU0fa5XmHIT6I7kSIex55+AUWfBEaY8/+oHqRviHvpYOGJHjEhhHHlCC+HbWj
9ClG4UwaP3dNCS4v8cErdN/toajilZLete7BPLqFCoCTtzXMdW8KjHVna65JKRUbsBXZE83cBUTp
07eNFr4MbEG8b7KcUz4d3y/FsiUJBV68P5CTmNqMBr9DzyQt+DV9CRf0HOJTINNM/idj1GzcFdad
Sw/J6lkS11cJ+CgjekIch/L/g95UXvA+9yvGIbw8FNZ4F7KaQf6bDEQCZ7ZRDqiRtIkT+yDY5scY
KXJRlFHh5lyyrL83ycAPXpS+kf6uIZcM2Z9x1lpgCA6I77lVzzVvJChqS3HJmNb9xS5fMDTjq1MX
0u5AVkYQDL6m0UShAXGp9dB9vOlBKAGDUnUbZgvvkTC6gEnve5lHM2Vqv9qe+hiunl99WNAqSxrR
4u0CL8+1DQsAymX8BFK8jxXo04mxeBnfleLtX19WngS2mTWDkrmblEWtAjy3LnG0fJIG8gzLcMvd
pRKEk2NZGksjTEv0R51vT6+xZqPNi/0k0WhVdEeMe3aBr/9SA6G6RNZVL9n0U9U9hecvaeJ0EbY4
G52+zJejAbUTcIgJwosiMi0K9V7cglrZhd0xZTnh4Y4lEsKW9L/ZEf7nD8ec+f60wv5JkB4f1w4w
MvmkzD5PW2BQP8Bt/AJU39QvVY+3UWpwwpvuqBIRSTyfOMaNx3QWVlcvlsTmHKCuZ9fHnqh1dZPW
pJklo96C8QPd9/EDhMiYjTl/h2PruO8Lroe7whLqPRRly7uRwxhfI18vts5LnyazCNMLZTfEfrir
pauBiE478JT6qNSiCIl/28RyqPPYwqdkjWT/IvR4wfcgKKdYjxBNaZ0cy8ipBETi8qWQc9lalfNY
8C4rUp9af2iv0exy6DtM9P74quia8UxsSMYISO3KEqIo+/uyA/PUm7/8PTiVHbqp5C1YTVtorQf8
AYnF+FkyY8iZPjk0uqZo144PxAmnKJi5sHZdP6UuViNitrdUKh7yCLw5COV3jF+ndy/2cfLzKBLE
SE1JlSNznY2VTzY/lqvvPOiUlQqGSZHWU13M6aec/Rdq3UtLzpGtwNENm3+un3kDzcMi0gMM0Kcv
XciBLSvjdyXHtj1Aib9J2XoQgx5qbcSWnMw/SmbZPsgG4BHet8OfAFqk6Bd3vZEi+sl6LUoddUvn
/UqHsLqfbwwPm5a9QWgPvxrvtJCU4DsuTkhWkce8j06oFltT1oJlLowmoKsTvrQLUZuyYZ3fWd73
8NsseRh0PLL44Fy2IAGJ74Q8UoTOOUO+REW1hV38Un6fPM2Ls+zLFIBTUoDN75tFfp0vKm3xZKsP
zLXBQ4dd7NmNiaIcZXKMQTU7WyXDI5OO6jrNNidMaImkg05dDukKyl3ke6V3QqqqqLDNNzoKxXbD
M8pZx3/ZPFyAD7egVGYTety5cjPjPO9wHob6XctLAF3tqgbRS+45TbxI+JCzZPJXYSeWz4DVCXhN
W5Dd10VfQaUYiASYxUaj5fa2aiGhaBB4DKvz0lgVm7tmVp0NmBgQSy6LE60NfTqnb9+G1MKJnFn2
en4dSyyfUve0R+GHNXloCWWN6ywsjOCqFENASCNvzZwtcYwSC/blngzhxzhkd83liTwRHtqNH9NY
PafYotUgUOEpABpCEXVRy4azOBSYlN/4ngypezxh5T+9dhIxKCpUzw7B0q45eSPjBGX8W+MumB2F
4Bg85gcXnerm5+oSVsD5Lu2hLQ/efpJujDlCN7gifIcRZrFrV1163jg88+66mXu1jIg5c/N7Fx9R
00Ma/4GKiQ4TkqmVaxTXFG4luOO80eto0eHnu+kmQGu5+HMphKuozFwmY84bG6V2ApIpVtduSdIe
pJIe1V4ReHRpMok8T+T+KZlolNEaUsjOMe8t7N7XLtuyHpOi1GuSrj3rsXCJjafoHuXEwJ0UmT65
4TVUbMEYjGQCR/6icjzbXarJ89u/6QF05Cs2diAG5ZbG9Zmpa3/TDql/0Adcki0rBIdWeounaVV3
htXpMcnVeQ0u/Kvnan+TcOTnOp+y4ezrkGcPFcotVfRMwij0Ymq6M5grUB1HI+9HuBJmE58vdl1c
GmbmdI9UmquXV/Ng+48u+6Gu1TJj5qTYtngW1mtlUKPi8eH+Z/YtIwjZbkP58s596+Tj5g+/bOUT
B1W7vyIMKQd2AbJXieyTdsuAavFruJNTzrd5/2kHWjzlDyS1Co4Q9UtXhk8wLkxoI1zg97Ov+npM
gkdCAL+7/nSjHNOUgFKbaQT96MBEhfy6yovW+zvEy9OuwewIziNI0DygEgAIrF84zx2vyjURMqy0
D6ARJsybcCxs2RSWph4UDXu9IqKetJ8c0gVv+zvPsp6P+D/6r+stHPiw7I5IXTxhZs9G5ZexsHeI
w1kvuTxbXbdlZMVYq2sMJ/jM5gNR/RdJWgC/DSRpEkFrdLXqA9R3A1BRrublTRq+QyOoZtJS+/GK
fAudyndL97ihv29xS8h8PwLWjbp+O+Cnk3Qkch1HJQIf9OJrcaCtqZtVdiI2+n9PcfiS+YAVIdP6
jXTxGcf/59p+AHY8IX13Cp9FPz80Yw4EprWBftprrjSY0U4hu8v12HEjn6tKN2UEQS5v1S+Cf7r9
nSQkAXxh1MbefYcIGBEb9jO1P9KzHJ+1LRVJRj+YOkCsx8Fp0ojIgJKs99+PWtYuqx6KPEdvl6QB
LL2rqLAFhHQiefPCx2w20Q1e491pD1YlWyFx8x+Qws5VoBkE+bWCYzunbKuNjHL+tlVlYk93HGzy
08FXy2VQtOdtt6JlThJPOd0fTZM8s7fkQVXWJSbC15rpUaVOl+BPTXJ9hufMycIxnJSWS/NYnvOm
7vIMNtMf3i7Qahi5wXC67OyWlJjrHrkTKdYhYwlbrHbm3r6EClY5Q2HmtpRiRNPy00hKUfOQN/np
EjILaILvMo7uhhsZEB35QwnyHXmMZkgAj2107Dv6DavfPXIuVFTEWChRvsDOKXPC/K8mA8MA/G2g
UDeTf6y8OYesW3dw/tm3jZiHMI88zdVNVGxU7s98+VdJ8R60ib/fBsxFyX8x3wiDlWNUbJpqd+DS
sEXbIcEXu8PXR2jkR42gmoK8ecQI/RvkZncWCAjskTwnDfsuzuVIO6y/Zn4ettcmNe/72VZ0BKb6
XOIBoWTbtUWo2C7n0Ksb332kC2D+aDzoOB43g8sFODFMX+IreQv8DeHYfLAtnCNlya2I1kmYer41
4hDYfbC7HZpNwKgmGDoa+p4MkhQjvd2Q5yOwHZ26m1Z09dwALgEk/gf4TxBmjMNONm0QtPZAgo6m
RWozdjei25xuav+s6rqAHHan57vCs+hf+TCKsTKBPWhscZIqukoi+9RDBfm8qaDnC1tu4m1D7qls
nVFPfAbHkf9yrsWdq/Ju1z1lHGwTAO0cQYVy0sbIoJ8f6gVeeZigUq4KpDCTDz+knUV3lDn3jari
fBe6BR3iTpm9feDAl4yQlAQPjI+d+TLiO+Lxxzqh2CP+j/BqH/E8H/Yo4XgChUlZBp//VIWuPAOM
EHnUv/RXO6yUAiogeOXWj/hsqgljSu/F9b2R0lDY5U6xh5wPYprLNtBFBOc4Bo/acuEKNyf+w33j
L221VCe5sROAoz9ACwddCkCnjRIpTce2Jmzcv0Ue+vvfZS/Nv17IsFuHG4V+YZGQM0PSNN0qJmGa
8+cZwda9GgkoHfszl5gNStOOo2jwDqvHwH/g39tIXAsWNX0KjXbYrBX9GOATMa7DUjdRbVJFxmyR
MzjVE994iVJdm/5BBFqA8gk6SOsZMu041Xmn3RG9O8GmfAkIdy/S5lKh39pWnr8iRPkKCPypo42g
+714sVnuld+867bfSGUDcs0M8D7xV6M+FbwiMOr53ZtjQF3NSAv4QCU+Iq+5+1KJkY3G5sn4GNi5
wexrF9hyPjfhfd1y/zlfW1sWaAMRzD7vuRUy+sJe6pgO2gkWcbt6kCjaixSOn6tnYKFYqCQKGa8V
eW4zlYhpInOn98Ek3fQYQVY7dcw66kK6FKrMKj8gDTpE3KXs4NzXpAJIl6sERkSemSSXBZF39tEz
V5a91pYJicnIPW7efbpVlwyy6Xk++KRzVCExCGCwwaEQSqy492JCXnF29GYcK0L67+3bl6GT1e0r
2hAR5hEK+EZr5TYJi6PEvPKureZHoHAGz7Xefo/9eYNjAed7N8w58oiIjd4k9J76MKN4DzD95Vfd
tcnrJswtomI/7Ibzd+PWH3Qa6CjjF4Cgo68gyG2taEa+r4Z8pnr16R7unIuOjrLjO/hSwSMfeHum
Ds7ZOSnkU9c73LSANcO8jW+/UhLUpBGxxFV8MCmypbKC1aOdDi00Nv7a5h4DwAblvctHpKc0+AUB
ttxLBa7jeQoey2mlwBHHlwjUkYzjQ7M9COT3Hd1sB71ABaMGcn74g7DRgvTxxM4zyROv8cdEJYgT
Huak/F66K2nicJN6iykmK18XrXlRL84x796n7wuPhDoZ3qmgCe06GBWZvcoH6V+ExKle7C4y/G58
7GYbgiEkTe7iQDJ7nf/zW9Ri8f/WGWa7surRS3yLocWqUWYNC+cFTygUYt9hzDjJmd82luQeK+3j
0cPkOtcOhtpec3NIOXLdBR28YS2NpVkbQVMbIBEoI4gAY/Nv8mUFBQmaMN52NK5amiEVgZGmbHLD
RCqoNAeTYbvqHv4aFidxhBZmq675wLoas4wQIJcfjPhLr6jVJ7XCddPireo/j3aVeU+URWEkCWev
nIYrNKZxxDcndaP70IQbGodHLmhg2SoFgcC3AEVN5laqdodRD/uKs1DBK55nR6O3OQRL0m9lF2F5
YDVRslw6ggxn1in9bwdisxRv634NnmVU0p4BBPCeWSHduv+nepu9YLFLAR1mCGSHUn168Zs1xqv1
fvFpV6tSaUm+/iLabSFvecmb2mQVhaqw7P+OSNfGw50a1eFBMveHrsFQdrUd91ATDLzG1nIVruSh
BWuNnMN7lwah2XVH4dHOao9yiv2zIQ8+cZZvpqxu34ySqcNebAmxb/qE2w/sXNvP7K1sOm+kdwpM
VWc4sONlkWT+2QxZkrPq2QwdjY3QsmfjHYH6j0cSn9yP52dH1JefnfM5awhAAV6zOnJ6edwfWsfv
FUDXHUGrYa2i1mwgoyDexZJJdJFe6aiJ1WPwImeHwPCB8/VqC2dqjHEvx6MQI6E29/wLJ5Yzt9Wa
QwrZ2tatNqAy46scksNz3fzzkobTkcUZGdR8hRNLvmc14oc/MinAPwlNlkS/84pyaNEA27qJ0Nwr
X1WnKFyzXPPee+oCKnHqg/66wFI48av+JBgoZJ+99xvCnAyXdaNUAF/t95f6eWP0v6hpo7gc0Fl+
aVtJ3q3Q2zMHtyb/6PNzuydi+nEknOf0SHzGxQN4owHLOm0H1LYorRfRisfjgWJTUSZ73u8ewGGX
5rBTEgu/JyAK77p5SpWsD2Dah3C+93P7uvUFVJtO0n2nP94FdkrvhDuU353kGOQ8Q64nv7VTg9ES
NJB0gx6j1vXtlPNPc0Ld85NTylUyyR13XKGuQVliT+MgMsvogmigslLiuaRXijB40WtynpvIGLk/
sKrbDuZvlswBZYCcFsm15nTv5c0REvt/zdjtGd/rP7JVoWR68goDFgXYPBOcJdBqCdXv86/P62uu
2YbP7JDSw+ifU1fIcRqy77kYFqVBLhv8mpYpFqE6B26g3N7fV2//v/WYZKWiQaI7KR4z38g+O1FV
/H3bbAW7msII7wwFB6Becf2bUkYbqxyq3q7+3TmlCbRghbtMpxEk3e2v9NiBF1BpVAuT1ToiD+Hb
C89Z5RcojYckSjm9RxZ/lOFpTNy5XIV9cI0BvvXPlMGExKa9fsOsIHfJLzFSVaKc2oVSBR8jFoNl
ZwUaZhg/P+ayxohq/eNB/mQpS0Xh5ZFWh9NiTCUChCKy8G8LMMKUjioHkeg5uqo4Q1bBu4h8RkE8
9skyNQC/xNj7hIQx/bbxiRdcDyjkb7RvLmeDHv57Slbg9NL37VZzjrFaV882zdm5535fUklnRDds
e1yBFKv9iYtt2yxGBZ5zvejk0NcV9PpjklMC7vBh78o0Cx6GYGYdbBdamgedFGQKck7Iwn23DfvL
NlFV2NXE6fHHZ+fcqGZL9mctD1EwrjejR2EPG91ViJ/ZY8ALeJGd2BlfORX9EgUcORtfKS6PSBXv
2c51jyvLmeAR+KRABPaGQ0nnEZbMAXcHDvFnJNJ4uq7APL5I+alEbxtdpecacO+37DL/Xyz7RRvv
/WW+M3CF71amwRevR+CCGouGy0jQKmzrYw3UVrxcGhVzLfA4AbyOjycO6C2mM6k6jZKYt4zpdk1Z
XGZPW1ciuW/Bu1i3H7d4hTa4/tVZwzaSLNUgYCbkJiXtAAbm4/GWCjgR+Viepo30jGlABaxnJk29
dHaC9DPHXpy/T6IwgTHVOjTP3RHyCrCnmovmiOTjqZP64QpOHPqUCPeq+7HnMK4BYHHsaA40P1pR
OBIiZD3KiHPlQX27xJayeuYzOkB32NiAUj1j0McM/WUbOkMhID+51bN09Dp6aUt3bKF24CNg4o1g
k3x8zx4ttE5hD+wcof62xXRR673tT9UreBinrAqZYs4rAWaB+Pt1T+Qn6ZeU74o0p6f/UXFTFoWX
IxKpZlSUbv+bO3RR78BlLAZmJO53ze5YphjSjwrhL5U2GTPO4/ZzBRyzMpywGulD+1MNxQdp1OgW
35c0c5R0pr/8CKEUOvDC2pi66tL4t69/Uw56HyiKPzjCrObEPkgY9kWg8iSj4gG1qX1p2Ih/dsdu
wCR50FxE4JfYBss51CgXn64lF83xET+hE+GakN86SwboKu36AKNgSE7evECcJyJ19JIob4C15Wfz
epb83+GZhId31NYRsHcz3fwTtfRwfTkuqr3z15pY1K9DB14jPk0MHL8J2OhfIxZvSDVhuvK8OxmQ
aIjpx66z6ps7AZVBx9B+UikSqYu0zKlgj69RKtDkCdlyP0NcyFrVZmbOVSGMAjT5h6JbDdfU6y3S
7b5V2Rbf9oys2nTbmS6MBpCDJVXeRB/1aAyrEXCyM2DfDAbVEy6/fyZUq3D9ytcMWZr6qxddgpK4
7rLf9tSBwRsN32BjGn9Hx5acdZxCr29VWecaIWzJZc58iecHgfdbcixMOomWSbPfrHNaC9XbRqRk
arzHaFp9bCSPiLyGaTpbbN8cV/j3KH+Tsdy8PJt/FZ5mVSGE6xgwFBs5ptFoUM/cknHEZH70jwmZ
A3QT9xHpWdsoptMKr3lCcorgx3rIX8Qf4NWNlXV5spJunCqgxekZxt+SFMBRH5ErTFDofJ1+cOWP
1441JgYAMc+ywOPRVAHscDWd3As2bd0/ofOHP9a5+606sPX+8f/al6pHLX5svBrAdCxYaCWPOBbA
fGyaBMPsommVKnhkn7L8W+z+6sHOFZc0d7A5XlNLqX/6OwOy5t0rK3WVh+3WjSIUw/4K10ax7s/3
HM0njBRCogFzCepPaLvvFfc5Tz/R7lWA5vHmadyI2dEb5MiKnKu+09+szR/oeSSiNPopyxhYUoXd
4NTS2YOcT+81w0oZWMjQLd6sJiTo0Z5U8SK82D2D5vDO+Bc2sh8DqxyZraDCrJeQztbvxLSWDyXj
y1xJF/1ihsT9Pmc9zO0W/+3MQM05+7+xSsdL587cAmfjiz+Ll3ekhWvPVNq3m5LUw7LO2Y46arXF
0Zkyfp/ZR+9lKiok0YbqZdD4RXeWNJwsnX7zE4h7gi08FUBwkniBzz2HuaXDK/wi++ObwVJB1wSP
1nL05N7qxHyqArBKzYPytfPATboV0rbiNJ9pBL+vv6Jlydr9oVRfQaXIt4WZ8bKqO5+GFMf3hed6
lqCE0oFVc3aQB3EFv3kDQGRSDtapiqbZmf1FexeWQhdMWXAR4fH3ByfJkQZ8yZDQ7XNyF4jSUhjv
v+rqr7V4k+8oPxHNqXL72RIuy7m33+Sjp/vkqbQ/uehmCsRLEeApYcv9rKPbA+jfVi0sAvboKfaU
SfBF5fwbRYEjak3RqgrcJ0AZb26EcSwSjbK4GMwkfJC9nTNhslMIMuzTiaJHmVkn9tD5o308zloa
31FUVjQ/oszdf6WgqSidFcGCrmHYWe4aVwnVCRmh2zWQhLnNJVmeGPJBNgg9vmEe1WJqIDReRBKj
xAAlTxVNS63IrvW7Ls4EgKFgeafC4QIUE7jYKYWCQrbyGldViCSV3tCXmx8zhliRpvrKOrpY1vMq
HEgbzDSnZvdLaZuinUwtYbhThC1J10eoXZ7Jh/0KILExFyk5+9EMRXOkEaen5Egr92miSxBshnmS
m8dXZCSHhhQezYpPsuIznvAMgIN1P5quHsrsj2QvZR4JPFvf/DD/cMtRXFRqVlR6lK3tcemwT5xQ
xqoES/5rbMXbulqVhFbTnVzyR9RuKr5lrZLekZKw+KQR2YP1+WElPOrZSIQXIaC/TUl3T94xlWu3
hXY+2uAG+qf6Fov/XhRXygt/3Dom/hT44zsZFVmzOdcryuDxkYqgq7hf1Lnnqhkbk4BOD9U/3KoJ
jRVKbiYt4eChqys11btISsxrwM+BlitR5CQhoFvVgxvKUpByrDAw+Vq/5cv86NwPgIPipexbN941
zjGyt7N+KuHGTg8ZkOw3S61EnIW4toJr8TdtOHVNq9xngbe29sGeye139reGrAa0Cob3Jr3H/G+c
rlVUrv5ZAIvnBOeMICc6VEPnVg0RwVcfBwC0fkp5QYAv5va26P7g9GSFVrGfxsTu0TCZdw6DU029
ZbLu/f15Ypfy8L194+yzYdNyxVWmCPIppe/hRqtlVVvhVle0eMl/ogfM7wMOmIezdnkH4GeH5Ur/
CVRmfwjuIeZqePTA3XfiC1KDY0jrzMPI6VXS/zYd+vYPDPR7DJIpxjIy8fjnfigtrne+Z3L+enbA
Wf3T4KFN2MqCTzX4c8JAP6WRgGoE+qaog6W9om27J/yiFU870joP5M8tb/t0LT2UIPC1iekDqkWM
oCQ2A7wBWHmbXDw3xEmJtI5ZOF4lI6+lzUQfTiz/LCLKtTwdzvGpf5Juw4hta7XuemgPdUtcpJBj
Y+ZSahqOHHWptCGi2/pINVvLuI9dQlOQC3/oWxU=
`protect end_protected
