XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{�|�����<r.��zg��,�9�!^��@���\^���3Be~՘�E��s�F�G��ˈ]8����!�:��{U�
`4�m�Kwh%�vX�09���K0Ⱦ�cv�tj�e|~19���$��o��h�����!p�Ǉ��a�;W�c��v��@.$=M#_.F*U�wDS�d���3HyMؘ\�'T��|d�,}����l����GS�?`��[�n�r�+E[A`'�l�Yfg�Sc�Kv��_^���}[I[��&A׃���a�>?�jSW�+�(�S��Z?� I)ܗ�{��)���F����o��c@{u��5����t�ڷ#��3ￆD�lE9��2���|�Ҏ�pF#�����8�<����-���a�w���(��ɀ����O�{YlD:�g�Z1"�!4[��7���������5C�o=�\4]�KQc�d1%ِ��r�]�}sx�E��q��d���/?�8��K�?���0"���G��Wɪ"��a�<i5<�("*���(����C�&�Ă;��D����!��ZR���N�&�_���Pf($V��!�牰�<�����n�b���Нu���/A���N����q��,��]�x��e���9�)m�,z���"]�~�ń7jc�>Ux''0�@�B� 
�����~��>��s��b�R��|T�q���iP�0?�C�A�}�N.be�9s�Д���fj$����L�C%G3��s���}�2��6}�z��T�t1�pW��
��O�kZ�ML�pB�XlxVHYEB     400     1d017_0/�e���uX�%�����)������QC�WN|Ƙ��C�z����F��Շ8�U~��D�R�E��ĺq����+��2?+��c����#���};�nÛ7_l�XR�W���o�߈�o�Z� �S�"5a=L�h���oD���-�}.��+<�0a9Ri
b���Y�;�	@7� �L��K���UxK�*�e��)�)�JHe �K�/.�ه)>dCK�����V7�"���&�gwJ�H�%�ą�7�]h��1�e�*��cJ�H���ْ!�R��n2�q�6�	R�ث����18���-�<��`���gL��/�OT�n�^ן�x��W{=�w����9ojr#�;��z�d�}
|ݙ��Fe|�և������7ӞG'v]����q��l7�݈q/E�zZ��~i�:�v�\���MQ+���Z������6k�*]����ED��>�MXlxVHYEB     400     130�J�Z�� �˿&
>܏����J�2��{�KuHr�?��X����3�SX���Gy'�j�W��:i�Ʌ<��!bCǫ��S����F)�������k+�l�z��TH���'䒰��wÈ�$[�� '��i�`0R��`�K�F�8*#p�,;9/Qٻ� ��O4�ujup��C��� utx,�.T��ɐ�{�%uC�@n��R�M�ڵG�A�v��8	A��hga���o����Ȁڊ��W�$&R�2�ٍ�Sڱ�&r��t�@Ќ�c��n�"){?L�����8_�_XlxVHYEB     121      90�)R=ViD<ڸ��9sЅJ;V�_\7Zo��?����፺?K�Ήг�����sn�Z� 0��髹�4Дx���-_*�\1¦�2���V��!�����-)�����L/Ǆ"��Z�LZk'�KG�2���WL�|�L