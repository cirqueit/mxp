XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1���S�������h`�H����`Gh�0�4U�i�3�K�:�!?�������$}0B�Yi@mg \5����Y��q>@�K�%E��u�H-�A�Q�iJE�Gi�CZ
	:�oV��< ��°��r��Î}Z\�A�������Z�Џ��>�e�I�2U��<��~�kY��s�Nb�9N�����~�\Y$�6��*�|���q�2$D�� =K5lv�]#^�
��{t�7}��)u<x����wD���\�Rq�xڜtF���?&��I��S���TGD�}��WL��i�C5T�>[��F"h��E�K��W���H3[g�]3�@)�z}�nE���ˉ��d����iZ�Q�9"�6i�	�ar�x8��� `Ã*}+�"��.ϳ�I"�-���~�����c��b�+H�a]�+�S.'�؟�H"���g/�{�ozj�A�U���rI��f����ơ��pK>V�ҡ�0���>O6�Tm��b�e������ �!���I號zkY��U���?�w��X���X 哕G!B�!Mv�
[��5�x�e�{��ec6���ƛ<-�7؎%P�������=K���qeĭh`��ڟ�H�U�J�ΉO���D��a��>R݂����̑�d/i�:6�!=d?Bb�~{~���J״-	.+a�wa�}�__i�B{]��a}��4:Gݪ�J�- �\NH~�BY}P��Cf����Nw|�E�"�o:�16�5�f����_�n�&H�\���⢄��O�XlxVHYEB     400     1b0�9�01�A=;��qf7�du�8� �tv�0G�n0
bªF���	��D��jC\$0�K�9�7�玁��y�%g�z՘u�N�����>h��ͳ�ħ����x�aN��$�^�ִ�ḍ��ְG!����I�X沦N�UN	�� �!ƹ�j��Ճ/Zf�y���E���S����9��g+ᷬn�΃w!�����}[��AbU;����䎻�\]�iŽ���-�dI���������=��"n7�,t2�0;Ŋ��A�di�V�_�]`u;'�����֤&������IAq[�O�*4������b��M�S������O�d��oL�'Aq��uC�b.*��JF�i�e�y����Q���&�G\
LM%r�G��O�]��Y�G�5��a��.���]O�X�r6Ŏ��#fH�9�P�����XlxVHYEB     400     130���*�
Q+bwˣ=��?]�%痝��K���b�, ��h7sVP%P;�j��v&�g0����	$��*�:���έ���X�?v�:�LO0��=����G�2E�Ȳ�������4Z�㒊��t��U+����^��!uB7��A�>���4g/w�L�D�h�H�����=#bp�� �)j|��vd�'#-�����ĵ%������N*�qݚSie`e��K�ě9�L	�Ғ��ZW#�������uy��f�o��W�\|/�����������ݼZ��Me�j2)͐�9lMXlxVHYEB     400     120����00i�4ʔ[�9eo0�[en���RW�:�2�@	��}���+��*b˦�}�|!����H<|h�s�o����}K��GT*����j8濑����87>����IY>"us�F��?�S���*v� ���D��T������K�~w{�l�j�㷿0毚D���#"����0�l�S�+ԉ���/�X�O /�lD��^�9X��X�[q�������{�O��;^�F���I���>1�PH����}�d�����s��CxT�Ep��O�:��޵&L��In�XlxVHYEB     400     170_��|�7�a�u��*[�sE��	r��$ю�|n{_�L��r�ɡ<T�w�K+�ys3�g��!?�-�j�]`���� �!o?[$�Tp���y���ۜ��8�/�T�s���l?��˄��Ys%��z]��fc�-- A�j�ڂVv����0�X���2��~�52��aZ�=Yk��%�P��L���?�\o!;���MxD4�h�$�bI�gGvìc�d��(��T���Άaŀ�����w�E!5`����z��W.�9��h�n��<;`�HA�˿�S��ã�Q*�jf�1�/&��	�b��^�3�`|0m;�q`�y�@$T�(XV������U[��� ����_��n��Q���B�a[K�g�Ҭ�~�YXlxVHYEB     400     1c0��R܀����fj�Tykc�����
�?g�����ط�j� u���vQ�0�/����{�Z8�gȝ?����%�=#�����S8_N���dC�Δ�2�8%�H*@�!rÝu��̼t��7F����m7G�7e����2J ����K�_��Y���;Nk^��uRT���6n�ъ��?�ՈnvLeo(��m<(�k�ت�<����5Ӝ����QYg�R��bf�͔l�#�W�%<��=���Eѥ�$CC�m�Z�'/P;��_T�TR��E�Ǚs<#S���3�A2 B?A��7@��
'��)�:����.C�F�k�0�t
��7?<���sB�X�9�9��t���P�_��gsG#	EV���q��br7eD^���`k�a=3+�g����:(�AR���}B�GϿx 0,�4c>�Б��5Qڐ�8�. �3XlxVHYEB     400     170�1��5k.��c��Ǜ�6��T�֟.kg��|�28���X�lk��w����$��r�1_q�t&^������9-çk�U��,
�������*�x�^���MW��:�X�h�4���p+�aUp�C�a�4c)rz�k�Q�0?�.�R�:Y/_�h������Mb�Xq���f�$-
�OL0d�+$�.E=aQ��n����8>7�{�N�`�B�쁫���3d=����
�d%�;*��I��;�b���p���0���2Ģ��$ڮ/�"5�~�����]v9��=V��G�i.Gqڷ��\�oe�\?�J|;�>�pV�T��K�H8^�w)r��|0d2x$�|�����q|XlxVHYEB      5a      50���XI��V��Y����+{t��[
r��ތcѽK�� �M@���(����ی�K�kK/��_5.�LH