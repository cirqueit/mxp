XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8�22���7��0(���.��ۥC�hh��ׅyyf��TR�>D�F��Z~QQ`�xZ��d�/��J���+z4��f���3^�i�࠙���=e@<�sF�%;c�Z+�j}�6�����z�΢��|#�L=]��xR����6L�b�*i�C�\���@��A�.��J�����}<g&���Z	�ܓ���O\��1�\����|{J�jΰ���]�
���賭�����Ŭv����)nj	A�٪
��{�ZD�4�^��n��l�^��6��B��O��z��jE�װ����h��!u|��z#�R���F*�t�h\3��q~:�X�����*�#7���b,?�蚱�����NQP��U*A~��s�AG�0M�<�Z��l?�����\���� ]�A/Z�P_��;aG�huj�r��N�`��$­7����wV@�m��-��b�X�A��Γ#OI�����4��|b(����a����.�ᜀ��R_�!�{	�0�("��P&����'d�!mS)*����V@ܹn�3b��ڇ'��̪W�Q�G�U�2H`V�����l5j`���5���[���:f�[�`7Mn��f;}��s)He����\*�o�������mz~!"�8�ӯ׈	�b�
.0�N�����B^Dկ��C+���n�f�d-x�A.+�o�!��!H�_�M��
JY�����*���;$�l� 5)��z�éCa���C�(-�8��ԉ�v���8xXlxVHYEB     400     1a0�5�vd�gK�%>�_���U�U�+���="	.mC�xb{~���N�tc!�:~+)����xnJg����3�ފL�����o_j��Q��`V�ZƧ�K���e���/U#���S�&,�Fm�2�O�V�r/B����ֿ���0+��e���fz�5����^��ꩈaT/�t)<��ӈIeF��c+�K�6�y�4/�s���l*�I'�󐰐��4��~�k�!��@榍��)X ���Zb!��K9�Hk�AE]��uń��e���4�]��c�ԜJ��6���a�R'�"�7�<��X��]�0�����m��ڰ.�$�
1LQ�6@.痧�R�؂fDx:��q=>�~ �*�K.���]K��}$���R����qpnZ<�3�N�.�n���ꯕ���MB!�XlxVHYEB     400     150G7�R^�P�Ԑ[�D�ZboWo;]�ݸ~ft�`&"i�\�Чw��s�x?\l��/&�ł9�{b�G�(�9dO��{a�FP*+y6M���P 
d�ƙPt�`}x��Җ�^�M[���O�R�8�+tX#��x̳Gr�&���xA�]�+�򸻡c�G� N���k-d�}��J��6�E^M���8�r3�[�ѱ�]����R����*Y���!������b6��R�%+K�6�m�߿���$�k��c��4�d��[fT������,]F�D�0��xV�����z 
�8����H=��%"���Rz���GOEj�XlxVHYEB     400     190w̥���:�"v��*�����
V� A�6G�
cN�z��HD��W;�'	�k)�#��<G�`P��ꃽ)}<5ũ��sTŕ-2��Z����:�X��}��h��M�w��-���8�٣I�1]�-VZ{ah���vk̛F��K��w�aۘ��{�hc��u��"aAh$�Hl!�ǎĻ�c�NEy B<Y�չ�l�����
��
��L)����Nc����F�?Ո8�ۖ��}��`�j}�!z���k0�F��(?a�<��c¯XOB��/O,
4)�A�Pf
+`��M�X��J�c�+j��eF����7�ˈ/���RT�&ƪ�2REٛE���ĽE��c���.]c)c#�zX�;&�wxi쓺���C,٨XlxVHYEB     400      f0�u� �h����0!zRB,�����|�`�-[���-����F��5����B|��8-Қ���8DW-t���]_�P�ۿ�-!�5N+;�H���j�<%͸����&�nM}i�L�Sv0������bܦ�~��0�ՄM���:�����Ck�l��<Ԉ�7��1E�a��
�܅D��&�%1�4�����,����I8T��
llD�Ԍ.ْrMn�mv���W7e�u�{�0
{���ʵ�NXlxVHYEB     400     120�����¥-؄h��oISV�����p��_�����_��[Ӝ���j�:a����3)�,�,��@�9��� ���F���s��{$���l��*�d�0#X!>��Nw��E��Ha����膯3���LwtY�o�xi��2�d!Ū��eZyRE�_�qռ3�u(dlU�'������N����^7�27
���u�����5f���Ò74D�f�]ϵ��P&Gf� �w%G�|	�`x��x��+�Ŭ�5?PS�67��ۮqM�c�#���lp�)b�]�-���%�f?XlxVHYEB     400     150�~�~���*�c�3��/���Ĝ>=<Vzל�:� ��o�e)���O�'�����"ŕ��Y�2mK�d�����4���֗��4Rv�����r�_�4廹��ϫZ��Rv�kF�l���b�CqJ�}�/S��d�O<,k���`��d���F�O���\��(������H���bK=2���4{n�y6c�\�oj��vZ+���*��gl� ۪��C3�~�~��j��wǥͺ��F�]����W�w�9	p:r҄��RD��o��l6��x��_�(��y��d�f�-����':E����:�u ��__�6����(��[�XlxVHYEB      ee      70����9��qB������X[�����܀��|��p$jse0���D�5��L�5��	.}i%�x����Ps����B��.�~��S۬쉘]�o�>�S�����̤��w