XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��͌���FCÐ����eh���%E2�۬ZW�<���������'��PS-R<K�q�����F{K�^��wrW�>��d>9{�0��/��e_�y��Vi�������-\B���r�I�IU��RnI0RA�H����s  ��9(2��d~���
Yy�;b�,��ٿ�c�*��$�¡9�����kn5ύ�zf����:�X����E��g��~9N��eNsՎ]5�P�8�A�!����h?8AT��Cr�{t��O�����k��2-�T��^.*}:�K���*i�8��oe����j�X�J�Yg�ɞ�&�nѸ�ny Dz���dC"N��)�N0n��cJe���6H�r=he����P}�=Uz��u�����Gآ,�v�`e(-͸�?q��y\����F?6MCw��(��]�H��NMx���s�͚�iQ,�@�B����g,L',\b�'�ˆ�K���i		�bQ�@IZ7���^��g\���,+x����l��(6`�S�dV�,C��X����s�'�[�����wJY��9���Z��g����<�-a������(Oٌ�)V�UN�2WQg�X������*�f��NN��X�Lל6�y-����9��*��w����x'�"�����E6!{�[i�}e�� 
�V���0�x��a2��+��Z(b�Om\b*�q�l��"�J`�ȺDsq��E=q\�|X��3we�L�;����ks���Z�"<��Fu���\A�X�p���XlxVHYEB     400     190v���rXB�p#�Bn�|U_5t+:��_-��~��{��5�f`+����[�:�n��y�f���m�ɒMTT�'[���y576?��>-ܽ�"'I����ַ��'Uo�]ɔ)�W�@^G���wD�f�T�L�/�XR��ƍ��άV>��Λ���������e������x8�����Yķ�'9���Ü��<��Peإ�ngp���(�W_�g	ĔWP�[�\prNy��$ f���5-���7����0��n���]��"�D,A�/��}-��D_y�M̝��V���N:�i�z�iR�i�j�������G�G@ohv�Ԓ�Ϊ@�[�C(Jcdo�#{`͗�f�.�;e>�J�刦��9~�@^��^Q8�ŭ��JXlxVHYEB     400      b0������j7��?���oN茶�2}�u�$�G�Ci��Ѽd7#���!�$�R��@�2�:~{.	�'��.�-J~����	�!���.�Sʰ��q���OEW�V�a��3��q3�N�Ь�u�.>���~��g�HWּXO�3�^����3����Y�ˇ�8|e(.V'G�XlxVHYEB     400      f0�f �v���2�W3�nBd�oHY�V5��b��񴏬@o!��P�'ݙN'j�n�R߂Du�:��r�� ]�s��O�]�K�����z�AqL&����,�_1�N�0X�Fu��g��f����n���9C#����E\�OV8�ɞ=��v)��"	!���!7�|�n����,8�Y.Ą˗��p�d��w�w�v�S��c��0}YX:��@eC�L�"��6V1]Pvk�"��h�<�m3XlxVHYEB     400     150�L�F�/�J�u�RX �������X�>���j���������ZF2��GP�*�@o�����������dlc�e$5����"�lGF���P�|T��\*�M��;9
��J&�7�¯s(%�@�pyF�����[�%c���Z�
��^پ哝���� <�/(�i �B.H{�*p��>J�ćy�����V;��+��A{�.N�y��u�ǹ�VY6�B�{�#��ҷ��e��?�v�����L$h�Ix\n}B8��O
�>���a�5mXg�1�$&� �>@�yA�b��,W𓂲F���:%��c��L)1E7��:eXlxVHYEB     400     160��:��Aw=*n�ql��ֽ?��(�=R$��g�|�	�ZV��wr:��>�O������60K_�~�B�N�v,����-��$�"aQD��cܜ %/�;Ƕ��稍­$\9�DN����ƭ.5Q�DɭzJ���۳ܧ3��,�,����lyS1�`�����/�0:W���_��#\���&�1��
N��7i6�u�i��!�{QǄ�K.��;F�{Hw�1���uF�OM��3N�8Al\�Yo̡uB���f}�t��&k��8��Q��(��D��T4�6@�Q�����Wz���o�V� �F�� m�g
B��f.��3�ӱ��4��h�XlxVHYEB     400     120s���ì��[6�^+��e�����T�T� ɕ	�J>� ?hPq|F��Ū�j�'A7j|������ߠX��AM�Q�z�L��|��yM�yZ���c	ɾI����f�E�5��(�6��T�'5���*��
2�Q����@č\���7����{������1��&��#*w,p֍��KY*�i=��!�H�0�����(��t��z4��9y���)�Bcz}�P�c���j�H���'�з���:�Yշ[���j,liH6v����h0m��Z|���k�mEE�&��`XlxVHYEB     400     110��P>�F(5��℔��f�nb�RP��\D�^빟�c���z�y�謧������/�U4����}0]&)HyF���ͫ��N��f�X^:9�KѶ���`�~�vg����9/V���y7&I���R��>_��	��V"���ݔY.Ws���#7# s�4�n=QG���a�m��[MU��Y�\����}m�����Eu�Yd��'9�K�l���!��P�L�J��v�� � _$�}q�V��t9��_A�&>�M� ϐ��2w��WKXlxVHYEB     400     110���T�c�Z��6\�S�}���
���&n�]�cq&FwJ�ġ��X��p�5���0ܮ����X�>e� �R��6�?�_�e��O����4����o�i�չ�7�9jbC��vo�x،>�VN�wG9d$q��)�_��^P�sRD��}��Z�Si�"r���~�ɵ �����b]{�-`N/����
(�g �j x���iA}��f�9Y�M!�p�9��KRr�x�㌭w�����J��>ϝb�����q�������9!�{`�J+X �)XlxVHYEB     400     130]J�6�G���A�[i]��
R:��*d���|��j"�t��G��Z�YTI��7V�f�fR���89�c;���I�ۥ��m�[b�W&	?|1o6|H%��,�d�T�5�%'�׀�f~Q�~���j'��՝eY8C g��N0$��N�b[����[	Go�W}�M���,(�=(��מ�ȴP�(�zU��&��(���dw���{U�d%���\�;�oΪ\Rx\���J@L]@�L����k�-�������10&�����oKW&����Z	)o��y.HLw?��T<���wXlxVHYEB     400     140��E4��8�}�ˎ��|�(L��A�����fi|�}�������^�����-��`0�	@���d:{�&�Z�pSǐ!!bεu�۬?6�t��u�"�ݙ����wE*��Q���4�Cah�j�[�?� c��I�<O�D\	`ɬ7(NE�i�������~݆��f�≜,����U�7Er�����r����e(�h���pJ|UK�uOBKw��A��e�Q"ᚺҋ�yl��/s+ ��^��V)^���ot����FJc�:]����yV%:G2��H07(�j�����|���d.T�c>kނ��oޫ��
�XlxVHYEB     400     100�X��9���w���y1��{�v����RS�I�(�3@6��>�?���Q��w
Xy
��B�b�*�\��8���I�1c�f�7z����j"����2˷	�p��q�����~>D0x㟷��yT���~{G����2u���ȞQ�U��tE+�X�_�/6��'�S~�e˃_
�t���=Xڦ��=��(��ZN�C.�;�P���-̯Jb�ૃ�ƨA�,�B�'~�HNK�"I��:��Ѯ���:J�<u���XlxVHYEB     37b     14088���1�ˏ�J��:6�d�o᥎�7aB�S����n�'�Ƹ���jf�Hq	�K	�)<*{�����i;;���"�Q]g�=�������/�$��&ۋ➘!���G�"��蹊#���'������9��u���ذ=��Y� ��A�"D0�'y�䷘ 	v��ء!�kt�(�j���~�so6J�����-�y��#;t��Kk��
�,X.��aҶ(Z�3Jjȴ0�'�{�s1� ��,��7�B���d/���`1a�g�~�۲q[ )������3��=<���HT݊r �O79	�
9B�d�E�	b�