`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11824)
`protect data_block
sxQAB/vsR3c84/YsuoI4QQ7yPbntAdoCLOjxrhwAMzmEQCzfZi7BqQJBHmvtdVJXXDYlxMcxJnzh
biSmvYCLEz/zCPIXnGSqdzod2DNmR7kGrS/KiVW5SQMRVNiUH6GsZSdlzmZgbaxBa19tNneoVpBd
9DUiSUx1IRgWcMO6CxDNndKZAr2T4ZBueSZoHApWReIdmTWYsri/YdxEgcMtMbLnZuCOfEla20mM
lm7IkPC6pcl5rX1POf4RjuksIcyl/mUvKpcDdGMJYs/YwKRqgGd7zww30JXGmcmeL2nmKJ7zWung
BYZuZG8x+O5qW/9SuN9nV2IZ3yCh9VIdPlRyAJhrDm6YkogKB+bYrZ60FGPIi2GN4X5cNlx9oNla
TgbH1ITCLeJl/i1Hpe1Li2tT5pXbR7SSENrmX2lglcpoeAp4gxgNsu8iRz7TgBBBfHWn7Gw7o2YK
S6AQiW4BDXUTpi/RxKMNBLV5jqSn5bz3Z7gPnUKnsBfKc7uL3S531xlzoPPcCkob2ftyKhTOhU3D
rrLf/BQ0k90SAND9Iz7D4sFsBKECr0NWK9OqT/ZLIBkx9dQR7ZtOaaRYzTzaZ25Rj5aSpXs72QlQ
HPw85Ca2Jig1htWLxEV61zZjzI5hss6O+K+GwzmGP/myMatr5eBK68QzAW23L4CNHwcOIT85jroM
745HwW0OYNbSQlyymfFL6kvG5MmuL/brUwWip+xfrNRIkAJKPoethkfCopVPIgFlMc3NiRjz5SQh
CwjEgo4Hd2xrxNup3LrpvywmcdfzK+CmTkR9faLiq6079oKdHgy50jL4OW5sUHWo1LLNbyf3xNqi
BrZWxAf08RmKiqr8NEWD9FOu0kmK9BVSfmp1iHJuUCKTpMBqMtKrjy5vTS3ovM3XAGpC8nu+zrq9
uHUfkApE73VDL+VDD9GQrJM3N1p56qLB+1OR2trqPQ09pq2aV5plcUDwetQzWTpHs7CKydrcaEf1
+Wtni4bBGsDNYiMbJERV6jio7rp/NWqUAuVJeVeBcrtTUlv0GCh5/1IsrIVzFbPbvHuIIaOnW5I2
WfcehHVT3a+I6NbTH0mD2mRJAQm4vEs/fNf8/rktXHsZHQ6yoF9JgGkAC7HrOsISSBnyOpuaamkN
ChgRzAiMWdEADIRLP8cHctIpoRW6jhVkxhzCiIogNTJxbsmFsxv+9IXcgZX7G4Itp3y1LhNkY6AI
euAY4LfyPTwvi+Tg/9qn1/mCu/6lALtqB+yB7FuNbVclBQCCheRMnP81Ccu4yB3KHZNjtJiWI++v
OX+rWdEdhKllqClwHcbi+uM/A5u3AqFItd5QbzM1a7/OwQZy/T9pQjEWA0ja622k4E7TxQAIgxFO
cSyfw2xmUnWKicofS7Bka6kLm24xQHbWqmBuyos9PKApDOKS73jjGhpjIORVWT2IQt0cHJlb7FZ9
PKRM13IEVhYNT6zv3MEQ9Ob+4Gz0jcMySEEwezqkYxRpyrrZEyov8AGLXTDa5XE94HXjvTT8+3fU
mESTzDrwDd/5jcG3brLZwGersThcbMSlw115yPTJYxKk01iLjfr+r32FOr89/e8lPun5AJF7FwvB
EPESRRLVPisTAozQUXtyc0laO0TemqMOMf19KEVx57J+cqz0QuG9V4m7oOrVZKKmC42oAxUN2om8
gDAbs+aZ/JbP5oPdr1Y5K1KNVxLfav2fYvhT3s1Xv5JwPHbPZzf6duX6xVxARfyC79DmAFKwIeQf
oBM2QZYtnIwpKW4L+NHnJXznh7jd8z8bL2mwsTwN/CeuWDsB4CrPm+M9levmU/kV2Q/yaATfYn74
ij2fVX9pcbvuelBhmoasleueiz2s/1SeRVZ1dInmA8A05cXK4E7BucoxFWSkhW+s5Sv6z9HcWw0v
ym5NLbTlHpO83F+j6/zo3vgj7EYv8u8UvORxkGH+kwCUSd86QNSX/XIvZRAOFVBlIZtOHsPTQocu
UicQipzNJfg3G31Jv/IZ8Dh/o0JX+NJ6yo/HKo9corV0N0Mjx7SwgrhVt64viCz/WFFGvLuV5ISV
oZHY+IVbpgYZ7yMQmoAIM0o36gWNRaQwcM2PdPPQl9jjrgeMwDtHt+yM+WfN152LvWHOGyLt7VpO
HYO+7nTOdPq8hPwWbjdsFE0OpGMdGSc64hACS3XiZLfblAZmPRd1ozfXymiDyIBK+v7tAdeweWWr
Y7wL/Dk2MkakHgdYaPOdBU7TQMyVJZKtPZJ2Uhg6u4fb/qlWx8HTkv2ntNb2qWhZqblFDVjoK8el
YxT3ZOIWOdZNaLpV+FIcXUJ3VdMf0XhNbuc+jV5H3twn2bnPCQRq66nuAcv9rGM6K4bptAGR1w2A
93jQYwn2UKp+DifPtQkNVB/qJsjtIsf0mnltse07aRCQwNteaA8Q6+xGia8tL4HcMZn7xHJauP3B
BycW7eozoAIfCPyh+mdhnysJ3NarnmtGz6ncLeInUJUqE126mFqBEM/72MFXop67lRhs3VTt4Qnk
ZOLxFP1YzXMAi87BN1RaoVtrvJPX26q7HnM1If/9Cicsr9nij4w/9KaxrelwCBwMvaMX1EMaJhL3
B9R9PF14N/EclN2JmRrrSxWM2g9KF9uhn9uHd+1H/SqXr55P2W9hqGP58KPSmiUu4IcfqvM+moGm
DENn602RzdvUhbrFQRLaTkcVCGVo5dryaSJPsUhD+ISHtXqQNc3GF7iODTUUwoFGp2zYda5teb4c
rHQjFIoGGN8zq/3GBc5FeLsTZKaF7eUX4sGrg0SGt5Ei8sXKSXfiBMENKCfPH9nBV9ohiqz8FiRY
Fm43GfCR+w6hiPKfXQ7nMSoW9r+jLqCJnsuWdozSSNi3vmkHOsfSpwZHpvv2t5kIKzzPPguJSCiL
jo0b8AZVWUtXDVaAQ93D3u8dVZnHyMpqK3To4xrhARiJGLf/qEp4uky2SmzZr3B+6HB8MimZfTxe
7VnUr+tVpnRG6uTCD48O7RKazWdNeC0dIS+RSL6pPp9NkTzQnfoGbLzPYADsUWmUKzN1D9bog8os
PZxVoI7FIrypUeS0V9Mo7vTW/JkMgsznRYHDsqh23eRs4oHov83CC+RP2vcuNe9JAHV8fowCqEAe
HxPvPFri4O6dRwDAL7GPMGO6CAc6rgyfLPaEeDzLWLw3SBCZzGLKqLjeAKrJpi+V/t9XZROj+XZq
RL/1bcNJAJObeO3hM0Wqe0Aw3lootOD0Hdq6EzhVzBBf5Xszue3TvZFiYqvquujrszA8BRrKue5g
ZQe77Rxmlu91wRZq8BOtMIM6Z+kuCTA7pJhGlwCeamzgfRPgJLcKC+8KqOh2rzGKHhVWuC0rY7jk
iO95xnDlibcItD6hEriZvcL4C3royOkfAHrKcJOF1vNYDsl+TmWJaVjAqIOO/FRc/4ij4zEp/bFo
FwEFwIRPk95czhkMeZQ7quYJrXKoBUBUQWGQ8dSNqeMVFfFDrlTrJ1BHqPaxnmYnEalinq8a7ckI
WfI9I8+WbUvSFaWlCsq/o3xY0W7hzczxsRR3IGjwvgRvLQxAg8lLlIfYK59aG5HdVrhXpyeppMrC
VWHxPd3sjD1RWl3qwf/aK1/dxZH4UvFujcnOUTEX19vXNXcDIMHSKbQl/gFGMbqaQ48UV4u0MFhZ
epQV+CbIwU3icM87A7wIyQtvFSNDLzhATTYvPoe/hqrtXPiM1uGvEk9UBdrtA1BPbjYqJFw0H9U6
JnhvTmojMuFWMiFwCOw9KKH7ARjCiFzF+5vziWipaA7ko5mgOgLEPQMqHFIqOIjVdkDagpjU2Dmt
ZUrKeO9+bbiS93nSXnqjEzPhN7xk+c/Ib3bkeugge6M5q5AP+kkt4t3yy5kezjpO86WGeLyJzox2
E1ADBmdEV186WYJ612kHY+jjUlsf1ncUcipVyJU8A41nOOw+An1FB34AvKwtS9hmufqM+rmdrrw1
chS7haKYMWwPKMjWRW3le8xeva7KZzWcf6A96QI95BsGkd/9f5MBEOgNMjAMellZ++7mwq7kHK/j
leHrNqLdv+Jj+6LojDYxF8ZvBTClzIM8o70RtWySg+6YXAR1Imi+jocK/wsy9RPb+VjgAJuudU1O
ULodfcRklBvF/rpxa7p7VQgenpBe16hMEzVm/52+XPSbhP2JyppEa4tZM0OcIe4Xivh6CPxW6XbR
y2jlMxxzyYBCs4BYRNQIiyy5jhKwqZN1CC2GrxvvyKsZiqwnkRmTdqAGaXAE+yoCXsik2THkA19x
uiYMzyVEWUR2DwbNycDmupfaP8QA1vVxL4o2ULMEZzbmmoLZa9u7kuC0AXfT3n7+MMH/knY1+/kt
6P6vJUQSxiV6qT+8VKs3sDlA7M4csp1VoTrDBMtzrpUfUFRoFC37eUQSDXsthfbDSTC+zJ2bn/TM
UADx3yiFfrmWY7pUpKTr33rK/kC1TFN1c8OzTTMS6uyej9voOt8dH9Vy+HVJlFQFe2vmwv9bp+Hg
NXUF9DcTRVTk88oQpY5LR+fq1+dqlu/MG3IpYmknX3HNklkIR5Lm7Tb7QYOy/YhpuK9ZUAgS59Mr
LEwBw4AnPDIAK3uoX2zQhEbyBsUC+OhKcLq41/7ccVXTBnmAlCvObxpB72HaZ21aTFjtArvP181K
dQZf7oiT+z5+eDVf/cp0xt49c9e38w+M/cdgjOLxsIcZvfWlapD9cNJ1x6JkowiaSss75uWJCrCR
45ZyA3Q8bliLHaQqHaMNOYvU9SUtlx7L+aupKRtuFm90J5Z9sVkROealNvA1hT484Jz6cfilzXIS
M6Iis/Hd8OULbI4yfZJiwfdjtjyEsd2O87YLxDs5SBpLH7r4cfKDSCK8ug7ZfzTQhgwkwmp3xMs7
o63PT8SZUah0oS4dsM042mWIb0lcZaS5cFGDxTj93pl38KiVkflErjkmVdE4d0TA9RJif81a7L/2
/wHvf6xX9EkrhujUJ41pgTdWTQO9plIxKjIduohwF/TVgdt3f795dKmKkJZ7uUzkAYWjA5Qg3zlI
juXbu6I4EOoz9NYL8AhNXYYe7UR0Raf+Q8UTW3Rxf9pbxbgv6XEnyLEFXri62TnZJoR1cqP6QkOe
/a+ur+8J4KsBbA39dt+tcDUpZb/YW4a3fvIuSDJ6Z6gAWb1sLCjHyUssRb/Bn4KZb3cDRVjEJOj3
dWzo+F30H2jXqUsDvtkVzD7ijWcaRHth9W7xTbrEDvpRiZX76osu0GwoV4btD7hBVGdw+AjJ6R1z
l9//x67mi3VvQbpwgucZ6/7UyT/bG0cm9hsNlytTFxvVfffc4qiNLl496TCLnS5hfzD2EGysfpEl
pietsmd8cU3LH6l2L8N6fBFLQx0L4Jxwl7yoLMXD7cmBpoy2jLqUlOXH7huHOvWcPZuYMOOheETm
KgqSjhVltFpn8bRo3cwJzW9HTfCyfNrvWvEcfr94NUnrgoKLUyOBeiMvI3MqdvYoFZ+Da5igoK8p
81/iYbxowvUGf85sR3wXC09fni+73XVI5QSRuHK7Z/nzORzMd3H3/q+O6lYkPBRY/v7lfKYTrbLg
EfAjK+4ZOQx7ZWP/QVBxzbLX03fWMFziDB6uEtoVe2WbXfo+mpETdRgwKApkOeW4XT8wxTSEILWV
G4+KQUR7fa0+5Dmwl9r0qJ1EVncDUe4NMvc0Blwv9FWqwjIzmwzunhig03wjMqJ6X9C+EXi6OBgD
6w9UyngrQlsx5LbfIzOIZNBXUqqgXKLA+g72qPDmATsc7TAlIgKaMtyR9bEKtMg5Y0Devv5N19Y3
rTGu9JKDTVxCw8h1RLMWGAV2yC211sjy3TArjvOzVAqAnkg4J4xRPIm6Qu1eQ/+iOya1QpWIp0jQ
7galklsu4VnPWa115jAFWFD+m4VrXXTOYHOoVeYPcRBun2Nyjtncsq1yXavv1D08SPmdTs6LIGEv
cKdeH+BghXZHLgRbfJ8NPU1BAx47+1g06ahitKU0oAsa4qRF9aUxqmSWL2cWdN7iPWIvrak5E9gR
TAKiPK+NPUN8TnDeNJ9wMOAW9RmhlC+6k1Z/IdrgEAoIr9A5zUOcIuTYr/P6VyZ2TQPqH8oPgWA1
YPTF5nKAQOdRpXdgYcH5XOx8jY7ZndFXyUYmaYCdlHQp0xSZ2Aj5kliDjR2ih+H7OjjHrkZ6taIi
Y3N6H/4eG52HLPpR8bsDorZdLzGnzU78iIfMycv5BKVFLxxIeTj8JZ5TXWHDbkZiZxNOAHv0tuzG
RYyWy950XYrkMJJ/NwX/fQX6MUauBHDD/KTGFC+QUmMiATAAYwCHS3fSlxpjQKcKwMYd2ySWA6gi
ME1RZObcJlFszuiXquqV6773pGVJ4nOidg/rN/u5kMyffovRNaG5KKAwkc9caG8XTT8omrbSA4NQ
kLyZV9eMfRRaFRHi4rJBSa5YSbhBGyYunViMW3hJP99UfSgc6EeUZxhoc/lumwbdeofd0wUM5H71
zmtDPQ+nRcV8bPje5poGjvNR6wcGQG3BW9BHL+EaCMwoclYMQn95H0fha3nNKMH2jWOjS+ImwtXm
CMsIQC2HSiIehyzV4G0f4cbmePRMVtKvXElmt0xi524L/QaRU4WAoSF78e1b2xZRCIX2Da0tcAFf
JWVdlucG8PMRoneQIE9u6Ucpn5ltlza6/+6mY4o1cK+HCmpl15Uhu1M+9PzNMBmFBhAU2vfApBan
w/Pw9BXu9T3vARRxDsvAwX8uao446gt9xGU1kIlLDVC40JE0wKA2zaWKLg0MlXCawcVb9VjbIJCd
PYADl5qH3upkJTGvHYkld6v0+CwUtPXwXqE+UW0Ae9CFjjSlW6pwRiSVeAP1kNTc+e7BamgYebFe
4vhZYwudHH0IS0pEaliQG4hSj0ePGFu3BbW/z1/CdSzaa1s9ydAeakexzjF0dqi2idj+2wMrbgjw
nyxPRREERAgdg7Ma4NA66WBYpiw4YMawE0kQKcUACWs9o6VC/0ItiFIH6KRiPMiyirucEY7K4aNv
TQcBOIpnkWYqr/gR0N4mqlcSUGXsK554tw9Pl5S5s2fefReWk4jchpZOXa9z42FSD3zJxkicTSsO
I3FcaZ8kgh9IvCeqd9ubH/EoUXd1YgmLgU48jDEAtG3DfafWqSnk30FepZsWt5nHMY/j8AbzYcPv
ehXk9AQmpaB+D6cbePjEoKzIMbn8MwxJ7efBbSEgnt6YjpJ/clUTanC1mLOncV6H7KfIIVX5EzSd
TjWBeETxi8CZFfXr9UwuCFnI7h2rxlO+IpDXuW6TM/l9mDIPiXS6gmrIvykbWM100nIADYcsWVMi
yWwlYsNvWNvZDrTE4dK39asKsx+7xIj08pLqhJJkASSNcZSOAfILJe1kbCgIWmGgF4r3o6N2V0qt
PooqrR/+UUHA5boG42H7ujH1fW9rXg6VLBmUyAmO0vU9RV5SvTg7xK20sJpE4PWEOHFPDS3x4HjY
8z8C8rn/sbs/6/oNFBNKI72uJORVgA2yE+yiewwE8gLkq9cifiBIhY7EsuiZLRq2VkBNTzh4CRRI
tn02nnl+hQD+ciJfDOVnMht79ZoixZvxeFLimLpManUur7nOXTM2XWDEnJ/3iuqKE8MAIgHDpbUQ
p/KRMFoZmaznXeINC9i1mrpHw2bKC+sSNZNr1rjNn6l5h9RAvNmXa3TWQAAKmX2bxPjF7hoqiNwR
Md9oGa6ix7BtkdtHBiNlSqYxEmsQY151MuqzAxD1HocBntwL09t+Csnh6/0anc+wqVOECr5QvzM1
bqKPMEBdBJz8aSf8YOD78P0lUH/8Pfq9wAQmUhLfFC3wfjWJOgwmCvFoAwNsz/dCQxH1qVjv2/xU
PHw3gO67gRqw/aKHpFRG1bH2b8m7qhxeH3Ehg+1KtiHtB61KVksd/9rWzqRP18qaOs9Mo+J3phTr
2B4nXApY2guXCynAjCov2QSalCxrQwnWT2VnznjOmUfqZLyuucf1wSTZqv5TKZ9BSfRx8S0Ge98G
7nIksPgZH6fmXaQW3gjtkgXQDhXo/EoOjCp0sHaHO3HJwbSJUsI/2qX+pncNCfijYwcD9MuHhBSg
sOMb6u/bXWkAPePqHV6WqLj1Wrh4cfVYP6hI6vcHu8ap3FwamfBS0uj5uVv6MEzAfxwfHOKoezXz
Ya1Bz7XbBVm6JzZ9gDGNTia/RmvA0TB7S93AJIj3xvTVQqCcczE2L3osJHAVT7CcodqHBEGThLqy
qW0aZFJ+cGRQYNr8/kU40cE9RKvSJN35kENjTEJo3n/gNAuyShzA5MZnVH0VnmUkc5FHDpVbdYdu
sGmcSHMUDuxRH4uPNP97nuU/pLVlr9Sfhab2xHjinGyX3hR5MHP0toDyVbmmVm/oVPJ0t9oWkegL
c2urvaCte4Y35nz/zzo3lXhjHYNi2aQWAT/b7pOYrOInagkS73EagQtpPmz2814GfrXtMbIb8hVD
sWR5l9U0pnHq+RPfZ1sMMQnoj8dn5gEZoeMwP7i4Mk2jNVG66fKr/ZFB5ef2LQiqufRlw08rLkzz
pPZvH7tlbVJtHErS54mtxVtyEz9m5qmEz6BI8vqpMu70cq4yMihx8DcS5LNL4NWoQ6pnpxDOf37h
vzN2Pvke7ryAMJ0U6ZXwu283riC+2WLQd7gmyssaA3RnAo9EEuU3a1CYUxmb1lWFfhn6IT83KVLZ
nHovO5NELQC2u9ccLj8HZOig7BgNmeYORvBJD7emtakO2Ly3fHcjE1lk1hsfuzQw2+nTH7dcqVQt
vyJX84nEvNXnoDHcwwNSX/MbN6faiP6HacaJAOfAP5CO7NIUSuRM5AeyWAidADy5eYTqUWFw31fB
1/b0RA8cpRjHu0j6ek5znOvM08JTTWBF8kcwuGeUYjkFkCe99ycDe0bKu1K+17Z2kn8TP1kYvCDK
QMiffu0XFbY6DIMQX5lCQz5Ewtiz92HVXlNQ+dpqyiBeYKbtvNkc1dnWPg2NI8Ws640mymgLcFgY
ZfBN23usWVxG/flJGgC7HQV0A9l5PzyDR9mslJwjo9f6fJ28xfobtwsqWy2Zc5paEgYhSpbuFZew
J3KJYCWFSfG1qtOGwQiCKmZCgiQYYLm8nG/fSFXCn+xrXo1NnofWhN3q3IjmSORAPjRM040wgS28
J4hhZbEKHECeOVLnM6XuA/QczRLMe2qycAg54dGK2KEv/qT3R8+Lr1sN1mHBV9lC20haPchw+k42
IPPQB59HGrTvfHoqGCs2P9OMpkY2R2H3ddGVeAtkRYviCYtd/mbpUbHMHq0CcahYm4i6DL4ecjOS
obtnn9BUGhQHAnQ+AkqozrlcVZSmoMZqypsQufZLasu2Dl7d61jrB0+cZcMFFbCxIOEjQqZDpZA1
srDIw1aZvegdPf/rW2rNC7FyNbWp5ngUbTykoTLFD7T8bdNtLy5Nktpfxehs8Z+k5eqrWg84OwZy
GJaoqElWiFCVsNr8GHYiLJJLnMrwdHyLMcGaD3azvhKuc2zkDmJGEQIq4XKMKM97lQ4GmMTaYWqD
z1VFzYI8X2AlS3eYHOygcc5hzqWmiZfjXE7NFp3qpgn5JsyeKQa4aEmUAqX3k1NwfTDzKiU/t/Zr
4qMhkAmm85ThmFtzRW4ilkZ1A8d7iuZbDar3feYFrVZ/5iWNfqLV9ieRIULjVF+mj3CRFfhPG3TF
7qPAsG3V+zYL5tRVhMCERiXlnAkKC4eJ5tnTsvaNEeuw5HSvuWphOnBTu8SQGZhrhVeDXua21tX6
UMuZY6rZ26RALWq0yNJaxkGLceXPa4+94o8mQVpsKIstb/G/z3AWWglQohLecDS1P25D9szUGsIs
ENqC1SeoiPqUyg2IulyQeciVqJhokPeTCwv0y2ezvETlfa1sKdfXWxakjtbQrga34imukJvNLiwe
r/9AXdkNoPM5C+f/QWrNu43vNkKZSJ9EmtmGjA9uss80Lp9iffsCjpLgRdxxwoHiKWqskDOJ9CZX
4AjsDIRToFqZKe0a7MJzQdU0G0+4l+A7C4YW0iKc4MX1Bw5hDtC70te5G0nQ59aRSc/9qizjjMRO
Ks3w7A+OLjA7fHh4Lh+4SmhfJwyakrmIhyXM+sIeRiWNg7OdsCd1F1j35UlJNBoZPdSGqQmw8oa4
8IJXT9lOF7bk1lMubKRA5FQqbes62vb8QMsW9IN5x0fEHj/t0CIJtCxIvoXvBHUXFCuYdk7MyqNE
/cBFNP7XU/8Al+Lbk3hQQgA6I/qYQaESaOj38eCKv3IczrHZCYg8UGyXmhZb9pgNh2whp6WknUl6
HLg5Kp2nSBwT7Qway4j8uE2M5d2bhrLYCwyvQTPPNBoPZZXEK6D9+Z2ogIGnYJNb/LVfvjHoVWBB
EDcH6u4swbMPnP23rs01NPUcf41i6G5KjD/+VsLQHcu/k+7nXaI+uDSkvjQB7iWvDmISYrDIRTqP
VA9UMLLX2bSh9vzWSXJ8WcJbE1TPm5BQ+BidB33IJPHc8AkzXL5QAT/M7qloegK9XwsNF6nOOZ7N
m/EPRse8wqSXiU04vR0qt4rN3gz73pFhHBiNvPO4XlKt6T5IEAHiGeiPU+7yiYgBGafeMxWXkh8U
+ZQ8miOJ2vTJ33jClwd2EFNvAPWjzF2GF1vX104BRayZb30OXsuZVA7mBd8+chb5jZsQ6wMr15nv
+ZyfEf2WGMyi5BUqsDZwwl6f/9v3KrqDglfANMbFxQdVTEE5bNK9fW0MUZWJrvGpe0BcXu64f1vK
4y3rcACdz+M6AchbHmCRSmxUdrOs4mO/y1llCPFeliQty7hTrXH3Ju86v8pWU6YMg5VXniojKCBw
9FAbFG2HG1sWEb/JcYZO3DxdFCpvo1QE3Tcp1+xdUfcZ4+trAEN+8x/OnUhREdc7G6XVTXspAgOh
FAEkmAMzPuztOHqTNHg3/WasDpQa7lODIAdMD1B+rLe3VyW60zToax+Ga9Uq0kTz6TSbxlpw1yyt
vz6SIeVrZe3fmNtzunXtZqB2esSZOxZhnUK4O0/V7g+gLc1UfXwDZ62UfR8t3AXe2wbSAjQn1A6f
88h+XKHscZXyuV/WZAOObVnlZX77vAr7DZXsto9KHcop9bpVGgf7nwDMKlKdA8E4VSvfgnS+6Yym
iZieoagK7oczMW6Hw40haKHmoPioBGFVvm9KpZ73jYxWDI5pQ+urEv4jbAf6Av9+AGpsscbhj3oN
prb7JlObr1mOEI55bHdyTvx/fErkhrkPpsGmWHvKU+RwN5sM7alqYPU6cfW5uNhC/t4qYFdy7h36
l8PPErwAOG4PNEXR32scdQAv9rZevlMvKt1Y1lnJLRLOyiredpM3a/zheGITep1k4K62+guulTyS
GQ7MojmxChh8SBHCA7h4tXPX+eeolUtVr4sIVagMnzPPkYZPTB/3thxqwKD/oiwTTQaqx/GMINqg
lsyTFCqu37vo3jvf+3omAniGeNVTlPCIVhjHBvfKfTko5J/A/PUghF/+NGq/gcQCl/IFs4wVn+Sj
K45ILni9z+F1yqOO9tYDGez17EwhXsXvkxnGlj8YsFPZcA7aoNWyt+eEJJ13GId9CvM+ePWcPjCR
m0v8L0Lk0WaPdysBNYryTW3CZKwdzgpNtu4IKZM0WZhIOLfk9FApl//mcmG8SAX1E+O10l+W2zZI
akDUo+yJBHYvZ5nlCf3JW6rp9zvF0hGriDImmG1jVrRrnz4B+0MGdaD5MX2Ga/LL5yhcc92SBsPh
m2f5Srk+f9J3xJvKmW74ZL2mIG4bT2NKEFzFQ8+7Am3B4HDvqu8fiaspCBJP9btAkHyH1SmRm0cS
GYmD6eg5t7LuWTD8ngGVVmMAO5pFO92smDzk8YVCwagqEFA9VCTIfV3XS2I5SlgBKyBFujxYjbuB
kEgBRRMaMg9DJK93Alt+F2KhbNUBiuZeTyNgA3tOUH4zxZ3vFE2pUtgB/lAVlsJVR2+Mu56YHEoY
kzD60ejGzdXuSznDR/avx+MdsobeTsMV07KvJOx3JkknU9D4zj1wsxf6veLYfzflpzCei8MQQzHC
39PRVsLoy5b+fJj3fd83MEgbFFOjYLxCaFt8dqna4EOEsXf4eGTSgYdiR91Dnt0NUsjuzHlHTFLV
xZGYcLshsE9Xd51JYF1WZj1JTgLFbIU9rDM5UBrnSkV+4vcVOuU9d8XXTPLhoU9XfZicFpgfTqeX
TKI5/Y6w1QY186XC29bLDKmbfWRH/hInaxsN7r/qhGanNr+kJsiQzNKNCgLCyI7kEMT/fzEf1HWy
4xuFdwjNZt93y/+9BCRH3Dn2IjMzDh836FS2232TdTY8kRWYCcaSolceDJm0W6s1S9p1pH20Oxqj
OahgE/9Noa/skg+TZhqx5eCOi/KSJSrOS6/kNf+SnYuDjiXfPC3PNeA/dBrcl6tpBMdq5Rm6XgN7
YV2W9Bfv3LCt/mJJlAuL5QvUu5ENTJditjzB/2UxJylcALhHcGB/0YFweZLmt3JV8rFkr0KXMsPU
EMw9AmY0Xjlo0knt4JB9jiXh4qtwygFv+dN230LmTjTu00G1icC6LJ7pKFcJsLPHZVU6RFbeG7NY
lJ58ld3BbprhvNQJdGVwXVgeq/oguA627gQidAfilvByMdaUdeUrZY3I7IoRCNeLcrhBdd5wNGtg
5PH1QoixKU33gD6eVaXFiG9repEDt97xFUVQO8RgZ1ffNVBzrn7SGD0MlDDnrpAL09U62wQ5tnvN
KNUZsZm3kwNmr177CG0btZBdM8xub21o6lTqT69VSvA3ty4y14AIxPQJJamDrvAA8nqPZl8bLiol
36JuBW1/VxwoNKBApweSh7TRMbiPwrqIGxRZvDSNaShW+ZO9eFg/QQ7EPsGc53xED0rwonl6bssL
vwZgLde1wnSDslNKrzT9AvB7UohSawncyfKRE5fuN0w0o+/aSy6Kdw9PoXXGuEvBcAxbO90xz1D9
DzQxJ86BhfpJXREDXPU9gS7yXXlvzSaykXdcjnTGKSHEmK8nYB+3dBkTDEbtGbQS9YPJWW0apLaF
ByLH0cZYidvX3bpmq1kvo8LF0Y1WVZb22wcBGIWxrRoqQK7nvFry4um3PJv5N2Y1zAp4jHiqJoKM
WRMe/e4ZC/1CGcfkOI9NJa7p9i64NEstTaGpTdf8NXOHBeZWyECv663tIJikY6PspqGdvNn0zk7G
+6aXWclM2zaMqQ6tJYaVNX3l4SHsFDGVLO+9wZK1bCpmMqtVwIBVLGHqGeia3f0zb/IQ5YfPld1H
578GZEQt5AL/MTDBAHNg+k3dm5qfxUSvCw44JfiwJpOGTzVkVqw/a8+Y7FQXmx5kl/GssNuf4trc
vqCQymY02WvGXG5/vQDkAtABZJeB4vGqdxRXVuT9zScCXQVtCDnc6ueedbzUUDmSxovokk5FqTDE
/mhVhm+pXt0jA5lU3pxl2Ucmo7zqAePfG2bpjjFpwltezKQ+ErS4tXq/1/jb3E9gLw/OnfuLrglf
lH+wu7HptTBZDoS/h7W0uEDXoXE48+srqg35hk6UDC1ClGqtwBOdjGIDZkMVGF8YZrRXtUjKH/82
D1O1Rv+MCXTi1VqWvIstzZy7GbjQUI7mEuEkoHgnh07MQc80HGH5y0OBr9cl5t+1bknGVqy6+rw3
TLnXvdPPl9S9jZbYbOeGK8iQZxzWR89M0nV3eOm5GPLBwXI6pkbyKnGNawOgX3xObQrzlOjtW62O
JoAsjDwzXjpuO2wn0l1LhrZECzMw/OWmGHNhAbZC9LDim+dbByhApu3WtRJKUz95UqyTUBZwtv/4
0sIQ+Pa7INYSdQOdrzNfn3MzxfzvHF19LhMiN9e6mn6VE1OqAn/bismwLp5GmNqIMen1Gas0MmQx
XqwyA2QfLtmmL4Q/v22ae6c+KZ5QmsL4YU7op2D2RCWpqi9s/DfQ+JPGm6N5aZJe6gFqUQPuWqTr
g3vfpEWU1c8MJTu5D34HbqvQgF7dUpAZApg+3+FdnNgGLDDXU6RPx1zfZqC5ORPJKpn2GOSJAiXo
5Xe+dQ3msLS0jB9nn8SudRMJtk64JcRqgZnMr7ZFGAJBT2mJuzmIlF/r35xNlr1QaOWTmb3JzCH3
XFxFTzF1R/INXQ/Ti1IMBuUS9zPyvnSqStaLRgHAb1P7U/MI50CetLvmZURyRPRnKqxtVBgtfl1E
c6hRc+iCvWtYnIDQMyBxPaUB71CgC7udIamMoe36EgCrQAp2MxjIWCp7km5hrr2qLtvsyU1+e49e
0PaJkTU1elNaHsnYAUzHkDrZXq175LbyupJSd9dUun2FzkcAq0hZ3ONT3SNRWirmdx6qt0a+YClV
f1u1F2ltc5fIXSFj+VeU/cLqvJQvm8PbyCzIpVbFM4qOq8t+BJdhFHKixUlPUX46m2PXl7XVtzqb
kljGeL6IL/U387F6AJurUJ2EHOedRWwD5yCusxwy/e9y46I+PFmhn5Am86TpEHFLvdgnnmXf/MOL
GDFyMV5gIQBYBadQ/BNveZlEAkDfmP33Mk8bJ0HqKmB1yGtBBv6xr+EN3FG+0t2X/HiwIskaX53A
QcJtmGA7YhRLt4CRRooPQowujeq5eqlxtWK+pHT0c07Dme/5ZjXSFv/Km2Jdoe7WAMofKLlXc+Ve
YFg/HTQg98J8ny1/9XuW0YZwr0XSDNDzBDYP70pBOi/TkEFMNM2R/sJwHH7MNRUxh9wZOSmGMEuZ
UqUQ0j/+gQwq9XokdhGM3oxkg5RxfKasqdZwkECdKriQfCoB0ZKL9jFg8/TQkRR26Cw9TbneVZz9
ffBecGHw4KhnpAdyN2ZEs8481e3fFSXDDNC4vdgLcx53N39LjRaksFahd3O71C9GLSg5yORAippi
6rG30B9Q7LMILYZuzs/Rj1zWWgnTmbKmM4w4tlWm7QuIiKGhgjee8YyxMf4nFhnIHn1dudMq+h6N
B0U1aVXh4nhq0IlDGACJq/8eBrVw6ydWiNhj8uvFmlGJR9lKHJvPJnKx6ZdR1YInCQEaHi8qoz/5
A2hXTfV4oR22P1n8E5uzAKqS4ZKcXwtfyKSA8YDHE7NGD+TT1WiXZkb0uptl7bm10EkjKdN3OVw2
hEMWYcHd741NdXB8bkXepvBseB39Nc+zUBm8OuLgnwfuAsZnKA0SKXaF4tX4eaOc4yBAcwMMc8tZ
DOu1zZcmIEzYAz2PG0Yv9hZNCi35546BQUqcy6a8CHIh7mwMhhNVjo//xQb2fwfCh5MiYwMY7dFk
YXH3fpYtJzlKZd+CXvK0MUzrjEyj+4XjbHKcDXzR4GeCQLVlOnDIN+h1w39FZL0BzGvmedmyUsLo
lXtwCql/TM4xysO3lCbpYDbiFlVnNiRgZ0/G2NpG8cwVLWDsoJLHWazR4i6Gac2FX5XFKLGyMFOy
1Ly7938KWsCmB1wfMohoDeNm68e4iRcT9KBBC3D9NRWwV1hhQjrhfQNSMLl3gFe1rAns18iHlOOf
hwrXB9kEmA54xvSQR+mZvR9Wc1ok9pF+9h7K9IZfX/0KlnAFDv9tjyBzYAVrgeEFGWkWgkagIAc7
0WSwWdaVUuHM/8vn+gN4z6aijUKoTyHwxYsmyIw6zqlrerep3smNflC6763HFUQjgHF1qaBZNpts
TMEYUCC/CmicCS4tPJJrIcMoLZVe2NaRZEI6Kf1CBRu5o0XhofzEGtXcmguGjInmsQ+oYr1hIjBe
Q5DZFZn5n0/VsmJoQO4pzfiujyvpYDr8r4Fw9Oj+YFV1pACV4/DEHDfCf+0Ke5QeDvrxemnVoIoM
4QbwfJyP0Q9Jyu7cftiJH9PaGtQCIluDDw==
`protect end_protected
