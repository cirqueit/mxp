XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#�l�x*7���<(=˷�ؒ�,��xt�>�G�Ӟ�$� �o�L���v�����)_�>C��u�e�Y3�ӹz�Y������9O�`:&
�K*����|�o:���5ESd�ҕG��I଍�o�8����@2T��)Ń����񄩗���3�Rj����گ��<�������x���t�TԤ&��gD�$,��
ς�5<����;΂ p�Rt��$�����eu�M���4>���s���&l�D�zJ+�1H*<1��e ���1�N��k��s탌SU�*����_��{ތ�=d��*j��Y�Rg7#��Z�S>�_�2U���������Đ����OY�a�m�~�d�9���kiP�@�f6�6h>����W����m��Un�u��v��'8":��Z��߱�>�~͔�~mW�B�IM��S�Tl���	����ۢ
�����R[=fI���e�J���\��!����"��6G�������]%������d
^T���\����ݍ�|X����Ԣ@��� ���$���΂Uh�F���ex�G���8'��@���]C�#H��Ԯ��i��� �v�:���5k���+��~>/�M̔��-MY.���-DY�&MOg��$kq!�JO���i%q�l��B
�bQk���}�B̯y"^�I�V��uDR3f�Ap�8��@a� }0L�!�m��8�2�xOf3���X�$���(�3��<HR�Ʊ@��D1��Տ�^XlxVHYEB     400     190��A`�27��D��	h'�L�Ҍ��q	�ɋ�y�M��eu�Q�.Y�U�%,��,S��VÖ��!,�Z�9"���M���S�~bK4��.�MA�}T�]��������1f�P]�U���sk�n��b�^�K��1k���y�"��4�r�gd�Z��y0�vޡUgk�[:+u:-���4��:T���se+�s'!�a�&�{L��W��G}���1���2p��Ek��]�ɧ�.���5x�gT��nH�w�z���Q8��8 u�t��g<]��O�K�:��Mk%e�[e�1ù�t{��(������e\��%�6��C�/�K���1ݞJ�0��i@6�D�K�G��Q��!I���vbvJm��3]m�ŷ�ci��B�?4�P���Z#�w��XlxVHYEB     400     140%��eW'�]z�LX��Ž��Ah���KB|y���J���:L)u�q�:ߞ�|�V}��0d�"SjY�K6�^�O�Z�$U�{Hd��g��t��A�ó�����*f��c��Z_�i*-΄H�<�ΐ�.�	v	�H�7W�&[�^>�y>���KcO��u� oI'<]�g�N t]P�|x�Zm�.N�<v�0`��˳Ļ�����읨ӌD�Xy�U��'��x�r�$F0�y�|h���:a`�]�cts�3\��5�ޟ���Z�M5��c��o��h���%t�V�ܓ,aצM�ޭ\��+NEa�.XlxVHYEB     400     130�����SYzlsV�uʜ"E�[�n�qֵK �����|^�*��B@�n�!�s�dH��+!*z�Lβs�#��T7Ak�GS�)K�G3�x�����`ΘeC��}yѶ������M��	���xr�]�T3��;W��x�_����v���NDS䛛5��$`���X���D��#L�Ť��P����q��C�C�����M|H.M_B^�d�]�k����=׃���]� ��D=u�N��?�`�i>y�l���4�ԣY3!�l�c�l8_�%L��|#vRU����G�;2��%�IsXlxVHYEB     232     110W [)N��{�e4�� ��@2rF��X�ǜ�g~��]>��'�	�3T�gN��%o�
�Q��U�q����N<(?`�1��?��!:'&D�������g��9�BǞ���H1�g�t"����|�Ԭ�E�eTR�B�:�����d}mUр4+����]���l�w�2^���<�*r��W��������mW�.8�y�Ѷ��,%+���t#�X��2�(Zd~L_�u`�6 rXB�W���2�Nl��w�BڰiqBcG�WCj Ur���