XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��kKf�"��}�$6|g`"�z��nVVGCE8 �.�9+��xq9�ݫb��AD�y6G��o={�5J�.���5��W@�=�y3����،"���K�`.q�
���x:�r�'��~�a
�AG"I*ޑ(�`��� ��^�4��������{���fGճ�Fj�箯�����s�8��3x�,��к5�!��x*�_S��qsp��|0���PK��DR�ns�$ �VA�$�#��-z�%!+	
���RC `ٞUfA�Ľg��e�<��a|��U��[~��%s
�Cp� ��l���Qj|�=�`�@h�ft2����O��h8���*B댑㴭��5�ArJڐ�	�F���a�\L��7���?W�o.4q�w�7�qc�66���m��:��{�w�.C�À��Yi��y��j������%{)zzdɘT�|�}�?F��%�A�_N�L@���~<]֍^�?�A���Jm�z���s�me��|�7v&!��Dp�p�g4'��AM!�6.Xҕ��u�ut����Lv9���o��>>�����r~ީ3xB-��({�޴q���lw�g ���bZ�c��T�-�N�!h�t1���JŔt(G�����[�2�&�-|�,D1z�/����x����5�șEϟ�L�J�1�TTLio-	���/I]��QB+I�g�P�(�Bw��(���\܀?m���"h_K@�9���4:#"ˋ���Rm!E6����nM��S)�<~w�u�`4�XlxVHYEB     400     180��nV%4	G���m�eM ���2��2 x��KeZUԡs~�_欆�~F��pu �����c�Qx�3�Ry�qQ�Vf�g\y�+��q���
�>�P�JXgz�����GS�dI�?��8rR��lX�� ��I��O�>��7(9zDjN�=oT���p�Z �@@���:`ώd��b�j�������bũKWc�YB&��d�1\�+��}�3<����1�Wv?{٪��$!r�~U�u����$�6�SaN��/������<vc�!/M���F\��&�W���l+K�	��n���)��s��w��pT@t�������[D�hB���:�X�(:s�s�Y���A@�^�!����r�ʮ����i��zXlxVHYEB     400     180�0�r�	v�r�{D�Ǎ�h����u��d&�l��?�H�T�.3$ԾX��Ξa�)��T���k�~p��N2�a�����\
�~���v}\̰�<�����j�f�lp���f�P�}�.4���z{U�7{���!��3O. '��52�W$І��.J8���Qy��Տ�~�v�P�$�";5��>�܆@uֆ{~���p�C:�5�(ԺX�`4-���ln?��sӦ�Ժ=��3��y'�'����|)�ii�q�@����K�w�U8����.��
9Z�I�\@v�\����������d�,�v�Ө4��JK�B�G� s��_��K�W� ݾ��&$^Z?�H�[�n��U
��>Ƙ9-XlxVHYEB     400     170m5����!��C���os>���#~�8׼�{�,oåL�_H�/
���� ��J��G 7�a܈ԅ0��6�7Ϙ�)Ї�&�8h���,��~��<Y5�7�p*�P����fa��汜��{���$u�OuO�{��tƭ��^�<-���o>06��{��/�r"%��^~G���}��*�5���,���w�m7�N���X�8�ע%b���[l�� [��↊/c�`�|�C���U ��P83����
���XL�� Sk��e��ޞ6��E��՝��������t�=HAKl6�)�$+<j)N]��%'D�t\��yL�-���˘?��:5���s��w�Sg�8un���l߄�XlxVHYEB     2e8     120�e��d�j*�Ϛ_]p����	�X�<�p��˼����v�4Ŋ�З�&roL�ۂ_7�h�n�vjR���Ө���z��5c���g�7@J3�(�W��혂�7m,�K����V���x�{U��D���z�o�ط[�+q�J(�[|lK������P5�O扳��.�;�bl])�Gu�t�7�Ȋ$�YҴ��`���H�e���ሺ�Į%\�I��S ��q��_to	��%�����#ޏ����d@u�.�c�0�ξ�������߂��M�F����x$���|&"��