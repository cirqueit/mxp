`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`protect data_block
8rF9izYALFa0gFH3Y1uqsuEqGMlnecW9W/+jC/hznKLloRHK9HMjKXvTgQsG3z3iEGELwzd5UacE
yjIkA19msJuaTYIagAiheCjKrWz72bWjQnDZAkDL0TAC5auZaDSU5zSwMbUwoSk41bMpENGwhPld
0tm5ltuGIwKkKjCNz58NJHpXSGbCNOYSQovBDgYAREwIIl2ZifCj87wT/eNDbKJ8664klJC7Dv7G
q3kVZ+ertQColZRucyNeqvhQNOYesA2Q24KT3oC1qNy1Hbr7/hiWF2//Z8xrdKOqJfSTOvTnssh8
YZdyhd8ILmUyK3h37NOvSOgkXih/lrP3AhMLINQV1RToV/d3KqsFK8EXMQAXHG/bU6TWS2lI4uKX
87/rsrvFKSt1SOkkaypDreiPFHYglYD+x6gReg0H/S8mz9cAnTEZ5mRzRme2Ei5iZVVntD9Rlryi
3Bb78kEnqFsPCsFkf35WzsjQJaR3W+FJiZ3LevojWAXXOimx2iRQRNDhceeG0E40e6Ko9GKBFh3n
iyeNnSmB7kIJI5p8k0PBLtw6IdwewMV7wR/XdO8TUI9ruw+ILmuYDoOZ7OyM32Lgo+2QGkHcrBD6
bRklLKf3Ofj9AO1fhZ75zzVoeAj/nEYnIj04prYv+XMugJjSgbpeMFjLw3clqiYK4dV/0CGn4SWH
pxKoalvWu4VnImUjxF3aJk01fcFh0WpJY1l8eOTcT5gATzYh2qHKJ9FZ/+H54NcjczBhWOGWXqZz
xPWLvdR2hFyLmNXc+XpyJ8lvQ3SqUGhwdy33LlDGBnDvEVzpztKljkPI8DjOyBrIVH0+kWeAMuGl
ajvesc7u91RCcK9O2oaCcw445TYpidPdgS+ehmrwzewuouUP/TFhVb1qIvtXRDZLF5MP9oA9j3It
q0nA4MWb3V47qWW17USdzWAYov9oWQ6eMspLvKg/IWC3NYoijD6StHAdgEIkrNXUz3E4rzN/Vu9C
1xJ5UtbDQF5KDC7Nqhx/i5kfzbdYqD5inxZhriyilSEb7FFW6VfJHTUtehCNL0w6qxkPHB5BvVqi
q1b2WCHrkaVGk7Z5oN/BX4IpboGoNKueel63TY2xJl/P6JoQcTSdmYFDB816xmEFQcJ2ROUV8hoW
FpuvMWxKecGK3ImLJQvbrcUPuuPlKOEePtyxEFdm4JUUKx4MlEPKjRknePzZW/4D+zwKvG5n2O//
480shjk56IDZ1F5LygS5pyATVHOjn/6yAB78Py2CjeWsg4iqFHrkL5JMbsFu7qzjd7BL71Y886df
dD4sy461agrzGckIXsKVyXNoisLz1VlrRazZCwnPv/JCBfAfvA/VVQ+gWjs/zxK56Ix7YpWVF1YN
TxFK3Ti3P9GmXC1AbVfhYJYHhZZ3UAFIbLGD+U30hGdLIjG4oNTqMmq8HVNTPAWM47KgzrrkdUV/
By0mn4pRCBZgUDbRe/WodAZPGeXYCt4wEoyaKZOLvoGEYSe2JAVW9vif5omEZs+PQ5KnCm6N/GEf
vr9Su1ekD6fOc0JdwFI+xBnERBrBkvGF9ezN/7gykg1gvmbjCKVBHC3dzsvFvpKg3sa3XuLAE1cg
+BCFALrkxcKcoy/u2/lw7TssUw7cdXEzHgEdwKSCVe09Ax5I4786zdPR50ZJucPI6Tn5ur1NtcQb
NW05os4ryDRSBrdsGBhRA7eFmlQ8/TVvTO8xLJW+ca8p/sC3ijs7OzoErQqGzPkuOg8vv8CtKfF5
RwUbmr2QPdATEyokUgz38XHk8uCPrIOhWJOsRqnqX5U/INNKmq7WTciDWnLFanpl/NiQRAkVwY9u
HVpPBCmJwn1CLJUmD1waRi13L/IlJMtvIH+cpuxnO2GAJ8OkkxrRePrrPb6czPcLXofQURI66ZYy
Ii5LSa9agfpaSbrn1Ayigsj7f1hr1lEoDuspqRSS4xXXA1ZVjCM0HCy+xF2HxVuz+S4AjaaWW/Wp
uRCe05fbkVwez0Kq2bqUtlPdwI/kc0m4aT6T1bBRyIRXG/cBqgXWdGHZ3mMul1rEbDSsfXeyyd6f
dXpSAfJ+9vsto4DYpRYNdxCn1DOYD1W05NS48c/Uwgq+R/wMnJvFDyAAFcuBHkWeWvdUYt6D6BLx
NFGRqlVlTAX3zmfid1pv8BjLjBOtbP9DkCY+IEqbc46yKy66slyZrrxulzUy/Xt/SO7/Y97hoboc
YUR/VffTPBhhgTpPzurYMaow9rfDJy7DWoffa5ogf/9Qyi9w/bNyV8a+qJu5h657/8GTOBzI7oMa
l7S1zw2/r/OSlsetmUxFsPsd/jrRiQhma3/WGwV1CA8GF7DcOJSnBWV2ESUixFg2IOgrXw6+VB+T
xxhGaTy09EEK90ai08GZ6UtTfrLekpOQgACJ/Px5WcqmrzgGonF7XzsmVjoKsQFOMGDuoRTsxATT
ykeNtSPMQa7C+yhe9bNgzyQV+QScVTyDMpiCVfEgEId+bgkR/f7XY/CXI0SkcfNsy+fL7CXYBG2e
+SeTmYWn6f0mtTq2u4c4UL8VEI9HblecyCSUaZNNEGxlj+EseaBho0RtwG6q93uNG2MYA8L25qUQ
rpfiGESVpzphIeQuAZG2YvfHarkXcQLEx3nHCNAAnbGFQZBBC7ZzxVvA4PAHjOUNWsP+XilApu6x
vTZJ0QY9WNfB3jE89RmQfa4nagy98x5YMr+OzJ3iTpbBGQPquRj9yyFAWktvvqKocGEg71Q3BUez
m4RrNPZsAvL9CyZGOKzJtXQmbwBLTVLFAcTyVeyvYpf004wA+l/ABDQwQfCkkZIcC9Zn2SJIhaES
FlROsOWdkZTJGFRIdMYEP0ydCQgd+vg6KvY7zShE9AfVTpcdmeXOziVYiFUOVAKVq9UOuDBSzHUf
CHB8gy9JGLjyaQR3bTlVgx1VTO86FhHh7sxmwuS0EycY5nmLpOcAFo4Y2e8PTm3CHAXnDZjJ2t12
PTFyfTz9xqQnguL8fh4wBzCHpurRrDyu8DeTLRV5dtXIZv0P5wo0oDVCpdYZYbRuGF0UO3DB5zzG
Y5ouoV4U47MeqeSs2098KP5Gbn+nx2B6kemO4Ro/FQKJRqtI9/lq/zeg3p1CZfSJ6AzeQrwDLgdo
1hQMxxuzHsnor8MJj1+m0sDNfpY1xuVVJlbMWQngvZks0wdk7PrwlpyfRedWPSGnvBlhmAo/T7N9
okWLBOPSSIlVnB2TzZx8VeY+NhE/kk4fB9Z/ljlISq6XIT51IP3kTnIs4Wipn4yb5HCEUcJwJGrg
cCLHscCGvRu7gDVxUP2eY73ZP5/rcOstwcd90WkJfLoHi1oTkkHysmUTCvIBpXAbqDA816RG1Xph
YuLAdkHU6g+tgLRTk0kbfmB/Wr4CJ4bvnKXWnuiEaMoyWfL+BirRQnH7aE1CEzsAfxYEVwYPJ0cS
u1tur3eKkmlohtOpCwgQkhVR6+MtdL6NXEdKh5Mq5aGZEZZzsMFU8N2jjgeL+RWgnXvayIRN8PuL
NCHphXS44vzfDnzCDlqoMJLwjy1nHKT7yn3F4qr8TipPpn56xtiL7LzX34IE2ZqI40az8j66ahSh
fz8FwJ0mWODa+yClrQdQh3qBfcfzST5ji2hSlsG20wjx/ckf/dXtXFWVjlISwkr6WO4lA+VUeyiB
yawe44MIWR7zlhrmeBGlqImlzFbgNhg8wat/tcRwP5RUR8WqKQcZd9EHwpaGykrCgkXWguzv0QVu
QhLzOZzPUENPkRZPUfFAu17GRwy5VgR61kdhJfHY023mw+SjKTP1V3O6uZn1gPzFWUijXsXdqR9B
UcZQD/+O+6oRY6Ld+mrt03+gT8G4/KR2WoRonmlsz/neuU+E9alD9roB153/ikedYIZGFmuWatGC
W87B3XAe1Hz60iMuCDbP+La7v+RI+3Gjx1AlNWoCn4jll+aJ46sujn58KzRqmpHtV8vXLzaUBZ/v
5GH06GKy7fnmeFXwV5nXnqeUhO1zI60T54vDfh79jY9znIAoA0ZnipdicjVVIoBxB89z+QwW+Xvj
6S7iaP3sJx8xc4TqFzYCXD8Kduz8ubEE2pXEqYaJFG2TB30ihi3GfUZVJuzeX00lID/XccBNm+Sb
lxqul57ITr+exUI2GMu61H02gtUDugMHfp4F87e5kmtdIgTSPjO9cnNA0rb7mQp2w60rF99REYW7
/zg3VCGPuAnv7P9zyvdVK7QaZhS5Is2/RF9lCCxKJSwwlctkdl1GlVC5gOiywlp7M2wv3Hurw4AA
fh+vARqczYu4nc8zgnqK9HNgHyx3Wys4J8pvAvzReLCRSf9QSL/ARpti5FvPeVVDvVLmdi1Qy+/8
WEPIk64yi8dI2Z+iUdyn9rG2VpmUEvdiVbuKe0Pntcf/l3piGEFZpmv9yXJaVh7Np8VI0xCMPyBP
gbprVHfzcSLemFFwUPd68nCxZoondmfQ0JcRnzKJVBnpLu/64p3nH3UhEVqmWL4ATCaGH8gldYXS
88dndnk7tFAOHON65t3dvPI0chxtkrWMKIEmn/QnU7+dapnHaBxKdQsmKROihHaN447IqYgcpoEp
cm2JY1VeK8xmVwPsj8Ne6vZ4AjYIJ15tt/ctKk9E/1uBeAs5tRINY24/mIf6CbgZmWLKbawdLThH
tgOiredYqxVA0EM=
`protect end_protected
