`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13920)
`protect data_block
FAyx+PMq3/GpLspoyvV1VQPxmsJ/VSe5cpI4ASJPJRtk+fT9oQ6ScH3KMIqY+4rsWuFJOUh7Y5yd
VThltxHYuf/nOX+vPXABAGudsP3Npl+rwsyI8DPjmXhk/LowwMrSHCyErrVPFolYZysJDbRwa7I1
0tsN6I/7xrtzpgCka3QmqmUAzmQKNNI8eJ+G+/450N8vLPcAdhAWRfzZpFmMIKifW5GHn4CZ6Xb4
1hohF11HvfRzMjm7Ez/CVVjFptDurBt+WVMN8DVJYGGaZpMXzTrlMgELQ8z0T+oHgol2cgIRMH9V
wPdGk6aXj4jhxNaMEfESG20F985dsBkpzTkofMBmzdkCBgmn/8yP5783+hErgL8Jk3bmIW9am/ru
8usg3Ru/sNwwpQ0wAEa+ARLC9ZrloJ4w9YY0fBVq5mdtZi7jvxZm0wOw3UGRpsbE28SQymMgzumI
pWz4yKYaiB+5akPNMm3yYHoDdrZn0IYvsN1bflrfJRMWXYJyz7vPJdvXK+P63AjkPzbH6bNAPLsJ
py7Z+sGZem4pCyQaF8wHQ0FYpdphE16e7rqO/+w6BVEUtQRhI54du5Hx/sxQ7WUYnxcC1Rweu29p
CYflmAw8Pur470OekaRucOL4z8ev1pTsPm9nCwcbFT8IEZDxMe/gY9bztTTqBu2w3FxQ0Yt9cX6p
l+YAnrjW9uSWvBJeLn4GrywTlz/9NE6oFvofEm6ZhYel9rXl+RerFkVkoUNeE4RcTPtvP6+rM5d3
FjbZYk1mK0re+giFwUwQLaA15avCmTrFVIlt1lR0SIJMvDY3eaBMH6PYbjrTObHYV9UXT+V+kNgm
ELsz0JWG2hCCvcs9ZBd1AG8vlqBgR7JbW2B94/bnrdKm6/j36OwIJAGwLMyPHZ+A9guWyLoppod7
U2mqhtkctQ/E0e4phi7I9JBDdA+uxYdf/6d50wWMcQOn9gZs4kfmeHU4or4jeNtHL6mYhKMQEIWJ
9ld0jGBc4IAQVy05amvrpqhrV/nTzyi+2QagkYjEPu6jhFiXs6j4mCKkSKGeGjXZ556aMO4TxtLV
s0wgIDsFuSSZdObW6bksNc50jszpHLY/32oLzkcQa/3UWZWH4Bxoraai8sqHgIAvkEqHnfjRPo30
dbaeIwJnL3zbmqY6o1xDzFPBoHP6f/3ImJRk6cDsULV6cX+TEmTGRb+2hZpQrwKKwTgB2BFs8rc4
GEuW24LaZV4JUIKpqV55Y2kT3XXkmw2Eya95koqA9FB5uZ+HqZTYbfchVPh8mb2tXXkWceW4ihdn
BBLuqGJlvRyGnI6i9yj3Sdj1tnPozpg3kTwNg3e0Lvz8gxQXf0IuKa+uDMhDhWz/CrRf2cIngeXC
VduX+2B7fj2ySglEYzJWviOlWOMyk11DRrh5x4WoSXdTPpy+JHbg9dhj6wvdAMaw1R9Yid610AVZ
02AFbF6D2lO+HyWWzsN19eShBYq7JcM1V2Ieuf/QnlfKQuubv6fZ+cIouqlcDwuSnhcsv+fG6IOL
UNZGTobu50vWEfaO7l8mXvc4w5tOeYnTFUA142CLubefkOJ+xeTOfxcHO6nxkisdwfslzanO0+eh
4YYEE/3mhiKjxSroqdiXYv4JFBlypY/lOWWigwSFhnLlvuBGrU9dqBHEiqTmYXdDcC4eKMM1tAnZ
au9Nj2FrmplxiJos6OnzCYutl4hz75MG2/ER7O/nn13wWRp3zZdE7aOEkXsOO5yeANgQydofmR1Y
hmgr/UwNlvtu1dNO1LqnXpykXgFcOL03Fp8Z6HlvRGFG311Ira541+L56kVPvHnHPs5m3PPqx7m0
0pGMp1ZypxIMvmZC9/R6ljrupJOs7Mo2AiXaMENeIogzILEbtImf55uuxIoXWQ5mBoYNNZ/RgjG6
aW2eO+nLcebCryzNumwApIIhySm7DXM1nIs37dIvVVNs/JJjumc/hKBcj3pdU0FNYW34ZQ3OmpBr
6N7WR9a4H0Rw7w9A/nGIEZZy57JhPDCqO+R4g7JqDJv5cOg1R64ho8fLNAmTSMerxpNDDZRN8IOx
8AcKF2R37fpqPVQegs+AIKErncjmFwBaByJLv+mKvNVYe3uN36AKTi6yoLoHZeb9Kv2mj/A49AXf
sGkhnMmnT2FPOZwDY1WrYPq756bWzTLJL3wRgRhKMDPlwVq7sE8UAc+AfkCmdJTuQq8MJd1VZHDl
1TDXTv52jzoNEQT7vQ7Fyw0YCxWI6OPn3AbLQ2cVST/dcey/Thf9l6reAO3S7opTrJZsnip+rcgA
GYBjMS/Wc4fBOk5WfjoydtpZq27ZcdEkLqZ6CASWLt9xIMSR04y/NIgpQa5I31TRsMKXP9FkELPm
gs1X8J8nukTIljioG+p3whaXEopP7SNOudHUkDbATJmlgXHTehhdRTBt0w1BMi1wtXIhxgDiYzqy
Kyr5/kqjrYH4vfvcl97+M5cDc7/a6cwSvV0vk9/OD6F14NDzSw9XXzDbXZmWnb6yHfFD9MbFB5MP
hkeNUUKOCiIqf+KUZkYgwkDBy242CRpv7oSx0fl7Ws3wEq2bfyaYDOkRG6LZv+fI232NuqbRFPwk
N5B8PLQI9U3FLe9x5qqqh0h6UYotHzAeifjvlsLi96Btmk0Zmmm4LdJb4l11iUvW5UMpALopPbp7
NIDlhKPoZFPyKohJhjsirRTq6Ew+xfTDres+q2Ka64TrCvB/iQl52QO67crqKAHC46wF3SxjTN3P
ygomVbd+273YMgpFqOJ5CQ420n4LFCNm3gAJd0DfSdRPpOvaX8ZFPUqlG4VzapcHRvEQodF3Rrav
9fZCqaZlt2x9EheOeOcJ2amzn0r0NVV17DEG32D6IZCnMK3DVe+yC6XNpQYcffR+3VGJfvFOp5N4
n2URin8VrYdmVBWtT6HVeKbrXsvv7JJDziNBi9EuZOxAKBW243MYtrlvgOmWw40bedRCwcg5nbaf
xMwzXzVSaJlJpCTiWvL/TZZN2MRLmhW064jIjpn80cgQ+HG0tdjvcnrTNKMu9IuwbhQn6WCVZOsT
YBtF0eCE3UHb8e7dZlE89oDCB0c9Uz+5e7undrA/ZhD+NIo7rjPuYKVL/H0/WgI+YdOPnBoeq5GB
x9VWyVeBRRx7Gmxuhf1ClyvPf0apGsbr7qyvh/5jAqW4wLmVwkJoE3oIijL4DBeb/Dn0RLQLRe2x
D7JlyIfgTiBd/QCHhJ8FHfDRRZztFt8FqLblGlseC7ucuCzfclbX4FsaySzDGtf/Tso+c3DxFsNe
yojeQo6n03khVGXz1MpZZ1KSVpPpx3+hU3RlivrOYQ+wt4D7K5T3N8Oiegov6H1bmgK/kLIWv/Wc
DbT9M9C5uRVzbTJ1BRlbws7hj9aMY2hUhCB5RmYsF1ptz7hcNBlECAYOesjmaiD9tVsm6YeVQyJo
Ys4szMdlIGkkVReWBYprfiH9k3LjSCV+cDGrpyzQmFOAY3zrQjwZYa9pXwrGxY5AzDe+qfJaVRu6
Xw+edxaaRNbMryXVfMg0Zj+Frco11xHHtCCrOF4vGUu10sT/+g7WjFZvZENRfY6u5IrAhz7vHmmf
L4jqdPKQnO1eCaS4qyKBzmwYJzS38zu1NJDFLN3Rn3kibsNEiWt6DpDQXJmPcrnoMXwBX1oFI6r/
GJrOZMeEb7MbPFL+MSBIotEVMXTXEq62gkSdGFjuxxi2YCZqKmn5YxnD5H9VpaDRTSzWwYh2KipJ
w+mXciYYUojjXiuC5Cn+F+RXXsQ23qk+oTd1Tp1zS4VhvWBe+FyogfrPn/Zbbf1iL46/ad6VzmP7
2HjVanyE/vwXZStMM/QWkBLJ7lkzGi5qcyT9fP3UaiMqduERKsZKSTBxMz/7Mzx7Eq7IxO0WuqWa
rEdLpr5RjW33pwSWyDObbvxr2CeKs66Fg6DrVy/FYwDIjUn25kHFGOf6wkvQudGmYSpfVzyVGOl9
SlS8WVIQC/kbOTijv9K9Eop3LawqoEhG0bTzyr9MSzGC6Vh/PNltAjihyL74Awe16j5Gha+fsHU5
q2DpQyVXjhTGQ+UxjUNi3preuhUgJLY689T7xzlgt+DrQdOZcvYCmqRcInZCaZtc4RaHx/jA91JG
kqQhRBb+szpyX6o4boue865jrNo6oPFzD9mJbuLa/ZZCJgzSarsz6OoNHlhed8w950PBEvA+I6y8
LImd3OCT+7CXBjlKWs7vqPhpH3nfo5+70Nv18qO0cHWvV/z8AmicYdFVqMqP2EcaerBHK+1e9xfI
owM/L5h+Uq2vXcisjTcvu5D5mU58WF2UOm8/waRZq8VRJhsNwISg1R1aWinKFsDRALB6AWqjCSxy
CXJqoYpUoeTFpLjT1yATeKmez4VqnWPtyb42+IPYvlEuoAcdSJFd/A1zvwl/YT9qI82hxOG4BhMX
ZvcZTtEpMdO1F6tH7wpCVpg7kpfRaToCPesMNfkIzueHO6RC2qOhrQZFaVkz49CvuaQIL2dbKezN
t6JkGviMDHr14ArroB7O06EDEO6vk3xjGH1Cxym/d2BZBhvRGbU8+cypeUyv7uo4QctN5h0+rTxa
G1r1aXcr2GU4t3np4e4k75PsuA1hyJi3nEkmuctB2aag1MP8qswdZQA/XRBT5vbKO6dLHWY6MroN
rWkUi6pQfeIgc5N4EXwFXOv3btf8C8CtH2VUXuvBI+SPttrTzOD/ngAyPU30ip7QNCvUDx+NxeIm
2Wy693jk4P6E96TMt8fC9C0XeeKEznP4atAA1vrNUsk8JW//IBe/3aJSE7dWWmJ6+C/F4PNk2k8i
5MYNA3M1B3scFjVEtT0OloIiOPuz8j3juHGxTEiz0f1txTMRHHgdVMoKQvraQwACkYx798mOi0WM
pCmmj/1ky6lKDuaI0DNtsbgt/SYdfYRdbPlqekdJi4qPfBJf0w5exMjX+N7zluZhCjLpKpXwNu24
SC7iXKBAiLBDh11xGFeEQtShF65eHGALnTmUGTpv1k3z3xJ5VcAmJj9ixjS86mK4R/9MPrcupzec
lqtn4qdlLuLcHwOmkAJ8JJ4tkAOp5zH9q2k5h8eR7VQCUOwD7phKbej/vawS0ZjkxIIs01b4PxJh
tstkRK0NcnM3wEbgCdDtappxRba3Gu2XgXSQ3zmuSLdyv/sdDgsxwVYUhSoe+LTxk4ahCyperk0K
okhi/ylyud0LekQYwVsrO7GXa/D6DqZ6p+dNmsXXvOt+iQRfU2x6H9keczmyqgq4QLMWHG2o2UEo
AwZHYhYhzADODv6I2q5iBENsh/MxsTB2suyYMafabp/tWR65yTWVSGJ2VbmmX5WSo3JS8MDufrNw
U8bB1mxCSN+3fyRd/jXjUAd6tU19WBXDyQAvbbwU7E4o2S2u4/a91KKQ5fEAt5XSLfY81GnfzEtt
i5ySX5rq5g1zoiqAwsEBwNF12GeyqIOEgfsamtmtmis76+UuGcI9ZZkkL+uhkQdLwW0FmB0iQZ0E
8pXT+AxuLCm5iPc3GFlFGKjHJJ33WqX/yeZcZj9vlCkjdNUg6IE4rtM5NoFx9Pn+kqyp0cAdRVtN
X8PzK+Ji0K8SMt9vI9Vj6KmGCVdxeYzwgzf16AcfSql5BNVp5p6k7Nl0Fj0YlEXPF+3ZAlNojBtX
qUZcRKRGIlwX64ZMkLwAUPXYI2bcOKQD2gwVm93usd6SuIqxTx9umXWVPSGethx0vkY6La1aN1hF
m/60TforXhwolC7Mu2rYLWfFetNX7QgHIykmINLKoCyIci/qrDMNXDqv/FlpDE1dXEu586bGJ8yP
eUyVQYH6T3vVDwmn8o0E2Hy8JbDMbEuItXDabe46rHVs7kMXQKvALH7VvPgieyce0GoOImqDHZF7
Lbj9q5oBSOWt+Q07IVbyxcBuhWtMnnliOYvMN051XWEcL4z4UEUYUi9M/TJyBR4UEQ4j7T3ra20q
d4pyJ+nUonwJmRYvCsEjmSoR1uu8ell+MEvMBg3eMWUECTyygsoZ/KzLitsf9oRv2Z1CxFMe4mMl
V8iIcbwWv973iu9SfE/xCJe01u+Lqv85olzVjImyfKYXIs7dbMjvoWS8i8TJUJoZ+nESdLb7pU16
YdHX+hcaLNyC+stFpqkh82brDQQ07rOzMlFJCQttGmihJVAijtGbaqzMWXO1o0u41ZDVeNZaxo4V
r7vUz0ZApc63AXs3D02klWglqpNmImQMeT/vbl0ZAr+a9l/rRnZpO7L1YRbKCARC2QY0qK0kooi4
V0we03SIirhoAiKFujHKqgELCE+pIXVtFFPp5VXhjEw/nC8s1ydgCJ3StaoYI27LzkVYjqmrTcyZ
k5KOECc1v4LsdVvqxVpPSEmVgUXKsQ6ZA9F+6mU2qgsQx/6pk4t4jHUA7Ak01ARh8pCAiAnL8AMh
QHJyH3X0NIYmPy8V5xFSTC24NTpF1uTbcb5hZlTVTPDEC5HARwz8Y7tKdBw7OTyxNb4K/qrleVkx
15BAYwjF6lQkan5HbzqSjXc29QFw8CPWfkMhyeejXUzcXc5PYSG62YXGhoho0PaFV7Oj4iFuaWxm
iS3TdAQpLfI7XrF2h9vV7PZ+5ppuO0flQdkLLyRXbQSnZpN6HURcjpsqbIl0/3NUpzYrSH1Xn+vq
wFdiW7GLlOibkUJzQkuazv7Vy250bVGzqd6O0og7eZ++NwIAKDIwyI/sWmrUF9qQOVBoNfAvfJBA
hWci08gmTWfDCR8Gox4MxNZqkIgTCTvALiI6Mw/E6v5OFNziAngM++2NyMbJsk/r1HXH9/2PY7vj
YAZOvtT5j/Tc4pq1TurqFeWX0Z+yEZ4YkaY4cVNoSTzMex+lPHnSm9Eq7BYZa2vfrVGxrr95MoNp
8U97fQGcmioqTRUr9we+8C3IgFntOsRgabFTflwy37PPYR7UkcxapWW/K8KLTNe5UswNdW+PlwLl
BbA/4NLLcBY8nV+u/tkVWRHwLie7Xd7L9zu8w0hqaJDJGu/3/1qiNX6D/4bB7jk9OlmGwxzRPSrn
gWNG1bcPa9Wvq2yE6tY5u8BTOU1KqqNDBnCcVmGF4EfK+EoW5tQBVQckCQMjsNBTsRRrElgZaHwX
LJO1i/VBR+adGkwhZT3X9JK7Od1FYlpJEQFM/XynWFZgQL5i5SHW+rs74qada494U8P9iKXaVeF2
ZcGrDYaq94SEwt1HRlcdugTM4VNWkMnTzmiUG5ljcq2Xs09rwUJ3GhKsY5MtmEDHUo2KO8Z3qUa1
ghgniw4udQdwOpu2unBU1WOrVsnZPT24b2KpljTqGCVjem9ts9bcyiCpTiN9WVXDLNtZAacA665z
kLxEO3rNULbgxS9AMcZpWAvTFI7gp9xV49dgDO5dVV5R6JY8k1Ug+ohOk/B0M7R3Lc3QTLMaHxKd
cITx/h8G1Xqb8rgvDmdW0KBioHIkcSZZSxuELkqcHKbmKpE/uDu0XExMEsi33slKAifKfMXHkCZ8
pxF0UGfDWOZN24PTQN4kwboLCqWOfwxcj8sZO+yAsxKGZI03MBgCftmhQnqh6aLpr1ocZMHYFnDN
2yCqxQ7WATmLgcyygrSogzWfTx/4xz0+3ZsnV21Wci6Wd/w4rOtPEk/My3Wz7Zg3l5PGqKqb8vwP
4WSSiYX7cY2ONZN8zitu8LTPsPuS5w1xAXlW3S3u0vdGUqQ4hHx3Lqf6FglhkqTcTLA45Ydt0EZW
O4zTBy6oTYeGGdAtSKw04NnQ4lkcXmMNKlWemWl03LfHi19+Rc+7nMtTc+Vo1mfY6jcWCEEcG9Zs
lux+MpDCJc9popSdFijD8MYm9ZiNk71k1cOAOiVZn/IFiaWPvwrODIY73fI3ZKBtak/laXTQBiMz
rtNGZuh0LA9LtKzlr0iUyHVxQYc5P/hlBh27Lw//YtsVmXRZT6jV2H7j/sDU8XubeVYkWIxCkKis
OSSs7s8PU19/2LfWon+IvjQLKLtPoMzhhmrpx8cdBwCl4Ah3OelAkzxv+J35VkN7Hea8KOOskq2i
asoZN4UTDhMX++Zb9BXLBzI5grwthBDOh6+vMzYvpYvKWsw1Iy0uOGpw+Q0WjhNwaXg1neuOrG1j
cCDEc9gHQPDYULdfFKiWMNeE5yhAj70+JavwtOzCqDm+Gs16AbldBzmuNqgfKnrW0x+fZyRlgZnv
s1p3JFVFV593fNDFvgU8Ttea3TJu2Q6DXhrf0HVDALgdhxVWF7+TegmWBM6n/yso9S1BKWs2spP2
wvFroznaQDn8pi+PTqyB56Vp/n7Cy71TbhGpuK65StJtK5017kwpIOlGJQmINOTDn+e6YJapCUpD
Fh0BVsroWqAyKNDHoEq3dZ1TD1hQc5I4Nl6aTfhLC7hwOMdiC14qumTeHFDLikHwkfsox2ZoOy55
81tAYLrKd7oZBBcOOHccaSX49JnbteGcJQJOl7n2hHEvOz49vT66enV4h0SOErkRy+1SwQrY5qTZ
Rz7gue3ypCHE7m1tzH41ZK8VT2Stqobznj0T0EJrmM+DZpxm1KhKbLd4xZ5FdkrVjpWQvCeQuDb5
/We7QXBzJH97fSrW4UY7MWXjXHsRfehF53cFKqNKclvmcDia0PwyC/zrIifut0EsAzPL7PCgJ6y+
6aCFmiHJIwZTaYos+ucmW3tsRl9xKpE98CESzAlV6aDH4KEZ0RRnW7308rVaRec9DVgfoXxDTlXg
6MV3LE5OGnF9PhNecMspeIAkXKkP0PtJtmn6F7xQ3TYlq4FgWAc1wTW639POiCYIFBuIkHw5+0ad
OmOaeEK6ZxRv0zyvXmr4fBwkRYiNVnYyapCHrpa42zEySOzQ+/FQRhH1jTJ4QcXLCU0mMz3G54Po
iaZmyDx7gChucmO1oRN38CrjGFPQjbYK0D2vHdq9sYw8DyGapbChhQeeloTAZ9qZyyQWa7iS6nLs
fEjbRQP0NcUYHgOl2Me9tzjAgWf5JNLSo+SoBVzHMOlIrR79I8dMaAtDlP3rI3N/IyS4rAAZVSfV
aAmF2K8DK0rJOABoGx6XtNACCbwE9KRRi0rNdLUaN9fQTOXBD/CJOsa8SwPYXJ1NXwA3ZqPkWLmB
pdZJKK590crzTUmOncOlzbD9w99lJtjhlCps9R7/anIFm4oAbczWRoR7IJoMTmmK0rEa3wsWBm4/
eBx93btHU1KaeY3ynExgnrAO/nmy6v+UBUGdOyNREZZjh6xYtKKs/VGtSuf4wiUvV3oSShv0P4t8
05cVy+HqnUZGzjONfEVfaO0z262ZTAVSVOsH1Ks0fk+PYUfNpfoIJyVgvaHfI8uaqUwhpD7lf8t4
pIYGY1zB3xH0ojasQnnWlBB4arwI2spyUpuWDdU95YP5aub9c7u0YmvIPZNXvjRD6w+Dbl//o1m7
guF2w+OqDrtiecsVmmiLbZw4MekaFrdYMXQA27ZvN5o7gnGhZw4xp20Wb4HC31RdibbVNV2K8YBQ
GkiStA+5fpLB4s0Gfebct1/9F2qXEvBPbitkXYKQHiilX/TpqMaI/ubPTpKJEG1bG0XhCEBQHbz+
8CqtIBfHz8wwjDWsQKUvma1l6C7g11/lIi8Rt7aRcSxeU9O6n7JR4LCBoHYaVmTAhB8T6DKC353x
9Epo920C5w2mCqDaYoU+5ss45SZX1I26pcuEcOb8AQV5HICLkiZF6IDbzF4ZccZHbt695g6lXY96
9NkodxbozZIv3dXqK64Np0Kig4LQvH0ovuQVKcKgdY75mLGjiJGpIh/6Dfwoy1IjE5kx+51MhR/+
Ehhd9sjjmcG5Huv4+dn7OPytJVFHO2G4KPjC8wdTyhlDhuiobTaQVT9qNWvbTY9prEdA9nYlLMcB
LL0nmlPg/ythgUQk7QG5fHa0mqmwOMyMYNYqFEfrLxZq7iwLxPDdotyoHut5kbliDfIHpn/Csvse
2TD/4cH4sPHin4c0Qj/c6HdqEMAQSYZEPmBugdJC6kM1Qg0Y/Tp3OJjaAs4MTbpIidRnhnV1H7h+
zBpv/FF4sshHuuQ6pLPfT8WOTdpEU9GySQejq6O2+DzLY1fKmLI8+4FKtg8FQOt6lnQ6ZWRYFxQe
PUOb+FZQgJMuk15LBX+iOwVfjbSh3rHkr32gMqyxRAL1FbKjr6zzY5gm/dAHknRvBmeqUqe8q+79
61+OsAAZxVg/PkvCzZYUBgoYtT4qadrQezHNp4QEy9qgQWmuSeEWYBHNj/VId+CqjaL09eE6GRWq
g2YOnt3opnfAmKBUIlYKW+lxBHR9oyDLpNEaQQrEVGNooUtukDf78upwxbaoKRV+EBmj6vP/wr+2
A79kzJE3qyZKn7M4LhI8tn7lkeYtxWVOnsAwDqEFAkKvctkDVIhJ2lSG84aRonM43R/GeBvnZgAL
Nvupjf2m3uTL4BsI1MjChLM3MjW65RYBQvTAKFejc/ey4f7q6+xM901FqykI6Chytmz/C8n877Ej
XnmyWA0g+f4EOj4XKt3gl1WRcR4WjSTyt3Z1JuVNButtVH2a4PFl/Uu/pIWnSbuTAWElSxOFU5wK
xtPsPTsNva8AqJyVqXV0Es4A7oTShUT0J26BmTN65DeSVtYdhlzUu2VdLSYMLCCyEeOoV0KfxFZh
uO69psare61Plti8geC7T1wYpG1LEXhbjZC1c0iWDhDz7FfajI5Gd5kpN9N0KSMx4K8mDoV/AnQ8
JzJO0Sa7E25cicJAFRjHFyJjkIHZ10by22/MXx+m56mHpFYyvSEDE/yH4keOn1wkE/Iv/7TNuom8
8+qMCrnK2DcEqAfFeUUv1Qc6xnCKTEohbaVEFnnhQ1wS6/fiNugD8CVXR6/SE+/q03FG9ShWP+cq
5NvqtUGptXp5s4UI7KiP423tZaMPAsvC7Btec7JARyD/bC4Z+grSKltJxLcJqJwTV4dKMRhXyniq
mNmwblWezEnbm4KUiTltwjSAJ3uYe5M8NBvoHa6T2bbNt3LOu+08J0mcZq1LlkcCFFPIpq3H5okP
aU7Qqnb//SIAQFXWoZl2dCYv46Wv/NR1UH/55alXYfQw2WM2FiLIbs9ObbGw7bP6s/gWhVskP7du
gEmuH/9PtH5TYLaTKWiBH6hGv/PZWS/i86dS3L1XnwAoOAOMpjrrZCU0bG7brZtFiznxdpb2Tg/d
3L3RqKfH6jXmICC86iSKcrYVAeXD1LjfpJcBUl8J+/lOUe7/F90Zs+lYazwNFY6O1k49qd4pFWt1
T9Q16SQRZfzPofpbj8WkPbRVt1v0fTcaEGyCRw0I0G0Qpex+rUzBOokZV09jZuS8Gjzl1DHPJ9cv
PeMGI33O3odqqbzbLKAdmcGX2PPLEwd2CIvaQuYD1iTX4veb5fs/9U7Eq90vG/g4xyZs4E7gCjW6
PBqZb8uzAB/3/YxCTZzu2U+E7/Ya05LjtVu3sgY3TvjS9qhYA2iohtihxRpt8jUmiC6KOkiTkNd/
xX/d3cKVHUTWRgYKn/OZr1WU6b91SqxkkLEccmItFkKT6kzaSTdoiQhKBmaV31MpN/KN6s+Ds59v
U2aLtKesnOUysuHrbOgASFG4L8tM9NITYD9sbHzlWAGC1/lObcT4ggOwcfjoHDix3sGUUd2EEes9
bbaritnEwe7+AH+Amuth5bLLJX+dFxOHVoVtTzDFF92OUD/xYPD3303ysUyEFT4sUsp1nbjBN4RF
HjzOITG32yD/piFzitKJz9Dga3oOgehZNkDaIQdI/p1f1Bs5hzHUPTZnnaF8Cp8I2ZxJZcSiUIeP
9yoFhz/CHNGPbR2js7itqWGbbvcMRMUdkxSdXY51rwlZzmEK4eirn8PuJsrCqRwhZgzzVfo4dLwe
OROZDIfXdxCc61jU/uLjpGNCvPvSkgzsOgD6LLZ5MFGP/DssF4myJtLWTJfbqoqZJoduse7gONxd
yik+/+f82QLdNLIb8etQ0RvUQ+IvY8CpMMBXt3TIG9hqplLsyg1TEQcMoQtjWD7ENB35g4WuNyaz
ECMOPaQp3gpc/1Y6Xkepaho4ULX7V6DuIA7Z5b77eWOXbHZ0FBxjniuS6WjT6XD8TJBXwqNhXC8r
zTkVnRWdtbWvNVuSx9wOYKcW5H4xbBy8af3bi82d27zlL3ET2YhFpjFWLRzyIRyfOMJtdIEEWs/A
SsDODY03HWRvlvEZDjyh9ZKj6+8ubNqY8CkND4KaZtJgk+69OStqeJE/2HG8xyC1D8xfvaex8rrO
NMFaBT0Nsd9OinL2vQ6OUf2j3rk2aY4YkH/h38uJLRATUQZ0snJ8RJVZ2UM+iPLVZlDJjMpkPbSv
anJNfEyKhU0xlJ98ZQ2exhaQIZr1pGoIoSl9kFEGvEHE7rE6CiuQzPFPCSY/I3wmFFbP7LwlN4LI
ILs0o6y/zklzRJ3u1xjmFHsOFdYL83f/WvCC+ZWwx1V+Y8BHyVBIRfQp+5hQZX9ULPcF70kAAMUE
7t8lswKSaF9e6apsba0AC5b8B/PqtgMrcLRjT/5/gVF8GhqquGogqMch3Wg4x1h26OYdRbhqOpRA
1D2FBtfdwYzHy5uyKQRpA1PnyJde+MH3fjIkqgOlfdLLazqEXzZlRmz1RE45v1qzvJl3NqgUJS48
rTDIN42S6GKwZcUpcUbgaLUkUiuGV8FmOtm4BGoE5BEF2zIIkGtuP9FUA1gWmJR91knRCISDXyt0
QHdlsCHSWqF033k9JcqSFrNfdlkBGHEJJSArgcBAcfcuWbDCHS3CP8cjRKNoG8azP/3P/Q9O6G2/
UxUuc+on50IXL7phpFXhB6LmJFems2zVposqzpvhMGX9bN2FJxEeVe77NIvRL0wBig9s3RWlub19
ayy1zL8UfnZd+VckKWl2Bmcz0L1lEXyeZ3s7pRKKYpi6p/nLOVmIhf+W/lN/aeGY1NppoJfFrKDd
0vq19LBtjo0c2D4cwcrb2r+Vs1sJ6K16zPTeoUGdA/MCiW73W8B+A9p3YVIJOkT0+nixuKcRjnsN
1j62LbESPJap5dXyHK4YV/vXTHcdG+2VBjjopjWBKyr9VCygGeZLtKbHCt6KIr7mJjHxILaUTlQY
ACkX9WlvQoYD/oH+HQLNhoVWFfcOVUFipu2xwg6TDUd+oepvro9TP/wFoiAxnvWPy0wnUiBM26fA
VbGRDWG3Hp7BvF4y+LM8BxmZoQCTgjMHsleIHrdYnaO0/DQaUZuDrU/Ixcy8GWtFZs2OYGExz/d1
PQH7n/r/Y1J9HtJtQYIdydb4nEFuY7ofp0zXKFkTDHQeN/qZOaKWUqINWz323Pdebf3RgS3CkJOG
c1SlDR7PqPFe77MGatter1oXvDCWMx+U0U5MtbJwAsyPpSxvE/SavXqwwCVJFo8CG1tbGhnTxeof
L5ABv0tjD9IiiShvCusbLl8oBEwU+JnRz4+jGEIzR0pk3UzNEY4Q437v79vEAIPI8GcaPyJx7Vt0
KPLdOY/bBmbu7hosgtxKXc7VybcuQa78OoLA0YYRxXg3egP/tqaGa++VZc38iAxBj/61xJsqr96A
UeuGEbHZPhVYa6HRdms8W8hw2eIytkOLJVXgF64pUFU7AuZEw4lzMGE9to7uLOn9woUEVHH6xszC
ZrJfJyDBmoT+FNoAZspiERyZYJdG3Ik0S7wFtXg/wQKB6OMHVbdlitKbvETeB1SAPsH/Hu66ciRW
ZgLXrLm+UHYvNej4kzgVIJ3WwLhtoXnwwblrLtkyqE+C0+UiJpeudE/LajeqMqWOef1s3ynUSQM6
DZYr03FfhXn96Y8u4vcfKsWwwwKKGT1sm6o+GhmVzxor9aM3ZIIfoelXXSwkF6imIU90Q/URWouY
73CHODJeu7TN18uV/XYUOyaUgOTEMq/frX5dA0FwKQdgB60b1wCKPFCEOdb6mi5Nn6lNEe0m2K2t
Zn3EW5ugtnibINJ9yROu2lxeyMaEonEBaNtSj8L/cXRRMxh22kYnQjkd0QFQdv198Tpfai6XckEz
gZZBqCyGZSpzs1gHe+44UxwrKGCBGcEnr5nF0o/langXopqhOeYrNW4KGyRKmsj+Y+1D9zkM5gv+
BxEtBdxY25PuTw0VT88OFBaoWB9KEUioxIFILgdeXEqLTIbE/DmS6hE3A/IZ4T6FkMKSn0O7caHc
biz+t5x2K+2PT3Bfp1Prmrej4kdVwG6mWMhYq32tarSUzKBX/1dOc3y5Kf2uiLFyeWDP5NG0ZDE0
wEqa1oPEBiMIvHa4Bj3LYMKk5L2pRYPSm2RgKUnFHciL914pgJeXk13y4tSDSy5FMCA+3myDF50v
LPLiCACB1GTOlu3aG9cHUGRnOvraRohsH+jiAIveKPLU9w9JBuwzwN59muYuPTrpNdASVSoGmCnh
oCvi3T8eFvELJ4kALf91GlDQRSg/9T8XZe4t4rkCIrAAPJBCrFtVhPeGRw/U6xMi3cixoSbUPt6m
hZ/ZzM4v16uuasNAxQucEp94wdp3g5B3lkZux1V5kOAStOThpzyMgrX1APPMBI3yqlJrr46pS0g2
K40l/Brai5P6fB/gif3nKnK8ndQ0In12Y5NIthxZ4JQMuRi5sxFBALbK38bdkRJP1VqQqqXoks6h
KzHYz1EcwJG0YPlz/R+mOeoiBtzOl9SQcn1tRYlH36D2iZXL2MPgpA0TNlS+Etu/lIKhu/beCQI7
BfPE8Fe17wTPTNYSKQVjw6z1A5GMdGM+FSsxRbmwxLl4zgoUPriWYXCtMaeY5CX2pqZPUQy/cMZQ
yKszL4Lu934VF0+hVNDHJEo6FDvA8WhRVb2ad0c4g6Iymjt3VHv1KWha62Uh38p/bh/6eR8w6rha
ZiIO0OnId/T5yA6GZfl153SiXCy488sdXvTQ0Ir3qBCBvHKkZL+RG1NkLWHKUYUYM0RKEUtVyI2x
m0B/IkAUzB4KRaQ87PpaqZaQjock1CTf71yNK8PDRPm1OsSe9BwhDFpj5Am8bcoeEny+/XOevK2k
8DDzS4RpUgR5Y7tB7A2cO/YU/Xf53OuoZep4VS3QLTZHdyv2ogRtKEnkzCwj8xT0+MQqAtXFMBjC
doLZWx8Ut73PhUMho6i/im1DIux9Mv3wbAdO1x8AV4Ey/+j7wnqKIeEm5dTSDq9llPuzSLZvQODd
tR7d/Bt6s5LLgxNMVOau2K5+1N1ujydTPGc12v7bR+Pjz2cOyxz4Pmo3a0QgNnOcciARK4bHzvZT
Naek0Ylxi4tnnG6L38UWXomwVNtSfZeKjxpkOXcBLiyxTUvmLARIKPssvghixWcY4/g8OotIWTu6
Y/CmzmhoQFko5todoIESxsM5uurujUE2LE7FeMb2QcIGDh3nQxYF+OMfxBpEQR1QRQWhtrjv/Gqp
FARAYl+x6qnCAVBpcmnObCaPTmw5bTJlXBrO0pMi/hYCEEGniPkpHiyweos+1nhidoIqyNqGWAtL
LYwz3TyuViDdomAgO9xa1xFfzHtWkTpucCjoAlluDrGGmodyttkrdhHD2+bSN15oo3cc1/9SATWp
A0xa6dXay1OJEptYlQaoXqK6KV6YQD+9S0CbmPgvc4xbooHmoUThJy7pwahcbW1iuN29CaK47Rna
hLz9dwZ4Vgjzb9gUvf5drMhclz5Ke7SxAWRac+qST5lzFje3b/2YBV4wkvA8HIDFQkIRJlkKhG8z
izEu1a6GS5BfE99m2M1IuZqOD9O4sHygqx1pAR5hOeWmf3lfpjtubVQSow4qBgRm6KKMFJV4UFru
b3Ri8MHl1vJCxtrOpTXMb+Bp8a+x0sbFiKFAfeq8r0VcxT4chWsG7yHlyo6PQ0784k/0rRjV0Bh/
TvohODX6BjIYNWVunrJSthYB7GWnn1ibB+rJqjNvEw/XLaECG8kUAIZxdsIjIsUvaKpJAOrOL376
83FYxhhJzYpQm3wdW9e0UHlFYA+XLM+icpHMBMgTXF6SjHYuRWn/UIubNkkK6jSVWuL7Ap/RE3tj
6ptylwtTmXgr52YdxbnAWIfjN3CmNZEW6hEqv65UMYgud6uw/IN9QJpULlS2H9SkhXmRMGS1Y7MR
LWnDFEKe3DFYSsJ8DsFkjEVQoriLmlR6XKhadYRFFmj+nEkCJMatFhLWBnHJUqluAgw1/BJH/51S
m29LcRPtSkl1tCbwQZ2uP8gLW/LNpMNisQSAHFlq1sHXAYwZG3CZKj6f5NfOmT7YzkPGv4xReTqi
kjeRN504fAxMn0U8OZqFb4xDQtX1rdZ98E/Lv2uj+m4Fu0qRwN5wBh32FQOK2HcXNiJp4VHEg/go
SFuhCtXL8yrgjFRCT+w7NQg1Pjq/R9q3tNjsbOtCj6nKcKyVGB+vYzT8jacKVv2qRpZhcaVUQkKc
VSL86giKwTmtXtMqemXzXovqlgi1VSSuEdRR1e5OONQy81MQPpVOjEjvmzKgLfS7rcbVE5HjxiMm
xg71+InrA3l7Wri9+83KJf67tjjuBNaZbAPkWWxEzVif2M6AyV/eSmE9le/fCCR8uLdQCTLyCeXj
DdvR40fQiMxcshKbKMXWL63UG9L2XX/vgfuQdNRuwNY+jUam65ytQOsvnIqN3wdVrbbI9vjv5Ybc
XX3MR4b75Gf7xexZrZR1XsE9cWrxjgCMLuJiTpGkBamt6li+4mrJsiKWCbXMJvOORXg1dcf3Iw2N
3P3wvcon7z+15vBiflyuSKLFG2QgLbLUyB8BKKe3WGmgE3Lqp2rOjkup7XWO1zFjr/KaFL22uX/9
BLMCtDxYGmLXGjf8yhrYwQR+ADrGQK/Ci5qSpuDLIiaaiQLhGnDci5l9o6cEy0thyVzS1EBOmv9Z
5qW2T6ttFMyLyMkvIBL1jKXfYJtHfo/qaXXuuQmgMa/Jx9cBI9e1I9Q1QN7mesgZrh0m3Inrx9QM
oHCClAFuYUQdBrDz81icgNIJkb60n2kbTW6MIPri1XCI2nhhBl1agPbjRXniWIsLskkEF4sCXnw5
pAebOEDu9704QLRT69Lcrkiec6mwfuxEm8rebhMAllXYgbZi1dak8FyzkTfNUvf2rKvr37gFCw/s
jksiKLjs65lI7Z9uf0WsCoEWZhoWb8vYHJcYpBu1NW9BGI2+zgXoOHX0860bq3ZZWpNVrbrDErz8
XwH8DnYH9NLLzUJpzolPeklFa8RMFoTDbr1Nvclx99kzub3hCqgjdxsSuZ1bzjeoZdj0cM4r9IJw
Jh7XrLcWHYDP0CnkXX6rrhbg7cY4qS36fbH8/l3aths+1hNeRRSv811RE73EQBTaxU3UogBTlne7
HEZ5/OS5F+0/UH++Av+TaQ4WZ0g6uZqN4eeWLTpDYsBf8uj+DNHgq4heNB9PXa2wgx2e6io4LknO
ucJ/J4sUbuLYpGQaX5pNwhHgni0yQilVdpKMFRxVBA5GfD77VId4ce3OSzJKNdFHmhDzFaKecK5W
ygVdPq526Lo8ma3thGgY76wHQXdB7FEwvxGcS07cbxvMvICWMA0sE5cgEmp82stJxsBMzccsr0vM
McYdj4ZnuglPPrnvCJhoLEh1dDiWgE5lY8nhN0Fo0mm/xoKBr/aLLuWn8le+ndEQccWfSN7oX5Xd
zNsswXVhrQUzvF+BR4SLfaJ1qfEl227wKByO651xfubMW+gfZy201REbGjbOvZGJ5OQQQBhj5jur
sWjXWHAAx62PSQ3I8WjevKIhepxZMWw1WNqmfRuBK+/vTp3g4/UJqbHxcS1jzNbnoaWrcKp7Zf2p
JvsuQVGbvoRhykjS/QHcB81O7dthfOQZ6CKpZ/LlcSNv29UJDPFhA4CzIaulZDqNMWjKOmigHNc7
q7WC9fEn2yxVPCiMJcwkAxYVB6NGdHn1R6rKLQEKUfu5JUaW/8dOzxy5KforewkOWFu+rqmD6W9l
rYwvMGt70Jbp+dEiuxenLUZ57FDMvrgCHza3TJFS3gYvROve2/rpbyP0ZTE0JseyUaWLZoZOHEa5
vuKPnBcTjlqSnY7VgAqz3H6ofhhfW5oovcl4MHVQNfUn/DEzKHAiFwe/HGq+JJNrFEAUmZTrwKPy
9g3lorypZL2gd65Yf2fsZAk4hZ+/pqBLxyvitDkirqJypt5AsXarA8CSv2A9WbKGyOpvclSy5B+9
S+V/0gNSe2uxmHsuhQte54e/YFVoyyIPCL4F2xaXCTK0JtdDghVnjgDyxJmxEZtEjPIBm4SYA3J9
aex2HXfuDdQjHt96a52Uyzw/SSvxtx6LI7fVAoHwesSq6eGwCugkohxOa5gOuNaf8s0zWttM/Kmi
KA3ynYdP3Z452v1KNtmYam0R77Kv644FHnswLxU7P/4gS845NPBbKlQmN/CwHjJoaBVx7pyvM1Uo
hQb5xVyew/F/7i7eGsYJwwAv9cREfendZNi2vKwwVKpHteAsdSI6SwDDHHEfzQ7o/UEOSOQdEURf
59UCHo5rv9PXr5WLms+xfrXH8iYS6uL2aFzPSbp7qtRHGWMjlb+OYAwLjGAHsT0iBNgG9VyxGz16
Vp0b1YFTtiGeSr/x4XVcsgJVt5L//pk3RNT+dTBpp4B5eg47gZGp6TS5hFuVD4vKkLFu0FgpxtXU
sDjw0VRXrXwW/KJAN0mMlpMCs3bUfZZD1SzV2XyJpxKOXLKemm4WXFfs7XCSsR29fybkEdLcO4W7
4+nJOJJatm1sOiwR
`protect end_protected
