XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���`�wD��X�F4
頟�Z��ؒ�U����s7���Ԕ�w����R����b,�	o��u��j��49�6ʡK+V��u��:-�7�F�2 �I:-�ol�}C��D��x�H�*�;�kH�n�`g/tm9��3B$J 3�>M�����B��9��H;�z���re�ŗWaOV��R0P�����<$���`?(>��"�;X}#���g
b�/��RΑ�.�g���"�iCv8/4�݌j�/'��	�� ���C��x���P&�^�}��V�]����q/2��7��eq�\�/l��T,�sj�Hd�x��` w�
~ʴ�}�(���v,k��X����9E��\�`AoC��>�1��F�^�P�F��io��虲�2��P�|W��oڬ�֣��?!,����sٷO��T������3p�Y.�%8��Dp �_�ya�c�Q�O���A�W8/��R��8m:�I�A";w�9*�]��ZX@>����j[�51ao5@��RM�Yd��f �N_D�f���۰K�I�a�C��LYڔ�X>�L�D/S)	�\B�X�}^���CA9c��4]�>*mL��鬇��=�}�G�V�j�4��䷓ߌ�A� ��?���!4�_g�;F����)���\fq?k�b���A�� ٿ]��L3_��:�?��Ԣ�m�n�*�d�_�R�;�ޜ�'Q�y$TH�M��A��C�J�vF�)u������w-ޒWJn~�œⵡ�\���:�%����)F��M<�h�J{XlxVHYEB     400     1d0��Z�d�1��,������$?ٳ����B���)��׭��~x�1Ƅx+���lf���Ȱ�����Mp0lA�gn���m ��~�$�~�^R1�>O��G��F~"P,+X�5w�W!��v�2����o�Ƃ�L�IV�G{���u��j>����y�&J1�X&g�'R<�����Ձ�$&�;Z�j��'v�/��=��`��+�~�{��	�r`�N7�@���(�������z�e�@5��Iv��S�1���yv���2��{�}��L}2U��l�p����l�ӱ��,tJJ��o���)FQl�'�R����/��lV���@� ��S�c�A[ʏn�$��«�b�v2H�k�p8������`]l[W�PT �����Y&�u
s`k�8�n����t[[^#>ʚ�K2�Ѵa�	�/Op�����$�	����A� ���g�)��Nc���u��}XlxVHYEB     400     130o461!�����#�.�r @V! �뎬-��	#�Qu�=�X<����)�}��{Z
��������0'��W�������b��P���IݶOu�V�Nn�����H'��W߲:4z�#[ѱdZ�h��x����Af�r�p@A�H>�^_u�y֣���&������f��	��ZaᦾC��,�U�ke4���ӱ��P����ٸ���YD�358����i�Y�A�!ѹ��{p�����:�̰7��`���rh�XNok@��1F����ĺ���O5ch/Ε"��7���XlxVHYEB     121      90NxY��cө��[!�\e�1(��en�a�� ��e�"�n����$:.��kM:�s���w�ܬW#
�Ρ9:�;{�.�����s�����a6s`�}41��=��S�d�~zu:[��j�Kh�}P����_d��g��\�.�iwlJy