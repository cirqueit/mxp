`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17984)
`protect data_block
Gyo7ENYd7g3jzbmS/9GN2iv27yLEZZGy8ELxstRZnkT5t1cHh7k1yb0OQiQoXqK/7A4kfIAIA9SX
3aYOxUthSHah8N0hHLKJniOjei8sO0TWTyE1GqhBBsAGaihmp+x59yVj4vDcKNtt3ZamBF9ii1UT
j6QH0xx8wTwR058JmOCUsCSwqsUS81YzgrtwfAYOsUmgChr3oroXJ48ADo9TMMW9dyRhzjosMjlD
lQpv8CE/79GlVSAAiFPPL6DhYclZ6jOsQ4Ujjdl+veExQ6kkEjq0GAQeWnETsHiklhnaxNMteDT+
PIYbTeLVfjK395mlZ1BLuNRNyWE3HDXIpduiY2QnnRs6+Xzu0gZQV3RMi9+47p7cZ3YCGNh/DTFW
Oq8x6lXDSSVIh4VizuClBesqh/duAQJ1UufdxcvoklyshRqCSZcfC/ADJPTIw0OdaVPVcxxjKjXf
wwiSsTwnUrbOs+9Bw5PWLgyOmCISpiJPfames/ZD1+oPt6NglKD1/smJKX3Z95/KggYOEZAe+4Qx
lxgi0riMR46WJP3WreJ5bDGlamP33t4zu9sesTHlp/cGeDoCPOv4ONejcnP1Z56MmB/nCzyqqGMb
ha0NeI+ZrTJVciBUSRqHNfA6Q2l3+cF6ms00EfzTrBGkecyKj2ULHqmcSkmuoTgU26OEXndi2PG+
062b6b8KF/2o7VVPFsMFfJvHnTORzABRGcs9GDnSzXiRx6jwSE5h1ya/7vtWzr3Zfw94aKUC1auh
enp5ETDILnidF7xH1+/ZUt7uQTjNI4ik4yH5Sv/ZUEB3XRFDUz56321KYwCRVqmtcl+R+RXr5Sbj
ITNLZWlk/1oMRhV2iicYM4VfRKeYGCLUlcxs0uCtcX8lFKZApZ6fPVgIu/V2oku54q6PT/KetZ36
HdkdHu5jOkDube4kQxVxEByqy3ZmCXLchkZynpi1HQfkwzIUJmP2rh3D1mlr2rc2LqSEQ/HOKxka
sJeZLcuiSqNG/d2pbCDceYZl7gfhO8Ny9Na72jmIrWuQdpUDEt4N9OL2Ay4p+uAANW4qO2CJbNyM
szdMG0y59TBoqLWGlrIZoO2DJyOiAgCaByxRw4FbLi3tJeF9pCP0fmoGscKGBu7e7wzadmHHGAGd
lEX5YqBtd+dXxM2UmJnBiwqi7hUl2sVaWeuI8RIbSQ822Jk8izIUMFUvtLF1mVTrlZEJfasyz5h4
w9I4TPcBZU+TabjmnAmjdjMY2qjcIK7hx6Zva85YDl48LAGTUqTSn4GFk5/ce4HDCKk2y29IaL4e
1UdMG+sTPF03G1Wx8It5zKKDJ5dZEXBVmntFqdEyS5KDPcKM6hLICG1hauYjaEsYlMPpf6Q2b43C
ag6OrhDhkR4NrL7w6e2HNM0vCXnxGDUhP6qENZS5TlN8faa5/L8b+RitqnFiRjV4u+LjBR9KZKR2
YXJtVoXbOKS5Xamj3Xjd72wXTKvQRUOuJ26uIGLirgGIZQRKvbOr/bu8kyRXPFOlS7cfjnF55fdP
8bVQrS9NGNb7QibRtxQLJP/bQWcrul7MAO8DoRsk9CoDbgWbVY2i0tb4CdG5p4eFQEKwfc7Tg+vd
UXL3L4ZHna6USWczM9kEzsNVVhJwuG7R/feWad11QaL85Og97xG9rrMXXh/NqnGYC+8q09R4n0yj
ov70HuBy87rLoIsCPvGgiA1aQad1zecfP7eId+LDz8VijBbVuDwmqW6WbSsPDqiVfSPYezDljDvt
IHaj8LhlQ37GzOLQIhdYeaIhRA9y0GGpzUjvbdh/NaMVRCNXxfqdjXq4NFQByxucWbDPEiYZD9Q4
xQxhPOp/5mOJ+Nr+3zZDwBfHjDZei/j6toD4O94KA6Kn/esCkEFAzHH0DygPXeTOjZD6A0YmuTrU
9Jr/RR2gvz4kma5nt0i+ilinm/TbukqvEU+kWMEnVx826kk7DSWsseNmE24Eys4FfkCSv0RKDcbC
nY3hXkg/UI+U+GNkhq0dbKQYvQZgQrFtffj2HvEeqtsVZiDg00CaEtyOJBSI+RDPlO77X48cNtjT
Wq2rrZHEk8NMTQW6I+ROpY3Xy6FV3asUMHjvA+cjpx40N4CoucPDvsCowFjL3h9oKeb1AVQEOnZz
rxOcOlZ5cCako97J1ijNx1anXePQ3+YNcOQJtGQAqfR9Nd7/JwolZO1jsRBa9MpUNc48Rrx2pSe1
qtyPKN6mYOBRi8LP3uQM3CiYt3flLSjrifY7zzHhBNOv6ch8v2KUjhSBY396vPr0Yg8JkhI3n1V5
yT1EnbJsCPbNKGwQX2k6kQA9O8jj8loOnEnzY1YzMF2pcg3i5D/IQb66eCvk7D/1XXFjfBnQsdep
VDaAnt41x2jUePlUbLMPxFIDdqMabe8livLd5Rb/tLLqyawmorljikPBrcgRxbtsJGmeAjDV+Br+
G0B7P3yFC6keydwvdbvompAg2bdSQJVH2uTV+WvtJhyNjwnwjNpS8v5MPkLbqF9nljRSlwjgk2GC
FySlzdzxPO8jtnSlMPQoDKaMu/rApMQkt7V5bS1Mcfor7HBdZAQdHvokEscnhH0O+mvOo4IEH0LH
oJv4TC16QWvE2yrUaH7Bz2dkzX0A0aNehKBkkU86U5YiS82Ez3TJjifndPaT03cijFTdtNPhBqdO
TiOfY1Ni+L/GWIMvy4dtgwNQa6f1QCGXhlmAvsrhezfifdz4+tZHcd5/4aCP279zMHQ0581tQ860
MBi5JEp/Fce9/t3I0YoiIF86w9Yf3c/D9vKjjczrkm5Stidtl1yxH5fTiiKksMlu6ZA2at4JWjcQ
coT3B8HOKezgRw5TzU7BwYaQX5YXcP4ThvTUx0GEsU+xDOrtQfp1apmbsiECCl9xXFy+d40xGTXc
A4wzPE5gqKtYEvP8xYaQSu8IJ+aHFB8Uq9J0gwOHsvFQ/c15R8HmjS9fm+DuQK6oZ4gag3sM+H39
iW4xNoFYh1qqLDImO5St3YEBvYWwPpuOwJybBN873D3YB4MCVS7pJkyT3kU+GSQBaRaAmZc1IQOs
pyeGSGtKm5QfGuPjX6u1OZCrNy8rQoJF8LubUV5KgCa3/pEbrMtSJnC+zDSyh6Jyvz/Yh81/BxfZ
9bR566MjKxf+2acZOjrUCZyCDl1L20r6vlSiGP12fZaw3wLza/KfvzqUEQJF+N5KvY8fiO6k5UXB
aRvQmvLDDmRbb+MhRWd1O6lrZdmdG4AnNRNibYkwH+hvU21uYtdhkLs7RaYKGjZsMjX+qVqaLO8/
6MGj9qmnv/CcE2f8MbH5Oq8G7Kgl8uoslqR+SLn+dRCPiOKp9o02VvEFtYiPG/L+OQa5oqF265pm
R1tJt3EBGdaNnGQ7HaiSPwrHZY1MC4tGeyJrKibp7piVSzIc9izSrw9rMFB4Y8+mwxDjvvAVR9M2
YFEUm2NlwMNvMQjUFSYKjZOieXQPjKM+nedeXiGx5xrSd4PU/phLKvBnvQ/t6xzJ/MvXrBfL7bha
nCNFBsFKxDlldGtpzQAUaPG+OWxQifEZLdw8/9jrtWHcBqjx7E/F/ADNa+EA3vrRcNsfhGVSvcoP
9/Sf9dOw0Kd2igkm+7DZd+lJIupaBrxwtJPcaC3f44jSmshkkzY46nalCBbPdxnA8QxgVzo9Sb4A
ekA0v/T5svkZEgvyWXIa/yKJrR0G9y9lx6zkOvMUQ2ZHfH0jz/jV3hkaFKxig5XWCeJGz6by/IF2
LCW6Gr/kzQsAvBxCbOwHXVGOcqFXEm4GZhOI8dlQKr6aiQ4WOlpBVHWds4LXFgyIXUh5O7RDBOrr
3kZI8Ik9NplyiZNEY3midoabj2grxQYavk3c5wqIwziej+gj6YqASK+e41zxfwWxm1lI455A8vrz
pt50P79xNvJWrLMWDuhW1RqbytFPi2103KJqMf0iNkchl4lcKCiclDG5LVKwNzxBs0I1TcxyVH0v
IJHq3USjjO+lThUOeeDhwJqEt3qHkm++2+oftR3HC3jGajcYXYqEF02jzFsc3HhQWuc3IpNH0l/I
6qNyfcnh627lajgqS630KVkFdvcpc7LFN0Gz1v+4RzOi6j5aJB8uPzNLCjjHjE/6zsRjbS/yBFtL
OBoHQ6eMzTsGuEQ9+hLCdFiRsFivyk737uOl1+0m6tSpCVbjUnGykqiSX97CI7x4O/w3gPO/3I5x
PNvIYge9wF81r7OySaIr9N3KnW0+VZardrFYDi97KdL1Y5ZRq2s/iiOhGmDIVQERCWLZJsaFokr9
phhLfg2wH4zzcDATN+1hTV19WyFOknUrv5Fxc+NSJYna2QjunFlpqZCrlPU/n47xyNm4w97yBQB4
fkqFJ+aDfNM6BWlnSH8YVFEsxaR00NPn8K91q9CtSvQiQzEKPj//9WdPoLy17NMJEHwsbylTquHT
7EwszrY8eDkgr7oOawp6p3TeTFMlyrDwakOStHNSxOnDFnQqkLyqhIaGGYoLGwAVYiSSVWcLi1iH
aKNHsnfQjvXIE5MOM1cV6m+LihZoaQ1KgxvXIlLB71L1i1vKKuH3ppuY9kF4TJWJG2QnvyiVtahz
gjHbvGS7Vb5+scDMlqEaGn4KDrd6rkzgGwlOzpVrsmLsfM9+EIbgwzkYA07a3RRHAsZo6GHGSPoJ
3+6uTyOEI1+7tZxiHsBgNuXr2l8tQ9M8Sp94TmN75B4CfertwrvbkZ0HIJ9ELbkJU063HVfyN3SM
tHPEaZwRhRgq2NcfGy85Pr7ce10sZmkLh92wUdaz4hvJm+ZoYdrqnBYn49PyPURGWOd6J71vfib6
1p7tDCyt7uuxhOiW65HkoEIKAyGDv5TksquuownMBa9zuWs0R7E1oiEwueLLLTca7yjSy+ey2elX
vzsB2vrhQEgQQk7HgttXHwwUI4dgX2kNe4ba2KqAkg3cF8dvyjB7goHb0mFvJ0GQxfg17qJlzmiF
j34EmOnrZb9O7lRZ7YR8F2v791K/wDpcSz35NsZlK/knfwjKkwYoYQ+Hkvj9xAopRrRSCl+g3q1A
hiIl0Q64PoikA94LSiccNUADkXmGx2B0HrmAQ2XVm1YssLdPsbX1z2yqQRMmRH7HZf3WcEyUzSqa
bgVB0alX7tzQpaYvdgWBJKQuniX96zcIukxhd3rBK9tF7MJjHdKaUidMicqiiqW+sPjZ66e17qUm
iSmD9OZRJpJBaJCFH+j3l1sdCH8dJL7VoL7DHrTBiTNKWZR3dcC9cahZAs76kqYeFtUIemeisV0M
vfoDrnfJRRLwtubSZ848evYnVjf4ohSvJedxpi8203yWnLNvkr0gWE1iT+BMwrhkYRC2xnaQp+E8
ELdYwMEQLTYIAebDygbkwa80khOFN5qYRFuV+zJBn7VIhKGCzYnuvDsD91j08b4qOAd7NTzf86eT
CESpaHPBaDLxC7twle+rZq58ZwzW25kHitqb6VRuPZTnRgk7kHez6/BmoojXJQODgRvFzvuvEIq5
J7NvCYz2oJD3QujSIOTfWadP33UGZGzhjL1Nf4RxUfS8XMbtXcISHOsNDJBESUZ0ByFdNKGgGBAp
zidxgoIHflZXGPGffr73+l6MkLcvZ3+o2QfQ+/cVjBer3drS+oVMDp5rK1PJbL4AlfwyvodJutzw
YaxeilhdW/kSTSlObVNR0NkqDg4L+t4p58dbyJY4ko6ruyVjGbLNbMWbAvcuVd62JmyFXL/i+p14
7RgOYKlF88BHRE3SkLbK9/poFDLgw2XDEosQ3ok1a4m/xpr6m0BZyV2Pn0OmzuGOq/Iuu1Zzc957
jAzrdij48rnyO58dw9Y7+DgJxh784k8C36ZJByzSXvuC2a13ixSYi82V70yQg0tWEI/NCzlQuE8U
xT+Kf2AN2liah5QG2EpLxMcAhfNd29BSUCvgRsnaNd0WMgLu9Uyfbsa0Rh3idQl83dRdQPOM+40U
8SpVuEoBVb0edaKEdIHBUfhcvub0P10S2LcFj3BKZbAGFLwLZYBiu09nvc/Wi7utFcgfWiDC5n32
zjAgj9RJYHr8SiKxUMjDD3m+zuHr536JwWc7gTrfAJT9p+4/olzQ3NjXAlB9iikTCst64zlryBzm
3vT3v10KyRuLoIDfspMHAabO2q2gJa6LtVNpg8Tr4nGmagyPWvPJrPhQo0IW3xhRIEB87gYIOYfY
xwOZ1We9O+Hzk+fmOq+smzLIsDsslGeCdpiiOUgJX47WeeAEWv45LQdLAOMre/6TO8ArDf2unvDp
6JGqDy/zYBcORhydktismZUTDg3MoVLGO2SQY1LTPZ9MjaR2H01Sx6G+caQQHY3LCSBhIOidyb/t
a3GKjzNSZGDEhaoldBv60YGmI4NujboiWYi9ehBqG16jjhoK+MaB+Zvl5wNyXdyNX1DnHqISG2ET
s0A254MLu3l7L1Ck4qMjpID80gJYMrCb5CJe1h5dTbW5IxRx37xuY6pSQbSTY/+ewmsT9f/c6of8
D552Z7zbIfCtwGqODtPHyabWQvmpqaoIkk/ouMTBA5ALquek2eWWEj8A4BUmeSmbIEMD5dfCMwtk
pfE8p9XK9W1J/ke72qhNb4xFBGsKOQX8+wXYmpK/KoPmPrFYIKKjsUnl/xSnjgQqyFMk9oyEWGM7
NMVoCX900n5Smj768XvJtmEXWMXz4KIjTlZvMpcUPVGQemHr7OgnAhKZOGfXsKPJwn+4MaMylOxA
uXJJG2GJTkVVfUfgFhGFWhHuYUFntIQow1TmBXLY7Hi5r3gnZKpbjTkCvcs7lBCgIxE9D33tdHRs
gMNwAl9lPTLlPDcl1jeBAI88ZzRAD8Cm+ntf9PwCOHYr0bl5cMKU3JuPfbubp4YpkPnpnRiGHkWK
y9Cc+1iEOrC7Lr5i/rwJ23C2D/xebvVVNmazz7DziZM848yRM0qr6EtPpipE8NmE0ShjDcT/2+dE
JjwDAEJr51Tdq+OQF6jp7ZVg6TOxR3787V0HaZvW7g9EaSLeu4lraSyB33OTQi/Uxz9n40COrzny
qQilLRlwFYyptxQEApeCwf+3EEiotKjIQYLOlZSpNDAuxvKur5P2PiErS5ZwdoGH62DKus9xOndn
MR85ol8Q461OtrbHo/zJHje4wavuzGRfOCRIRLfsGGjkk9Esq+6vHLCBcPtGEdV0I3eHyHdryfYd
50+VB5L0jkIizPT2ftLLBRgw01FBl5nGMD6HHtEy13xD1OcNtrNhxTS1+BKPjU/RNCFOd+9Cs1Mi
XUMTq4XuIRyLU6+IeltTjMf6U435D7cZi6NfUTS+IpfATqs510RN/VqsXl4LhSsLmMk49xnO8h1Y
xoZyIuukDSrdRDaWAcnXnR7JHfrVrlrwAULdqqwWy2/mTKqnuKhqH8719Loyqb/znbT9SgHKJqOM
Nn+wf0sJe677ulCt1xrujqkNXrPihIvM51HHl8M+/DG/VOv9vVGvRkO/EYxLurzTbzhi5o5J62fe
0fC6CsTE6a4yN3l74hvOonHJq1oaNU7zQE1M8ke6GT4MpRNTur32kiMsozm+F4TfnQxBE5xuGkzS
7NOE8YfA+whguC121XaDfdZzY4Mo/NipKq8WW8oWnedLhKfh2jhjX4YlZ6p4gsUcgC7ppARwFMbw
Dc/jhh/5uXXK6WyQuBpgynr8rb7lg1hsJMvboCTThJW1emX+RJbybzDxIvNbZhn2v59dgbrb+d3W
/UpajZTphAq8uR1XzgMVpXxcjk01pjnpZdUXHz+lQyRakp05lKsCedMQgaFnghJnQpO5g1FZs/Bw
0ZuLKGxJKMuKA2mDV031po0pUiPcc7hB3we4f+MQMQ5gH6DLPFu+wQWfz9p70cOwZeQhEqSed8D5
N11YWMovFuwMXNdq087ZjIBD9ov9M44hOmpDdr1C4te7Vc6+Ci5Xwg3MY0UJovign7nEYvtTAj/0
0zHsYcEekuArM91YWzOWOgxJTtKG0KgzUn0WznP3yInA4O0Rqy3lpb516e5OGif0C/bPFTaBCeQw
tgPboIlaY03FOXBBpYWNH/zAv7zn/ya/cjNUk2yOl9X+00EOfIqDE/RcPVW4OA8pAnRjZq+WOF/Q
oGbPXZbHVLkea8NU2JovswFcK2h/wzxZtwYva7zqlYi4eIwvUdunoyYEGf6E+FMsvE0ZvdKUrRiX
ZS4GokW3nTaLcIbPHuAf/0SLP8Wsmamg4kvPlHjwV7Ow5WFFcoZpEw2dM6gUPFn2Qg+t96pWsBYm
8DeT6mRPUN84zBAf92fLm5zYjj8pZV+zdf91S+j7Pu/SjQTxC+cgyGn35fBwW0QKlRwhlDKW3/WD
MgeW8jxeJ6CDTDWE5evulfcHUuEVOOYHhBBg0UQSR3tAhee2Z5ZaZX3WUi1S+fjkslGBWYxnbczR
2rwq6R3V9TIZsApXjOdTIsrF7y+ZIvaEBgIgY6Nz7JqYOgKNrtFNUDn/LQ3c+XR7PL9zxsKEMj3y
nVgViVkzR0Q8iAU6iHRUVfxcUwQhFG22YGccH2csxq+d+PqF2NhJfKAB1GLjxyqvL1KVpXvQZUSA
VHMgtI3Ha2KBDNKy6y0iQDzL+qAd52h9blnET8OOc661MbX/QWDnNXRH31zT9Rjw1L/Wze5/GxqF
NPrNksqdPgVECCE4Lbti5KhuJqtopN4NxhL3y8abz1XdLRfskl0G8Y/EOyhe4PkM68ppjNXyEJ7v
GZDBVghXe3QS/if+gSpgiY3bdssJZlTdWAkq4EAPCrnNPS4/DP1f4Fl9/3ufhixQpuu7yZ9zlSpS
c2xKbf/cuzmdRpRC6EqpKvLQB9PIJg0h9gRctw9fBBla76TgTymFLZDXXqgC1Qm+3AaMan2jXJa1
cd2TVqE7yQTnQyemyYDAAr1gGUxiApFuB92ovPTVcd+KQUAdozj9SdmrOdw5INfFsTSOZSGVx4HY
5RcDh3OUv6Ld0hbXzut4CZjOvY9rTtnNMGegR7Z7BuJtLA8Vn2rmRJsEukulgbrauzD77NlF6171
S11zrJkVNMnhSufcoWv2soBWoJzgT7IZdZzJEeE3pMEaIyltPnGY8rAcqnrLfguvKD2NKKqZwjxO
Wo3gLX3luCWcj9r9KOIPc3gyxMg9+6M8+gjTeWY2ltJ4kwu0cwCfb84LYTiVNFYvLDe3VrJ5kkwe
ykzTmzYqQiGBHBmJ2ozodV5xNPEyfGzF0/mHSYMfM/s5UfJ5lX5uHvl7klRWTqpfveAt3L6kLHaI
mHCsSOoYhaXS9sk7pM+zyZ9qfASVgXtOYaWMq2ORL/XlF5uCNU3CP7bS2EytxuKv0T7tuiaSK9Hc
CUKqIpIJ8eSEmSVDJ30xFYDDHy1IdhTjRZ/IVv+1w33w5TiwVjwE2erHUYY6g2kOROpwFZbWj6wD
ljzFZPSHvjScptOuQEHV7z3d6EjZaUw3DlZPDdWbkla/gK8NjlR04mGgrhTNqVb/EqGQAe4sLky4
t1SoYfdZ3bMfRAE0IvSpsiEvSbsKZX+KsPxAxtgsIN6YY6FqPTYoRgfJ41NQ2/oRBp5x40hjNNMs
7lxjdcC0krtQzGJrt1dx+YRLFO/WvVVzldXc6hJmZEZRbqO7cdOH1gB+KtEx2nglYANOCxVDWGDk
kECl7rxRxEQqlCCA5+Kb0kwaQiz2YLmdVmCSVuBCmOLw6rfE80SZY1N9Pqhrx6lLke0tIeeuEyGS
CPJ9b7Ck+ahPnY5/X9JLDCs5J29aByncrFDi31Hl9EEE5ztXkMGJo+2+ba/c3/YJ+XPtNaENpz2b
dXs7sQJy9Oy2z2CnlSjcXeyT8Z3suxYNRuEvZKwKU9X8h2oAcoNBGUi+qNlpDmzs3gNGA693I637
ASuBrgEjaRbJfBRgznFWa8g0wC/Oo86/W/1LVjdrGRwlT++TbzqV34dG/Vo/kEfPXDTRwNd1FcTb
Mj6Llx8cR3I5nkWuiQyv0assd//r+uZmla6N6ZNJ0IAILIvRKdA8nFw/DzxoftbB48Hlpwp/RU03
451YgVjg741m6AzOV0W02nrznPihrxc6uGTGzXvJv0znjeUFfARmiv6ZV9nkLTAHKswxv+MW5Jnz
GeR0eKnD0QE6RBISyvHkzjCT/u+pkURw4BPp74cKT8F1tXf7a2wdgQ7D70JpXkb6770hbmAvGF4R
nN/EU0AfMV+yHWDg6NrT0YO3T6hgB0IRaidWVYfDfbZ/2Ri20hi3x7Lp5dXUgM+B3ryv30KZvqtx
uMsWue1dBN3QsMEMQLNq5R+mSr9KmUppg/l8bNeDZq2hgas7CvqqM207bh2o7mqjivWoy1UTZeTv
IhKz+tkR6xS9s34sS27pqARHXdnGwAUb2ZkBgrq8/XvSA6ntaI7fz2kVjDFORapfxxVhIfySKxba
BOIztpj4kHgaBucmpql0s076k+me5/qFeG+ehUknM6fAaZ3/590NWr0S+hX66Mqt8XwgHMBPcuyL
9DOO81KlI1e9Lxn4Ku2epcdJ8IwJuU5eOj6m+dyhRUfgfy9cPauj6hipDM2oXUKIFdZTyfIf/+Td
b0iWEpcImnxbxQy8eEfFgbH9GQcpxOIPPBCJA60Y55H3Ws71rgBQhUSsFJzJCGxg6iqm/qrC8B68
D6XpDOKigeMdKZ5rU25qhk4kX+klsYV+Ajb2B3zCtmMFq/8UIY3rhK+t+4EUbdFT9CCSLLexe4fs
7X5Ud8nX3Lvl+d3oBtXzGw1xDKDFG1h1rkNZAp0mlUsuLafsRlF0LfvqoNjY0LP6igJC05N5BfZg
N1PD6UzjZZdN2BFJWUVB9Ay6+k4KpEpNxw708Yep8dt0tr46qYgg02ULhw64rdjqQNc3Rhxiu/Sc
iDmeYHrkwk8z+reX4OhLOF1qlrpGjsMC5KeOR1BAQ7rwI7vMgEIsdY5rFOx6u2i0H4nljSMtZDuv
bY4/r1vBWBRDbE73HIaxqDwMbxftGPozlWhsS3UffL4EKCY6r5Hb+7ZrWZ+IuhyheHLhwitxMrt+
hFlzlBNHtgUJD8YLnyoCqQjt+CtSYrvao70EQ211ZK29Nitr8Z0Vi+45vnjxR6J/c/M4NNit3JbP
dg8SnGnROJF7URBo6fhHle22stq4dtwPtLjkl+yPgqkDJRBAHRg2+1scHcnmmZjhDRX47/HumxB9
D4Hnf1THn3F0AcOYpazp+/5OS5BLxY0Hdz8JkzCiItVyagEaBNj4t6zBBt85t9Ys9KA8FgZIt+T3
28d4utpqNiTGsdMO7MM56fvXmsnCSofrM/zHG3rVMybxKRD4ktzeO5CfUuoV/tFT151TtOgCoWGu
RjhQV4oA1tWJNSd/GlIYmR0Nf4XIuzY96OFvh7wu/QP8UDFsg1d4V3IzE8zBewa3ucNAhUmjp4W9
Mz9MIGL4Vv2AyZfqignRbdYnoaTuj9VJR2w3khKqPbW4ifkC5ODCBsbPLe1woclqvg/qz8hL8oHU
okZhdtlAldG0KJ0VGE/b6MklgUVtivR2bl8+zmkQ2fTFQhmd1ctjEY0zohEpe0PwLkZa9iM5x8l7
qY/SyYugo+9c41zUnMMR9YDHPwTg38KFtlthDiK19oXC3CcQnhw/yP1hRNR8nCt1VjNGpW5u9hd/
CJ6J8JNNPcwrOo/cvk+zShzp8Edp3+yLGgPyx8vQRAee4CAlg/JbthUhYSujqQtDOg1fn2S7FQey
Lt43WkGOtcG0jENm+kJmROSnrskG3AfnPFeX8AGMCTcN8ip5h9e/0jN0SNWrNTr4+x7QQGqCIEn0
iVunzsnO2HRBw7PS/ERY4A7JgVVPIXU9MMlKelVrU5XGPCvgG2buMl0ZgMR23sJqG6qlKL93twEb
2u4gzlykNP2/XJy5JShXGRuBNHoiCVAjCDRXcdAXWADCXepQxuoAb3sx8FFKzr0A5jyxqLCCTF29
kEsyI7715XwZBi0Q9gl9n9HCyuRRo4tmF2FJSQzwS5PNlt5vcpOGRTuWkzjb7vlTr0dnW7t77InS
qOcftki/TU8RVcFpUis2pctGDN3l8bg9XXBywERGfIQkghgRdCCwQcziM5HOEumtevGvumeBepxE
SXvIoSA3s6QSFI80slXJkuKzVuizOJYWYmJwiHz+d8S7w2gv5JtSwRjaItbVE4jumRiLRn97HVBK
gJomoLOS0lDRMtHhmJfdj6f5T0Vwx2K1ybYUS0s81Zh8gRPQvo5vGU0nAu+4nSxrPcUvBV7AmK78
EOGbYP0V+3JwJo9jeTLlBm//+J9XmpjupYAwkB/xwnvPr7wn800PER0NA5zqyRWU6hPPA7zQEa1F
zyCo/le0aS4YLtCqcONL5sjBqvs0YSSeec3P55KBO2EKdwPIWNoU7OWdEE+uJSgpwtr8PWyJe3tS
jb2eiNfTdTWRCoi8A9yxn5OI+W7KIET8HvzASiY6/vmoSczsei+IcAgtqLW4mRmodd78omV3YK3p
U/NuUxJlhEafKfH2w2GKKVSx3/fAMVZuhkkd12DpDIQFGt0mrEmBzeHx6uFenLLk6+H1164TmH8c
9zsVLpHA/rTUYaJ3FOreFtLNy9XdkgGvAPLLC+SLu/2a8Cha5D37aBcy8OnypCQwEX/VsEtgVO6z
IgU2Gf6nLvJiZYw69x7I9Tgk8z/wc0Pyo6MLBe8J5Nzc5HF83m1xtrki3f6DD9t59a+jaCGXzP/g
8XOm2xa2JSLC/3Q5fUFdonJaVNhjUdt84MyJVBZreVjItqkqu2S+/8zqN1KbmBOqhhL4C/lPDurb
ZvKdGMMLCvZqDx+d2EALY9Xqs8+4M1SSCmka5vQqyGWWWSf5L9JVhlzIUtnjczv7nXPwsr8M1H5P
gS8xBQi34ig9ZBoR7ZGnHTLuEkwoDbBh0TuLyeFm46Y6GR3XtbgEUM5GunpkamhX4Jv+L3Lfkbjf
CPIbIhx5xxjRU/pxSDZqBdV8WMFKcgZ845iDPtS1TTI4fcuBNDfMySny3NUbwX5Ke6fF8wq9DcgZ
98qJruuiLdfBSPGPWrlWUP0lUhGuK1F/XdUOBHwIqeD82ueeNTAvkyBn/eUk7wuI/L6U9mFBz6S3
Y2Ghz3U04NAMgDoCE3VuMYleWb/O/fCJs+rAZ71bRzPA1Bf7/Mwjj8OvoMxwsDKXH5mdfhuWGMRA
BusY2yqLmBq0RrtqQ5J2TaynJZ4tnbKwXMR+XDPLGXnnl5Y+6uHcjCCNCU/n2GOIL5qCAvbVsOuj
1589cvJ7kvBXSNM3K3YQU3ayL4CbuM8bN19c6b8HDVLozkDd55hDhtqOo0al8+v41BMZlBdtRFXD
m4Hdjlk4D+mX67mvw9JnkndAmX+NYSHl/SAziIZ6O6/QFrtS/+/46H4NWL73TOmEBeyltra1pKN2
eghtHIDY6ck3E9WhYps1/68ciYXhUvfJxTKKBNMlK2c/oP/RaRuE4Xhy1yjquccbn98X0mvz0kCc
RjrCmyn7W14RFsiQSDbbnljguFYggKtCjgckUgd+DOBoz2kJvBJPsKrT0Q7Q72FSedkf3+sEHhMP
alDaaqsrGvHO1RoxIzeUKqUoo5vWwdGbo8RwsiaIdHV0/Oz5gsaRBwbn5g5BHmTu78nikdTEUIxM
gT78a2vfbXE4Zm19pxpJlxvPBZQ8WJN0tViHp12SedG6KfqgKqVY+WoX9FjCzGbCAfE5nD50WjIk
jbSKfFFNIbBE5+6Dti+tkqA7ARa3Tu571G2AOUOJMGSpOPw+vucorkfUTc0NMJWqjSxz4MGANh3Y
brdEwD29JTKaNhoZDr0UEFdbHT59q8azRU3MIlI5gnHJ/HsHQg90Zt9LV0owy5sGs3DChVEzvUGZ
jX2Z7TMsnqoLrtmAOOt/q7fqvb9bOjCwn0uSkNC5N1NAIpY3Yu5KQ4LztB/tOFaE2J32PFhprd55
TebY9uIbllsIQEbGNTiRDh0nprmKWeyXBk+FTW9Qi5vwa9m5txwSYbyL/Tb7UOWGos1jtjHCoRPW
8v4pmpA3p+rJxqGskgno+PeKXJI2qfPSO4BcFCGmpRlfdQ5uObL7R2ZRmJgiKKjYmtY3aJrt55Ux
te95NyHyHiQUQv04259FkySa+6c2zuPYWhKbkBX+IuspZK8ja03GY6qK3nLfunejnfYY4tkqrFQE
TYzuljVnchRAVwc+PibwJa2G1jcvXe9oyf3p97IZ71QsbZ9gYlFb315TOdD70zQ6FIPqrv2JSK/4
xTz42x2LB6I4KkYkc/KW07eOOYtXQ+bf/PLa6VhZ2ILuNK3e1l4wrjrw3sNruQi/4oorp1Sr408c
GtGrV5hMns8hNzzrO4lthFkkvraLO9MkegAVR7TRWVlyAx/j8fyLd1uLwwlJOaIjeTL3hYv62E7a
9m4KL1nQeqk0r2qHlH25JUJiVpj50POqSXi1yo/hSmh37s4W1dLURiTyxi6+sWnONEPP3/ScRego
aQaTwiBpG9ebP/3k0GUWVSwcBO/oKbzBOv9na6yZ0veR2VTJx88I9NfuHyuNxTM+eOLkulHZIcTw
cTcIfFOmUf/jr89MltPvauhC2gsnYJFSPgUttng5z40ZbDUnuwkQXK7+NLRxsVmWjFlTsUNV6PQH
0G4y8AwTdH6Aiznrv7gH/IbLtLUdqNH2rqxklO456Z8+9z7vnag86GOr0EeUXiUXPup9anWkdQA0
vR717dMvd5gEuB+Q5bBKDR5xbq0GU1lqUtv57WmHxv6Tj1jjZ0tRSoUoQoZy9V/eINZQUTlDgnfp
qoc6Ym/brcPXH38/bJhdrPOIB1g+fpwJE6IDk9jHgsdV8FvQ0Ye2JDAwKKQVnlkjeD8LxRdccgAD
C1jw+z1wf4459hdJiBKK8id7aubqgmdBRqijf7whZ/GdWjlJAZrB032KPJOlCqskAtw4BFdDQUBi
IvWbMkK/BoFyE09wHn5L+lNu9EGssCGC662RwezhAhXLhy3IWC04e0s4zLE0amDorDp3NtxIT+Uy
M7B/m6p4mh0wgU0pNecxei+3qRParJYBeM5B0OWi6mPu+LhUNU6bbngtM005f09+Tk9kMnGyRsMY
eV6AnCMI0m7AEUwXKVNL6t1wzJeOf/k9iNQPacimFURWEI0wben5wGG1S2N4PYCNPzpBDjynVdCv
MYh7kyqQqsA9qIkq7KPVtksz1xSer1Xp3AlAzbxNgg3gdU5A+ZygH5F/RV3YDGJcrLOF+PRZmfGl
028osYV004eUr4z4cw4GOkdjRb++EfcE0mK9p7w4d1SOv4AkpMcWkNjieO1zbxHc08DgAPvxz+y7
g3v49/l8sEJ+Wq99rNaozYbjJ8XdPzFvS2OOyLyz+/IRy/X+xWo38zEM7Exy3ak61BI0PvZnlL4y
EfsRWUQzWYnlJLzytcjO12s40dDTMR141JnEfVXczwcg57YJ10lOkD/s/9PL8v0IEBCDuQhbZGBG
zpB0A7FARrANM9v/HZYOXX8YxGGT8ltENbxWP/PnGT+7vmZ3caxzkm3Yh6Luu4IDI2VLz+bV3N9M
qIZc6yzGY1yJNPDssijZc3gtpW7itcYEJrT78eS4jLUnAa8hxQxJU2wpxT/Ehp9WogEafKRkphO1
Mpp3PCv5J0xBmX4o4Kz+50Yj0qVkRRKEIkwoin3MO1fessoyQSqCGLhxD34Q5X6WO2HfBFGu3Fqy
5g5voKspBnUKh3dKPUyzrU4cv7KIsq7pZ89QONucgHTa0TjsXkKmove7nQYij+aUf5jxOpJ77CQR
HaSVTdb4v4D48wmKGwCENAI/nKf+uCjq0ImVVkP624FtUN9kRi8hjawUvvW1n6d7QAHGsEwMEEpW
o5z6gQhx2gRr4Hyg8M+f4GsE3TU+oFFH8yGJ7RZ/j6UpC4jQpe5MrVMl804ucoXB4A9wCIus8ZzA
kblQ8k9308jS7R71C6Z9e4Tiyc1Z+dQ0rq8mzpE4XJGUbohS4BPP8klBVIA6zEtrSS1jPesfmpJL
ZhB/hBP2qLnk9UlATIPgATrP8/kuQM+y6jI7bHIIZ39VRJRgY4zj1yhUHsVh+hsEpqT+q8Tz+cAl
6zsZQbxJEOb2x/evma1EFNtFLrXgtu0og8RhwZG17eUkZZGuo95GM4T8vxIlLCyFHrDEIM9ASHlo
tXFD+hJf/BD7zgjrsYh50HoKx1jljhv2pO97RpahurOoHzgQ2q9BZEatqUSqXtad/zwx6rZ9ti0O
onN1dDMcNK4J05MPXuBrUk4CqWLwBl1rIMxvi6wPb697rtrUW3R/UdEbbDf3oSEJ/DP0/j06D4Os
/M3mOsXpZnVtcMGye8/7kH8h2rdnyD6AyhBaM3P4YVw5lsQ8AOEYazGUXZESbok+YvY1UbAudZOQ
QY7Flu89l1msdlil5yV4gPeWcop8orNTDMLKcRrh+ytmA8c1hMFEN1oB75h4uPE1dSOGV7qalnqt
xyOH57pZwkhRu/mO0IL4F1FLP1ixAyLuy0MXvervK4bWh1VlVvOaVZIhqvk05BrY0oYXXVnbJlCJ
QmZJnkhrmVC/7sAOCKh8VDyoE89L27kFEQCPUS28wjGsHQnvNXT+tN5wn7biK/qGprWQE/118i9R
UmN59isnGsmCdZSiOtGFKbxFjKK4dMV0js20/yomMalsqYRSKmrvjm0OU2i1sNjqddMkFdb6TBMe
POycLew/dqMEk0zFZr5yvGTUMQ4uhri2lWwO5gidFJVPrbbGrau65tK5tHklpHnxlR+8fJDS+wa6
TUCFc/Fx21QRZmQO1ZrSikjeXAHq6g84H0Ar8ExVq4Bfd5dOHqF6ul8q9OpN0h+Y8avornUbzleo
cexRa9DZ8TkLsRqTV2Hk/rdZbQBB+wcpmhDZ8ycLFcWxdOiFklC0X9/j4i+p9TUJEeZUEtAEw0lZ
7eFSn1r6O2mcPWHaWSzJM6huOZbqj2N+thk5ggiyLsPVf/KS9nIjfyhAXJGWVDyHs2YsC23pJd6T
3BWnZW5D3CBjDIiwNsyXTp6HdYcHDP+xAbGNqhrxgBe2EUlufOeCMtn4hUOSzum6BQPE9SdmNRJz
IJKFCammSnFPqSdbMjP5loXi+J0QAXOsni4zdRrkSp/atFafWE9TuPvA4Qs7WMfcFdWAp8zHqOj6
if8s9vG77paa25OtuDPFeHB9o1F6W7AP187rgxcoPQRlqVjQOUYYiy42fDAFk7/hwlm7AnU0k6lf
6mcGTZLgUcUadMTauW+Jv7tl5z/ormAw/ggHrKgZWsCOzjmD0Su6ndFL9Jh6YQWy/miaPtMYqbzm
aAnd+/se9EF7wKfU66s6+EDvd+RlTttQ/YG87q7VKiCsppppqCS0/hwDwu5buOcyhvahFRG4+RS1
lH5bwgUYFsRpQweG+kwkkhBTo4KWs5QRlU+5mIbRGCB7k+mBlhfN0C8tObCxbXXz5ahHp/QLIFZr
+EOCtJReYfqi25O1udsbS4Ml5ZqqvcR1BCLcpfIHTNGCbn2ecV7kEDhkxp8Jl5Hfg+blqf4UdhIP
JX121j3NnC5f/+znmd3HguaqLWexVQv26w3l9BxgS06f2jp2MajvDEcGBTUNFY0FQTiWDD7fREN3
mMoPOcGmFqMYz5dk+1OjQCeGi1E8areFeoZyQR01zdXJB66tAgGmJdGoloUGHrJdifZ3lT3izWew
ZyT+HqLhBKDjJXsR6pzNjkO/jypDwcfgTzOy/tOvPSjG4GpUTJi9nDhe6vwyoP0JK3XyfhVHLxy/
B4nOwD7C5AccNVL4RvOxzic55+VBdfYxbSkIxgghSs4dMET5w7dfm2L1WKR5RO1DleJtv0ms176G
f9ayxR9lrLJH9JJVAN8fZRj1l9Iz6CoxujzBidehN+EYfpZvEVuuQpqp4vNfItfiCSYlt6ZfuhC3
F/FrYisZQjSu92hOwp0UlJdHNDfI4OPTzNXOBjMeRUaPH0sRLtFlGcxU2dPVxL1o7wXxoUSvIZMA
f3W63THJrJSlbSJoBO7rxhYJJ3BlT/0YWGae5M6WzxrjGOSanR1ZBfn+zzGg5RwLQbJSpSexjd5/
1AD9B6kZlG4cuOvpBalJAaZ3FXGmR/xQjL6BxhOOqzLp3pGJifbYP6dRE2Y6fsd/IFmnO4AAgtlb
I+Li/Dmea/xTkV+qZ+4514HRdvnq/wLWntStaWGp0e3c6d6mAUqoemdRvkzju+ufsYkBW4KYpLVG
wI+W/FgkXg8n2QoPjP9vFWu0C0VwQeOQpECBkZcL45tSJxQBmio5VIzO64Sr6OSIpicVzXSVwrlW
M75xTqw3SJ+uWE96Bv3FULvlVe6W9RGNW5qBnnJRAAxsd5XBAsAarxwFRe+x9cJkQ2coiiiJwPOO
I7KuVzqcNqq2VtF6NDhJ3BvS60bqe5bA3VIz/eLCgPq2xTyC3bCy2xKqBd8Pm6TudaWAzYLYt6q5
GrBvmhztx+0NmFlSTzpgiZw38OwLyliFIZCXtrMATywhI5Fu/ZO7rZAvaBP3L1xQ3qociWPFxU6g
9+nD5fzUEfKNPzEd4RElkp4QcyejLrBEFtnIHI4KZCnCGdI5UiKdSAovND1B+Pdl1CJ0tcGnRyvP
lNWIKbWjFHY+IDK2jfueNjo4dDY95y47QLtBg0HeEvEdT7SBJ84YeGrjZHjecgEcaoeBqvWMoUTI
JsTwjGhqj1s8P4ZPOUvL5pVX9fZs5KXnjA5/CEXsRXFdFoSK16ZISEVcNLxKNmIhdL4J79It9AdU
ePbzh9DM3NyMfkZNzyV5h8XH7PfR8U2f6Pg/oHLqn2jvMmb5zDI11BXKcgd5CoYf68Bjb1Q8m8aP
PmeAQ80uyW2be4/rGura1S/NAdfzlrVk2advlLcieYq3v4KNrVA9R84LflDpszSQS2CYQUKXEFs6
uHmClO4N/NcwExYUdgxX9E3sVMxQBMx3ZqsrpVMgoEBMsXOu2tjyLpUGdTEuZ9/tl1PQ1RGJsxNj
iQcXZsbIVuy3MHl1V9SWau1OCu1Fdxv64Jn7gMQiqYNg9Rx+6FJmpvab3cPL5VO5/qHCZyNwaFHa
gHS9W82PLm6xqgmQ0l5lSQaLuAYwHCgz9eUOxDjlCi2CaZNiZ8Wp5Rct0CrDjPPM9F8ugDAVeZTR
QS6wwR/+tRBkq/z5gVJYH6s+nErcTzMWx8Y5rV+1CVRhEE0ae0oWK6RduZ4u6aVrxgO2JosHw03H
ayQ89IQBIfKbnXWjsb5rbKLvQeIe0GLNyyU84WeHOLwiZaLV7K5O3592qwJAivD2qvzzgdtrKI2A
rNhv9u8Q1C0oRUOMM8JPoUTJkdJL5JOLRrwJO+9ydHCIrCp1n+iEc/lQdA1u2jR2LcgAzPer3BoY
y2iGn1tymp4vwaAa6RFTNSMnZ0mT19EL6q/FXhxY++QzWgEMegHWgkcHyXCDRg/SKdfYrk1MhIwt
g8+pT1cVPIsPb9o5z/Fh7e6+42g+VP9fi+AYuQ0cbRQgXtTXCzK0OB34/Pb3duvLXNOrPDJA0nNG
EPbJfa5GAoBpqakRyzaMN1o3arJNOhQdNXizDKfqLCnHfkRbLXrTvuazBy1bH1fiqztwZUHFEMpl
To9SFYIluwd/AAP1pD9HRcMhyZIB1VCF1l/AnvmBU8zj3Jn/UboWf6seaeTUxNSqQwwb1G/JQapu
iI/VraOLeuWHBha8I+QPkpKsMm7ns4B7Kby1PUAR2HGz81coYOuStLp9YkIKF4SCKCODqJBfzS94
PCfQIV30A0tLCM4vOOIAsmoV+xg6vdC/BJmXSdl5Vq2kINN1FTpYvSCCdvVpqOzJwVIO2hwRgyRL
X8T98r+JdQCw9+Wx2OlbMHZds88xCwl+9VpiJAGATyPuTPfQWxP4rANSihklu6L6XffPDidAUBhP
6xIMWHW0lFZI3++y/6hsguxVwOHvc3rgW5JbsKYKBsFkUwbE12pgBPocC+5dBiGWvQ2AeQjWmVm3
cXU/UCNSf43uZ4/uNFjVL7Tsw8GlhCwYrZgZ5074gLgDoYvRF3i+d9h/rBV36cPL1SYH7W0PuKYS
yeufq1qHEK7FrHcEqihVfbadXuCSwbmrZcBH24kmamWW46PN8VmPXV/YMOpHlTbDBmwJ2sOQJgY1
wtVNsYsLLLpcBJH6tXLqCzqI0WUavUMZR8iYWlehqYTT+G2slaOsduH6AokU81nUakeiUJB7AcOG
S6qNnzD2qzE8nUg/O6Spw7YOp+fRPJwqmDxjlEDLVNC2Q5RQn++TtJBJIdXrWn7istQFAj///rgY
QSUB3PD9rVO00q/wkqQBx4v24zNuWWRaDYOY6jXFG8vYVAPulOs8h+is9rDbdpOc0byJKzkaeOlo
D+lCvlK73tduZC1PhK/nXTFd1ylwwWlZKCzORiey/NMkYItdYimy4hz2YKrzOnRs9U510twpbaYd
TNndsT+Hg79eJSXHm25pOiV+djNot6Ya1c5lgz6pdTCDYw+E3q18zSV5UjDHWxN9ypXMpu6sQ6Sp
y8IDg8qNxROgi8VdEYXodmo8U3VXW7cJTD3s9pVcTIG6GyV2d4msi6TYan1kotgda5ZfivziVUnk
Nn+pT7Hsoa9x4pGncRpLXMDbXnp7rpb+3cGIPjSHEEZZ7030FeueUIkV2xacCg6w1+ArLPCICwQ+
AoIyKuWLpD2LqT/OCfui00OBD9C4S5m5dcDcEsazODHchibfGHeiMbFdrCQ44elw1pbUViqAJEQM
DN/1dWkY++p9Rc6O4+ghJa6WfdnRkIljrAmX2XyPdy93MsiGDGcGvUW413ZebPbVm3XfYdtHzG/L
JTS8P2wsKQO5vrTsO9827+Wz88ehHPGUOx0ydjkfUeWU711GcmulYBI6an8M+e4WfSHb9iNUqnWj
c5puCdWKr60nxgk52ZoUm2AhM9N9DQxTrznv8X4aKPSrAuXyzxltIS1kW5p8p8ByeLqRERhqhGXd
60fl0qhqEBH5v984XWq5E8/BCnBCcoTK2wRS0+wR9WsYt63T/WuCY+HfOmLmGfXGQVDnpQ6BbPh7
xPTN5k+yIhoBTRC568Qbl6uEuEB+AAb5Q7YbQUbiiD66bxO9zc/Cx+E8uKs6Kk1a0eaNaGOuUaxG
zMWj/z0sjoYWUsK+72N41E4F2ZaK95Al+nwnXeO1jeq7jTu5LOTj3sSS593pMYM5NM/wCy0n0TtQ
xGFtiQc6WiPzCL91HvOKsW9JiROG7p6FrF/Tuux5ithxjoAXwsRNubJJkvt6ft0Ole2TDUjHKkWI
jmKrXfmDeolkbrUAtLbMrX52Rl7z29ZrZQzgyi0yqMWlajAGwXTLodvBYBpbVbYlGJn/Yeem9yc0
cXOluEUenCw/AsSmsgGVpe/IyFh5X+lrVKwXpbSi+M4WKgJOYP4nay5t5UGAbYggLqkUhQ/qBgfF
l8RCYZir2OY4vWCShVHSiyj65ZwLM8s35Zd/Qqxwut30oL4FFBNKLOP2PCqkSriLt+ajuhDuehpi
OYywIB/mHqruHYNxUF5Cktzqn7u+RHfsV3JKUMafOxNLFvRX6dXFBvOyFmkMGnMICBxfxR6396da
XnG7GlHn6DkROviiG/kIreiJQaV70mQuanQDYx3U5/uxG5Z/+R9ntZ56w2hAF99Uyx2C5rhd5Quh
nFthp+LiBaHtzk5Gr9DdvQRGBrjalE8eEFapbS7jZWwo6FgEB8PUE4HMTPWOzTZEbYXvWwWG8izR
vGPNF5bfxshCRDF37KlmWfC/BW9QBofp2gVbw4WY+v4BQo2pYxWUgaO+XXIKB/VTGfI4JhXKGFJL
8GfwgKp/xZjyb9+FJUNq3WSGwP9FM8Q/SQHq0NCYYrCoqX4/pHXN5Lr6LC/jdF8S1t9X1BzLAF1F
a4fuM4ZgIUVJH0a3ymU9DpUMpALgeR+H8jtMvzVURZ/Iuz5QB9JEKukOSbS1uBdUSZmZlEz0wHck
ExXQ2DJ8ErWiEgGz4adF+yuWFmwY0rTBbGZYKTuN39ne/Y1ARO30zBHqyeK4ibJq9ah8kN+sZqi9
VBpS1clzXKNFQ2mWpi5sahHe/LeznHFLWDJsXzQX9h8cc/jjrDKGeKjIbtDbFe9oKtsrg7twST5k
xXNqZ2voE6nCia4IxLvfiSKK21Ti/A7nXkgm2GKES9SWpadFUrHk9uy+3fvYASCMw7L5Y7okGP6R
Vwtj4Lbq1ILGntYk7yVfQlONEmiEPbth/bFBeMpuk6IWiFcvKLXq/ELYS7Qe0gX5igHEBLvNtgjH
iyn+gZc08nksrLLFWhQqCXFr+/oUWsrVmASOdU8ILwmjhQ5sg/GS5aPVDZCeV9S1ULSOnQgnrI8n
QaaALzmJ0OwaxqwhvINDYonzTm/IBzCzSu83zrmy/aOgq9K8rgNLNBzZhRmRyRD+/L2CaoU/y7jO
DzY9rXHm5f0NVEoBQ52v7wCdl8tPkMWUfREdaMX2H1xnsduw/sOayfF0bzoYBi5C6KZer7V47N9u
ALOhEon+7sQpTtWr9IT6JQw6F9z4liglUsaVxcqssK+BCLxGRN9uNaSnivcQcbSgENZXxMGE+qed
0rjasx2PZu1qroLJpJJAhN9fUx4u2RrdeHPUtWT5WuhGhO4ATA7sirqCbPbcwXYV48b9TgQ2f8U5
8+RM+a2fUE6ucXgtsctmpjDwNCR8CAFv6UyXmu7MspWPI42lS3QBvPogSp1mEOgDlX0+kuhF/V1S
b6xbLtXs4epJ5MUnkMpKps+u/64zBRRTJkt6D9372quv7wCwLP4IPbTJgpw4RGR9iXZCmIM0UAmZ
0isBlU2cQDs1/CLGm+CdEZAJHRWR6OhJa57d9MrwCHpk4bJ2OoVlgCx3mLsaNUj8KRvkZfYK1Yab
+lm/xKNmFXoRcgpf7gRLgjTLk7Z+XIxu3gyS45golhCt861+gQUwPDUSZ/BLrSXlhJaOZs0mAc3q
p9A/KvNC6EoEVZBAPLgUYk6Lm2Iz4CU0Lfpqy5bZsinBacEzYPEZnCld7TRTKAA0N8Bpkgzlak76
08iOnxIBZjEHjwRESyRpu/Q7lPxNBPEJN0O4Th5nsJfX/IpUF6PnilBmKpTiomfh7F671Nvo1e+6
ocjJgM+OuXlZgCPV4TK6Egzci53cb+CbQVDP/K31wDvgr1zzozapHWevUQFhDaMedqjxsF+u8eyk
iwqD9XWac5EZ134Kz7Q6PKbdYOK3TgRNqEIKv02Z4pZWbCbjql+1DsJnc0SBdO0FD0wUJLT6oOav
pFxaA7yVB/coyyOYIKMNlF1c8QpEWiUrWrBNHk50XxDHmOoUqQ1D0CRtdaL4Cwz1rA2XUnT1uxpg
JMCnEwn0VxnwydHzYknRqn0oD+1nae1aBEkm2Y0uDQ0aQfHIHESa0Et4usou2G1M/oD0qBAOqaq4
yMvTb/L2Mo+kC6b2QZJ1fBhCRSLn7IknDxzEYa+xwGf9SdJkMZqXROf5F0QItg0fAhYM9BmwvVcI
DkKL4xdZQMBReI5fbeIOOPxKHAsclCExWPLdBgBapSKre6N3rRbqVb/S5lkmBfYPyPXxPU1akP85
zTmSw4jQx+9Ep8HkQ46Li8o5mWU+QSMTPKnvNbPqcwMcleTTSOZhhyrQtjVH/TiNxq4REIYUMenN
Q5pRXHFXIGBZNihfwOr39b1deDcIygWRjJzMaxQ9F/mAZuRGFgYK6vyFSCWfc4w1yLrIiezoiZ37
T+uA2d31/J4sR6LVZW1dFEKD4l9dYg4WPOZzKFqgcdeOrsh9kwcymmzHCDRhjAprygRwojNC2ToB
Ep4YksiHa8vb2rf++O5mHuBjyAwh5wB87AhQKwx3LPVQTFumAGIriVe1kijunLWUauIIjM2CmH69
GpT88iX7SkhKoOl/I004AV3Ok6oZuE3u1Yvrwuxb0TfA4SOeReJhxP79IgLI7fTLTotYcRF6yj7L
uu/ZwWIMdCy5FVPvmeYjLTV+LxyQYE9363DCq0+Q8H9MwGYSetpNEhDoa7jlvE87yROESSd81bdK
C4jejkz5qAbqJSJ58D51I5CSh2JsFt7gD4DgC82bqxwuDNGRFjcDbQEy19ps019tS3/yj8bEzX/m
ctm7pp4DJ/AqGRMm3mwZg3WOeIjmizd3iBB3y+w=
`protect end_protected
