XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���0x����T�=������44(!�|H�n��[}���fcV�G�x�ZǿE�^�f���8Ɇ��;���0��6�Z� J��O\�c �����>� X{ߥ���E⑍� �|kP#h��i,?�����?S�2zp?�{���d4gf_>�-�FkϯF�Tu-X7\�@
m������ς�k�i?V�v]ơ�i�D*?9z6�'�7Z̓�4c�]�hS���6U�wp5{o�1"�~#%ۉ�z�ׁ���J��Xט�����U��=�*��b� �����AB. ���b{���%r��Ǝ_��
%#�*>^YK'1�R�J�[��B�OOY~���@�\�挦bjY�_�`k.��٢�4��脍�0�s�5�'�ǰ�R�Z_�K"*��d�#��p��z�.]T��̫֘�;�6�S\�͆Ϭ�W�d�þ%�7�t�Iߩ(�&��67��Wn�pJ�8J��5~7"��L�eiʳjuS(��V���1����`�	^���r� ������fUi����#�^W�ե�D6Q���̜�W�S���J�*!8߱eY��G�?~A��S�&��K���>��(�:���_!�X�K}��f�,�^���� �eF��� 
G�Q�Q=���1$o��D`�c��WS	�t4�x�ߞ�!w��g�����w�6ir\���GM�<�|����S����O:�G�5{��{�-lL!��>nC���+3`�T�ck6_�B@?�ȁ���^.WZ���~=N�'�XLQ1�ĂXlxVHYEB     400     220g	��P�������n��^2�m0vԉٖͪ��VbQ��ECg���p�u#�'(��U��0������
B������+�a|� ��3�@w;dI*�6->2��I�u"tI��������O�r��bN���j��mlӒ��0������:�hm�_�l���PP�q{'��X_�E�����X����L�T>�@�;
�5f� ������F��]���j���<�P驰Rl�/������
<+Y��@�|p��L�]��6�I#��+.�49����Ċ��I{�)\���.���0�w/���>���/v����t�D�D8:����F���:{L�tN����H9Y~F���3�ڢ�C��q���=V�YnT��Zt�� zW�z�1]_���@j�!3�&k���<�ė.v�}�K]M=���ic4	QFQ@��no��[&�||����'k�8��fai�޵2x��4�\�(Q��
r7�����vz�s��$q��{��H���G�"�Y=k�"�j�L����0�a'�����XlxVHYEB     400      d0{�4�RY��Z�|��>���1ۭ�Fd�EѺ2���%EI��{����=*�p��쿄�*^6n�\˸�i%�Q�=kl<C��uޙ_�Rh]@54���!�Q�|d�m�v����׶q^"ޫ;h��n�W��fcmἂS�ni��+<�%�C`� UA�H�^'���T!�a佒�
�wA/5A�!v�02��vn�G��`_<OfXlxVHYEB     400      c0Dp.�b����9k��mG�S����_��SQ�{���]�[��pOT2[��-<�h�S	���_G��i7�W��� W�]�^ضVg2d�.BF�$���?n�22��D����v�®��x��		8	<��0t��r�;a9Nsa��s��쭕�@�m��u�>/�q�xJ�v9OJ���񎡀Wa�9T�XlxVHYEB     400      c0˻:��w�&ax�%g��5	/�q��kj����PΈ����ҹ��^-	�(nP�K��?�H�<8�H��?���;	(�4���,�'�#�aJ+�p�{�h{�&=H��W8��K�R�f������b�¿𡾁��G%���S��2-���j��D$e�P��՞���c#�)h�:�	���#Ynką����&$�XlxVHYEB     400      d02��Yյ̬���T�kLb�� �׋驇�:l��Q �NfA����#���l&�P��̴n���O���L�qy���u,�h�hŧ�6Q�i&��o�7�И��h��d?� gH<�t0b� GV��xh<��#o!^p��(�A�S��z�-����R�/CD`����ꪱ�eȔL��Њ�n6}���jXlxVHYEB     400      d0�>�]�jw���ɶ=�ں̓n�G@ck�C���-��Ԑ��A(�ݵ>�WƦ}������_;������S���01ʔ�Y�� n��i�i�sCG�nI��<o�2˗R(̇�43��F����6$Ҿ�x6;��*f��ۉ�i�tk*\p J
~FD�!ؠr��+U��-���b�^�#�������M�b��07Q�1�CXlxVHYEB     400      d0���ڴ�N�x �$�lq����x�I�6����_d��aZJ�lf&H<���+B��h�ճf�E�#�
op�v�6{�����8:4��%�U$T��7�Z��0���y%A��xhD�;��m\X�ǌ��Ř(8�JU�����/Ae'�n+ FTwL�`9!�3�Y���J���(ߌ�?� �]�1R�+�y�qwZZ
a떩L�XlxVHYEB     400     170{Y�1���k�[y�vW�7�#q޹gc���-��A��r���'*3�ѳT�:J�g�����ƙ�ˠ),�����+v;��$���$��~�K�x݁���^�j�Fxb��A��UܕoPli�`�
 '�zp����b=�9tk���[!��GE����z��+�� .S_�WUx�wU3Ͷc��PK�)�����Y�#'nH6(�];\4�u���2�7y%"!I`<����pѨ�>y���̋(�GK�lޭ�F8�/"ݍ�N�4!m+M||�A�2s�N���k=][����9�!i��*K�,�W�Q��)t��V�<�z��`�+i��i�{�ؘO�Q{�^(���'6<W�XlxVHYEB     400     140�O�I�Ƨ��L���P�%�,�+����Ļ�W�@�NL���Zr]øKL���&b*�L����̛G׃�q�M{�_�	}��<pۗ[�q.�&��L�S.<�����:e-R�3z�h�8@�\��s��3�A�ӱͨ6.��`����i�QŜD���G�R���n�õ�c�q�S��X��7흆]8�z~���}h�gOӫ�)g �No��O/�����շ�=y��^EC兾ZP�}��mS�����T%J�4%|��{�ϝ� |���QC;��$��x	A�pg�:vi���I��y꓎��.���=6�,I>\�XlxVHYEB     400      f0W_�P� ��Lf�K�̓��J�vt���/��3�]�/ϒ+c���08ś���,����gS�k<}#[1�/
,;�'I�A���R!T�J'ɝ ��Tρ\B��h^�1�l�t �E�� 7�G�+k��c��e������}�Q�g���[�l�Ő��6�y�Tf5��	��%�C�h����M~Rݨ���W�1� �'`tj9ZyB1]&��O�9
k�����s��&a��Js�cb���XlxVHYEB     400     100+��݄T�S5x0�{�(�l�P�������R��;x��R�"*;���%J�j�7������52�=�~s��lR�Q��/���Z��T��!��]��0����H�b�h�)5������U�eϪ7��y� FF)�����Ƿ��Ԯ�@(<��A�>vqLVwPC�p���G5c*�>��V��8��"���.��HdoF DޘqJ0�ŋx)�81�Z�����L�;Km٥���T-�J��ӽ���.>��XlxVHYEB     400     110n��-�v��u�w3֦��6k¹W�j����+é-�ǽ�c���K��X�_�^�e/���!��W�Thp�QF�&�=�N��B��laz0g|�,1ӻ���w�`B���>?�^�!z�[lgV�����I\��8&N\��YSp�F�m9e���X��w��Ѽ�ܛi
`�/?G�S
�=trĐ���]ը�̤��h�D<>[���O�b�MH�&y����� 9����N�V�#!��v��d �J�~:=�e�ps$c�XlxVHYEB     400     110��@��/31$I�}@��|k�A�Z�Ht�=�XX$�	։wV;ٛ�G�����Q,�*8JجI�<P�c}��h;aL����6*=���'�50�p�WGi�&`�n�4C'ˮ�?]2�Hz|��7�;x�����)Q�-��E�:�
F�8�sQ2�3����:w���d?
�o8��G�;���O\�Z�mz%��/��Z�� ���I�����fS�!X�-pd��1����ҿ�$
�^�71�W�K�V���Uv������lW�s�͖B�XlxVHYEB     400     130���Q���&��@��k�6���I�%�����`<WI����=��fY3#�c�*({��j9���~A/��U頽���p��ο��]���|�M�x �9���s�;�r�^���E[���%��5�g�W?9>�_|Kr���є*��R�N�ٶ��]^ �(���PIX�W�s�X�_�Utp�����S��Ce�Z�o�q�j
�֩��JI�$H�J��K�O!�mbA?1��ʊ{�.��׿,q�0|�-f�
�J$�S���>���z���i�_ ꟞ �=����K�,������$�B���XlxVHYEB     400     100��*���M�^-6
ƛrDj�{���a�P�����4��w5T��:���|S��`l�N���*R���߸�^��Pl��;�IP2c�=;�8�Q��{�ղ��9v���D���D�Z5Ұr�p@�p傢<*Ɋum��j�r��Ty�1�E��WS�)�^���Y_��ⴞ�e;�X�m�<�ݶ$�k�A�*���#���~@muʦ�3m=��=Y�H[�2��T�3Yf'>o�h����5=��m�w��	SA�XlxVHYEB     400     100U�UJ���Y\�� L��Y0n>@�ǜE"�itF5�S�l/���{�RM��@h�L�I�6e���FT�2Z#\#��J?n{V���f$x�(���nP��5�{計��V��^��
%u�^�K�(w���3�����5	Zx�-#Մ+����^�uX䳎��}9�6KU�&}p]�ަ�xb3Z��.�+�a�py)�]�������H@Ԙ�� %�5Z�Q�#d֦F�YTQ�%2�����0�U醤��dˬ'S��j�XlxVHYEB     400     1009��8hD�(_��0�������P��xk�w�"�3k��`��էbg��ogd���S�>��g��,z�ؐ��P���FHo���;0(5a]��p>%_x��:��w$����6V���E|Bb�'C�������yN����?��g��G+����|�i
����I�:�Ӱ*>���eMFu���ɚ����4/m!+�)������Z�V}�iʅe��X�����ds)�}��b�ܲ����2�XlxVHYEB     400     100ߐL��@��z���vfQo�QzF�NJ�i� T�����.��	���֗�l�tR�$�ƓTb�UjG��<c��Ձ-�j"���V�j��	�r�s�c�`a^/ �y]��ս�>��r����:���9L`�g�9��,���Cwrw-n�`8��}fI[��B	�OK�R�Ѩ8�A�&�z��)�+�QVD�v,{��H.��OS�aK�Wc��^=�t�X��=�ᢒ�0e�C��SH"�X3m_�;��P�S���6����p��0XlxVHYEB     400     100膦�`��O��q�cϚiƔ�<N���^�/H�Û^���k�0D!�'ϝ�_�9�#�4�e���I�S���ۇy"���>����qL9�ݴa����+���Lu�bȣ��ز���$F
�ωW[���qA'd>�f/������i�
�=�+Luy)�b���Z5cP�Ql!���]���z�Q7�I�m\,g�s�$��Mq�-C�C�	�QQD��	�Zm����%)VF��8r�!b*Ȣ���}�*[AҾ�XlxVHYEB     400     100[S��Tn�  �S�HXg�s�*�8g��$l!J
[��J��fc��e�8�R�;�,;6U�uq����|)a�=�ٓ�?K�УU8Q*��[��K���g+��Vq���\�?�~�an�.�j8��Ƅ��<=���@cu�B�C�nYaB�>�'����̛6����萞i�\�M:q�/+�>�A�I�@�ƶF�����'�ߨiMo��Ϫ�]�mQ*��P$�w�����.W�ߙ���_��L��m���*����d��XlxVHYEB     400     100A��<�����WT!�id:����>H>N���|H���pM' ��YF5li�mg���`���M]�;76�_���j{��I��ͭ�]��^^�-�zV�4�<�3b0��0'���ߏ0����hxq�?̶�
Q��ɘ�o��m��Q�z0�e��vl�7�E$�%��ĝ��hC��x�i��Ig�Z�ׁ3KC�6�9���#��|����kaw��Zn�lCo�(aj_�LT{>��uY)���銢��g��N������XlxVHYEB     400     100,�N2�����Nd�Q��H�[��<��*�?��o�g�WL�˹W�t�P{_�I�dp̏�S�ÂQ`�
� �Z��<w�^xX�=���|�O�6���78㩮B&����d�pH��O^��ۃc�=D"a��eb��i&}�}iĆ�s���TfyE)�cqH#�+�z��5a�&q����y��1��m}�7Q��0lC4�_�0&�$S�@w�%Fgt�d��<"�Hm!�c�����ϊ���J�XlxVHYEB     400     100|����ȧ���_��Bi��+��*~��GU�m��
�i�����BN��l����]p4�4�-x�P��eA�L��C�Q���-)��@M����R߾AkL�����
)ܺ_~�����7�p�����I��!��F�?���4�W]���VۦF0O��8j���k��ӕྡ��:_����p��C�Q`�Rg��2]R	�ۣaJ ��>y�@f*f�3�S˨�4���N��c6e��;�̝A�����XlxVHYEB     400     100�r�<�-��w��	����:�m���3-!<Q��X�ܒt�,������OC5�35�3:Q"A���fO�W�8cE��v�����瘢�į�NV�|`���R�7GZ��^S�d��ɴP�ld<����4�#��9B�ⶨL�UZ"�e�:j��#���Kr�B�2D�0xE�rWI��;�3���|[�m�\nҕ�	]A�W{��;�p��㪨 �Ǩ(�u���T��{���h���R�IVWXlxVHYEB     400     100k��![:�S�n�����HF��s�H]Π�*�XЇNGKBQ*q��d��A�;�����͠�PBGX��4���Ѭ���Gg�8}��XkۿB-�u��:)�L%�@?
�T�/i����
[��jۚܔ��Z���K�ۿ�Zn>_��<d�9�2�/�>�HS��ftض)z ��*ʳ'9x#�����2��2Oo�i9R[�����ed�ߡ�'0��T�?���N0?�Q�:x؞� L��ATd�5�p�c�=��v5��XlxVHYEB     400     100n�(s��ߕ��j�06��Tc$+�O �u1�)7\�U],�Vm��#� �W�ŕq���KQ�����Y�r�Y�HL����7j����5��Fx����l)�g5���ԎMՇ��b�����緵{O���s�R�1�{�Q�ݵ�����M����J���(��Q���$M�g?V5) ~ ��u3���Lʇ%
~�(��=��y�o���Yviæ�,��
`�[vtV��{����B�Ė0ZKR�v߀�_XlxVHYEB     400     100M�a����/`@v�����q�^	��G�mmE�'�]�8��;�*�n��:ma<�|���dTPa�O}*(��0$Z�ķJ�y��S�m:~�2�G���R�5_+�xC�	�#\tɈ��8 �N�}�s���;��b�xDg �,����Y�uIK�Kl��q��;F7��XNd<8���u��D���o�5b"�\��}��x���J�yC��[`5Vb�����W8/�5c���B/����1�vW�*�XlxVHYEB     400     100��}���|��%��s�����~����~�i.Yo\K�'���\c����DP���M����:x�ƶK���D}�p%s��q���'i�U	W����}�[
G \��6�Ǭ#�Cx��	����*��JyJK��=�p�$Jg���K8�&|���7{�Ӵk��f3G�r�F�ベY�A��H�&r�����_j�2AĂСS�L~��7p9�������jA�u֗j	��m����y��#r��/��	�:�XlxVHYEB     400     100�
���$��ZʵX�c�E����8��l4���i�O̬��}�=�������?_ �8�SN�J����$:PNg��t��[�V�#�4V�G!�b�Q@�dd�{���\*����^�"=師�{��|��UD��#bv��כLk�7-���Bdϕ�W~�6_�q:Ϣ��X�4�Xщ6�3�>�5[�&����(H�Ê���ꇕ݌�DQ@S��z֏�B������R�WI��;�����;$�"Z��DpXlxVHYEB     400     170Y�3K�tD�NlB_?�ggt��@;�O��\�-U�%K�K�ג�\:1×�GS���$i���PJ�}��� (&�ڗh��<W����,�7��7���u(���`t�*�К;��PE�DS~z�loH�E���Q��L��nѾ���/��߹� \g����GV�9ґ��=��߼rT	�#��i��XQpV������Egq�P��.\���3�M�֬8\2͇H&$��д�4QjM�f��U�� kv?�0٩��1��vc��i߁�q`y??TՏ64�����-\��`�`�l��Q�6��ã��pb���8���/����:�c�}l�'}�عp00W���V�|9���6�cx8XlxVHYEB     400     100���ղ8�/W�Z��f��~���En��0��k"PO�I���۾��ڌ�qcz6��&B���I������Jc�|'j��њ]U�<%�,-<���^+w^o
��S]|�1����Lg~��?��eϻ2�������v.�c���	�`s�:��	1d�`rg7y;p�|���m΄o;�)N�?����3(Kǜ�&k�h�����N__0U�HK޳��\ ܃?څh�6�?o�i�BG$�
Utm�?���W��*XlxVHYEB     400      c0����S:�C�CiRk��n�囐��c��'�}
��t}�(:C��CJp��Tl������U�g��
��nG��� +�ƒ����l�Y�WA��~.�Nk�C�*�<bw@\-�+ݖZ��!B�I����h8���A�{/L���~�c��@�2��+�"��#X���F�>ݯ�ґ��/�ʣF[D=��u�XXlxVHYEB     400      b0p�C��}3�Ǒ3��-����L.%���E�=oU���y���9����(���� 3
�ԓ܁=ܐ�6i�r�,1O+޳~_ek��w�aF������!�>VT�p-&�Y�<S��Y�,fG�u�0�ݥ��u�� ]���*Ś�P�yJl�<��܆`�E���l�BdRd4�XlxVHYEB     400      90nI�ݵ���g���&���O^+E^�Y�ٿq�Ε�Q�\ڈ<��p��l鄰@ַ��!Pl��/��x�)��:������/Ajr-3Ϛ��Y��Vg�з��E~���q�l�C���f�F�럒�RZ�ťN#:Z,/޾g9CXlxVHYEB     400      90i�a_*���y '����̋.�����*����̻����k*/��xfgt&�v'`ꖜR�&��Ōy�w�m�K�U���~)�	VmKn�T�Y ��܀{ �k�<��w^iAX`��Z��/N�O�A�i!��/�Ė^JXlxVHYEB     400      90<o*#����N]���HTn�"s,y�J�@��7�뷖�<��\�&Yu.6�Rw�"z���p�zX���<�º54��n�2Wk��&p!ґ'��3��� ˻��r��&?�F�q�߷`5W�(�O��?:T�!XlxVHYEB     400      90�b����d�I�Vm�w�'���NVnJL/�ܵ �=�uq��9K��b��sP��s�����=����B��,񒀲��w$-� W�S�=����M<�#f`<�V-ǚ�&�eF�r����4�ﺶ|t5[?����aO{���!uXlxVHYEB     400      90o��
Ņ�=�#Q{v�p$H������O��ѹ�To�ɔ��M�9����]<��EX۶aWgi"Θ9~9�<�[1�]ᓾ�Y�X��& ���J��r4��6�����^[�����_�{B�g��k�t/+,5]�����4:�fb�XlxVHYEB     400      d0d���t��(�>̺����q�(fC�W5ɻ��R���+Y��S�7T���Z�H;n��x���&��p�~�:���J��0��&) +%�k讑%��N$6����g̲��p��A!V�����X��K�M�ƈ�Wp*�1�Q�����3sp����z5�x�E$@g����	���E��71�� g����.�x`(�sO���׹��
�XlxVHYEB     400      e0s�۱dp��g����������H�^��:q���,SuI/B�D�on�#����)���*��ʗ�S���&���N`p(�b�I$���dkj��xϜ���|���*��L�<��3M�ЋG#�y�( �Y�i{7��o����|`���� R�r�Lᐞ�� �'-ZSr�2 �+Ұ5�kP:�(���5� c��T��($Z�wj���CøpXlxVHYEB     400     100�DC�{� >D=���ч���y]N�ï�:��������K�[f����{M��K��l�B� 4%�8B���1��
z�����K�������:���5#���1�{uߐ>��a���rtp}����c"�8��>[Q$�[��`��Y�.����(����30 V�_�����6�BL�r�`�jO�V�Rr��8�Ex�d����]����Lc�]ۊN<��̃׽�����eȿ����[i�X{nXlxVHYEB     400     160��ճ�10��y�X�C��m@�$s�Q��ɖ�w%6���V�zC�E@��]�y$��g�}� -2f��n;$U���I��?�C[�k��x��n?̍*!����9�j�m\S@�e��e�V2�``;|@�g%s�6������*US,bo�+*�N�8Y@`�@֛�e;�eN���ȋƋ �'�R�<���#�r���E��]����?��X��� �Z�[f�AËÁ�.}��2G$��%	*�Gs̡����9�pJ�`�˿�t򐀏�U�R砐)-̓�}�F�/`��ZCj�<+Cmڙ]J5:O��b�@
䧎�l���(Yk�o���Y��2�XlxVHYEB     400     160U��a��޼�,�&O����>���D����)	�]l`�O
�yc��wL#)�YL"B�=��*�)�����8spۦHf��2�:C(�vJp�RMP����ǫQ�p�z*��� �����Jn|��d|k3Q!�,*�O/�G�NT�2&!�� [n0�&�<�2���_\vj�U����@����
�<Oº�	���E��ec��V���3�=J/_�����	���Z�����Ђ����h�l�b��iZ�Ґʩ�o]�l.Xfa��?��%x�Y��e}G�S�a|1g;2D�_ٜ�&X��Vf\��)�y����(q�/�)|"9��%�i	L���V�a9�8�^B��MXlxVHYEB     400     140�#��b.�Q�R5�����D�5x�D���6�8O�?���v=�1�sA$4`Zn���yN�ؽ0�`�1	��t��悡�$�b�Ho�ì"��&� 2�B��z%���P���_um���'P>w�j�z��x,���]���}�0> �!�jZf^6O�6a�SN�כ�NQ�#-_��)ަ��3(������%�o�b� \]T���U�6������6�ʴ ���_#���3S����b}�P69�|��\|�Ia�p�;&�;����?�*�0^4�ŉgՙ��~����orÊ�5����XlxVHYEB     400     170��0P�LhOz�xm�?\V7Ĝ�|��w�>g5�g����n����E>��@�2��[o���2a�L�9�O�>��
�ahٴ���J�(��JB�@��d�y=�Y�����s�-�t3c��ߵ�E^�&�}�����1!t�EU������c�Ѵ�+\���^�����E��*�r��ϵ]n��;)�.�0��NT�&K�t-�؟(�l,'���\������X&��j��+H'01�w�,�A�ߘP�~|�T�B�kh�l�km�M)S�4���aW,��W����=�\e��7d�(I�e��i� O�?�LG���$�VT�E����F�W���KJ�Sk�I�,* }�/pd�v�+mz<u�!�����jXlxVHYEB     400     150h�s7ٚ+J`q�L�}��˝� �������NWOk�㘹�] o�i�36���3��`���d|iA\jS,+4Q2V��w��o$���V��� ����q �871U�vK��֐�@��F�����"��V�K������HT�f���?�����u3U~�
�(tx1���x(�i�Iȯ��n+T����hr@��տ+bD��ȞpM�������G�B��z3f��s[DU�'�O�2���S�Ь%�u����vu)z���
	����=U��\��ג��m%�s���2�_[[��N��]��A@�2+�;P59O����݅YevU<���XlxVHYEB     400     190�6��]�����AI)*vK�k�?Ā(��q��t�{�C6U� ��.�07�w�����
�b9\R}ч�Z�Ô������B/��1�ՉU�-X	������4h񊀌����ِ�O��D�NG.�[�O
+�7|V��4��
*9���LMx�[��w�X��A`-�I�SZ]��Y��M����E�:%���y�z"��3�#m��aU�JeՕ��B��7�ÝL���߅��1+�}С˧��/@g��V�H�H�m	8�16�bRCޛ�2�yy�ID�����E��#�V���U�/oԩ��f	�"MC�˲@cO)�:�]�FZP�a$�/nv���y���T��`���J���C����G,�e��$pz����[��`M~�Q&�qʡ/|���XlxVHYEB     400     150�B�Z0k�fN {.�]�y���)?'���P����"���@�������>�W�č���F��5�F��`�}U&@S� Bl�����TV�B��
�z^������OX�.[���̍F���L�ǵh<���<�������9�)5�C���'��g5g��4�^�捿�(�tj���M*��a����<��5��mͨ�C�ϥ;���Ͷ�|d�z���+Iԏ��bf\UF�<-�͘�>���e�������,���T�i3��|J(��W<D��g�œ};S�s΢����^�=��Ғ��*�tߪ��'���ķ�N�5 �L/#�:
�OJ�XlxVHYEB     400     100�)���q�9��Yh�E���M2zT&n��7w��H:R!_&�TKb�a\�FX�%ډn�J@�F�6��/�ڴ�h����JD�"�t���Ge�(F���1��f�S7��������Y]�aVwǣ��t(�F���Яcvm��4R��k/u���6A����q��֬���p��Y [3rH�C|Pk}r~ؒ�4��`>��惾���lqr2خ�,ut���L��[7~�0���zG���XlxVHYEB     400     190�c�_�����|�����f"^o}6���7W�vn{b~��Ja�`1�i�<�f��J�_\4�j_W���u/��Mhԭh_�-wk�:���V���c���S�Ӓ����"o�����$�_K���"�E}��H��Wf˙IECo�QlXJA���y����(���{�d��d��䑬�q$�������&�1/������K#IM{������P��:"�Q���y�<��q�!k���}B�
}���D6�����t,]��i$�z���⊲�bڇ��@ߌ�a��\b�`�9;�[��1E&/6��t�v�
��1MWγ�d��rE�Dgo�w�[�!C_]t%%j"It��,U]xOkLyx�*ǿ�U�`GL��Bz霘��G��;�ϸ�kJ%]?ZXlxVHYEB     400     140�t+_���^T������-U�z�,��|su@m�DRD֚)J�����|��Y�5��L�PP���NU3��́L�%�p7��,������Cݍ9�1��I�+Y{x�.C���y���+�?7BKݗU9`fUZ����j+�߀��`�CB��)M?��k����3G]LڛA	�wjL�s.@:�E{*E",��`)mO26v����g2��Q`�[L
t�Ҁ#����r0����O`O�+*A���r���o�X���N}��G�a������L���l��N�'�o: �#�l���%��M�鏌�G!�[��X�K�)��XlxVHYEB     400     150���)�* vܣ^3n%�8"����X��S�J��+�cH}���h�ݧx!5xF��@ӳM4��z�e6t����f^�	�6���]�b7��.}�Dn~�}HH�����(�C
�������E[�&m��3$��O��x~bP�k}�f��&ۢ��-�h3��uw�&hPĄ�_~M���i�R�R�>�eC���֙���wY�4A��ɉ�fs׮�SA��6)
]6����y��RC�j�j�TO9��%Imlܬ�s���l[S�����FJ/�/BLH��ˢ���J?�IyI� Zpo�ff�*�v~�j�t��g��7�~OXlxVHYEB     400     110�A1�ژ�?\'�À<M�T
@�^q�,�+a.?6��k���u��'�MX����y7=�7�t�a?��-�-K,g��x	����q��JA����N���|H�q�p�=�t���������@bI_2ʲz�w�N�s-��V}R�p�T�V0������H�ߐ_9��Mv�u?`�J]O�{�I��^m,NR/X���JK �#TQ����E�}>�6;4��T@fǏb�9���}�ԥ���D���Nlq���|�bH�R27�c'q�XlxVHYEB     400     160���f���u��u�;m���8T~��XO&GX�c9�~];6���.{�k�j�䪓�}ۡ��8<?��q�-��i��9�9�ၘ�R0cǌo� �J���T�eG��d �����c�1)��h���@�j�X���L��*J��>
��"O}ٓ�&�����HT[gb�ˣ�6�L�e�T�6��AԚ��l��3��kdj�b����!�%Ă����[E�Q�S�{L���7`�3x���	���mGR�
�G�}�vG�������Y@�S`O�ƍ&��~���w�$A������F2S ��nŐkg��i�%�F_\H-�7Ŝ'��b�p
����F��7�T�7#�����]��p��I�XlxVHYEB     400     160BakP�dh��rp>�,#��8�R=!O{B��%��/UQ4��W�L@�q�|Ezq���"Bn@-I�4�[�
�H/��,�5K���fV�PH�ǘ�4�]P�(D+��N]��vFks���	0�(�n�9븛v)Eλ,���u}%H_t�d��J@y7�$E}{�E���}�hȻzw8<� ;�g2�P]��SS�++���׭�a�tz~FC��X��у8�^�^b�Q+�4[��ns��ml��!�tv�\����yM�S��pΩ�"�Hc���F�����A�#�.	v'8fv�f����R\_��o��MvI�k��[�����|*'M�*�Q�A�����6=`���� h�XlxVHYEB     400     150UyhN+�~�	���ix��-Ak^�L�os�z̰^Ն�{^U�'N�'kt��)���	o�I���{���[3r�<�:6[Qx�A!�>G�w@�P����Sʊe��h�| ����ɡ�ha.���3�=�S�3���.T�3j\Ӣtf�(�>�p�$P���O:�qA�+��]��AnT��3Rg��g�����0|��`�r���@^d���,
˵������P��(���jI��N���~��9ݻ7�Cլ�/��,����/�90��ם��5:�o{��ڏ�Rc����%3��"��G6�@:�hG}C �?���ч�0�B�XlxVHYEB     400     150�y;;�I���`�Onˏ2�g��Q$�NL��b�S��!'Z�D����Fx��>D[�b\`� +,v-���\����!����f��M���.3*}N"�D:Hŗ���4�~�,�K,5�&|$�m/��̪�Կ�"q���jq��A��(J��a�M�q���JuW[�X���1�築5��}ԁU8�j�L{��Q�I��w���5���3��ۡN�N-;O�4�gǃ�/��[�H��tCy���v�L�y���!��n��D�ێ�D#^�/�?K�q>M��~�#zR��?x�$9V!r�sF�+<��xB�	Ǚ6cWl�����B'>��W��XlxVHYEB     400      d0���[G uBm"XD�	��q�����ќ�o[V蝱"|�#ql���Z����/{�����`�R��>��0�H���0?���Vw�:�{����s䜲�*�������]���X[$���2��u^�吰����S�YlW��vXt��"��E���Di�]��*�?��zAM*;����I���^P��lK��#�o=wnZ.��Z�2jI���XlxVHYEB     400      c09v�<�ma�_�^وz��B m�n*�m��l_||q�s�.��`�X�q7�n�d�e먠�EF(,��`
�eP(�u�n�j�=b{�$q݂�pzt����dV�w���q�M��4>��RU�V\ g���\[�30���-�O��6+8F����fB¹K ]94-U<����ڹh-�l�?���a�jXlxVHYEB     400      c0��5�d|�V�}-�Blw��:x��ڑ���jl� �Yb{'vzAo z��K9oi(�9NR,-->�rG��j���	����n�ԁ4f��s�y�����H;-	Au�M����|�1����L��)�8�-o�W�hy�>:�f�0{��1�!�"��/���H��m����T$;6F^?�� ��$��jB#XlxVHYEB     400      c0�7�FR�T3�=׾�O5�CA�C)]�*dl5J����-������b�t��+j)��oQAPf*A�|����H�m|iY� ����T^z<Q�����L1���$u������������b%[�#�N�k��-��=�l��׬��K0N8�;�?��І�2@.�B(�;��ǅ�.s��4���Q�2�Kǈ7MXlxVHYEB     400     100:��0��h����	��_�:��B���rġ��eqVa:/&Q#�P��o��WاnQL�1�Ѽ�A��O�I^�cց"R�Ҡ�i(^*�d����Gp�AT�+Og�A���+�}Hz��Ea�nd�f��y���io���ʍ��28��c���0�_.u������c�Ă-�˯.���~;�^���.��b� <u!Tfd�z;��6��M��B
��f
���
�k��b��'Je�>����6(�p���I���y�XlxVHYEB     400      f0r�c�Tq�8�Xu?��_"�x���ȷ��ٌ0?���V���_v���� ��
��Q��
�ܛ�6��-���Ek�&�-h� �^��WC�j�쟶�PT��ZǄ��`*��py>gqrLi̽� �q���-/2�B.U�HX��2��W�Y*��>O�o\��Y��(�m3������7�u�ʱ>kJ���,��j)<�S�D�T�c����?�$�-ڃ�t��_�YJ��ImǏXlxVHYEB     400      f0�SU���:#Ar@�6O��p{͛�Ҡ"TQ���n�<<��x`��C|J>�X�]�F������DB-vB���4(�1����0��M9�$k���x�U�s�Ȇr�1~��7+�v��2m:�	�K�k'��&�N��ji��p��Tۀ�X\t�^�=,�޵XL^X��S�Ou��{��ev����>Z�N�0��(�;�3����W���"̀A�|��.�pm�XdJ&�?N������h�R��MXlxVHYEB     400      f0ޅ+c
Wy 4n�B}l	h�A�u���B�LHgD�p�m�݅�$�K���P��o�}�j��V�"G�~�^��5 �G�a�5��)ģ9�H
p��O��: ��/�/3&lZ��!4��?�D�3?�=�����w�J�8���Bl���������׸\��D.?���]�[Fk�&��%@~O�`�S�c�o�1�-���d��?�;��0KI��j��`,�kbĕ�f6�n�ULu�W��J��XlxVHYEB     400      f0�j.?��d�B�]*9��)��	����F?{�[9�i�K�i��F{ �Vhe�9G����J�8�R减|Hjv�Σ�X��-
�b��e*���xi�N�/TE��*�uH�;�W�wY
��%I��!����1>ȡ]��鬵nF�m�L��B��4��x|�C<��<@�Qp[���u������(o�4�{N�\S:�8!*���8M�u2��k�Z���޵�b�~y�����h�(::|��XlxVHYEB     400      f0�h�'��'��=��|����_0h`L�],W1�yBm-*Y���ׂO2�wG�Kd6�=�����`G��7�``<���)|�C[-���j �P�w��j��駇'8) �.��D���ܞ�ur�\6'� d��V�r�'�sٔ�d������pMߋ���BT�g��k�g���~�x�*�J�%�?�A�"�|����@g�i%�J����.����z�Z7��X��jA0���&XlxVHYEB     400      e0�/�y�H��TI�ʛCm���$ޫ���s��ل��}�-^��Ur���v�@���C��d��=�e�ZX�|���tlB��Ҕ�~�u��^��f�T0$}�/��m)`���r��/H��ʟ�y���4'?Ͽ�j�,�1�m$���xiVb�a:�����*����DJ�L�*3��5��6�mLC"�X)���`{�����՚���E|��T}��W��XlxVHYEB     400      f0�mrtcD6�H{��%��Y2C����87r2I�>���U*�o��G�(���W�^ʨF���w%�4C�������"��,�6��k�\����!�r���Dn�D��H�nj?��p@�����ʵ�k���p�'z[�W���{3��r�����L�ir�q���f��hm�oO������cE����c�G��|�V@�6Zn��MK7Vg5ӧ?����p��>R�W�4����{���B�XlxVHYEB     400     150A��/6a+���v��ƞ��C�z �T����k�Zh�!d]\	���U|�uJ��Z��Z�AiJ9��#����L�Y��,PE��)d��l��i�d���Շǫ�L��R�^v+U�Q�ǈY��b\�h��$
�I������ ��J��w,Z߲y�<r w�7kd��p^ɋ8x�v��ˤ���!*�1|�#��a�OK	��V1o�Y��ഷ��e7)��=��n�9��d��x��C���Z����[�"�>TAY��E�����$�}�hB�T&����ے�F������͎g��A�����}�S�\XlxVHYEB     400     1a0#���ݧl
��R5C�	�������ة|#@����n3�t�̈́G��Z�����{�J�EAŽ���s]���w����T��_�_�ʝ�rh�]��0�Y?��LP:w8�R��K���%�ו�ѣ�mB
��o "�\�OR��T���U07�k�/!DǦ��ԝ���܌�KVL'p����u���,������5
�/|���3c�]����L�S����|����c�.�2�`��L�8�1�(�+;`<��OT����)ٝ��?�F)�$I���2����o9>��T1��F��0�����H[\ʰ��;':W���&(�rb)g�S��zhq�~�����'��I�@.:i� �T����J�f2g�j��cڊJ��y?j��e��MOO�.^DW�����IcXlxVHYEB     400     150$A�wR��A<�)�vR{w��}cd:�G7����ť��R�bQ-��GZCL���	�Hy�
3#q������L��샘�0�9{.n*��E��5U�!W ��Ƨ
�ι�-M
��*{��v�qsZ/w=�z5k����|�52�>sC�*ۢ�2p��PF�ۜ��
���dU�	4]n�gv���A���%�UV��>�m�6C���CӦ�r�M�K"(�>QD)����oOE���z�v�;�:4�"�Tპ�\�a>���ߛ�YBh������]4P�B�$�\�+�v�`|2�]��=w9uy�(����}r��%������3��*;ֹXlxVHYEB     227      f08��t�R���_X��3��ryv������~��̷�������	f]zB��HHB^�E+*�޹5�Ȇ�v���?��3�H�;�#����SB+��������;�)	���(c,!���3���BJ;o�Z�9%����fH	M�,kxsѿ�\�q(��t�m��������\�G�;O��j	��q>�(�*����������,
DD=�I��[Fyޣ�D{#���
�|�4����}EH�@