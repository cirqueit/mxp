`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50720)
`protect data_block
TwqvliIhF1ew/jQxLAvnLPG16GOkn57jfmXwd4FQU5EQPuUf2xCt9bJLMAwiqe2FnZwHD8xy1qVl
F5MY0g/EBa6JmV5eW9w2jEHNGkvofAh1GF2eoVkICABsryiwoxGlfOWnV/g7PQ3JgPjKiVBJi4g3
xVo8SR+VbpAaDQlOkFlyJTjdHOiF46oHmb67D6A2jHjmrU7tum+rvBnO7n9432U8OGBswsBOZCm6
/u1gRFyo8rln3H5HNxzVQfPCU/7Hww5NYPA9uGLtKatAtWVUqr9XBIxL5CICcL7FCeNQANO08bvG
d3UNMyms6yUDqoDsP41xXoUKzCYWZPKTdabFla0IUxi4lI36DzMUX9eO7+YmOgZHCO4W4PZrtwOj
0YKwvrQKVlUNi9pORIAg/r26wKIxBrMDwtHnRMPiwqw3DdfvjgT70sbhFqaDQmtFryH8ATt0uUwB
IUs+e5aya7IIGWN4RqALSwDKkWJZhROb2xtTcJXUlz15ZVRbsIIVoow0+5NPIhnImrufXfOPjOyx
10rF1kKo+R19wc0LCIUSSTREdCi47oq65QAv2wPVJqly8rYfv6bzUcziWDcLFVzaeAmkm+vCwrRl
TURW1tZ3dLbrLvfFhznXzTkH3TBWAhaxAZh79PiJ4h3bW7mElhiQPrpai6tIH9rTufc+26gwZ8xp
Tx+y/SohNMAwfsM9lKHfUbSeZVXREpLW98bWQaePhu2hnWqUWfKdwUT4TrZzYtIwWfo/gPaVaQsa
IvqlP8d400l6qWGVFLG9hhja1V8gBaLMnjehXLrsS98WnfF0GlahjrRFpfRgsloe5lSscy4dOTgR
BaDFianuk01D/cQ9Ed6F/vJAfRslUmFFy2TUFbU5ezinQUAS0JOMfSaIiVvAChohlBVTXx6fvA3+
w0XSknq9LHDFefssTYOCz+cC5f9mVW528uNSJxH2fmx8czbv81pkS9YjLC3sFeY1udzxB1gtynpF
GjfkK7+LVomswNpIZ25mv/MCeLjY3WA+N+l3Z1CDNhQuDcYv+5WU3IT0HgSkeBCYt0r4Tgcyi0JP
kG2TvZySve5WI9CeP1cJGCUDQNvMtBEMBokS2B4vxaG3KJFbQ8w9j9SAIVjkDK4uDniFrfBkOlj5
zWf0keSlXSBj5bFcLbXKp83tF+m7veI9QXnwpDZSJUW/cfXD4GtFfTUvo2aM9XCBwDj5LuLaYJns
P9/iXMrenl4cTPD9E8P8unLCjjMklJd1S+UzBYg3g5KiBhe31x8lsrVT6FGVn7FQJvrB9F8+Dr+T
5TXfl89TqkGJk2JCXcyqmDKKF8f94w6TmeI8AzUCu3oaF7VDGyiD9mJJoWASOHdd94MnEtx1A+63
5WGuv7sRVj9TEu2bsXZPPy5dzi+Nh4/qGy1lv20AwMMBiW3knidX3ltzFzKoZC5mi1AaISj5aZbw
BclZuvlE6mIrRFfRZaHhWY9i7Im83jPpcFUDBMWmI6QJ/J3aBSYV0YDiZ5WEjjgCYt2MtqFg6BQb
2DQWAprphXVUceFs0fUL2tPbVVhfTc6tiavuwVyY/dlwrsxW/AsVm/+xK8WCXVOkfb64P+qWogfv
HLXIxanm23+o/gmDA8cLbty8fX+KwPHXQudibuwBm3TBRl3U4gII62HDe8m7uio67K4Ib6t+R1qg
4yy7pygn8yRiZdhD7W6d9kKS0Bi+FMZYiFatBAqwBEcV+9jCQsr9gk+AB6yCda2003rEzQq5TL8W
RsSztemaLvyAvHuehPGqmk7hgNd92x8FXdZ45w+jpJ0/ApfBWFOSQEcoU9wFKfZXUfwTLeFaJ/dc
mLqxGyI7mcD5yz3YSs9xxX7Y4HBtZR6kcVdnJkPJGUFhgC6E4U3XHOKNfAqfODvHAMGFc0kjrayB
VuZn2pwwYe/4XdM7ZN2S8t9MY80FLqgJ3rG3ElRH7P74dcXNiNfulaHYodB+ioEVz1rV2G3h4xqm
8WCc5DW/4MPignzlmFL9YgSGmEkC9yHzl5zXdRE+NjXbm2Bs1lfsQazYN6kA59knGSYUpagrTO+h
0bLfcHleueXi6oqpu/OMbNTUg9bbqnvpSdfv88NvIOqraD5yarCm++nYWW+VVHXA9D2X8gFTzqUy
59mObc4YbhY2OMRrPLzgfjNz78sAFLEQRahUqryXkq9D9dyOtu70ah5xzyuQu0HZpwow8xNKSykv
FQ/5IxkNMjouK6FWYFSjp9FaLvcq0XbdLB+cj8irscnnRgbRKf8KH7+hSa2NS2hJNhQH5s2bM8Np
JModoXDw0s/A0dkE+/qFPNp7aNHxmT+va9B1buXqwHzq3iR1OqdhJh6wfxV7u0RoZ+2uHVVW4woy
wvWRRt0VcKNKvL6Vbw/MKwsf/gM0m2Le72JJbDa/4ntcXylMbvTYcfiWHm8KtlYwdkhvFDJna+b4
KziV0kyvo7JVzWw/FhR2ksbv+wgKM7MNjimDzZtWUKungvJv3w+iMDLDlE+SOpniAKvHsQyTm8Tj
aRocBfSW1flqSzCnUFUkyPElToERZ9imTKlArtPkNa+vdMy6NBT7k2oxz0RHQeuIAAlyIAlWf2X8
etNdh9SUk8ysDDy5yHv2jnqtaqXNwHA5XBEii/+tGcUMUmwNHz9bfM3j1wbbDTEUCaDpQBHpSHi/
PsJSZ33larJQXdWTk5MYo8WCO69Sv/u+cQBdUzskF9pzVlq5QRNxLVGnbdxHUNCHl0aTOCOMvdo0
QvF9IGoV4VrvvYLJrM3lKe3wo9f9s8qZqFPh62Of11KipFMkzsJXyDm0CNfUZKK24tXRrbYbtInk
13Hs3TIR+tdTY2F0+QOqZQW2TjL2Q53se5axg5K2lF/E4qg9/+ImHdSN04jOIckJAYIWpoUaz+av
yS4rtvi0f1Ir7UefzhrdyvNd2IftwP/LKX8MUgUA+7SZSvTES6+qBqVrk9Z0IHyYK9U9Q/593/O5
K8UImAhjoHVptKQODklAOxD6ISHh9qYoSH3azhxVBRWk0k/k7zifELsx/Yc5rgFjPFTHkzu/ucmm
bnzaFHECdGYeodCv7EDqY+lqwbH/fe3Sdo983Dyu5XGAf72x49UWDBllYSJKSNeJuWzqxeOJmAVl
MYk6480J5+5i3LfQIGsYl2xLzuk/DwqwH+CxEMDWY218gVOoz4iwdaM78PV1iX2qX0wApvPXpi2X
4WGhfGGhOMuQlqbXlpSD95I3VSBrCuLZ9l4rsDO/M8WR8RpVOTGOWsTvLfFEvJSeSyE2gppprdnd
VRYWH5YrLLOjBawqVjeFZooZLKZ39lZaBN/sHc9X+h6CUkhwdxEPWVQk44Lcdi/6R/sfGte/hlfM
4vKGke2Fe/EtuuNIfC8tBcJDgODqKDvtMucVEjX33Mb1q5ylNNsuN/gbuT6dYPOB65DBwYUqQkVO
h25NRrUR4K4V77oE4bxJv+YL/OXIAqjdJy+EqNVATEz2V2BjbBQ0K84EA0THJlaPwGe4kWVJtIJD
ouLzaG+xppgr5vzC/1ynMshG2qes/5TTegca0V6S8JLA9ijRO8ykH7G3isc+u/qQ3G01i+NtngaF
0VX9xTYfkbevV0pK5mhxshscpHRnByCUz2YcNrvDQq9wWOsaX1CgbmTt6BrpoU4/g5k68x31e3hk
Kpd3r1uvlBUkDkBrUJlMfU7R/wnIr851DwwXo/aaNE5QwbixbyHEthpijSm2QCwMzsgbkNWc7Rzy
XBVl4j4yDY/FrU9hnknvhltwwkc4kJ0IdH9s8xrobZZNyCuF6BLhejgrKDUbAs5A0j86W7v9X1WW
RCVB93Sfa+EU4qQ/JQNyH2O2WIxOYTzZzjKqvgA4Q+WcbccpuYpNy+E/yho17B4IO6GFsN47CQVF
eCplf26wlauMVK/SvcXqEMXjiK0E3CON8KZqw/w6IbjVWiMtuejemgzB4be/ESFeLAxqjPGbqs2o
a5acMaQAG6VwQ5hCKd9thKOeJPDrf5n09tYm166z6XXQbqKbg2Fa4HfYNuj5vSoXHR3cFTVZHYPv
jArD4E/9gJCYgbqndlcxqKGH1QPTs5FbajpJo9Tu1p5Ylg8y6p1ToMuFvvmaHx3aPVNcgbABP41e
EnirxsjFFr/rNVe6VUcSalneJd0DpePwfzktUW53Am5VCSRFB8pX3bsLcVwbHC15OOkXWVCrrjqJ
4yuAr/BAsg4SgTs6GIT9AQVn+cIsIbV7ZMCutas1yQUsGfgfq7VGxnfl3ERGBxUywXBvQDy9scoj
Z2PoVhSf1I1+BFe524GfnPp8W/gt5s3AIii10GUi+kVc9aGLHjMjGhvT4gL/o3IQnSFIGNXff/wu
MfeFiQfwhb9o+rygF/9S4o4E28HXD+tuiMo3UfVa+cYJS4zaEiCDgrg/GJdvpSYdqZLS4k+yB0MW
8FGjctvazW2rIz+yhGWrvXiRB6Dd0sWKvLiHSr430sNJjgFZmXOCY93LBifRwNo/u97sSKnfc5C4
nePONiXVnvkhd5LvVSkKYPghnrfKjEFlaDwOn+vot6ytkYYh2V5NIeOpVPRx1x0ZYtr/9qADpn9M
YM0VDYdlerLIzgRQU/Zghj2zsj5nWUVigxZJYnGcVbbCo1ziCt5OzEhMWw+PqykEPLeBbSLaLYA8
DKIP4wRFpwGRdb8SGK1C/o0nAYlNUcbJW0ux/3075p63I6a9wbwBnV199Bl9JJw/j3/oc8xW+GKs
qeJRtkCykGWYilTIF0j8mucTHSZbCqZ3+OOD80N3RuAMgEj99evVB1BB2NilnT2p/2AqB1VfReGe
8LHo9qnHlEU1++rqYV7JxDVJdNE4CKf4A2fA5l5TVGNNvwKShVX2MaTMRUWaIfibmg+Pwj54QzUx
M5Yf/8dvjVchY4QJPbpyj0F3wU5pjUTG9W3eVnGiVXPNNDKNQuN4v0QoxRTHHZIx5k3WsCcIlFM3
ui7cjaZiKKuyirv9qWbLmOjHDgIViS4IuTlPwf5utUIGwqakrS2x1oyMndEh/nPyzia45gklaJ0J
vz58QfWITAhN86DyprVq41VU7nBkjoxSHSlh2D6QJstfqeT8EZyng6TLDkfNtqXr59wNpjZjxnkJ
rqQGQLYbVLhCdYbQTvCQuzySQfWRpA8vh4IO9HrrwBn4VDNdN+6O7brESuGbjbVGzod5wuD/Us7x
gBB6JCgQy//Y/vUOIkjFRZVkngib0FnjDoHW1nUWKSO1kmoSmlIOVVP/bpP770W78D7NEqPr5WpP
ttWNxU1TPSJX83/T39ekV/GfWwBRCZFmqKpaAQziXzecRlKQXxUu1PrG32mMcide4mzR7lp5WA9N
oHHTFVi2vFEojR35BI7LGeqNnfsVkV4WMOEKoAUx39VmMZ+9UzlPELoh12Ecs2IJux7NPqAmPVuP
JJx/3rNAzZIa9mAoE2j4Rz6Rd0VsRSdRaejWCG4sXSehg+ikUcSFNEy5FAx+u/WgP72XVHaPY7ur
b8xbAaD6RzDQYdsNnMT3cAPnYM8MkrSKMy2DwhliBbKMYVKyKWzvXbRjsWZhvRs8zzs0bsjBVlY4
bpPKLbhpzWKWFH6lSJLsQOhW7UGBz1CuDmyXQz/HvuXllbZ+PjwvYDthxtsRJ0HrpUHHQUK6jvxS
4qoVPSy/dhMznT+3viPuGtS0Aoclml1Bs0FuJLekqt0Yij71t7FMOMoqJfNpU9yX5md5ZBmzWA3N
rD8u4TVztAfOJt5j/BGq8P0/1QJYpOgENVKYKHUYDMI9O9FP5Zi/koVsPL8UVvAK44mp1dn+x5DD
LD9zDJMxn3G3gSYhHLcBbI4kLUmf3e318NUBpNjOm8ktE1EBe2sMtrH7WRnh6yZTWmPHX7d9siup
fWkyGgtZwEfZwOtWTK4nlnKkTq01i20dZvpwbjtSVai0M967othKz7SMxTnkJyW9NH5jR5K9wbr5
bv56EWaSZa4U8lGo3Vb5doFM6McU7fDgRNrsS0ME2d3g7WIwsTB+yVN+jjCzWw8YICjm9uX6VOw/
9T7DC+6bLTzGdvgHMuxYe50wwDgTjW/umOoMKWc81QpJ3ITYgySReTXhIJTji2WkCpZHTT59AgOx
5/75icdjRNenapzOnf9lYNR5ka9gGps+GWBFAoqmA6jojMTXTswN5P8/ID2B4//VDHisTIRWy+Kl
qTCYQqXfRzeqqPleDyCWIqtEXe4AvbGtEJR6iagFkMszU+ZyiYzbZF1KQROYbMjMW3JlHoXFAyKm
1XQvWtY9MaF851exZfQ2kU0W8f6j3pNzP8LSioen1/JNY1FW+42vAewACtqP/1WN62KXEJWKXpfa
9bSyzxs07y/XwSNt34MGkiV/60Y4e9vz7D4zm5rgydkQgBg62NdrHc1mSdoqxn/ZlSgI6v0yljOm
XUHEFXUAqYj3fUBjL9basFwfFvFaevS7+JAsAP5B+olqssB5FppmIkrYrwkJcLhQgsCuH1FByGX8
kCeYtN0mSav6tgyDe1whGkyw9NGVG9vDy76RqnsevHbhokUn5wNGLdVHgiYk7CjXddJX8nZB6Mu/
6Zb5Bt2l0MhaKx0WHAsI+6orQ6QCWgqfvSnhLK05eCRao5EbZAGDYv57kX35T1CQAHe8EH53WClJ
j1uRltVpWxxkAs+xpVq5TDv7/lfbbS8h316lGZXc5dnHDWPbmGwouxkWLV5ks7OYPtA/xADAngpg
wBK++MSBt5SdGBeoOWCr4EV9MgB6XMoseKtnvG8WDfgefa/zY3DLr9oaFiwi+fH72gKQhS+8tffd
GGP5UHmeh1YK6q4m3xqX2hgmqLgUsUDw+zkCNVegz9uyv9UdcAdEPIw8f48soqw2y5S2cJfuN0S8
7gVtorh67F1fiIY7SF/zvLTr2frZginINTxMt1PLLfUeb2qOOv/alOyengD/U3Z44A0Byfu9Rcp8
vPNGDe7Pnt3e0JSvhQ6QXY7D98WsKgdHP75JzJ6YMrqul81FIFrfSn/PePu/3S+8iLAmhSoHOvEY
vwyur184WtxAzTPO2+Vw20TsRrZH9QpYuLAirIDBIRVnzljkYILrm3rQ4qZPUHH5VCbigDuE0Afl
/iDtOilmqtRLxwHkrTTj7un2NnjsAWFpZ9Al4HrzyRktcEYzSbaLz++/uiLeh/D1jlpEu6kCp1cq
1tUS8LWwnwfGjGW0W5seHqEIorv1dmZKENVmpTFza7boMn6sy6abALwSFEaIjp3+SN8hAoc1zTjv
Pug8HAiWYU60MQf2uBVi+lCKOpozfl7TGU36khXzBXq5qAgh+/zkPc+1sGNbjwQgmk0Jj0iCMcqk
/7tA1xu8CkbvUYqV479RV2KQTGj/Eeht+7/M5HLEW+sTluAxkUW8EVlJQpWJ1ncH7FUWlSatqsBA
0MlxlUNNnOuKMTF+//qMscFn61zaVh7X03xQQ1xnaHbGUpkaPEZetuEI/gFTqez0fYIWPSV/4oPW
zUA+DROQ5SWtqrMEENVDskr/R+oZZMwsjxk9MSy43k90tuMIED4VAOeNHqrj2fRwLTkWDIVcRtma
w17V+J8vuF4tXSlg4aUklSmVObMJhWKIpLl/xQwpTHk7oksqJhRWPsZIAbGMZImPM0Hzei7XRaFk
z8W/k58dMSizceTiFH9UQzj3Tdd8WVGqOdA2faesz6dEMz/9yajbmEAxylWuyi0gA4lkaK+0DENr
sKBj9NoyrGuINIikPgucY2SmQ0Km71yYs/FVNtOBNQxDrf0s3/0OPAoWPFYT0HarItIZgc4MBMA+
1SDv8H4h+kJFbskjItLzMe6VMjj2Cp4HTRoRZJG0Jg+INCp47cHNKd53UuOsVHDiQR2+HgiMvqy0
qbPmQuyvFSrfDV370I702zGK63YBWm/Iqqgz2qRyJIwESArJaapQJJLjcTlw5aj3MDHXR5novyMs
hDCiiFT+9jAKrIRFDZ4zmL3K3xLItgDJYgCPAMLFe3m8XF3SNvlAbd8/P59NEAfiiYGDg5MxDqW7
qrP4KL1xcvhysQEdvSoYBrR3hjcEmgTOZWx7Q+CoF4PIsemB5cKrvjiCP3Bl+AhsOjNGrWNLzVB8
yU7nrR/MDXMs7QSLhxRJqdIPONTGip0AeK0u5g9bTP72ueBJtfTf5VAkZEEsi6AHI4wdzpMdikmH
RZO16qhEM8UNHwL5TsTvMPN9xHxiL56v537AnjLZ7T0ck1T6iOn92kvIs5gMxEAj5plQIT+H/PPO
KhJRl99W15fyZ8zWBmm2LQZ1/GwhEFEXYyNGch1yAKr3YK1Ki2KggxPzo3bC8ExlGO1Oin1IQD37
xx8xuMULBdeGwnGyu+leU6+PkHKmzUsMqZtqCcbIhVmFT+Nli+QD0Qn2VlhxlcjxSGqnf17HWkF3
RRLa2mzW2PawnhQ09k6yUnsl+PbhKsilrPujoF9ZpT/KAGrrOgr5y8boTfguN5x/RrsXrfxWY54a
4JHBdxm2guQYTCkFQGPkQ7NyT6oSWRm1rc2CTuul3s9+pnxbe6eEBFoLAwAtIL6wnUH2PZgeqPVW
ql6ZNDE9eOEsLhQ/yhJyzUTcT1bUxkj6NE8AvTPYbHUjagWd193meseZ1uYDf/XKg8NRt2urE2t4
0fVeKtVbG7AbquvWxI7h7yhFTLgy/bF7Wysq2f+ero77QGff9Glye1GwybyxKN49ylOx/GTpVcs4
25nlIccdYJxuAyc8tmtc+8yanLI9WYafr50EjGYYH/63WKf3gnWcxy7/me9x8KR/LGQoACbYXL88
zGr25LJ5d88I3TLc/b+ATRqa1iAGipFEtRJwwmacPCHPyYUSXpQsyIIeXsvKeTmJPxN73iksVkT0
LBwqCJq6XtoOmflDevLDXR1F9udB4R5xzI61ReMaOSEnEaYnY53ZwLiSK99G8kp2M+lrR0Ont1v9
U5at1jK1BoiixaLU3h3fmmQPuioa3hExoPjx9Z87sdq8aZ/G5NwNR4/bGFh+3DQA+VVl6LGKZLgw
XzB0czPn9Cld9hD3AFcL9jP2JTs47lTMq2OKe+RQnnSeAY+AyWsum6g10V8g46TpqqQsz0LPSz5Q
NKyaTP3kid/shfyg/ngoEowK4pGehxnHJZIkZBsZ714g1ZNi29/Zy9HjbvZSfXz9sHJG6N2Qpa/k
9A0RH6OzvnHShuFnt+pT/TJbvd7JGk/ixII82kK7JPrq7yFtiVFKK748l9rQB6qA5uOAnSxxrRjD
Pub4VYJiLkjANSN/fXLlTcMyubYfCEu1JFT9D4HYAcSN/grLCVJ7wDR+AtpquTEcPTBKpAjDFYij
RpWEDJHEYX41RH+/UMOW+b2IkZkDoLpPpckcSLs8Tvr5mRidE4WjZQH1O5AG/zr1Wia5mzOMpEkQ
Lm0Oxw3JBnkkrs+raK5xjebvlkWHelDK13lqbLceRUfdxR7OeKgKKz1w6km7VsmQyXNSnid7Jq9f
7sDHGzTO8SduhhWPsm3ayBPpZ9+KK7DWckTLlUxIVnhnjmu2j9SSb9Gi000rv/YVrfP7xcwmCMei
B6iOG7RuZk8t6Ogh5AY/faIDk9ypmTa+/Ht1sTfO7d5+ZB8FEfewzmCei+oMkuaJxpemQNCpysB8
cGJCcNaWiW8spRtn2tCZj4Y70sOrN8WXCO766nVPTny4d/yCSQf3gKlxj7orF5IvZNOZvkefmm0y
23U+5PJ50h7Yx4xVup4iVD7TE/Npeur5XevRAsrq/JkbwFIZ/DpOreojGn5V6+0PocGRoKeWvDz/
DISEl78iVQgKpY6ZruOHOhNMr4PbK+DtqYFxKwkFRAvXiEF5hhpOj3u+qI9BFO+yI7fog7n1Tdgo
MIfOTbDOar3cTsnt8a8bJPcY/W2noi6ymux6f2f4dLDxKHa32sbjXMY4EwWiSLvUXw7Rw96cSdRM
g/ELURaJDEEmDDhY/QiwOYErydEbtYoFUI2P+3dYRUrtAhyOzYNvu/kIxW6YeNYJhXw3/ZDMplbU
ElEkMdy7mLk+MDQDkxV5UBxL6iiFam9ZR6RRe6efAzt3Cq5qcevUGeEGps2FwxMsEOJfNST3IuPD
Duo7SgpPFE3VmYlEgAA2hLiHbv9WiY2AwA0NBD3SqLQgO6+UwyISjhOupdjnBBzSDPtz6Iv8AoJM
Xv/PjfadV4hI9VNClGuEm+7MPnlQ5GCk7DI4If4CrBbFNUO+3pPrwZG/398+QdtByGEjKM35DSkz
GHHK4sGKk3iUSPPMECq4k/meiq/0qEOUwLo+oNfsBx5ah8eVs8jfTpiswWnXZBHXCbzEFx2kJYLw
Qw53vNI93kQ3SCsxchM9gOV480BHNpGhf3nkc9g37D16yUD9fqp0a+IwYLlMs2/f68mBKqh42LJM
kOJQTDoQUoZyxERP6wGBkdhFpFZryJCgwryMzmhc3gEUnTynbmbLqntJFA8/1JHjdLwF/g5xDSXT
8UqWQOQ0FPKNAZBOWAsL8/fk3nenvo03BFkwn1cVGhDppxs3LwGWp5KSzoetq5s8ZehiOS3zNx/N
H+seEHvIb3PJjeBJCdynsuXsbEU11dMd8G6+ex8E9qRE5IZwlEibFErW6SXAodFcN2LaVaRmoVW/
GdB4DJkRD65Rry2Y19ClfDpcgwz8xQGHPVui40XTydgHzCisiumifHQoI+c//B8icppSGCafI/d/
x/qVKF6CzvzMp4nCBa7zaV8ZGO4zUF63akYcxkm/osDP6jhgh1m+3p7fTICyOwLo5lMiTgBSDcoA
d3UKckz6h5bHClyK6dhK9UHfIHBUz3x05558bW5C0hbvxP36zvOkrnsmbTXklt+y83A6Z/LLG7OJ
12P6WLVnPRiOJ4dSrc1eBAMULLI9ir3Fik7trTAXYjPm0YdmtrbUzy6KaYvC816RlWVqu9y8p1yV
k5vzXNXGFqAcuydYO4cYr9X2wPA87fPx5vWGwE6wGF0+vwKYUFJRaCk1+BQc9Y2oNCJeq6V5wuSZ
FoRFnxtAj+oat3cLX7ZrdeLyz7ZhKi4rdyG6ZoYlAmUaTpHp3x2fsCc2qo70lC35cUEmmrjPK/VP
zxth1CxayuB87fqyJRU5Ih+2gAHUzqbLIcFZ8oakZvOp+QzdbVdZ0FoeBRB+Y2JQHK5+LAzhuOfq
ZukoI/DL4EZobO1rk3H8ROWpxx197iPPXR+pqqXzKfjaAdgzrhAzNxArkfOisKGH0UUPJ9Ui7Pzp
eUBYfLSgxiZWchY6AhmdGonzRsm6A0b69UuHgJCSyg3RZSMFsoHY1fjtiOSK6ja15k0ydu/JagdP
jwDlJvGWWcrc/28jYJuznWp0OXcdV+tRRXMQZH7QqVMi9UrF04UFNTKsYh9qJhk8kuLHlx2KRm3D
NvWonN4Mwti7bQ82pUyIWtkdhj6cAgsnrqw2w1FSJYQApHbWc04HBZL+Dnjjzg4Hrbum+JvrPEFW
MlB9qtu01SmUFFJfkL17O1u7/lv/VPp+26xEhZl9RC0CEL2OSKDUQeNODRqR/t+UQ6waqTEzQkdE
ZgwS77i41S2n7vSjXuRov+4kHYRtHzyPDwgFiAA6MEPmvB7PQ0XEleqfTzgjIr9PFm0/vOBFBeU0
vgXH+OaWOeYCcXWv1TK4xLvugomrDS+vItowEKrMHxvDBMSTOWe7PsIQ5M/oRS/pmfkSDz5LLA4o
nxLxwchv0/XO5lukxo5C3lNW0vRl55kQqg18lDgEL5xy0Qx7EgSNpCAn8ufAHffQXY5RSebHxXgC
+oOd+/9NdVcIcqExZ3oTYfUBrJh3oEJszm+3eh+o5v+j9rje60CN5s+RDRgHdwySfWo7NI2Vapne
Ap1Hg39uvzLSvquwxDFvXJGKk3HhA2QWPktzbaNWO9CpIwNV+OceZ5TX9fEauJ/BTdIsBoS5fU5P
39BMiNyCnj3xytxmWr0YX5YGsVEttasxPs0OzOpcTgIqgGTh/LKGFh5CAyC3BCYZVsdSFJIsXVKA
7r6XTAcuTn8YzO986DiMJitvPjFPeut5NMQKlKDsF35/nD3ncT3Dxr8lZPoJRc02ZpZE3V1+c7s0
bFDf+9U3P8kOknkHGzz7ARdH6tJ/EJOWeal5rQ48IiV+PiNTl0YWvqt+epjyaj6FXArXDkrnmSiK
r0M1bYIkYAUQBrldpLARHRQYz/txoKGtB4z47i73UJ/Wr/N2p5GbGO9trjlzSrIiScUm8SDcLnT4
Vbc4NxY5VsWjU6lGbj2N0yyT08WzdIR5aL89FO+tYibjLSgzArq889Gbep5O79sQ0K2EbiTb9Qst
2kpNfUYsp8scqqNJoflazqxAwDuthLSqj4aQhmqi8zfrB7xuC403TfNsPxhUasImC0hZQISz8Yv0
Cn64+shQNRSwSHPz9cUgLK4ITt27NULxsjJPbQVv+hxgU8+S3G4wvJ5PXpddJC4Tdfj3Q/m99wF9
Ajk54+3ObqMxTa5BLpSiupOfFzM5TJNOZIM/hfLHwU5M+KAiYC78liM05Es3sC/ozmRrrnCEpsTM
QqZlCvz0fcNtUODRtkU9l/ALSC8fVPa1SLtLBuKG/qRv3Ur++f/rv0aZ0iRntNjN1CG8/ObPUy/L
YQWFXP9SIyypMcWq1yM6sIreSTwYj04XRWVQ9dmZJVx/snW2AZObsFnORJG9vhUhy78LD7QI8+St
oCBhOxdgVUu5EzWUqjbH5FjoJnhE+exPt2ndZ6z/YSePDgJdZB5JEkKNfATn13sj73EuW5SuMaQ9
r2iH4aeGrP5KRug8lzybX2W+7vP4409sFGUN24JOcYfEIrWoucM/+nOOOw1Km1yGskQLVdC9Wnqs
dVRkfKOIHbBblat/dkhWOMAHEhGPeuFmc54r2rnI3r5QZQl+lOoi+HEdyIuJyyNbRqTTj0oZCLbZ
b8qoHjkZUtIRZvp3WDIT79FG7vZh6Zvnx6T323A9Itc820NvwntZCB+xtiyfqfy8EdDWyql6ATLg
cVJkCarAEhu5+FcDyMcjDNG01KGbd9gg647gGYOfgxq34Fz582SwiTuCO38unTQKF+lA2hMM2VmH
r8HyLqSsz8BalEpO/Yn++xy+u+b1HZaSBP3xWTqA+H9TKejs8GzcVy8v5Lyl1tCnBluXVGVv6KZX
T1NJrxjS4PR8YUnapxORMVzDwUS3afNCl/K5tUdlASuCOba1Ijbg7neagYJIlkWDAJ8/Q8SQl4yM
hGHKMQKJzwstIlK6mkuI1XeaWVNvg1DmcIdSJYD+z0s5Gm9nKLvmcgkmPyB6mrYlQsZh/1r3IYS1
5InpMe0oa3e4egqdVa18Xjn2KuSmHDRWF7rHF0jakLmQuj1NWSRM/aFqcNd0d4xier1To2gpuTJ7
1yZkjXP3GjRZ35alk4aSLUC9+ZTckkLmoBqN+ddL9trsL3qO0NGDtZmMSy+TgRiePSsh8iY8I3fV
8808T8BaC5ztv7VjLEP2KLG1Fhy8BJsp9xyHZKgozGQmQA0N8zswZGB6IhJ4sKPobn7zF+HzIUhM
Hj4EVwMFbSWL+7fjEIW/XHtNeK6EBeoqWvgiFdV7zLWodylib0PSb4ASEV1ROqpp34rPf8z6HMx/
sRCViDu6vb/6W1nELE74fSE+Q8VznV+RD80PFFaJ+gfSXT/Ffh9Vvic5cOGIPOgGSRLaOYRWKHiL
3NNwJd/Ah+yvyxH+ZBjPqhyLGti7n7MyYL5Awb0JcKhN+xvBeb1PX4rwoKNdjg+oTEY5nAUe69r1
/iKIgWB7Udg7kk5yIgxNff6QyCbvEFcwOfUjkHIaa6liSjFxIQ5RHyG43PLs6zd93EJF2r80VQ3m
EKWEAmQaoVsfpvobE/GvDP0J78Yxi2h4bx5//lwJXELk4Ftkx3MzabpLhKHcsMHDu3QYvv4Bb9E6
YkblPZhmFn/PBYiVQIjwTsP4IBMRU6o7eM2l1jPsd3Cf3iIZd64bJfNYARHyI2SkC1Zprb+C8L0T
c4njlwoQI8d4VRRqm410tpY/IfZBvX3y2Y3tnSII8jJBKWtkx4EpzyrL0/8Xj7UuOqrH1insFkl7
tyWknWPXYDhiNbwDolSycLb4PslCpIsPysSHskohJjmMItOhWf9YKOOHZbNKtEGYpRsnFpjT67vj
ASGC87DGdBJXCy9LaOUyoO/519yQdXhKCKteTJNnzxb0nO3t75rGTqmgYwCV5zIPI+pVFtAQJR/Y
VBT4UpKwNJW9YQXzRpvonl6a/QZkpLy67h07YsHfL94Marzq+4Da+VQVOXQVloFYPCodz33a84tt
2+aidmfslnb2dHU4w62yMJ2TESHBcrsaTRfWcnREybnjdYEjERvIiyym9/tYEJSp4yN4IyU9vpBW
hXRWenS9jmdBCamR6nYzdRliMIXhpcQBWcC8e8CbkZr9qaaVaWFyESuQQ73+xnkm7wNql2icALWn
3V6hkb0+SyLp/Xe/63EEkYLo1eV5MEf7bd1QnD4kMVSyDsLP7q6hMPvmMKNZRz0Z1ktscSVJuwp1
9n7QBNCAWtzQRCkdnZ5TXLKxYxcA1nsWUcq821fpB+cR20VhCyyWt2ho7CRvX12xgmV+umfKvmpZ
EOjxxGRCrrs2IeD8zW2cmZXCcHeQcTIH9v7wx6ciHFZLG20nC1IZcwQKSefYX59IT2PK5xK/1Bgs
OhpLt1BjTQ+6g/5vkxeWH56zQwLAXvbw4BC03uIb8BhjtminL/4T/B+MK8pPbXxpAApTDCbejMIM
2bcCr0HudHgXl2ORQGKuGY4lSV2pJ9NZXX3vwftP6/XliLNPGazR1vTdLi/5Q1fnlua/0lrol/4u
W7jx/RvVL5d+IkkHZfn8NS7/UAxB0lLmoZ73ZF4XTcBmn0cqVJAObQrgtYSn90q++fsmDkJfX40d
BeVi9lkvIXH2HmAC2+t7tKoS0FAYnIBSoyC+6sKFFuCkBlhmnBNpYzAGrX+Aqj0fUC7QfK9xbJ9C
6H0cZqMt+S1kD6tkjs6jod5y97pEqtihwG4qnTCKXbs1Q2v6JqJ9v+8rufK0Ees4BYrLhCx1ebgA
VqpKJX9gogyTOFvpOGwXKIO+bHusMknpkzS1k/uglz/A4ptveacEZbuOWeooQRUFeVSfAf2zCpnU
y3TqbLZdZT1eTwuu9mCQNsMjQjXjoG+k9weYiwbjXAKzS6GA9AZ7AHrgVG4PBMR6D2L2RhLvcnVN
1eRuDOf961bO+NRlhspJbM45oNgacAiLxEplKwSZV0UKP59pp0FyzibBu/WBc3dWtFe1pUL2sT57
aZpmRrNdkeO0LNr/pxIbnJxqjNggvB7HFtd0T1osS98jWm9awtgzr4+JoZGPM6KHzhZ+7dMG+TtQ
q/9x4x/RhJlLPPIfO2Si6t1aeY0cwk3/8v3V+NvzbQwvMnKn6Yk1K55PF9x5HagZimu7ykzvPBD2
KY8s1/1kHS0pt+5jucMhA45n/e/i+ItwJycthVcSPMcjXxE6fgNm87B+AnmfH0flXoIgGdFjkZ07
yME8X/d7rGXQsXY21vHWSEOxQITh9xZZnFe28LZuKs/V9JmDbJsXuDV2ixVqOLKLF88aANJ1+3Bn
ok1AGjo7MvAnnnXnmc5XMKgaWoUZndl/2ORjJy6j3OlWnSyuv6PAFX2S1Az0lynj/mvfnnk3qcLI
09y2lg92LOzaOKz3nh6eW1SMUGpoPa1fY6gf1XYIo2RBJshRCG2z/SOUo5PSpp1KYY2nUTpjxapE
FEmP1XxWjhyD4LpesG5hGLNq+Dpv9dzVWviRYrlmWesBZASTsKxa2VPlDlaCISqp9ZAKDgK4s2ET
N1sjD7Lx7kbNb9dtBmCli/rMhzU9dRG2xVdcSa46ur6KUwKRSryHWAI92Oa+iFsb/OlZL1FKjfdv
D/0EUkgIjGKOAykLt/H3nzOf3gfG9NH0oWHEEPyexZswQ1dyu/Cd87KxG3e6ktVV0klFc2fgMaWv
k9EJSNLv/TnNF09KQjEt/N+tk5o5rs5Xea5zD3VGqgZzyhbk4W+dKmmbvzCR/z3tKQQbUTCuyXcG
iBqpBj2Z+yDgklxUJbcdQqec9g/WlS1hcXgukAbodF2gvzgNF0Cf1lbUOhXUG4W3ID082A0NndpF
5fazZ9yVloVr460+laRhJ37NIkcPhuU3+4lXAWWWy4i1a5hDnseSduOkvqAu/exprEdTlDh7jkoR
Ahp2rN0UMa2O5dRJy2W2VXxwVKXntx/8IDgIeNMe5M3jai76nOXTcpZP4ai9lqM4Ds/3dU/L3AoU
DmIJ3edMcJzCR9WWE1J12ApcfCWFXweDVcQeuGMIIJbXnfWj8WH2inftXTVCSLMn+UAwwlbKpLfG
WzotkgP1uIw4O42vfgJkNJgilw48G3grg6LXSnVLnM83+nM8vkMgKX3LbeVBSFEV5LyZXp7p8HJS
aXli7WZBmETSOgGryqHCovv46ucqbehsvp9FgSR/2lHhqS8Y9zIG2TQdL+KFOKQIrLxRgshgdg3E
FF+qfz3Yy0qvjlma8QokV01iZVTuIWa7DhiQxIL7VLUpwNqcJS+zAaIWleJmAAGSA+Gp11qa+q2M
MycuoSk+XJ93ZQUzCSfeKhSnfMf0UQkAG2uvMOwSTFs5HH1rpM7SB8hFX0uz3TssnAyjUgoShccQ
4HHSv05bTInr+xPVSQFqsVSfbaQqoI+xjyjwEYbxLZ+R+mWbb8ubSlztCIxM1YR4f0Qs8ud2GpEY
B6TxK42oA7gl6RV1R9+/OJ/L10TdYFXBzrrF9NE4u5SCen3XNys/RjAW70Rx9oG/feueXmcO8+MK
KEskcy4qP0pam3T1PPFgLjlYy1tuGEXct+bpdZ8tO4zKDp4R/NQGJR6OEk2fjF+TWonjhB1yMDXS
efwr/BorFWmpynutEx5y49sJiB0rldPzAgJQGAw4zCxnqbfUGTggR0Sv5KMBScwR0rIb6BZKGxX9
ftWZodsgOGc8YKHLcekbQAqtkceL7l4EXNIPdXYeCH9jJVua8AEfwfgewjGV/POry6Bo/KjptKRn
2OlSbSjhbtByZd15VcFZm4iuAEoCr772ryM2tjHvGk6HQtptJ6ybToaGn3Ukhq223W4mxS4uKJE3
XfTtqyyLbtBKnqPpnElF6HBtouaWreqqXJV+Pc1pV5614rXrYWsOuzPusNiI5yD4tomh5Ju6uhL1
n42LswYGBxATJMCcGBVrH60E3JnR/1hCu4F44lLFhS9kPR6N79dTqe3xnuMgpIzIzOY+mg2n1nOh
onkLWafyhbtJmQAaNMEnRgLSmb7sMg2wbW3YzvGW3Id9cwIPyJ1hvFwENQq4u8s2lpqSSVygguyS
UTpQenugvcAMNdi2w+PzaoHtuSOWMdpxRFVwJSfZbVEzfr8WHLJnIbWTZYz5cmUl3udlZ2aViPOt
f2Rx70NZG+YprNnecvx74H5lzBPQ0FJMuDuvOlXlMOI/WGH33RCkuxHsXljTbRylca+DLkvItfCv
3D21jM47ZYUDXEsWbBhc6w9VUt09nPrYIC3guNcd9tz8cfC9YQw57WzOG5yqP8/7XoFDIqSC5mxq
a/w+mPXAkIw+uN6pVl53fBTC01hHp8wq+o15JSBw2zDp4Aa1WKukglFB8EegNFGA5YuxL8NtRpC0
RJMBpTbE3FhKfcb4hmJWBswTfhdyZK05j1WJQd/IWtzJzmWGjoaR3fjzNbSfZV1QevZfTx65eNNf
1DoeCATGquv6GhKnxIxCrqmQvl4NkAt60soA7vkPv4w+X3X11QQElXtBkybNLgLFS4dK/eE0P7dF
EbX0EkEN7YWFsuspc0Arl444vopxpETMhCRiRPMqkGtrSsxraqvNCe/np0Lt9GnZ8HxR/HRPJwqr
kZkUgV7NxmdDjmZoQ+bTGrDPpzyQ6pn77y1vmtSQz9BgvzrQWe3zXTn3+G55oyqKFOjYgqLMrSx9
ssodGd7wRb3eSZ1qAmbMoIgR0Ch8gCcqzbTFpfg2oo4PQn3PG70xWIhSkX/0OXeqJSgIEoQsJ32x
JrRKN4EcrZ5ReGcATbnXm1BdrNoNquNiJOf2QVeGFO+hJHoG/CPpiDbfghnk0in6hm5qpottVdF4
rx8wSl0BXGcagR7OiH6+dkiKrNjyk8z5gd4T7y6lp9PIWzZTcN/4MjJGHvYapwAp/i5ze4Qnb7nm
pJo08JpkGx3EDKoLGMnodLHzOIW4o9wREvqhas/PQh3jv8FkMjuHx/7z2DLM2WyIrnRrDuTx62ls
dQEQIyYks9QLR3Mt+n0J+MjxO73WPI8BbG9GkgewCjK7kjjQYvgbr8lx2OM+aSrjfOxkq8i0lapj
JFmYmaQ8MlGGVlsE6VcujYXrZIt4qA7ImoNz1i8egTd04gs6BKbO++gh9aCi7ByqTvr9BXy6Hwts
PoB7mmQAOTodTpQTItsLVwNx4FXMMPbeDiU7VDCRwmAp55x+Ibsmgh0vaGDGC/flbz7vNNjz7knv
DRemXlIXVT5DCMj7vz7BlwhF1fSp/jyPVpG93XxFymIPLG2pemi1LJlVC6TXjI0D3EFVJkpPg/cM
sutiuIaKNLfdO0SvCteNKDdr34akudC4Bjb8uAtJNcJ6fF3jxOiRviyhBRlwH8viSzDMmN4AMn5d
ENlYmJ4pOOdIK7iH65iHJnxpw8SQ512f2x3XHHThk4R+pc9+oUKvB9gyUCEAsVt0T3X4MvtumoGC
1VZ698Fb5dJQ/58u8xwFcj9XhxkaFPVWuevuw41oupZ4kIAdy4DEvb0ty7sptIr5iLop/KhiSkpu
arVot+SxlT0XhI8W5rybWN9Mh2//8qhqIeVy4chIn6h+DZhs9Kd/syOWTIla+MhXoovtNVKvDlrI
Qq2s0IQh/RbL3xrIO4XOhmkUp9xuJZH9+cEtnFC+o0n91wCjlH1NYdCBOqHyfv6htsRHoD5xQfe1
OyQGqmZtdtVV0hPrBfqPF/q6Sb5EA+h8peuiEFY3a++Ik1UfO8v/q/sK6d7YgnR8IWNP7hyewhdC
WyC0ECIjy9yMZQslBQ+YgFqAUN30HAbNf2Db/RypMMffyinPrlbT4dkjNRVIU+d102E8GQ9rYein
qUmOUzA3dipSIzjX17cwvExyn2FyLbeMuTxFQIbS2jyIhlIO6ksqqaX0VF4B6IzWldTm7PKaJ3tF
dYIy3a9UbxEIBki3uQJstgvZY9cWNcZWKOGt+zV1mD1pjROVKPf7MooNmmxLDjF2b225Pkq0WjBS
Of52ahK2o64nK7hb4jDF0/LOZJ1dMHGa++ltcOjIxsZhFqDSto0voOp/VKbHqfb/EL5FuOtEHEEq
6CJDCxbWmAEPbs2MYx8GaDBCvAwSr2BNv8u7te2MTHexCTEjl5KWkQiNOrV7mG0f8ZhPjGH65pc5
w8GyIQLrky33Mq5pkfrNmsMjW0tyXFfcvUZm2A9fPzhVCIxO8Kf6tK85D5LRT7KRSWmJn8uxORa9
KGyPYXkftRiQwLHhab5GaZQf190yAqhD8QA5IPHeSIa6za2U4rDp3iDeAlgcR75/UpQieBYYpZKY
+cZIaucFCWOwAwAXlVReYAM75qbexM53k8T2uBQ3//L2j2qvbw8zRuSZMTirNtUCWRvh1Caq1T83
aeo1bVdSjEWivjRG6EPFaxckFupg8HXX6/vlriR/VeoqCSGEy9sAhQw89ZnrX04NQYxDmTwjLDeD
4Zd6pRHU5MMLNDae3C+8yU44TLTjYbHFybYIRE+fGalHwbc5MQURH5mpKUM2xkWu4ufHFCLFWN9x
Nh4siM/G2c9xPi0v0nDe96j6zgr4SIZSlRxjRWUBlYBi/nzegscL/cPD0BpjFIEi/rQw8ZfJAfXt
Od7SOgpB47jItAqpE8HC6Sur7RW0dLAkvmO0Ktbv1N/giP5E4E4Lv4mzeu1oEIuW3KkG++oagASD
16oXyn0YlkX9t/1yh0qlofyuuh2CuYTs5Ml0oJPzav9RuC+R8QkE9SgdIr8QDQdwF9qg2cObOyOW
vs3SErjiFQPFTMjRdoU3DxedxyCTIkk4+gQSFnEapzBSRhma8uvR/coZdW29ycCnk2+gPRIQdQxU
FrhEsr17RAypG8FQbtVfqP73/hBbCpS5gPOWuTLmLc1xfSsy2VR4yxhIpHuU7aAUv6y8e89p85sI
1or0zhBr3IuTl7Tp6zKyGusL4U+SrJIsUOF/rPqEWfjlwvfy5giDTwbX6kwvyrXPcUFQforFENf2
KoeCzmq4U28336WTgIqJUJuwG27on2h0vyeqBL4MHzQBvrpObAB8j6WDwXUHeUsjCEFJOkydeEtu
jk4XN2sp1PhwDR324EJGDCx9vUyImhTL3239SgaK5Nvl5+6nJ3Xq+DZuz5QyoyV/uh4TSvNIckQM
42QxaehEEmN059GqW/fk6MbkiL0d1jws4qUuheGmsE2y3ydJoU8EM6fx5nJlA+oOoDNms8GpqamK
HgdjH3JeUNR2Nrp//YvF7P9JI8KJZglehdWRgPKJDfVBJK2a9wRduvmPeTmCooYZoaae+S9Y05s2
/wqev/8Q5BH88rRpdzHie9Assz2ZB4nA/ZiGDkSyOsszxVfwOsRKCtEy986NLQ5SdUWUhXntGblI
bqizYsDtmsJ0oKy0RKCGQIvGu/jdbH+x2xEPbfRkX2b7bSKB0wwsQ+tAR0N9MYePaeOG1p2tKbns
E7uZcqvNqnCQ7+ZuNLgIjbOV4qt2T4XsEL63Ni4TfkLfy62Mu92jFkLo65isii/84YnOYqlUNC1s
01sH8nT5D9cXz4v5Nd65aWNcONDpRrl9tTYVsOAJ541BfXWIIJKg8pXfg/1wCG94g0WRrm4T3rMx
avILsKH642x1q1tiTiT3J1GtzBIzetvsVPe9CO/UeZ9abSyGjGRtasFJMU1JkR2fs9CgAXReqz0g
93fvGtMOJVcz0qaNJ9llrr8284JlNKdo3fstsy2PjAWvSPhfNbqD+mrDt6MTNL4E4mOJj9TfcktA
NB66QCE0UTEEWMYF7XnwSmkmijRoXoDbXL6M8HCt12j3F2v/5ta7L39aDGMuzOReawEsuEBeBsEl
rIR3wkR15iNgOozX6CrtizXzpCkofh8ueiE40eRDs/xu7HdYhgZMaLCxlxF/mLGrURvEqVazLkpw
faQWvC3r6PZYNPxksprH6GV0a0XsURAZVHIiQ50IxO3gsJnpm2T7yh5OgbyuOsLSzhwrbYnItEuB
85aZ7bLS8VE6Y1eda9b71sJc6iWyZT1+LK/IUnRpFos53xXS44vNLXUBD19rsNTKwOOufPVm+jSy
stsnP33JpoeocCxx1y7ikmR7kNffjQM7pJIOQrSq4bN32ylvSUx38yXGgLwImx+CJZQf4lenXSrN
MMP2gCnjtd7hDe2P1vCjgBrxeK2ZbbKrKZS6e6znUcpwDzkY4jJhVsySOUb5Y2pQN3/GV+blswuf
e3BXpB3NQ82ZeMyIjO3VsG/+CHudmszyeBnyOaoIlGAoTspZ6pp/QcvD4QG0YcDfrsqkGw9VpUge
R61Vz7FRg3FaWcTrZ5CzRvGukI6K4k2jYvAkfZBt387BUwXYpqV5YWEHXcGUQq0sG7W2TWwJfOi2
2waD/yPNIBo0vbY0DXFys8XEPvP1JE7utBE0JLag4MG59qmhG9eMAHQzvRUOpm9C/oa5Tv4I7Uv0
KCVrgo+JVa1Kh2yyeq/NadEvtviSJTs9TW9Z2PsUdZr4Mhbopfn063WKlcHRnPXnlUsV6wQGgAIN
GGq/vgNAAvMtrnCc0Ic//gzWnbnT0x66O7i3ZIxO30HoRT4CQBPwQ4mLk5Xj4ZWP0z5EGKFp2BI1
onGy5NTRpkv9QW/fFG8lQYTNIWRqPODZWrF93IWBUM34pwrjnPQDYTTvM7I9u1uZb0Uet1QMczWb
7f2z5KomwEOnA/SPDB4eQAuZBG1Dw5P1NxWj6fqUATRlLHio0Rv0AkmR419wRfpfQD7D3llUyYE6
Jg3GxKJ1MJI4hhe5HaHVAddmki+pAbQEfZscFzQVIPjeqpQ/+6SGLG2ADQenRsUaK9IvLzOSGep6
zYR3XbQVyzxnZzDee7HIhUUUp2ekiIrw11ZDtAj/28zVmlJ+icdOLb2a2OZPFe6e2hsxXSkMlcXH
ZDtuZtH1L9Iuy8HWNVPbuZE2i9IsP0W2tSvlh/hD+dQkP8KzLd7TmfPXcPUcSx52HpxLCicYljxj
H7JX/qJj8+3iMrj4QrT+neNA0YgmivgnNeEptRuf6ZuRz3lX59QbfIQw0Xy93Bca2oCDrikb3+HS
c/1PlH+Qjo6Ut6cxc6+Tpu3SDDdVZimE2HLVWBRWhC1h0E0ydA4J9/X4Sbqpck/PvWn70vHmWIsD
KdZiVNqekfS7v4jkPdTVqeZf7p8VU5nlqTheaEKqYmXwwWOv4GEtjvM2rCpKcgBOj1XwaCgqFZ9a
g7le5Ii5bWB0eQYis7QRBswPP1VDueng3gP96k9ltVLIRB7o1WEi0OwovSwodU79ok8zpb/fws5l
x2X0qqxBMxZ+TBZ4mx0r7Opb7UXBswU++GUegnJgjDLOFLj0G8MZJYaS2HCFJ4ZwZYAY/ph1xe4y
a9GeWLsHJ6Qvt69nH1erVRWCelLGxk3Ar6OFOyoXVqoCT81d974Cxy9Oe+7JiNarkTRVG2QVpiuA
C6IsY0mfL3kDIzOrwqeMag5p2qyofjT5zfYXX3NwrVgp8/zEK/wUEOKxEU0w3BHxOswatpJ7xW4/
uBtygg7jt02gOlr+NFL5DSVDVrin2g60XfSXybKiBUm/d/UMQeD4ArRLOPf7bicgb6ND9k6g82xH
tD5HnsiiW4qnc0i6x5sABvRHjEgdiz78hXnmroK9NCVeweujW+KLlkgvQ0JMv0uAlEysgEXKQy/2
mrEgNWa5qF28+53HzmFD9zuEFI3lzH++JyoZL3NM+fYe5lxp1k1JgfeGGMUDyCPzfDxg3fZKD8Mm
GYLtJfDEyYWis+lbfhigNEydYBSXJPhomCTt7kRcBknjOZPvr3rloHGwZRJsK6i1qL1N+oIsVq4j
6LfGOaxkZV4tzgHUPTGuJJqDX2JAray5ER7Rxwxxyr6jXsUQiJOhqXE1UCqWkpavygb1gr/z7+1B
xjHGqv1ZWsJTozJUzmOh7OTvRrKDeO/cUgCmf9CWNTMYrRE41sOOEqglOO3pW7rvy7EqABy9c5zN
QvdnnpNDWT1OywPNBB5fbnEBx9oOCT2gnkQwNfxCOQ7KH259HO+UGJ4LBkb+mClwmDWzT8mO7k7L
ufJqvwk4OeMFwBzQs0u+z8wf264LxysmSQHtLY4TijCElY7N2WJ0ReGstItqqHDsUHVHZwFWwr0/
Tt0304W0ZNjEBFjMGFENVDpZHYoDhPy9b6WF0UpnKFEAB6sbAn5hD+vnnQqhFEf/qltrpNJo8Nob
m6BBQ0mjHAMaGJiuA3KUYbEmKqzGeeQ8LJudGkwTKFwLC1DebcSfRoNqE+d5CAyEe8JQGrKWlSeV
zD3Pzc1814NRlN7HmqG9I++/3Nn+no9Qlau1uKGOe7nnyvyQ5TAk4b1HcGcQCzEPJttwOv5MslwO
+w1s59GoqUFKrNabX94JuQEhejiBcJ621egMcLyXIKo+K+1Zvl/iyKafSR3Yujy0ykQLm3RlZ9yN
5GLo3xCjlbFtBNetuO8Nhm5gns5v8C3KTfvN04H94aJs63X3mWt5zcqZppcAfbFgo+4XlWJKz3CH
MhVS9dsms9dybl9gbcTvFTBycMef4XWnpRwh2/HKi4gxnng3AP2J8xQF7T09SRRCnrToodEaYNZh
05rwvJDStY7h8jRKQ6uFJkfR5CNJc+IlgZpOS1evNhqOmQLRaZJd3gW4j1P0JClRAGwdE0hZXy94
2bbO69LeO2wEjIOo1841ijG3/7mbNPOIbzpO+WFJtRfM9VmlWWmQGK0gzMuPhTmnvy++XflMZSBq
O5ppemEnP50LL2Cs39GajfbvQ2oBxfmIN/Bw5gaeSZa2C9vGTPTLKhtGJDnoNWCBKvdn1Xd7gRUx
aIngfNi4CB9F+OG/Y1LgeUZ4WKGfPAo4Ld0fy2WsK/zqX2W5+/1QnPJsRLmpgJtmiYUnZOdV5HPy
YOOCpsskaH9aM794JT2WTc4KM/QG9boouzVyUlT+lYPIMH9H1qTRt4VwyRUP5WzKuDSMc1hRzD0h
KT7izHPKUXSxmQyNOeGDnErSOVsVVbu9znfe6XNytmY0vaykwn8pYd0tf5O8vBDa6fvj0vOmaaOQ
MJ65AXqJgo0Oja5q3FqVY5KhQG//S9jskeIRKkyfgIn1WFWLPRHqv8DNATzHWS0WThGLz4+G0xq7
e6Sb4bI61x7mc86PCKFcY9ME8O3GLDtgyHpvfMmybEGxDS3ye17v8De4H1QJL+BrRtyJJqwZqTjd
p/lY/knSTrv7Kimn7r8LG99PrjpBm/UGACOI54ecdSQeRtd+2nL9f8LeAutuWgy5p83uHy58GH0x
WCmqtDvMzMep2AAk8PKNWcPTFJKgbW9n2CqfptzcDkFmYtQyFLhdGofjaPSMnJq+EQNg0K0W182o
Pet1iHYUa5j1XAorJa4aKca+DtLDR9n4MnSIZ5zvvFlHm2EIh+TrbM4lEJfx7zuZi96TJ3R8K0RM
3/ruEG12uehvmL8JyYlY7T8uyf/eVoZ6VHJCKJvwTVdqPupotFlOGcuw9WZXZgKpPtXj0G/2583P
KHag3GJ6bjbhkJOlalVlzsltVe/lwAPxA/cZWQbIBzFH9t3YJghaQoGupUtsmjDv4owaMoeRq5Ti
KCpgp567XmBMctcw8M/PoWlPi6nXLWatTfCZGbbHSOhI2odDyFGeQTOwwddltxvjEBztKEttUdWT
sMnqTN5cz4kIu0uVIXfoWXc5H5CBEa+bxBzfi1JzvbuEolsb07RLMrNk2xAWVbHzfnjDyrxtc2ua
rD00ZDbX2dAdKwpVg2r7s30lF6VwVxcerK8Bxx+QjvV2usnjR4FDMDiUFSsteAFTqfhXE/EPwtaF
cjoxfrwR1rPsASKYmLfWi6CDoyKJhOWnqUCbk5XNCwI2nU/cWB/79whHY7/x6TNEedIDDuKFyE/b
to+KLhV78kkbjD6DieCirJPavh1YLbfJayFK2QgNyFVliKZexlOgKcgvPwU5wTLWb+fBAO6jN2LH
YWtQxCvgu4elBVOYOhSt4NvhoOo9d+dibI49qaXiZSgRZvGdm3j85c0wqLY4+UsOGzO0ZjeYRYXe
0CmGrPhNjAT8YP7f1JFCNzxI+VRhPgXIAF4acbGSOjVOHFtT4l0yXWye31QQskLxClr4oix3Haa2
17zgky0ZsfaiFHURom0m1VfACefL8uLHPkG9SHd+BHcdXCrbyMcMk0n6jr30B80zRQ1Un9Ujvhc4
CvAmRU5n6MNSrbUs7ie3IXCVHjSls9ck0ojpDKWRNyeRf/pPh5uyuM6YvntYoiUEMib1tg7NEi3/
hucnMMTMGwsAEOAEAGNwh/6hgKCKk3DpF5D/TX7szNDL0JIorFCtIdX6rGvL9wNibxCWtTwlN/RJ
ey+ljko6FCXL+sc7ac1hDl5VTf3BYBYg1I0kRZsQEeTLXrHYVc50bODDsFrz4kxKC7UXOIuAJtPB
MOieXhN5oFbjUyNwAC5B8DjNPbtQfD0NhC/3sdBE4F20OIC1Ra/mYhK2c3ZATPStUZSMpSVVo+Cr
80S4jSJWHCWV7TfaItuvRdc4KX5jCkpyGetjL9aRe4f45JF+h/fYDp6MDaUhhtQRIcYlngRFtkl9
E1FPtWrPYbjwQqQ/j4aqTn6htdzznU5XVUcXMydHoXKnOlhbBWrFwyuhHFlHlajdVoxdS1HzKOWy
RgY60AM2rIP8a67Xwyrk5jaWb29xfVpf/zondw8C6rfsMm9uEtFI+zmfqol3nbyRTL/2ThcB4hIg
g5B33E/6hdbHSOThiUAkVYmcld2Bbb6L+8eCFGSWwNlK55CVLxFRIEZfOSaOfru0U3C5d3l+33Ws
G5tVrnNMNJAQsq/JL4WurywFUf5Vu4X4ZGcKvyEERg5JIzn/XCKCvd9mMwb+pfX79p+TnjGjfi4B
lDFRGMIKRYyO3y/6305lZ7nMFzwG/ihGHVz0ltfaOgHsnFsDpKWYXsuG5V0nz243f76blU0kuPz3
ECKW+kfdntMLvIqzEmGajsaoNKv0K2Q/00RrfPsHpfAYPWx9HjryUHWzaLrYKp8cnL8of2vuDkTv
fuD7pkIjpniBIwIjxr6QOsgX90hjb4r7oasHnNYFPCDmjRsfBZboVLeYXd4p7ZwJt2vqGyIEagNy
FMi66sbWR22rluCYuBXXYAOC7JtAkqE0rBSy4GcH6RTp9CCBlcUP1WJ1zQPNvzRsBiM81euj96Pf
hIY9yfuLR+iy2pa4CGTcp6k45WAQLEufwFL+gxZ8xaxxFqctF2136RMTneihTb+LdsSMWMgxfJUo
McqPggZGMo1ikqQqYCaCm41Fi4LSwcdvrX54erp0PPFfxWaQEG615iEw2NAnUm7WH/gd7mjIlR3b
KPDMLWtzNcbwsEpGZmkXS7tMTWU65SK6By+mays0qtVHDki/y0XDz2HpoSgGtbgGnHrnqvqz7jf5
w1k1zZVDsEbvL08wYUfyezZUveDCls2PFUDCVh30LpwQdMrm0mKnm6rXRWEeDSi1ztep09otyis3
Q2eodkc/KjWYAqV1cDVC5YR5oOAhW8Rt+Ho7fso76fqEtucUUAqY5C89kwfF44+ibPHoCunkmrn1
ZHumbEHf8806BYBJDC9bK7UQ7HT3W6d+VtYRUDYQTlyFkAyjYTW/uRkT9a4wEFp9BALaIAQ4VMgQ
3PnFmZsQFxQlTQkKGdXgL4zsaYbr73IIfVCi80bpKDzpvj3zUn5UA1fO5iMLSXrkhK6J1QqKQJ1y
YFF/4HrtH+QfMdoGsUvhfYmCMuwIQAVMiK5O9RxCuDIzbfoFgrcn6RGqcDjHMJQ/+qucdB7uYvrQ
+n90X1LuLPXAa0WfzHZEYIEVSlC4mmyj3K43YydKpjEFqzjAWiM1YVvVeu80wlKGnMzDTF65DF4c
sxTupBuC8hNv57GommM45YIACUfgp27qbLBaHZ1hfmH5XtT4TFfPYMIe3Nq7ifyp2PNmDNZH80CR
f+nNtibdY3Jv+jefmY9QpuaNHn+ZKA50guiteKqcPsai2/bxzEIXVZNNCdIOtLhJEPoFX7cwHUJc
q8HbWuiC/gGu9yDd1cyT2IXvVsW/lXYt0qYHwpJ6Li3+jknbe/tGxk1kcVWO6yvTgGcG6mMZk4Wk
IYQPPn5mCQi0h8OFFpTd24OaTISuEPqTRFotbLrmB6NH1AuFs8RXbISogaF+8Lug/uVbPWfWlman
nggE7IOaFnxCfysJp4atmTCf5ianjtezsCVsVVsQMVuQiQmyEbQe/1Wm9ZKHH8QwDY36Rezmrqbk
YPkJmYA23s1AEZPwjSXAyJxrxPSpOvvf3Eg0z2hIt+sxSBvwnRz1JzO7SLvJ6UJrBWfPi9qRvtB/
OxGlwwnEmDlzXsz5yE9jYp8KZYXNscg7QReGlscBqZshp3Gy327KhXCoPRx/zIdZgZiiIZ/bwYPa
+mdhoeFgowdMVp60VHYL6ZrTj/j8U0mEzI1Eb+rRkno2PeH5Rc/SRJuS3/ovD4DeMqAIVQXaR7vI
Ob+j2e3fEayQ83eEqhAiCQjm5gxEqvyMgfra/O19f+KlEtJqaW13XJtLojt/Bto9ABWFB+kICIg5
XCFK3mVWAGR2mvA7PKLWS/HZPkK9SwXkPs/zl5uLpgbAq0NQMiDZVHP/NIbKrcp8DZ4qT5XBZdzq
//2nNz9lSeDmhbo8g7tonHnbGLfyHXdhifQrNoMPqwHgUar34CGt1Ooz+sXUCaj2OUWnGz7gIwO0
8v13tYgZ5oEUyiNnnw2yFifGXpWWpxiIVxNtwtrl3P4mRwSXU0+80ndi8fOiRTzwKRo/WHsvCHtQ
08ATgWkpu1TysRDOJlxq1LtTEfmCDK+NoIpZ9RIng+JlzqnWb6Dz4NIe/DfxcVuCUKZ0EXc0rOLg
icwUoYPJclnzOedftGCW6hug9LmoiyIvUIuZDsYN758ESFbthCdG5rFkC2P5EVgXxtuIMtAVxedQ
r6Ox3gT3vbBY8z5Xo1RUUS4IIY9SD2RbAWNuLZVYfmhxEDlnYv/r6o+n0NJc/blWUAp3F5nNVd7i
TLLUM7sz29K7QX91HLZkJEjsVUm0Excg2vmLeRkFYOfkAEDqa0EA8sXquZLTG9qSPudYYXC0S2aS
SuY5exT9XiSgj9krLOtv6CuqLH5vgblDPe7F+rYp+i7fXOJTctvP6QCFsPqy7GlznloMxfi4snFT
OcVr4h74NIEblAFKmSVH6UjbNnu36B34lQdSOdRoNfNUbCPsvG4jili4mRapGV34cQF/n81b3T6p
CLtS/NlT7VpUMVvgItPi1TXCijX6JN1HMjy7sTEJ5J++MWtBKXpeHIDiFA97c8ZPCOsoP9xH9JAy
9P/pPjfPRMD/+PNjO09C1NcQvJm52AGQXlbPaO76g1DqiPiAB8soH29abDRcS0HR/fRWULwrJwui
/it4Gee/8iSEgksBUmRVFAmXb8ryjtdICmcUFzw+kMp1PDGat4xuArjpaASlQGbyIeCtpfQcSvC8
CRxh72qmHDvNV1BOBErokbzUGqO1N0ItEY/3WZaVNjiBE86btPXBiCpMzZcqj/qVYrxfR32NbyU7
fPkTHIS0seTxIPet5kLCCQK7vYjzFVk2D12H6TKlCAzn4bnsJMadZNKc+T31Wth6NgQxNX3n+Gqt
5mFb8LBaA2EEA2bcleXXQLLxn54U5uaPeJqmuPvK9QuHjXxWnV+D3E5ZOE9IFRrQw9ltZXfQci5L
K6K5lV67XPyWBd0hAw8QAxYs3KZ/pgh1gNi3cxF6X0VLegJHGp9RZ2biV1qioGDdgGUgK/owY1Qv
tV/kQFudU1PVPoElLmNzBR3Z8WHFu79HD2yITH0dFgZTw9GUh9hM0JJwHx76I5KE+eFASVcBzeTp
O3ACPk7EE4KmjYiq9jYYnPqYKjZoeE0TwMjVaDE06UBtk7ZjRzow2loH6CV5Q3SiNRbN5F7aii33
QHHE+F2qatDoUCcN7KqcqA1v7ZBGkt1LyTAJlEa5e1ZZuPd5b1Um6gzBV0ADGdlbXV6hDXVm4/4J
khhq2B2pcPWCCbBUglsp4E2UFAdGgFTGethfmgqzKvS/TPgmXYaQ9BWycoRf34ygMOJ8gIFKuhmF
U4lMAWVM6QbdyI55Mv2t1ZY7EBaaCT2U7jHuK9n293mw9cix4vwnhuCtYtrTXRXTNaWI7F5EUMrO
kcsoMQqo9Lij1M/Hu405hyXsmuOLyaesheurQ4EkxQWQJlARvTlLLAPNZNHdw2c0M3dFOUk7FuxP
LNJTjYE+7lkQO0m/BTmOSy9zd7FvtWeHf24PnTKsInRDCDHm42chEY6YQshy+2T2cDJMEklyVh7l
YWoS6cCYmsj5Rkh6LguDywHDX4CzzHuPP5fXzR8hiBtriynaLqBvK3UanQLPueIbZ16k14BJ7HOd
Av93WDfdk3diiPu4g/tPhONZ4L1QACp94GlhGSuthMkvJvIiPHyohQPLo4lGv6Ddvf2ry8pRXIbm
9JxhRqyUhjKf//DQs+mEeiP/Mfg3nygPpR0J3SAefLaVjSfDht3RVUtyWk4TiSr46JFRogbOHW3g
eAAEcBHFB9xa5sXnNMh/8eiR0lX0YjKdsLyu777thd0qPxNeqRX2lzSoO/KJGfYTDxLKcJ/gOP+v
hITQ5DITYxkYWZHyBaMIohhQtn7WW2m/Ai2KGTUENZLOvjuISyLmhvkt3BCUmsZe24MYirxXXOvN
0xKEktqwxs5x3p+Tj0N3gPxj+9kjp1ZYXdkk581QRvRyuL2vuR5t7i407T/MkDMZPUk31rGy67GP
9lGNM8za2mBG8buoQJepBGbabfBRxi5+luT9i9edQsUWIe5P/BJg2AuiKz3C79B3dHUxBNhdHM6Z
rhkGnLMCvTgyGzQfdQKGv49Yjlk8g3KrWfrypHniXz5ExrDTXDFrn4n2qe2L87VDMNdglKv1Q+mA
WuS0TapywduJliqxLFFsdv902TXIf3QlM1+kuIMCa0BxmwNkbXYoWAFsZrK9S/3f7O56Madg280p
0eceQPe1pEpsajwE/RAD4sBJ8W/9lm2LiOij5FO8yb1ty6nIxgJYzBxfYErLic+LsM4HdB3mgcUU
/OJOViUfqF6mqQUqbYzA+6sYwivyVu6If0x5mswVv0Vvr1y6kFlVaqbEAsYtGTC+rwPDGAe5HAUW
MRLM/QkJw2hIF+Aa3paPSrntkm8yDIkWlYgjtxOsmUVamDGRPBaO/37bJ/r7Zq4V0NoUce/g2rGi
G8NVJrvujyaztA+PtqMSrj/NQRwP+opyQn1XyQRcEwUAkwQ5jHdk7L9bhmM5KBJqzSdrBx4bjsMG
FjAhZyPgcG/6h6PISg1hS9bcNhTSLhZ79/y1gzE74Y8ig2govdh7U7HAbE+eY7gAmmyUe9U+REnq
mohdZKJtuqAlRAvS5dAtX1gakynasYprx0xbpA7w3mxUfEFczvy4SXLnR5rMSFhXnhFoXOTWV36D
7IXk86va+G3SyqF1OjxfjgvQM4TY3rzgDtJfrg+krB+epNPWJVzQAjWhWSAONcqjyZ3XobjzGDNW
IEFJzyL+HXpG6F3mEYd2/NgC1HI6Ksi6XXeOWlhH+omAg6bHQEl36s0nFOIWpBhkja+nFrJv+5o+
dc9Q60pblB0lqtMcnrgF63Ku7gBYNuStNHfKApArLSugpcOJHEInacUcdrxU/ai5j5k0oOv8qEbj
pt4JBehADQDdM1w37+sMmx41lzjL1DoqjAzJGq+KcG0ZEoOk/ALW1shiar2Jldj8DGSy3ddV9CF/
4rudKjo2mfeBRELBSxqbQdXYzlcl/PeJtjeD3ELm2foCxYK+4QtmgzorknU4jzUGYC8cMrTmyGe6
iQuoZMuBUL8stWENMJ0bUXmD1msj7GHhPPBHFRCoCO921YQuyeJeIOx+bcDY8igcaaHDZkyeQr9Y
LVU/NXd5HRSvMi7TI3QwgLjV8NTFlNVh8LaKMFqMgNdZnuxzaIFxAi11JAmIala1ar9wItdmdP4V
uOomSChoDlGe8e2wh1PAj90sq8wKFT2txPHcuq15jzeiDGZrj3EmmzWcAzbTkX8nOrpOBXe+FYPl
w1dXGO6n5beRXkPfWwE/aFfDATVJR6pOrcO4bjI2x6sl1NPDENrG4uuO+n0GLmqMv0ssK1tQnEJV
k0WAq4JxFWG5AIaRphdlD6wUt78MCxeCxbICf5YK1Uq2ot09cOhpJA00rr2JlYMuBBybTJGONisi
R2H1VuCPZT5Y7kGF/4pOsu0oVoKyfLTeokKOTcvFFL98yzmrk9khx/icZ8VehDZvEeZHiK7Zq6qb
AKzMaiK7n/J1v7gTO/gJ9UvlS94JxM9NVy+6iHQVizSRRjrHme/CW4pO2iMqQDVwF5hi+OvtOl2z
ZRmwGGhkOK6mKIdk6gYWfAPh4NDLeMjheH6yD2wYkd0+73d6fSiP/g40TLMKr0oZ1G/xTIp8g/YS
MBTKPTNZ5nmKflX3SJQfU1lCcJFnI5415H10OVFZNX2FJjKm2WlrMI8YioMTAzDs+XC03vn2YA6V
ox61E0TEwRRMR1KU8VLpg2KYf0isgehgVNBcHnpIt2Y3Xx49Es8e8nP22hYuYfY186QiiCCO30yw
n1p2zNtIJv/l9+ZP9okeF3bI0XuPJKbG++7T/jfbglhoJSMgtSn8Th9dWfvm2Y7TiasdLHHs1e/C
c1+BPjoIG8bqVaFoBQGujzJaHNg56Aqw0W8PmEtqoa4O5Jq6w1wCik509JJOKL1HO7Y4mI5fZqcQ
St6QGwkivvAabE12Uv3JlSq5ldUq0RQGYUKvmunr1KzG14tLuHlsjJRFxH2IcwfQWuv0taIv+0Bf
k8/13R8nAKQ31qhgwhn0M7Dhfz0d/T0UI8WfxWzJwKtggzZyG6XDRuTEa8snlW6nHKo8K0IyaliD
wgUWzxVk8SYspSrptqVg76hx4XF+wAmEkBJm7OhMLqXdwpJ38es6vOlsbtQUw6tonCJL/+X75AEg
iEl2NEPVd7n80GhWpuJpWy1kjoC2vN+BFxcoI4Pysb52kzZ/Ce+OYdLzW9+iQ0HeVhGOVWJ1svlI
OZxc/GHCxNIic1X38rno9nvV/xZotOE1S7E0HG5F5OJTBplkzCeXjL7hcimDEgCvIqBUrRsCmLxD
hgjB5H5NCzv+783I8661Shw71bS4SqWiRib6ER3pFQR0zUaRAxH05hhUDKR9pk7CYn+gf8/UShkO
apZjttoIMmVyPtgJ70vGQWfEZ1fxKvzSq0G5LH4Zry4/ANc0phdyVYTeLW8zoIAYs5KpdrSf132k
F9JVe3T305Mo1lFcQ20YW123XlhlbXMdy+e4SZGihBkiD7WjV4zTDe7NKSoMjlgrCtvlb968mHEZ
mJ8TZ6jRIWOjTaFzAhQ7Y1thEBNsQ+tZbpe6W21CA62ka9utVjtXFW4s3zraBI9xdzEIa46j/He8
3aru+l2okA9k9tOgk2GvpSqED/B52OCIH1zBaM8sDJ0KwdGQ4TMja1NK0haTk2UYUcpaqGUo9Rll
/vCIUzK3GfAR8Rt9nZxZ01ho19YLbKeKzETE+V54lHx4zJQFSzrpSemD0WuOm+P9KHiyDxcm1d64
Zc8p41+XhvpaWzOs9lbycVQDDDWcCWDFaCaiPc6e4Jz4+dD/qwhqlRq1gcOb3NIWSpZ4y8kW6fs/
kELh3KoE3wg4b1j6Ery3/LXwrlwXilz+ZkvvVfBk8dlgapSWCtO/j+AwFxZ8EGILQvT+uZp7Rjd+
r67pxboDWi9KUsgOI1wmHiqNsL8SX3w5REYYoAja+5pUKMuOpEeGCeJIMf7DIv3sMuEOpcg5gKOt
5Bn26H85fxrs2xWthqiVnL59xaMDhiVRt1VgXbsU6NrzZjVflrhZ5e7NGRtQmLtxa+V3cnC6xxdn
CNR4ifkKtrpsQCL3J1zJp/llyO/JzpbpjB3G4sSH6EkBVE81bPXGVJYe5WJAkG2eX1nob8k6UTB6
Xs8nuN2I/jed04Nr48J0nmmZvi8cAo+MErctIZ0TceV/+KpNJFfqRK+pXNEAp9nWnqQZ/vwjgLMW
ecc3WRo9e58a64cLnlP/mxCXFW/WiUJUywzhqlc6mQZgDQgQtmWeNiuDJdkkGnORIdgk+XnV7gWk
+GDADWGe5M8ULxhiAT7kQ7MFMDoCdDXNEW502M5jPnD0cg9Sxs9HioXvWkzVZQWAvNNmK+8r2Kuu
3t2cYerIHwBHeZyVwF8Slb7LAPrUGGbxo/rHASMlB5G37PitceWAAB6g1PZYcL5UcI2uhlN5rLs+
xINMa9tO85773w8k85zdKqy2n+HP7HUafuqqHqQCufpXNOyvwPawceFhFo5q2RumNQhruYNTAQpN
b29UTxVSmmoNSd797miGw3ZjBtDPuFoEyNUCak9r6PjnfYwpMNABYpp/zKUgWm5pUbjpfF4v2wD+
yq0MePGOcX3SpcsJaKuapOsOF4aLzBZvwUvtOjJ6+7LWG+Za1aVqYcDDXeeKdp/UyldakHZap+xK
rJz7rTth2Tu+gXsBN44nuVBU2sEsvW3qWrniqQjVN2vx/k+g5O4TmDD/kMUvR1mDrp3v9+6eanJL
eltGYA14RAZiHjF8x891lNp1lkJRXRzcCTGOljzwd1kpRshwNyWy7jUShn0YX1QhFBISr2t20O/f
QY81V4/PZBaDqWrtSLzsdZh9kdtAWN5JkZQzmLQCLWpq7EAAH7kaEunwGWN/IoUiOHDXxOZGGoqP
I0gulBPUZtF3tUky9bImWarVfAoUfMd7uy45RZssT4oR3U2wnDz2oVnxOTvVcewCZr3E08QDTBRf
ts2BVbpTAHOlaRBEih1lTh1+roH6KQXTaXDAerCoJnzjIvfirZwM5/nYXZ+l4D3uxrmrXTWAXxLt
sHqljQPdYpHi/+QjLDfsrcNwxOGjDtOCWNJvBmAIuv/FrCsHR6eBP57wvkdVNO3NKZgw9u7wFSWi
TU7Axrk7vAiV1mfSQ5e1Yher2AFhc7iJudfIRo1xTGQxltPjgS0AXnxtwWEseVzpL5PPQE0SlBoI
Mzf0eHTAwQJU55YMgL6F0SDcj2LYMUL+0pU2wGDHJd5x6xIQQHH8URKGjFz9igHRFwZ8ENLquT3G
sIQDZNoRuVim05wBwhNvGL9FBEik8OcAYOocwAaBK7juER3ORkjTU+UwZctin2U+bmS1TyOwjTFA
0EAF8UYCxBN6/jJF6Z70wW1erZi+kPcolUu+B+XVWZClZf/nJLyZ0T5tGL9Xh75Nk6cttC1vfAxE
n2ReXQTBzwYjFcKtGhvB2nSBXX2YeicjA6WdIx8lZL6XYxkdzqmUtHiisuMkW/V5F94TTNL2qDYH
Hpmsc/koCnomq+ebTQ0ozqM/AzFZCv55kNftaH75bo6qHo/4QZUunICiH6XSf+DGVhzUq5c+7uWJ
Ei3R5lJFZruHXsWyT10B5Z4WRxtYlyIVC51ehUo0jTGXi1DhY61Sj7/WGE15+ABDrg9zAJhqBsOH
KnuLCZk58mhoN7Ocb0sJKyVmqOTXze0M6o/w/iM1bCs0DUoaDX/1G4TUFqt6AAsUOZPn3Gm5xXoG
4g9P1o83rGu68U0SqdoTUWejyTmzTU4M+BREWICgMVv4AYaKliS2I38ZhCZhfyIdNvAtrjawr9mG
mcjvsTQlxV4pgNpEm4ZHCXmS94lCUMmJ+tonf7DRumd0Ku4glUAJI1ZQ4X0mG/HN9TZZQdkfkhxt
2swiCV4aGLW1bQWqp02uusfZ+p2zl87dZggyLru1sDG7dQS1R2uF88/nUHxaI/vpKcUmnS/WnXbz
lLPbp0oJSghHV8YITN22JJC5lGlyrRnjQ/07g+23Z/grttY9U9b//ELRPBJFk5do37mFmTJpOb35
oahLfPPKxnUJl21kwCXIwV/mJnKkcwwKGrQWxQc/WjPyLGnKxvJuyEwYxb5kvGm6nP9nAfhLV7XQ
92bqTdZzHmf5qMSK+pUw67bDUE+c3gDwusPdJhW96BzT6qZIgXGzl81SOXYnYnN1OswN6AwDuge1
9k1DnwOvpR+LjL8lFWSnreRggM3d5JT1DdJh5EISdxRveC1DuzvqichT625DM8l4SosvYyAoigfw
jSv15Hu+geiUYZmgkRPpL4MrE5PfyM9q8vUyxcsbgUD6xVX9bJsOKFRV93nH/9hjMyLJCfIa8kdi
q1kWKlsLZquYiNbbG2vGTJULdnYQAY5b259cAe1cyTSwBycLVYoPWGjbHondKpShh8wApfKKu2x3
1xy3/u5ru/r51H6Dy0hE7ZgXm8CBzS8GzM9b3hRsfuiTLVc8AQxiR7RVTHCoWebK9S4GTdJcgLxZ
3y8AChNWK5PrtOrTR6DXhGhOX/zMXUxbkDcL0N3whXSnghGCNmh3XFV37MfvIFsiP8vnQdc58m0T
lYGmMqL9Z1CbA8JJWJAGyFiUHdwNTPwYOB95jZBJiWtdt4wQCxYhbV8zLRxwj8mymkKnGVtYk6wj
SFaYMUhiWcbizBeCvLg73GxqGSmU5wYeWesyxJLqx+G/hh6TxK7IgGzIb8L6P7EO5zJn7NsD/0da
sS0Ee5XqmMWHs7QRm9WAjRHN4tMo9CLPHyQ1zr/yM3gd6FuF9YNsQDo+mfs98yTFbD//LUPG0SIl
AI80pvEisoykPY4uAQki/QBaJXhlzT/cK3EOj7e7ZQZBzrUjk3rrraiuJ85XItlklOlgUMKBQiqH
WY9SW3bbI1Gp7YsHGG/N5SLADIcWJNDHF+RngRgbii4z6SQhuC+argKLejZFMd1UJMPs4xtCYgWe
ye2pCnU0KU5xh9JwG/Zvo/qobbHbZIfZx/P0Cufuz8r00rGZs64NSsZzHC5mnR/ya/vKlTzOa+DQ
EX/VmFLGsOltatgFVsQx488f6NHzphi/qhJJscr/MA0SoIXRFFWBoA42b1gYj1q5czkkAbDdfOcQ
yjJXDVhVnbgCM7XJGdeJ9J9gHlm45AZM67EnEtOSSb9F+scX1qQ30FROhSpBwF9jMzD/dQBvlvdN
wesCDuQlNh2H65LHflOtlsf0OlyaveTlniTqGWPFCHbX18i+bwO7cwr10V4BXEf85sXxp6atIMN8
Zat9jaUzU5aOeE7cIB+s2F0VkiyV6oLejyVqnpNaqoNNyequZECxclAdTBCJ3ehEl1wxQNRJ7Kte
ZHZ3M17Cd70ohXwsXUai5BwRhnfoqzJu+D/ug5fSNR6TPTLZdhytFuB8n5PInV1BFjka19+ERNND
xFR5K3EhXdogJGp3JMj9od9uxr4TOEEG1lwQxCDr7PQ4mmjht0w/aC8VHZvscyVKvcGrLozsaqM4
rCX6NDg1D2qDkrPChXslrCRg3HCCvEn4iDgsV7rbc/XQ3Pn/LPOSO1nSDtGHsmxbeblfu8QpGrBu
fdC/8oKlWzrswk19JL55/mWFZ4q+nnmjyvAsv5jhPoQDBbdCmnQLicmUbcY8a/27ABLSBCyb1JtO
bj1c3bu26wa+seKXW/HpHTrAdc815p3aemYFduwKQ0z+RN6iqawKvIylEmilFjLyEuW5LUwhk7ri
4ldeBuiHRC0mhWzFJmfVFTqQT10BR5ERlbkSLDbYBmxt+N+p9dUzGAIuXDsVTKEKKmgi8zyu51qM
x6pv4DQI+acUs+5pDiqpENWxroVK1Nk5/zn7YIOwqNMoraluLFQSTLS4t7Gp4xW5T6GrM2j19jgI
bxtdYqYBDoSzrtl9PXtBDZLKEz2RsyRXKu7ucO6VStAJfZISi2jghbWOVfnhijOEj/MoymQ+K1Yk
nc953cbIstduQ5a21sZ14ToZjA5Z5kThu1d07FrTrsrwYX07l5xrVZfPUAME9+chwfuxvnj3/vbr
vjWohbQ072E6glI9jKTW00n7alJQave601Tk0ju/adkESQHyR3L/2CUqGO6Ojl7vZcmSsrAOYFMi
wVtGsWWIM7jtKcfzNo+e4C+dUak1ftNrmA0SYXkn6qxZalyeXaA1E4Gvhm/kH88hRt9fnCcBzvMt
V3/bi6jcwD+UVac6GdHl0gjzP3nvIO0g61bCxcJ8IXKZh3v076KzSaQwNuaONzH7wxG/mIkc+h4k
X2NKk9FAPpsvRumDOxfdb+gTZTgASlQljMrvhTz8vqdcR4EzhQMwvvFtkOgjv0TXdUdh0jLmXDmj
n4coOygCzyJu3g1Ni8L+5dw1IOB1dCZc7iZlOMQaUIIM9OHsQWwZPzd0T8vatjffIkqe+JZG6stZ
IFxx9q2rp8C0aYazzh8YbnK7Lzglr2WQuqxNmvv4Eoj/qsh6VEodZTNM4H6AzuCSSNTH8UxNPxrq
Ybxl0ddZT0Hg0/J3G8Dg1NC0ufH4aPWsUHwX5ROfUB6UfEUZuM4u6D3iwXuJvPb2cozAMaJo/wNH
iAvewr+okoX1HxbDDidp/bSXS4YeoHNGgoPzFEv/i2cvxYhIG5i3hlrUIQWCF6BqNBs1PTVVfET0
TCePC5Q1sCGd7whw20pLDSjbqtNeYHCyphHatY0gVpuMT+n+DkPahs/55uMKCyeoLwC6vm6rQaEs
4VcvJkxhIS53CGFxCdCZcYZBGKAsiX1QejEiSXIa+qYDL9Lt+lYWVgwm20Aq+HnQdiKvchZ6repG
82J3WoFoBj+s2n6MV6YYqnBFHtQjewYL/u9x/EMgNjlvV4/u4j/ac/qb8WnMIZieIbB/qOJR5IuV
8U/nyXiviJ0bXRhaVJLdwYBGZffgzOGBy6dgb205fFJubIMTHuymQ2UoreIC+XMqnepEkDE4YMMp
XEKahZp72nBWb8c93UhE7RagtqAtrcbgItOrXzZla9/LMgFErpdC44JmOtDKZrlVDKq+9+EZkFdR
1NMqzw4mc9QJVX7oDNnblezEvO2At9ZTfRyrDUTPsi0ip8bbDTkbbO0LULP3JFg4Phio0RuTGzxH
VqH60BDaR0FlpeXafIBBsLgBqGi/mqVDu7Xidl4iXKZoLjRt17nycts6ySKZgePQ1zLojGDwAAi4
uuURx6f6cBenGf/IoueS79WsGHtP5D+jn4kkzfZ6y8Hf5KtRfSu8uFaaqkUvWJXPxNZ+GQxkR2d7
RrKEjI/xIwX4TmpMaZX1hskinOppUa/8uSd4k0DcYfIwtYIWrlXgeKSD1ILb9k4MeLfxVwTaq+fv
wHdl71Fvxv9NfHfqVtplW2XtK8T8UTSI+9n+/3NfqRvRSNvBdNetcL9PEnUHSVBsN0uu7Xef3FAp
hmRaYRjpxbkpMu5PvE6Ol2sL0zmFvIKpGDBn3VW0r4JP6A2KnTus8tqqmsOSbzG0RNQJX8ZBJ6qh
kuxyW8fH8xSSW2DtoRExYjArP6v51LfFNrQ280lBJBizJDIw5MarZz8xzprMgrOLgpqNmUUj0VzQ
a4Ww8c4dy33BRjemMH3LlBtEb+z9jjFhqtiL4oaPHBQBtkrJiz2rpr+msHBfN37k2kzkY1NikFfW
FilD19r72+kUpfkhZMpltNMT0T57U3hIPLcirOZ5PsH2wH3EECSgACHg3tKZ0K2MuZCo0mt/zQED
+k6TUXe/fbDQBGobwy6ytB9RV59qsvliT6T+XOuLCfB/EdMw2uiR9GCgr+4Y4edcWgkeJbzQ/vQb
zV7vmjJIk37mN943NFLBqxXH/fFc8xYTleSFRXbGqheAV1g+i5qiza0+6aF2OTagIkW59s0WtNeq
8YPhLjpeFs3SC9sSJhYRQrxQbQlTkGtZUtsS2fdHIf8NduXIUe225hJITMAdn6prBkOKU26JENIN
CosHyJD0FcFNwnXIMfTLTbSKKN1LOI7HGBVfQ9o8katmPccXGr8yiuIJZLPSml3EDr8Bk5gb3WWJ
KZJXYR8GXoTC0gW1iERH8Fw2DrWbfyzYjOes+z4tk++db8lA6m/o74bCWbBt3sJouY8mAmyjl5TQ
3e8PZvAXcUTMOZSdxq7PLWElUWdIi+ejzAbUUED0w3QEmz9dldRBT4MPwtpW9yUMJjgYz8JyvjMk
5ZInpYTLG38CpqGq4NeqGxG6kqEc58xPOs3eyzIg7ptIAjkTTnLocx4WobsIE8EMXlIStCQTUAAd
hatLnkHJBNQ7flC14CpQU1WZ9W71bksFFOPQVSWXjIVq9YC44MjrNs170/jBesw+SuNrbCHnr2ws
9nS9tKdBqCsDiJXVebhd7p/5oz5AAt0NF5CxuuVjY+L3IluB7mBXrkppbfwqr1kkbjnizhTLt2IE
YC+gTVckvkxg1B43fYziEX351/FVGBCMrIqVvUBsx1+fOxuIwk8QXPf31xqDNyF50A6VrixExmsJ
Gu6mfYzUO4lLnF0rHXrxPpEOyxV9u7jb2NndOd79uHfjnbfRdfDBHhgAPkQqRQe7xBBuLWiYTLTX
Eq23zFfHdiEpTiEV3BkSdlndVBc8P2qxQoo2lzgLtV2zPq29Y0E+HbZhyEtY+KCB4RicMh32t6mm
ItrFSh3ZN1vvnKaA84QLe41NoEuiGkYBo7iD7jygctJbtI5bTR+w2XtjGnROEw/s8DTVXKWdXZGr
hDGlkmmf5+IUHpXoAezrEtpqrhh607vwTRnciaEbXU0XYcvdDd50wW2O/ZIGmBSzzzEEeM6UUxCe
MMjWmHWTDYe5MBo5CcJE62J1ZpcAqn7xCeSlyUa6a9BYhdo6tt8v/+eHbJ7ynF1CQiLBEog/4B8J
OyDZeruELimCWLk0lOBoKWNPVQB83zfAMfxM9663brttGHXOzNQMU0X37dzcSCNOoRkuXTwrJhCm
e2aafgugHfND+mDMa0idwJqTGcx6iXCLiOehPEqlhI9HW8jPpzidAHd7IQWC53ygI5Tosrb5Bieq
EgO4Lqo50olaQzdcdUNj/IUm+hJmBBoLCKDJuZFRAEAVgWzGMVa8VUbnGC89r097QdOdIUnQqfuK
XGJqOcj7k+LgNf7zAuDixartVnCZQGKvIFthDsGO9HtFcVeYtttZLicR22Yg/HSFICP/08JlsUyZ
uKwQclSCIb+pMRhziGYepZdXXJMi8/qKLbMX923xGJ1oV2r34+sy8cROpm8CuabyHBDmtc77K0NP
AKzbMajGxeyw8iBs5kYBZ29IDBJDKglcnKOMXM4LsTWav4j30fC+Sp+iAwR4tLhtjSVKJjdPGS99
6k6BZ6XsOIVfdOLT0g1SttxvUcW1QvZnJeVU4CtzCwLoExs6CusrnzINcsnNnsaPSdSkd6Mvkq1W
SMACXP0DWkVRUtN+RRmvLQJ2BFRKLYm3TVh+wPUwo7H6otDlC/TKHJQWMjJrdI/8YtnlFjYWScfP
0CgMSj0DrD90W1G4CGWZvTaGVE+DOHlby0EztCD/0tJnpoDaAfxYDdX7oWzHkfZE0TmU+0KgJI+7
eWmoOKULKL2TO/QmspfNmd2Nj8CB56B4fY672t1YZYKqs4Vv9pw4K6ALNpjDtjfx/1GIfXsNM/g/
iyMWCzlrgFrxewWwLegQlNmRlxZutZ6a+jLFQb4ZS3wfj/I8cjwkPzY8QW7OgRaFWOcrVzXY0CPw
UTa2W2iBmYBvzGtcXL3FHFRlHLmWudHHVFHFjrg9DVQL9q98qg/r+Gqp4blz71ra+InW9gTRhRzq
slrSICxIYYyIb4KG1CVeDBNp3KajGb5LjIqo3GYMjK82x6b/GxIz4mXNGCSuadTDeMcx5ulV9FKF
Tc2msMJ9By6ZFNYjB0qB5dM8G85vxm9ch7I3sgq6MYf1Lu/rk3QJ6GHmlnBMGnHzAi5y4h3xODEt
LrHQ/WtszFUHxrnU+k4TvoSwCwG+TfIzRJejbj7QTsb0/Zdj3CZY45wRaPVxgIg2kMBXo7k5uIyB
l+dEH0o6bIaHxuxdtuf4rGO+E096GJqwUVwgENXjWg9+3Hm7m8w02RIM201dHmEb3FVWJ7t0TJHY
QJjVLEWJAkX4lcvI+JCtcj1RpW+lv6JXXOyVAnySRKCk/rTRCytewxQUyf0M2u0Au3RuLZkq2L6u
b0yXQZkTXxMtlcOnHfZdRVnwWBpiext4VitITWDUpJFG6fjvlrpRZGAylTZCTcs9Egnf2Lj49KCD
sEXwrhVqNT92ekBrhU+X7XnZHCtyXV+LBMC0RCOl3Tioq0ses+5RGw02uAQLY9KkXwi9lf/26n6R
Kg9jqP5ZXq0euKuswApe1/diD4LjFTVJBsGUAQN67YVZnlcMLPCUSkxCYeEE33/ESkGydLuX1WSR
8hnOsH8/nRWGKKyjVRIuv9/DvAppZ7a+iZVdsBcKKr8mw3rQkBuqBlHaOJJBL1nxhCvGG3yibtvd
YLdzhy1mY2f9RvzyQW9K4hyJrLlRjjdHv9FwVuPH/Rd56KuJs51voeSjLoOcMPFveajU84rVI0xw
jUuuImViAbu9+yciI48R1Vi9mA3shlTaqA9FMuEYWvYq1hJ0rndopzhYMHF/z3keOT6FRLAIjE8K
37IhgB1yBlCTXwOqFcMDad6i3dXSrPz+qN+XXK9dnBKg68RiwuxGJmXz2tsz+4qi6IHZ5YkCyaBy
IRngtqasR6wJKJx0BoNws6O77voXMEqVTkRtG76V/BZlNgTokzQ7Po7OM0KWPgvrzgI7WZjSOMno
7pGevxGPqrywAC4ibLFhxIMuwskAgDNlgR469Lb+ToBV2RkHnsIeQ6TTLqmpb2DxZtGcpHmopbmO
8dD+7hUq07hipsbilAhHJYOSaFT/wCNTqXh0f/UpveFRSghICqwxbWDr8QyGfcMuGzamzX6YZYaS
OznMtAMAErM4l1fZYdvMsnLchAb/bawkbVgI29g+H9bnLBwQ6vfO850Bp5fj0YlNn39c1V3NZdst
zY/sHaPeipB02b0AMEb5dh+2t3P/MvjnVrFotS3gWBfmKg+qIE9buBj1iLG6zQegnQZg4TnrNoxI
mK84HfcLx2yfIi/VL0nYahzEyxCqcaiZmNQ0HWWa/hl8GcrQsYs9b+dxQ5L9E9T8Hwt4PhuRfDxD
5JxUcCcPjQ0TAa7UQewYFLKCIz66Qn1s9kwobgmEJrNrZ/60iARAb7ZQxLH5iF17lw1R0nbR1mWb
wwj65q4hI7NUagVjOxETjKD4ndImjYbfUh87b7l37OXR73hRwKd8YZKhl5JcKKyrp+4DbVFjwZae
ryQsVIi6LK9NrVOxDbSukMQ3OAaI6053q0UMGMHCKxfQxWx6dvlp8FY7kovV8EZ+c6X5raxS9a6Y
POD8ViEuUOBNj2cnR6uHYqXIpNLG8i67hLBVLM+dFem1wj2l7HaEj8wv3UVZkPliytQGMpb6nyyR
4TKX+x/y/KGsfeFdaXO1O1oePrDzZWdAeZblyBSKRXIq8ixQUn2KHKcoCtp9BfS2Qmd3JugvatYv
T9XEMdWDrzCYasNxgHvGebQc2oSX7ugZA5frZcCn90QAIf2gM5/AzPln3kbAskj7FRwmw910XOm1
tj51Ep+HsMsVjh8D1gjWgrT9xCWQGMjqXkPMDz5lEOuX+sL0UE04khimT6nhLlwOscD4OlECAnS3
IUCDrWoeykB6wppqw9fHwNF+ssA67QMEfyP1ksNg9BHH++AVTBiz3PDg5wTZz+Obe7/GSI9HiWa5
hoqhcJw+IdsGnnN4ic6y+QoWDRmDhqWd7tzAxkHY3YeizGuXmOXarXxGh3t7l8udoa1NheRnmTkL
4tyd8qvqvXjAj20ABEg8FZVK6Tn+Wy4745kceXezmXwkuPR/wKr8sWXTkoJtmW7IEVn5u/URBNGY
/AzS+nEGWCFCJ5SdFiJLUIvgq+nVOpIQZwHk9JZKzPmDnXlA8CME1jJSEanVFHpFhdZ08o2rzQC5
TZ0+EuOTMqjtKdmNU7DgRO3fSigh2EYjHVviSd1R0NsmvgTUJmgU1xWvdwYH1jgJODeaMVGZqkHb
5EFbiQNO2idIXky/EMSfKo+LAypSmy3VO45oEX6K7FL5ThZJxKGkrfcjM4/wT4H1Xcyvl1VClMJF
w3njz+t3+8jQJbCvEnusqzId11d2xHKvXIXvHb4yknJEfazMdPWAA8A8d2oMoekeQQuka2sQ34Xw
MZOzi7+xuEm+HpjRK2YcuwQ2cLKiGJjBADsU9dO2hMZ/6/xEOUj9wM4uvl7yl1bVy9pyMH9orxKD
AIlE5AdtxrGgBTFEQrWPy1chv4lU7Fk7XOcxedddXua2R4otvSx8cy1nvF0PHCRk4x8vumZpNCAi
H31Jfm+hNG8Fw10wEqwbuFjUeRGLys2COfYhddg/rOXjSIkbWNTQYW7AL3mjPEHyFiK5oElelw+Y
2bsz5yU1BBiYdv0T6PcKymw+skH2ClanCOQu9BQJH+Jg2EzE3TcVWqXdjxIRUTDsVZpCkoOml3Yn
NAoKlRvd7m2g1H4S30A71hGgfQv+3if+Xf+TzOmrV6soJe8wefqc9nY6rp9HcHVUSyYDhigDCPnm
UZ92bc8T0HFn5b0n/QiM2FA9xHpjE7H556eMogHsJDB2ZC6YWEgRP5JEfgD/mdOR5rj2m4wBSsF4
RhYNliUNQAJ+JUzmVaeP6H8gqpQl1tKXXsCHWHZZ6kci1Ny87/0PoEPS3GDsfIhsGybdKTYuevxu
UpltXZYaFOKmTnH1a+ZvxWF6y6cz1R/NIfhGUsDy3FRlqBNMgncV9srRd0JPw2Ks4afGhLUOmljP
EjVgo5nxud2Q8cZsnNPjs98Dyk6bYPSxuk93aIuFN4Pz/hmXVxOAHeYjBut1hkn3QvO2IYzqvAjs
sqY03sCcbt+Ai8qlhideKBXE65jlkMHu+hG8A6q12ISEy2pP6UYOHBaWlXz6mbW/ORERqC9RNt0n
RX84wWX8xXjHk8OKDnuELt780M4Q5ajRnBQZ8LGV6oaQ1qfB+OjgM1iPe46+bsN+eDx0sM6Ilrlz
FtTV3Kavm1onLgOOnu8Gkq/3rmgezvriYcH/cW1WhUxORvdEN/dN5ohmOUoKIVBimToVVGrLewYp
+3pBob+2ARhfPxsa4InyAtXJTrrsECO/RdkXYyFlX799saIWc19yFmnaY7silYaWcwGATnVVycMW
upxpnxhJsM3mNW5Zm4d+e0kk4xu86yO434g6C3k17X2cMERlt/mlLAeGEwzoirUCeNcB0lYo8a2p
/hO71asKTyWX7f8hyV5XwV/gQY6OjdfZBlo13kCcczLVipQh3AODxNWCarrN9LYKGExH2wrq7zOm
sDt/qXqhK6yhUZNXMYqk97KKQq45Suz+h1IrX7J6gAnsfuRuMHahk1ivO8Ssc/XLaWfHlBdNz5rw
s+HTLbsOxXQegYBfE555UL71+jcozlEWANzUN2dZwa6szEOy1QaS3m7rJYvrvMLMSdcHVRyEshcO
9AIJKUO1SR4woNHUd93QNosqt6v4gLKj/nsmxQ0wTK2ghKRnymDzNsSpQsGtJDiBJGHIjj+gFdR+
DA9Aa5kTlypvHLPtafT4QTZQVReBlWVgz5JnVxkDB6jPjHnSEHhRevVHaSfycbjybO50NlveShFy
xoG1bv4Vlg9yqfxyvy349DPs1dLj8GoHrVNIzST+VDEG6zTfWkYzxJKLrEsfPocfOsd9lw5Um4Ig
l5zYAhH2Q/YGcCdPSIeOs3y7PJ+r3lf3ZyUKKbbpiyUW6UcHhKAjRP7QjDPgzOGjikbUwum4c4P3
fBW3jVM7sOrU+/ddBKQpkG4SMgWCt4pVj8OsTei7A/cEgZ857uGVokbTrNvnc+RKG8rS82213xZU
O1q9f04PkBow+83G8yksnTkujbWAUlaYATtSABLgYPb5xmPB8KlRjNf+wQKwOmK40DCv7MJUV+FC
B38Rc8gBAP5UFVVEfOnDJ9qiu2lgrD+ERxbYHvaWsAgNID9/Us/lWY7y3lHCR8dGCACkuJr6hFHl
mVuKQwlV5i5wzQv4yQyk1/Z9XQs6TT4E6bmxkhGMgGMNecXIJAqKOGCgDXGA5vw4CPcjjMN981wb
yB51P3u8xx7Rd6pm5oRfXxNSM1toq10s5OH5nvYvIwJEq9F0jtgDUd26otCHryd6S7mazl5EdkRm
jNuoDHUcb1jOcPsZQn7yQY9vWD3uFxnTxCSmr3xmBtsCIw+p/s0K/f4vl7lIdBshfDZWDjc4lP4u
km+zCnEFQlw64v1PFvLQ3bJO6AoAZSfDu6Zhh+6iO1Q55HFu09xt7AeAuOOXjW46hHKR6HWbqefU
/X2f/47qthrL/5iK5HjdVDnf6gb1v4PjwHSg6y+Lun6nTIS0GaRomjQm2frqWTWgjbBZzv+HakGQ
R2HKi3dy2ZeDK3Gq3VlhB7FqKv7GSvWoPmzWBnEkU2QTlKUkuhjUul3XgUgl0wwYTTFMjEmBRHjC
fYud+mXLgvGlZOR7Qnov91NGdVVUkGYkPV7ZkeWdZeSMWkx56M8VuCFja75oYmXVCsAY/BwJgOeL
fKUeEDxALvtFuA5LqAZ61zAqgssfvQg5xXtHeFI8xQ4jq4iVXSG7df+MH8fn9zPAg4C0gtRnbx2R
gEdJIVwphl+bLjglsAhZl7ROHzbNr3VfIeq2SHCfYZv+nMMb50Km9DJ+IYSoFpAIscx3l75mX4Sm
HlW2+HycWsskmAX6riZiN5aIv9Kdh2fH9Bdd1IueyT0FRQjB86Yg7TYfUZAZMdGDePKG5+BjqueE
uFfQb5q/BnFHL6W5RgvelqR6Excs15AXOfz5utXPMg/1UMe+3R+NIu0UlW98YXuhsIYpmGjnfqcz
uACpRSPw2Nf+ipIsnhPok5FVQJsi3oTURTCr1aS4CDPeBmZw29L0vRwtnxHv4I6gyUrBo1ab4k4J
f9lQOsewg5T1WKmujMKzQmwOr8MYNbKGP8C/vPz2IJo5Et/bKWgowzkBt4LO8jG458t69EWjwGnZ
JmeGHd5cHyKARl1pn3J7iVLd80DXbNw4YeuwSUxcGSCiGz2fM5UlvqDbJDp6pl5P+oP/6TJ17Wsc
IlwiO6jolylueNhLKtIKHmLPwTwvthtiw2Ls9x7MLhfeN9whGt+juUb27FQqFoB6ralbHdq7EGFN
cBhSnPPZ9HEN+MtXMxQ1/czh84frLASNeo0Uba9fv5LdWvjbUbLwKSASSFtbr4IkFdfRtJe77fZQ
myV06FA2TpOsHjuDC+W6N/Vb+JkRkpJlRdsZYSZrIdDmGS2XGBL4s4SeOEDHMnUnBc4oAzJMEXhE
fiJnS33jyP3M1vbSsJRFxiAvnZbXyqUv9YZmg51M7MPHBkRcKfDkQd+HW3aQDj5kVwkOOUCIXhV6
UlpY0axg7EWDpjQUblNck7s2/v8BCA703vtfgdHI/AsleU2xy/M7mcCjhweeyfHBRm05QRgy/Y1b
Gu4EPWC+8uFUkLijU/pU/HouHYyDyHq/12mNjc/K4DiFHjYOIZ5CpYnmQJiqB8pgjVIkXVg/sCxp
6ByZNC8p4LtD1AROKBiZ4ToMvMjTu+vnudNAwwoo8GtyGfcr2yhoxDcpVPhccJgpuyJhAQKaMXCq
PKUiq0FvC5GmAKP8eHetw8DsX/9Oa+vUnY9M7LW828GO/uOjsJN3cNqbFAjKtk2FVlf7xJaWLD7s
jT4vaA1ho2NQTO4jYN2orf7bgcyNVNhvVqOeE/qQYfMJsSuOw8lID91iIltzSd/sOwW8tHFV4Kg3
xBSTp3daEtJ9JpeAkpzHM/oJLXxoXECUXwJL6CEwMakk/Ek1g6++dSHhcP2hIxefQ/MEKnaKXTRe
JQryFABkByt//fpZFRdxrNjhmS3azStU+tIorEgSPZqpHXmuDN/l2hONEgQ19ADDEg0X8Q26L79l
dv4NZSjzdjO0vcux9X36SmOzpA/lQj2pfKyAnhbuoJN/oq6FONMKrn4HTg9zHLq17HvYBeFBtN1a
fcHLK6T/ph6np5sX3ZaOiB7x/bxkRVb6rCaPzvXxAEu7h1UxpjLAxWLR76blQIot6y6RDpzVoUmz
jNfLe1s64XfuT8g61j7THkfeJqIGVKBskvDuuiO9NwmL2mXfEaS9ylG5YcrInnq38R2sR8VrSXhG
diRWhoaWJhVjaWxeeoHwLlEoum2BtlLb0zL5ZY8MsNpAdcC+JkCVcu0/vmDPGsTWX2fs7dWK4hzB
d+F2MGLwO7OODADebrkt9jJAN5roa2igpkQQGWbGuyFD6ZBpyg5+P4Umb4SipXYJCfKiiM85ztd8
x9ycaCyOffwlO2PjSFMQ0uBnAsk7ytX+JJcKMehBZP8cZLgu43MyTkgFi3hG0xl9xcUL/2KLL4e+
ayMhauakPXtKtWpM+bm3mWOsfRxjwZLU+vbYmdRJXHNKZCSn6lJbbVeH6rjdA9z0HrkNhH7Tq40T
su84yGp1AmcJg0GB8Mfc1qC4HOpwdiehchKnmohf9mcTsD7UD4H84ZOF41KQgFphiT3AePUj/lNk
QC2bENirBNUCuk/M+9abTj3zE141gXhKaNVDcBstdcaQV9KcYAT8CrwxSyL8pJ27WNPvnu1FLt21
mFfPX5vJdmH46dGWsYHehVxhU/yeYtle8ahbNCCc+ZSHTs6v1kgWJ1cHnhJb/PXQRIcaXDkgWQR4
brtJFJB8YC1WoHdaFnITEVw7aLAHlHDpL+TuptWFnXKmsx4fQkfg/QP9fxG4V27NLP4FjzmAU80Z
OTI7t/eBws4mlRgTUaD35p1Ma5YeC2TFtP68tcJFQFaIoSUGXahXHTjTb9tIG41flSBHUXhms/nG
teVNOhQXQTGJ727BDg0lmkO01A3xDeB8sAPn2M9M00ulkK3JOk5Yfk1Zz0ZRPgIn5r1no5VcOviu
3qkro8kWKk8qEOFz+lYDmivOSyHAsM0rHkkha96FdhsQydZ5fTO3nHaTdajg/3vBEPdmHXQ2j3Bv
P61aTMjlJj8G3xHlJeod1BcO/QUgX3E1aifBbaJsE5vzHseChBr+lvFejl0T/JIAcz2xtuS2lLMk
4/6mBmuCFcY6ESxFxINuZeEnUQHfTB2j4QlAk09B3v+AjDJZRAcLuCQQewxnvqUeQER0J+kshewA
ztzmtU1F8U1Ughpq8OR5177WevVORm6bLJk+s6rpJYkLhYv5UPKPYZwUVmv5yMe/IRv8sUsywzxJ
nCVEAc/EqqGzeMUrw3aeYrzBBhkbQjA88iWslp+4pq4gYiYFpUOzKOX5OEWCEkmIWMMsiTiNQ7AH
H3LP2aJGLB/u6Vom/hkg3h6c4GrF5vqEa2c3nb0JEmgY1sXu3nQglyZx6LvA5jUIgXy++TdfHavS
A8Cu8Gb9TmGfRMeIbHqER8SJpXGYCFOD4CnTOzeQBN3U4qWkWkhm09BCJlj4+HUto8uVrbCSL2T+
08+tFtuXWAFsFI+nGdjgFfRY7DU8B8bzHMEt0MSuK+RMmfl1UNR9/jSv4eBCz+Z7FuELogfrCGfm
7GHE1GOhBWrAD4yc2oVO9wBDjyXUmBxAiMW2ysDMKxU3mTqYnWq6ZJw8sMlilf1sCSfUfNSRszeR
AWAlRfcr6fBEz/O1Aa77eqI6CfOvXhigig7Fbh05kKM7LqELBBSZ/DWYAsV89sSGOxHa/dogAvYQ
BlQNBcRaPJPCx7EoaFG5375z/CKmGsoxXlbIwg709PRloUO4vGGbixduFmNR2didoMLqA7Hvfw5/
vnA2Q4i6eXCYgOgDwhQt/3BsS2+bHwfxwGGKGUE7SOEOdB/mMPdBCXMbM13a6Vd7geY8t+VeEpJ2
nABwqs2frC13hFQatpByBtCertUdrhcAgP22lZWLzg0gJ14Q3rtHTWu1nl5psG5W2HMYuNkoNpZz
EQc1XHReniMbnAV6EjoPd0sf4/w1/stOhgRnuufnWY9gdfzJShNvz0gT8JvCqjY74Ce87Ml8YUaP
+DQWBwZEMbGvXwiRLrl+kJjiOkSzej5q0Ugg5BcuMI+ZQGw4ZRDn4+7LKDv33zL0VJzhml9dfLG1
qmcNJs8fCH5lq1UDFyCVZswmuU/d9yG98c6atLSNZapMAbvKOWgP71L4Vi7szaYSDjxgRUjCQUgi
4f3+Jbpzc+qEoN33yM9rRkiEzOAN2Ph5xrgpoByw+STeSWIpFoz8VTPh1W2BMSZpMZRhiuA9cutn
Z5L9cmFFRCsvLZ6F/Enfw4TaSgjBacJRk2oGqfiHoTnD1Xom0pQik6J4spU7hmMmqDYWI9MUe5Ry
nX8nRSQvPsAlZjk8UQZxAM9XZI2bef2LgnNyznEAXjG4vOYKhDQasDxds0si/LstsCdhV9s6hk5X
fZP6cy4OuEGLm43CkB2ADMJEyNgTuwxTMG4oQjyoFNG2KoTipmJvmwnw5gjO3h7PewlgaXD03HnN
u5I6FlZfhbfYBfC1DA51E+Hq+MRSwdv34wiPA824pDh/gs9Qw6bTtJX8Gcn54eE+HlIWJIi3OXSN
27qvfjjDbWy6dWC/Wj0twrYNlKbjWMjZWIU+Xv+97Znh7sM8Mr7XsxJT0Xrc95NPQuAjSsPcbsnX
1NzAheCGODKuanWk+CGun0YlBtLmYsLkAqYSazSqH9F8n+c1yzs9NZizP+RkwfK+ZPDFyQX9VXJg
hAv0NAlG3xZTTMukybgpG8lFOPsHE0JMI4LSQNfrWGHUGYBdWDKBX77xn8noFl5C+rKDSrJBCrD/
RtglovFUDgpZ14ZAw45BjGg6V9jHZ4KBg+qF+9gxqgEn4LDr3GfmWabixEvUTBYYFXbfDl1B/dhV
OqSRp6n7ZrvMqRKmlCznWlb2g0oE2v6z2d/mnjufM6xD/zAwPwoHumRQAgvkTw/gzFhYKYDUqt1k
TJ5QntCzrNHPsa4jBNmzxoHLp2ZLYV/SYdbsNGbSkfL03Np0A7GxWzBnKvQTOdkwavo3MSfiRwyn
ZnqMurLuRNQ/K0zcvxN+F1yflDF15R28p7yxw4vJN7AbMuQ0bRQgbZEThhm8IqCFEfigqHiCy+nW
mlcioURAeH46FBAVuENh9gLykv8+ELT5taIiSgiZlAl3TyxONZcflvFotr49oP5dM1LOrLydpe8b
yt6yPyyefVzboEH2kV2uUMdF99q2lZwfgLgH+bHw/qnuUAuR/NebycYSK7sVteihHAvhiWMgRA6i
GO5O5OXCES77sR+VaFMBX1KFDzZvnbGSrlh+RfxGe3ITATXElyhg96WM1PSZ0Qg7Y7/FJfUg/KuN
wup4jUNw5v05g6Bw05Rgnho0oQPmgDIwqVJaMgy9Si+ZnaxV9Bb3ysv7IbnE/uyPgZcT3Man26wb
wR8Uas9yo9t748W2pxVFBYunA0X2r+2FcurzUx0FAwRim34P9nXDz158fhxTFjOyNEigEq9Rfp6C
qqJiwIX0LoJDEE7V/p1r5AmZLXtJnKdEB13BUi0/wIlHJjb1v6gHgxWBd9GqUtH7nQcKWb+QRKz/
ld5WSf++o2WvturL+B+RMBHg80RevvmlSTyzpEhCZCcHBS/lo95BaHOQe+pfPVprBXwqY5JzvypA
/uDttui/u1JYO61dxtj3RVlE942JfXcZyGzG74tY5dYsiNIn1i30Wg9Lmz+0kPPIt52s6Cy2q6z4
yxqfE1Pqe589j6T04eCg0gXnvSVLpS87JtOSoerp1mus+tGIjRrqkYRtYZuiBx9lU+7NV/DV2Wrj
OBtywuLXn0a9YhL6wfZ85bCIETSztfwmVs9YMDcjE07cLaSTnYK70MLhxAJYyTC9sCZPyRJg75Tn
cQYubMf/KwffCWEGl+e12TqAXhjYV4a03nnhZQPydfK6DU0JggG4BDzKSSR+0nSmxpMZDllKaVbV
RIkdHxdtovSz5cJ+8OSxluTimRXQkfLg+Xm3M7O91NE+jcMUFsAen/EmJAm6HAdqCN2nu0BJ/lcg
GEi6EcUvq39RTh79MjHjy6ljYmij1Zb2tzNolXSvmiRKmutftyK/FKP2I6292zIMp0URlSpOVmgD
rrRQ/X3Ni/JFHk7G3GX6+5piZV2aesvOqfC1MbJ4LJTnzP/r+9WP96f1MfSYEpzGeHn5EzzprrYu
vq2gOVL2SSiJ45ty5rg0Jxo9/BxbdzKJAnssyjrjjM4BVzmL+e442wuGRzX+pZ8gYixrtvRFctXj
fnODMJB1Ge2yX7LzBc4TGnFYkHVStFlx4rL3drwT4UOPiDK3K2eCGXcPU1h1NCtTwxq3r7993zcY
hw1CUhjCSdUBG0e7/Vk5da/aFtESmbnmfX8fu/5yg8U/6o41XKtZ0KGIF2G9XapCn84Q3/hsUjeL
PIGzo749Qu6IwnlUbTUC6aU2vXLJNRD13gHWlswc8N5K6Sxb+TEDPefkGG+myWej4LpfIdPyg00g
TJ2CgNWQpTAIqrGACPb6AbAc7cRVUvjLMTM73tQSIVz62NXfShiI8pslI0FUjnN+jT2tX+mwHVvV
cqemOPq7y2n1GWRS4YlLJzE2BMU60wR8wblKoFGplsvkdvzZ+z5sX70dHBfJUISPQoyhc4IR4/jn
z3/dj9/QHPPPw9DNSDyMKtgATKuvSbj23bE0nytrrQsYpU1GFVO0i8TZ/UNtuaEO+6gR9ejQM38Q
kWINJdI88b3H2bki1hPHt/Fizt83Cz9naIORmI7BU6QryWjwabLA9IYDMpwH6th+ff4IVblyOF2Q
dIC3+ez64ki1ZBkw5vdr8egTlXrxo1/Cm2r0cBysg8geQfRRV14c5gfkyWfhcJdjqbFZVGJ2nDvD
Z0Y1ylSJhYIvmt038jdiItjGizAS+d3UtCqWR1j5Kx0j8fWf/RLLGVMO1uGdmoUTM2gBPWXqjOcl
Ed3jiJ83Cs8KulrrhwxhlQB9l8m/ajutZ/JP1dwBCWQR/LrtIwb+7/C32Z9JtbdNeIqfLECH4Y3U
3jmtaJM2hqQJ5wCvlKzBT1pa0XG8L+lWxEe1aEBOZG+Ozt7WBW/viEdOJlG5QyglyGEaEna4Or47
ZFAXjn9+k/CkEdIyMxQWfHmaNkA3Uo0YjQDaRGOIt5Uhv1wifdblyuOglYBypQB9IUsC2VOdlW6I
jw10FReFw549MYbjIIY5yzb4UIR5I3NNbeChyO5YS6L3XujSVd4NoijCZQRJl1OlMswEOHNanuzK
JV74UnFr6QUSCnYU7MANapm4dtnF+EEm/wP8PygBSMeh+yJtHuacxXgIq1SuvyJfQYr4ZBXkdc5l
6onrV1Hy1+tAKBnlTo973OoVv8pmyGG/0H848OJRQ+wldd+6jRQo3/M/xMnZnUFArgfobMBruSzC
FfQhQ0ejJLSh+3zwZzbrqVc6ti9mmZDsExpHSzV/TJALbAC5SC0EQkXWEbyZjALuEU9dNUpFp6V5
CCPLUFf7APjGx4Q1SvxOGs8y5F681QBfz5J8EFjSE/q8M3Hn1JyWnXpwb0P4BQ06EddhvFp1vhHe
Am5TwPkMMlcID+uD+WYZwe7OKd0XnwP7iUJJO4Njvp8iBO45XVTE/7jy48fPEpVZetwM0YU/DMjB
tmU3AgR2NxKUIfPN99B5K1hf2lE5UZwiLY41b8SZEgGKf7u3rXj/a/JlMzhvnXSo/4iDxJK2SOst
3qwZIhGWvvlfDxoCCz7v8tfp0OYyZUFqTXpQ+/1TEiH0BmWPTWAxy3BsiF9an7fUSWgw4/MmgMe7
QO7DwOJdeJ1RLHLYEOXqJayimbrpRa3aDVVHvBMgFkf6hqMd1F79SngtoO1nDp6OKZcg3XnlRtsb
hb4toeta4PMM/PrKwSlUnGOtS9BY34iEzvGhs+yex1TRMc12SnchOb2pXZk4Jq+88QYigft87K7C
ddfJ63KVEN1eQO+6TP/uqbr9xJs8u7NG/fa3efFFz0wed17jMjetAA2CUiBc1uo/K/PTaY+DF7+E
JEyO29apAGTabdNWI+nGKz+zWBjyWLXgm+en3UEFwSyyl0jcJTUFzwVEL6sOITNBex24cMZwg1Ve
EB4MAc+Xx/Uqi4Ck5aIZoFhXh3iE7Tr4loLPZ/iHa1GH6mVDv0L+Vl4xF3esaBHSeYPuLI92mfjj
/7/HJpZdRzcDMkAD8WMVN1U1l6qRBo75ocMfKrsc6gCVANJT4LIvvCRKYFX3bESfBuXu4L7AG5D+
UMvC64rseMYkSc1YY7YTKwXaUQ8Ac74UJfcxKdWsMKPn/mQ/F7KGa83H0Drm/cpKVfPhGmVbSAHp
wpLGvnysfMGt6JiigXsnrOcepz+CGcIp3NihzIUvz65J7JEUBYcWm+Xi6WpvQDQxSEzM/XteiszF
ycAUJKIHOzjgh6iMAF5XfyHCUDA54rg5QXg9uy2eoa+y2KZqGLegCyTEnHlfDWD58A6v1kmrJdW3
zi+2AVR5fK/hy/lBuFqWkbQTFv+0ttZXJk/9gQQIYidbPcb3D2rqFgySSLDnxErVohODx+PzjNqC
/VnXpR6e3LI1JP+tCnn/OxZrBLGEchlN1RNSW9YL5GIKfbp8vuZaxAKw0diByibTosEn3cVthNaG
5TM+eosTcZHHiv6SM1P7OF2bPoV06HBo6y9T6+B2CzqgIIK1Lrm9vXC6i5Uu2CCkjh/DEI//edj/
lcA/ULRazxAuU7l6x7qPRstBXJNWgPv/0Fn/0aODvzlbE3A00ayZvTQgWFjOx8gR9okoT7psmbkq
kQJiUxIy+00rYO6n+tp0nEKSWPpWZeSSEr6wSKOa5y9utBiPsfopGHMgLsTU1ArzuZ2ZPm7ybO1l
DJjpOUIhR0D1IVNU7oQ25OM+jQbmHKoBoKh+1VvxKlsRUNsl6wFJ4DCsBTfp09HqKy6cH8y+6InX
WquEJqmX/Huj9wUEH5kqVqudYpOlX0cAk9ehH5W0/RJ/gxObA8iGuEawDemX4r8iPg8J91aHVr3q
AMKXGoZAT7or27FySTAyvVxjCrLUai/alK/O1pkglySk0WWOr7KZ4X1jUZq4WtzjljNyttym2tC8
dWBy3RdgQLE/PVy9rEOX0u9mxOYTAdu08zHn7sEvtyWCttrk8hiPlgILWw6tjC0pU/KiE3rDH9Ha
zkVKp4fP9JLacM3RNzq/68iwWsGmLdD8UFNHyJltHk2oaqqjPoT5FwrYuWZwvyCKFQQfNeHHd3lf
WQmRM3bBoh0wAoVKUex/8Y8Bl1z4CEkBJqEAj7zAZAF6erB1bTGa/YHP3t8MkbzpxuEYk0Bzwo7U
59M/BqYXJDIF/1rvfeZXyMflxIsYP0IgZ03mwJTC0Ut8HZXg/ekBXPLDGD2EnEdxD/KGPBDlr+uQ
BLBgMy9u+6RX5SSC4gbL78bFWH8BF1SdghExca1yVWY57Fz8c3gtLF1iX16+Ep3TwAtuB7mDI2fm
QmJb0UrzzZjflHbaFZraSnRE/xywvxPtcXDwYwiGBEyswdJuHmXQ2JOvuMBfOj01C/H9EAdetcvz
gDgChlm1x5qi5FfeEy4t/9tiEt+tqma3MANAbzUerZmqI5ySKsuaSgM4eni6yeuP9HQ5TTyH7fv0
2ymuG53+LIllklSqKmQjPURI/DBlQLFj35xoMMrUAgKkmoDHsul6dzJUXYy64lFMqyU4o6AMMOIl
netgF4MGn54spFzc6+3FHfCBEg7EfHfj0r/G9Mr/APVMa84XpN+Gv+51s3RGjPKW/nYKoZqKP3ak
0IPdCC6HnnRVTUCC8PXzoNKaPXr3yRKXc1A76gIfu47MiA0yk4rYg+1+KQHhL/OGArbEC/ITq063
TUHGTTMIzEDzg0zdl2nUuSLn9vaqa+d7qUc56EPlQmB/mTsRgyZLJT6IhLrjyB0qBkc0kIwA6B9U
ESW1xJFrLfrHZbK1fWsciaOoiJITLhJt/rg1bg9C5MYG97jc+7iDz/dS2Ek4g6HjKIeVCa+uByDc
FpuDqghuus4Xk7XICHNVFn4jHvVo7fZJ+rXNUHzgNqJCxfAFAc3nK1RcXKCnL+eszu9h5Udqk1eO
t4sI/LNOcyYXblzE+pD4OzpHrMusT3OSVob6H6l9ZPC97c7jW5sJjrji9yqFBySeIf8eUUSrgcus
4vmSrhYskVH3Fys4ak1SsqZ63AjDCydbZlRRV0xZxTpQX8lSdhSJsLz3kQCvibrLk07xWwmnGCCL
LPECZlG1ihiVUfEFy0L2bzWTaVmMK+MMIYYlYs7xKQqizMoHPR5CYnYzD7wzyJNfzdcaBDDUHQ+T
tQVGfNnOtaQbkXOYQf6PbLgZtM8n7k2H/s+ekev/D1m5jY31dnUcj9+WAP1DujTG6gv87UsG6KIx
duNgZsPj/9y0VGCP25eblP6cc9JQBjgYKJdGratXVVKPTr2q6zJ900u2Evk1QCXE160ROmCdDU1R
Wgkrt0OBz2rN6Q6o8Ea0sicHtBr72DezPgS5GaD5GPxfLCczKyCFdSdRqfHgMOJRCunmKGfhRNtJ
DhHr49cAnWLQqx8OfQNvidOVzvRKnqRWf3bCCfA99MGuVhwFrjNM2+O6nTwJOkX1rZ/Gi51yWP0t
ZEn14zWeA74taY2LA1f8kIvyABgZmHD0T9iTRYi9OB9xHHZqO2lj2Hti6bpWxrdb38GfFNCGHkhE
7J5nS2jQo2Np7jEuOJc+2FMhfig7I5sBhSAAlEJ39JJkFouvmx5abVPv+MqdSZG6poCXpo7AN1Tb
zQOwTsNNKdDTjUASLaETKOBNdKq3iRjgFh65e9YADEX45/JES8DvYsJ2LLgC67xWbfUa3pxnmPe5
9w0JKpFQoPSZQBfpCBjxTpUE6RY1h4owTOEaVFwIsaDuoteiErbxFnZPg1/r2OMc22Yz9VmxV8xG
hqBkZGedh4+VxrpaHJKzXzH4f1aWx4wl5uGD9M+xKPdmf+ZXVdQNK83ucq87ZQpMcqgf8LWdERZ2
ODVyngRJZLscO18T5PKiff7PcqPDFj5nO31FaKaDjrnvAh8Ab5O2z75zWbghHPo0xNGvB5vRF9zB
tlBnc49kKwIBWRzdcYxIWNHDIKktcfsn4+nGITl+xUcB2dO+JxZUxDqkA4m2Uh+bjQFt8TEcDjzy
4CxtnB0TB3V8xcUUDYbifS60426+94ZuKjUFYpyWeChLBmutPdp/v44zKqdKXvoPwQOkDryiX+FN
ihJXR05dg3wGtUYxPreaBV1HiXpfITvHKIY/G/xy+zQP2yBdqUVt24cUZlO3S5lCBnMAJ6OxFD1e
vsls+kg74sNhib0ZdRKPqeifVou1EYadfDVRDJ3pyTyGfT0mCc6f+EoX2vjm8NAKwclYQSXwfQyG
3ZvATB71TC/usW6TFuTujdSd6aQoy4ppu41EtSilSKjXEVv4IRK69ZznqXZHB3fxMBHbjKpb0bDk
Ro4tGe5tcLaDMlJmYww2dqya5NtoUzCyEHe3ECZb5A0oYwuujPJ66hqg7Qtb63QoPGelbSRRr9sc
1rccOxNoePlZRYxeJA8PzZpkV+ePQvYGmwPr4QkiUlRphiQ5ihKIUgn/H6nhbHbgHiI4tvr7SaB2
LTH7kMy5WXrUIiqp92JiE4XZV7rIO2rCMiE2jy4tjWlPYl8JXTSrBFt/mbBmGa+pH9aUL2Qw4pBs
Ad3LaUjNU9JpNfs6VSpZRxGj7XTu1KsEhAZwdDdoNnzp42w/SnnuHnXrj7P/0VhD40d7SS5QO3sf
Jhiu6kK4BzYhBQJ2Lrm/Zzq3Eph3TyboDc4cm2udhP3zj+0zH0gzsg2g2kSVIdPXQSXOaEM40E7I
7I7pkHHVW0ky4JJKjPzFxvP/rZ1M9OT8izmLooidy9KNq3QKkZOR7IIawrTRgghA6JjgT9d4dNz3
UyKHPwLzWt7vZzpp5l1Gruwmobu2cwn+27QWqrXQ0oo+ArDKe7kULeNsO0KBBy3XAWxOBK9OeoJ2
SC450wsXjZwgW8MuGHZcMdRlZhxx58Z3OkXhUXNZpfpIcWRI6aO/4AAUDYzSUo9bY2mYT2dB3e5M
oVPoOXvyVANAxwEw8HSjtsPcZaIPrUV3GbV5Q5iiwF0gtiGV/HgRZ05xTZdFYjs9u09YnHKHylAc
m6chNkGU48HsvQ+/6jE8GLZYg2tdACDiSCvAkO1kU+niQUSP27ydaeegCbGS7xTaozLKA4gIfniN
eXTdeA4KIEoJ2wOuob2n6pr0yXhB43dofQkVaw7cWSBSsEtnOIJySy5hbndQIJ/ptoH65gkCwgaH
IfUVb8WC4FQwgCG0ZMrHaZvx0I4kwUKCKC3XH89wVXWUzRprOEZlDre6+M13odqHYZ9BkGTHw7TQ
qzu8TO+ze6PB+07dcXziekHxHFZ7dkurNaH5z9XAHKoo9oFB0M9MAqkjlYeQd8MH/59q/W3Hcg6D
DV8k+kq9pM4zyLedhKd0heDkWvUiAyabefxXAIRpBML6fXTQ4DTR6tzEyQiMLXVNvzcGRNqnSddf
OekpYnHyMhXBh5o52N/tAootD3Zp8V9bD0WOXGcz1ZxgKyZwMwc0iaoeQXULtUjSFmDpPHfPXSjW
aGoTcsP5BafeE5cHGn5UMq/nLn+7M0ia9kREVgpgOqJiVckM0zddvLAc3mTmTsH+xI/MOfLtfP/d
W4Ug0GbILhj+KfyGpxtuxX+swnlQXUCTR8AE02AZ0m6hAL7GdUUp0GEsqQKSdG34hgMkUcO0wN8N
3w69OIt/ph/LQKV3UYNtRs87Npymo6csxle7rZRDsMG+hNxDwWwlbDllcbCTNXw/IXPoSxhwOZCs
haipqfV5UUEwzGsxJ3gUaGQfiEdCOZ4mwUr3uJ82VBOevX4ywLKYxsqQz9cGrc+MICGqeB43pirk
ox0Il8UudRvsU8P+A6PV5OMAJWg03XBM4YZJU7IeL6cI9Ws3lAeTnGkwXk58/qayDzssJrzExzuD
g4vVGeBp8x0gP5ot5Y1usafHBDiEGeIQOX+nYUhFD6OO1Znr9f6/z4UdIFd7AiBRXzezxMpsLcUD
AhiIE7JR5jBXm5vbZR/8zF1Tgl1tBMmnRJqsgjMrX+vu2bJgtN1z7JNP/Clb20YEXyaIPGpi9MsO
9HJ1tjwK8yD9UfQlBr/YZpC58nCNRqt7/tm+G3IiWhp/aCQCVnP7MrlQPUl5E2d+Jah6EoFousPt
T79/SsSAYYtpMqIregNZUqn28okIsVwgDDdIt32aF7qcmbUQkirU4rIKtELY3cfiXB8TD80OjsRv
TnFB69XV+K+tT7rcM+GZj6e8cpBMSX+gyw7RawV8Vu23fJIOgBS4fI/27FI4giCcM/TIQkPhIYfL
wWRnWh8Lpv/G49ZreTZdnh1cw61TAn3oGrDfpHVv0MMoYq5/lOPhzp94qM3dprp9XmXvyF+jenIv
/p2PA4u3ZljzVElJqbXiDfmgZPbq2YJi/MslxlxKFYNxBMm3fMYYG4L0NGvvzKyOMUR355QMnFW0
2qxBC3vdoRhBETMhh6j+uczX8UeMLkIWFx3HzR6vZMnjzrybqIJmZvIJnH8btI5DdJSFLAR7W//J
FXBAkVejNFaKsbXyvrlqJ9p2az3B/zgOtasNufQzCj4TS2bfCP0yRroBE5d3XYbvHk7UwtWgY5zQ
2VLIH+eWunmE63IX5xsTvs86mVKVFGGs4YVD9zuQy7kmpP/lPYcOINqIIctsp38s8PHUuteUv0+W
DIMw0G33vBCZUXeeqXm3C2mb2en+4CFVLBuzAdSisC3sgkTL+5iC0MQ7MpT/sw3kV7wvS6x9nH/G
nc+HCQHOMSG3smsQcw2AODIEQKe0NX9INhU8jPOevowTO5gN4ODyTYDeR+0BmJRSjp2WTWPIS2bZ
QEkoXvvgCSey8oJ++ncDHcx2lys7Ju7NaxCbnb8x1p0ZWZN/m4c0XSvcicyFHnJXbB0eSybFBlB4
T8oMieeM5OlYofNnXXFFEYPhg3EOwBTkSnVhiFOMQp4x+E4HJhe0+r6iEOTgBHO5j+NiC2xXJgG8
BNNXIwOtLfv9YkK/GsJG9FgmAnLDCxPEtgzFOTPPQy3KBFq/tboGSQUXep+Gsn8JcM/b3Q5J5SlW
VRB67pWc2pVXMdP/szmCSidnseAp9N9wVv4d5Tg/aVPWZASxOIufb15r+naz7st5Ge+LgEPWSdK8
IU4CHK9+f/jdm358sMwnVkIMlqQXxhG/mSvCHGQ5VBk6TU2uMhUp2qnp2QU7AB8jDEd8EF3fW0vH
+20VA4vONtwG0FBiOTBJL1g2ROga4AOSA13a3FdTK9GjmwgOCfWy6tiZ87KwbrpIdQ+cS6clGADy
lejvU6493QumJmhzL5RFMOm7GCyyfvspj3EW3lS4i6IuXv5rL4jFVHplFj8Yi+BEScyB8AsZ3znW
6X1adGj6qn/xWPYFHt3/AmlOzJHV8iv+poxaGb2nPm2Iwmev2kqg79ZYSDU+B9F6MCCtDs3rF10A
EL5RjrbRVPxywzDLl1hcQ5+5DyjjzwRoQnhacDGzMOyP+gpMsLIi8XjmF0gAsQCT6doWQvUsfuL9
H+hVq9lOvUUlG1aHp4AK9+b6yr2PDdru3bkNHKWB7xINXMAnXdXiH96DOLnLJN60g31eXPn9Sl2N
8JsImPy2yeSBlL0E4zMtimUlt43YJhjWrrVoxfV+AEU6JWLTTuI3KVsQg5nkT086SNijj6gLDhyi
Tyk96cEngmcqov2GMHo6dAph63OLNHi4Wtg70ouxTyfXm7jg16+KTTfoRqPTbXkRw/VvjGtRl3M3
NnUPfjncUrw74ubfCo/W+wCIe1Hgvdoq+G+891z09k3K2xX5VT5874r7XHDY5XBz7hKnrLw+0cyf
txdZgXyUjasrG61RfUDDb9fAvbecXChThMo79gsaBlXECgQINFoHtmVitQ3UUjmUc8VWDtxkW+bo
fWPDIp4CSOsTjK55GC7asNkioUih/TpAjM2RInbuvcwdr1ZFQnZTmDrvVbO/yM8tqsS2pTBb1cAG
nio6HJDDZX4HqyuDWKf+G8JWc3jVhGJ6uEhKDW3aMOnxXDS5zWrx0fCAJGzxQwdRV9CadaH25LIf
VpbZMtB6f7TTs2jjo9fdSdNe0FLyAImuYGPhhSOFp0ehGa9wqdWLKRC1jdg0+wXYlDEPY0SYmQ1d
izeJuvemXITruilAE0qhlmXtOEA3zTccS1Aw1sWeKcK4bsyD0bla0IMWSK/qmPVWCOZh8xckDYiM
g3XzcmhN5Fv/ibXe9UtkBKOYals5YVeKl50UyCCRf2OPnrdip3joxglp5s4A9V2Wx+JjEc1u7akY
ga9p33OYsb7qwGAHxw/+5hKGaWM947e7CuRerU5NMLS9b7iMHVqLNQcuKIxSS5wLAiyJRjnX7oMz
Yqs93c/8m8JwFLIRI4ds5nwBypXPQxpn4Fzf7vtGDaZdJemkoYskS3a2elxHlwhhVV7EaQMKPxkZ
BFakkxBOnCz6ICCqDS4r9hZaO4/6srIaK+Foo5Puc9ppOJEL6JL39/7ZqZTtd5vFFuvwP7srPCeX
0XLel3NXxsLZWeSdYJz4zmmOcVDjShBQpYxtPOnuPxkpfH3BFRzuAJsK1gZ38WxWLFZKL20+Gv4y
2RXLxSyzrOP8H00m3lH9mwsNexOnMweJ/90jXWw/0cMgP0x/so9QVhwItYxoArdFDLqULHrYQlP6
F2qtgbmLwY5TWZ27N3mdvfxR9UysdS5ZTftM9P00tweVphHSMM4h+wosx3jOJoUVSRpk28fnYnr3
/8PaoD+6XFXldFGpZ5N4yQhEIBi9qJB8bTzhC4cpgtmccPsHmGMMyCkJic46OR5Xd3LCBR3lnzXh
nfrOvCh/FLxZTMr/EW2rAqIgrNk9ouAvvV68U0vo9MM6WlV5Ti4dLlt2BYdhbUwlMZHtwsEaEV9S
c7A833EaBUyfeHyhYL71GmE392HKyDmBOyYTbFHxsf54MOk01uTZjjS+wb+b2zt/vCPYWILuba/b
weeTe3FPSN29Fe+j+KPOo/8kJM8t9dDcDO3n2b7hKw0YwewimtOSnucQyfhkKTh7cn6jzHwECiI5
32Y9OQl2bIzIuXrz5xv3EeTDfxVdaak9TlL3FNgjjRppjT/vSVG6JmaPmwT+P0HLwG4ZuHg02aJh
y9CIdNwzIoz/OiurL05pwPjcwqAIauY9DoO53fnTPBSOpbk8yxOCqfzpcDqgE645R47vi/cWtu8Z
qFQV7oJ220CfTjhjM2CgGXerwc5MLs2sldI+hZeZxlnCTrgLVVJaNBFWXu4eVrDh1N530EEW3mQS
AbDDjTg8xOhoMg+9KtU2enVKe8/dc102IHE5yvKIS2V/Mn5acWeaew3drXHMlZ5A329PYoGfFwju
vcJbJokoxkmVhASvOw8OF9zlUBQuWSHA5XI9tfqwWRkyhC99EgwYxSjzsp34B3LWXflM258QVazA
wekg05nJhtK1g6zx/y9ePwXeER4SlYwuZLIb6fiE+AFGGERCFHm/4AaReTPTKHG79PliIvD9jv16
LapGA/NeHoY9bis1TjExj6RP+IzBOQPCzTKaXr81sVGw/xjXSU9EXddJF52Aa/6gOfkbPugf9Rut
Vj/zeAVoX9DbaAI7DTm5dzdIV8vBCToLyZGCKwAz5TD0Gi0JDqjVijAe/yDiRJfAQKfR66NC2ZUL
/HroMAt2iv6Xrpa1DBKTmkVU66xFB7Z3jhUZReF/zxw8Zmm5HCMFKCsrtQI0uF35xiWo/mzzQtEC
UQ5pBgFYspH9FXebPtRFGeLav8SgRra8xETc3FGqbE2O5mgPpOhtJEehoGUYCwGOTZ/VvF13Z47P
QC1aPNJFlXl7zN4H6sxRA75faXLmAT8PCDDTKd4anYdFL3Oa89HJOJc7GYaRRJ3HipGvfEd+yENs
3pyuIpfTNMsN4RIImrGdSbEE4qXEFNp5vIYS3rUeff5hT0ITm0auMCrb45admLQWdJvhRBok4YYx
SAt+jrxDvRwWBvbaYDalh/k96p8//Hok1Z1mU4D4NdpOOHCRHrm68pUNnECDJt5MvTjr/wHyVjWy
12IM1pdducuizhZRUhdUCJbDxNWfoHkpJXnuOaREG0vQJlzY6Exkf1n0V2ZvKP6DBiPR3nF6Fbjb
vYy3wC7xDkvj9ctQsCVQL37PlVT//+ksW21QuTXKr+qi77Xasx2teDy9oU6vznj8Dk8TXepF6hJ0
KHBP8wZa5YuLupe4yUl2o2jPbnOwSLnnIsxAge+0PE5p/yDSYQnOpXOsX4JkH50+t/z+SckSzRId
SXthya55PKYKjD3eBI702q4yvdVMnmOIX3KzgGC01AQxT3tB+oD4vol+Q+fmmJ8YNVXBRN64FuqB
bdCw0fH6wludDwWqpfOQWpyfmvbKd1V9Hhi3s5iPVVAwLdubagmS3ldJUHLmF89z/xVGCG3al3x4
dNqJUCkVog03jCIts+l4XRrBCuq7lll9vo5VrmKYFitDk0mapi632GAbmdGFYWRSXcicGoudzj0p
E6jvZfxJ+hlMsI2HJPmtWQIeJBBrmqIFUCauQMJtItGcqaaGfebJHqkndKr8R0WNyKnW8eW6k39W
iyKumq2luZAvBb8B4O+0ix20v8Q3JZUjV6zXhaUPHOxrYsKpgGwL7T2VIAOgNeE3oJ7hJnL8We0m
PPJvaABp46QV+O72bWFtlc8xTIfEkVPljMw1dMOCWv9+eWLzdruS3HWnia2tXhk2Id2CaRr9TNBW
U+KlmysBM7eBflIxaAJ5ZaIkwrA+NcXOX1hI9AQh3eANUcfaxcXkfZClLKvKiEjQUIJ2IwjxwXbW
Th5LXGgz1UabX0ACh0M7bj2Jl7HmR8yULWa534Pz+D2Qqy1YJotpWRt99wkEBnWuGyPFzHFumVIr
fNXiAJ5x48O0Mx4Z9jPNvQPpbV05aMs/UxU0z8/jegsQTzVKB9mt+MZhq+9p33n8ETp9D3F82Pkv
3o5PkV71PXpMr3K4PE6tvOQHsTWBiR8An/XTAOgFD9oxbwOTxOA1SZW58de4CZRdp4WeeQIsq8ql
sB0/kD6xU6ELXDJ8qDuAYVwDdOGM/jloPsoNZsQRDLO4iS93g5Ye+FfRGmnu1eP5wVXwJcHx9G4q
ndbczWo/SPWbQ0L2xuRFd0Z2rWES3tF7GzJmZI+mQDvNrifIoOqetXK4fKWhRpPQF0gswNtXWWKR
hsKCL76j9cukfVojOePcDPbfPT13SVW8Ceyu0ouK8FDP6i2F+uWr7tNN4YFGZrg/ZKUxbPcGjpOy
J31EjvvdTIvXqLiPCXme0wbUzp4OLS+/ZyGF0bfwrgCOV35e84xQwcvz2gsucKTF1qpKsJ0JER+C
isR8YgBqobNoI55NyXA4J+Sb6rWjsgwssM5cK+5d6DZ9wFdnioGZezUaMagyWJ8HcTeTUlo0ivrg
MjRGCeee4xE4qvcFky8W2PiARPQhRHIVkm+HrnvBG2Ek/k8C9BPMda02ozr8LqIEfePIAkVH42qD
9HCmaxYD1FEmI6RAFN6/1oNvzhAIWKHA1QVb+lriV1QKSI3lvFs8XOitv5uZ09vGDO6E9j+cc7B3
Zv2fL1VWyqinuAuWQLr8XyVeIiZRCtMaYX6xA8bsL1KxiOZi53Cjsqbh8lh8mvKc6KKmAa0YLa/c
8xWQsNyRFMAos00HvR8H8lBgMSSn4OqQInvDFisO0KcBDRVv8UZm2U5J5FP96hocQCfjziPWyOOb
opE7TttlXA2bFf33m0YMr4P8Qu7fikEDgkdrERZUMoGmshgkjQy9arLCR9vcNUSI5CgnZ+orjpOH
iKrksFBmQSGiPMZdYlNiMlW/Y164Uq9DFnyv5ujsW1I+pYaeloTDOjVBkEd5XrP2SUhYx0Xjbnpg
/q9oElZ/psxEUmISxLGYSXs525FrqKI0fUmIjoQQF/1nJZy/kr94y/felkslQpJtPleHTohld+m3
1HMb1ZmgzS1LR2IFBO9GO5QOveDCDN10WwbtmCHsn+8tcklAusCP8vpbg/ajPAZV+Rca7uwe4lhD
AMtIVNWTK27i2K9Bfdro39QfJxGKRhMHao6rlAn+c+nOQXkiXNyK6e47VuSQ6JaaPRE0o7HziOL/
mb82ChxjlzrfRwDgKb+fqVNYt0+QcavW9xpOEhoFexGKqdBJPuUtYOFML+9BzD026+9Cx/Yz9Swd
76Yj5QKfiisywRaaUaFsmlunM26fP0LdPVhPUBwiMHx+aeFbF1Xotv08Y81Ue+WBalFdr9wpbF1K
FGY7vZ8wFR24KMQXCXyX0GzMKdfHhPlAp+JRp3lsjzf9KtEuR/86/hdwzTSD4NvJ5oSoT/WPR6Sj
/uN/s+n9j4/sIhqMaUBOZACfMp/3JOahPia+8wIkosIc/BEYN4vkGJH2Lh/0y7RFSFwnHNiDFCil
9o1J5PjWMMM6HIzAUzDOVUatXphpb4v4YOXNokMdc8FxkaNXivUZSmVeenSHdQwfvBTvcEs/0A/w
fT8YCoSGGjYCSTBPnEHj6t54QbFMnLLTjnAAYRUMKzxykHCkhhMLOn66VcDbVkKamioqcMs7Xcih
DrQH5RQ5twaQZeB7ShLF27LvWzGmHglNHlx+ejkD+ER9lV8Nv6ZVfSxkH5C7HUQNhjYYSYvAZFTt
NwFUHEn0JdYlc1D1IfG/cG7yJfhBg34QKADafK+W9QvUqgaWFhNAW/rq8Ht66SQShflBRIFX/J17
Jv/J94gNnUdxzUvOLV5peLqQ/EIm67hUJ2BmE0kdRXGz7OHdXd1v83JqOu4IRbmN2sdOdL9YudNf
eeN3NJ3ya/1l4E48kD+3zpjcC6eH+a7EOoaRoYRHZqd8Uigm5Y5Y4K6AkRCIWVlv2pyyGxEuNNyJ
YlJ+MkQh+KLz/ROqPmVj/64xL31OOGuLT5/3kEgqmAX2BnSXNQ4raCqwTX9BQHDuLaRsoV8nQR7B
DmBiuDrXDhvsB5WOKGfULQ0eWbSz5kx+NnqO+vRB7z4S7rFwZc4D7vrSn+HfqtxJHWzK0CZwDKW6
jHD2N7VkUSuPwsPix1FIG3beU/TdbYUria6OFphpWTkBzrQjukYCVogxxI9cWtyOreXa26LE4V3o
oP58OHEKEPsmJMRUHgQWK+pEuzp3evwdxcHeltPYZ/llOak9PsWIT6VD9Z/fHVTnUZQfgfaH1QtJ
a+UgBAe2+3niBOzB5RY41Zb9omwBQCWQoRaeZVPeGS9RZflK2pbz+ARRTuXdkF5t+CG6SrqNifU9
u81YY3Xn9ICH0VGAKvv5zgiet1E5YKAe6ye/hcrSh96RDSB7kZUjfPgMYTgrl/mpxJsOlxYnZo0p
cSeC4hF2k3HnDxKRAX/B3cqK1jFbW6ub5+Fy9ATzh+CzyXOl9ftFwjKiUlOPYIHpDfqKsUt3qRi4
2OCZxyAZpQ4FglXZ4o7oSlgAazpdjidlMJWY6PPzvIlBT1XELWzcoFNXAi6U4SX4at1uTD8oRfBz
af3Bn15AQviKDL9OgA7x9X84c7b/hj7psIouUgjZD6GKyC0qeoTGe9FVJ5MhvVA7t00pRpNA0+6P
gtqpQYLpobOHD5/J898rmgwnKPoverPLm9o2qcLRhOfw8gVHjtrrMtI4iRH1Zjft1I61fQgbmaTo
yhxO8cVz2jqrr+gpzDGto4wtsLd+ZZ7Zxhw4jpMuMONkq+PX0jiSckqywkupjmrizf7huwLjNGOj
UHf6yhqqOkO4nbiuinnEY2Di9DKafHCHxBURL+ib5ziZIi4Ru4t1wKvZw7aKjY55NiZ6HD5yvrz9
JC0yC0y7rBRKN4TPhMksR0zjUplG6I8sbqR/KPPvemeoX/wfkX5S2kKwGVLjEYEYwYwK5rf+SLXz
YNUw5VYbW7dV0jrRwDPIHlaKYkS4Ak04TCyg6YmLU6OWwKOhb0VmPQH+uzAJ6LJAPi63YOkXnuEz
kqEmgWjiw6w/riZPdJY+m8kYlmG+5B4lIPSCHX0NeYm3RDKoJtvcoLrBhFCYYG09F5usZUdhCX2p
wbGUt7RHVr53Zm+YjcqakMg/wnUPp9kiAJdYBm0tM8mcd7eVxkSK9bVfOHPqgwjHe5U3ILCfEKqk
s62pvALtZ0ozD9AfYGyPb4JQzkSwa3tj8Yb4BOj1tkrolaG6qkU1xod5jXguPGQXbxaCuhc4VQL0
gsSKX4T92jijK8B8L9DN0sSNGPBT+iPuEEO4FjcWpYcUgU0MaInQEE+JH0Diss2STd64Ntont0Hn
OODP7+bJxW0kSft3DU6u2PhielMi/GoPIe+iz/CCs8CtK1M6UbgcCrUhV+hU50r3Ne1Zm4KObcas
/f9kspKXy2VDSS48H4/2UQOESoPF3K/eEUAtnAV5vfwE8lJqeKSZjHLs1QbbMbEITDIEHQ/EXN/P
Oq+Y2Pu8uaA/pIrj8CW6I0+zon44d5fwlV1KM9gt0a+sUxTFvwukzibUBqAl5B2h5Kz7V/e+zw+V
xn3MJD22c/ZJTAm+S0RufPIQt6uAlyaXxM4qUSYj9EN/EftTIFqnKoBX+zBi1YWPe8NNCg+fJaQc
KbljHszG4VmhhhG+GwIOubELXzoSbLfd5ZnpUaU0pB40cC+myJyrej+09fYUOel5FsN7L8o5Hxhb
Zds8gx/0eY5pbBldvcV1RyNZwnXlPSVk773ahMwNLLfQBQ2zjft+BP/AIY7x89TedBNZNw6618rW
yL51KCS1uth80vi5H0i8pcGKn997p2gPAM3iaB1hMtLbLudRxEx2zWOD4Q4weHpOdAemm+i6FX3D
Wt3O/DiBTnljmQGQb5X/RSj3S0U6PerfXBGgDk/aVSTeEHzMum9oKgkVj9YIr/1DuSvwq7nQajjp
q2YkP4LI2tWGTuWjpZTF8bZg2997Tfin5CiWtoVIOq5yxdrtf5kcsrU+a8nIPP4Pmjb9WQiv+yXs
in+XEIhCFRWIr4ZO1dzkAoZmNx+nirMY+ikUYXbZJrUPNBSkhjJ0zhEMA4iWzlpkRKkLFvI2qYU4
2lWv/S7Y2q52TJFSbWKtp+k5irFor3t8LUSBrBfCWQD5087m6jqRk0iQcN7c4jaCyYIPD04PDqLK
qdPyx14nbasqt2HTHN8Y0kMj+6UAsbBGC1+VETl8FEDF/P548bNfdbptuU9g39xs5yhM/pU0oLvZ
ZpVMOe4OVIwTcTwivlqI250nY2xi9a6J8e7vGjphYTJNiHR+uDBtSevSt54mRYKcImQdOdwOQlBp
5ePNjBy0FU+ct75FRa9WigQgu8y/F5Tx89MtXEx/nWKmhoU1mIybRLnDjhAq8V3MyWGzZU+d+bNS
b5NebEFpHL32ZGCpT8XqAbMU4Nnr4tXj9r5GKmU2nUAHucp4HMLkSMvy1nqiBWuvH0aoxxetfgvr
1tpMJAdeUOqEXDRo4qNrQuTVLdoNGmATys0LpvzxrNztQrLaM0+c1nG1TdT9llPScXC4FRAaMkvp
E+skKodHZD6WdVjntxizMuNyqu7GUGxsyxT0d5sdyKM+dMnw0HxYqc9lDsPdkN+DLF0UTZXLKD5K
252Zk2/Ln5tPEYR6K2BQCuGZ2kZgRt+NpbUbUu6T1cNwIOA9Ey2xgBvne8VfFIZezN2xJ9kWUy+F
JDO0fu1sHxlD84smqV68CI7PH2olDPVyXXqJDKbSZdCPBsynVUHWT+0Vb5pznvpogjoFiBb8gbej
47nnxteO3ve9Yva+gDR+BM7aJP1kWsOM5Vz4ebmli4NmzA5ken8f9Gj+dlrJohi/mz4FJAWktv6a
3g1LfKu8l0SEsjUvRXs5S/+4KqEbvwOTLhoTVbncHW2jcpdZQUCwAnZmRlMflT8=
`protect end_protected
