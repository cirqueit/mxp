XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g�����J�{���}k�#":=ҟ0��@��λ\ؐ���x5��l`5�~��Ѡ-Q��Н�+����>:��s��L��m��5���Q�{~]�ca	+�Tu�#�'�}NGn�T��X��گ�������2t�P��� �%�(�4u��Ѫ���i���H�A����|��~��H���.N�S�RX]*�<�3me�\C|��|n#(BG踼�]�$�o���s�@j4ˌ�V�7�3�X������x����t��ڼDi�P��03h!'��Q)6��ƪFT�=E�xh�g�h�I�סP����I��	��,@m�J��&��=?"�)��u�K÷��P�����V�n��󝲑���!ހpI"�_�ZnI|}��h�N�4���Y��-��QV�C�ō�.�S�+��M�������0V��fIF���--�&��z|�Gj��	Z��V�ন�:SC�L�]���:+�A��a�xc͏
��Љ���2ވ:�^s����">፹� b�G�ŝ��)QtT���G�bFź@A�k�ُ�ApPf���5��4�&��R�lΎu�W�L527��@p���>Th��r����A"��vL��6������l�R�d��|�z�8:��C��6��ī�Y,�1р��CK��kA�����y-�RMn����.� �ʞ4���E
��	ޫ
�}u'�s	a�ȡ2A�$	l��N�D��Վ_�+Gt��M˫l��i�XlxVHYEB     400     1c0��ޚ+#a��l��,��I+V���00��MUJ��a��qUq�ü|���p�voqS���9*H�}9��=	���k�,�'SbR>��|t 
����Ĩ�N�܆���=���40�}.��HL{~�{<��ǲ���$�lS�u�G�~���'l��^�̈L��I�x�*����[����þhD��`q�s88_f�VTl��UŊ��ǘ^W]�9��0�PCar��jʀ���2�Wx!�֫���]46�JX��ڃ�bm��^���erଵVOk��Hd�3���=�����(7�6pf��5A@M�@!�e*?�u�w�S����~�u1����8܂���:�|��~.�� ��++}`�b`�_��A*P�������w�ƛ?�q�v�L�Z��R�_2î����d��U�D4G��^��V�)�Ϗa���XlxVHYEB     400     180+��
�M��Ƙ������w ͚w>�!!Y�g��}�٤�~V�.�P���_���l����`'�=7��uݱ���E��t[���+����m��c暊`�0,�ۉY,�ˡa�O�f��dfν��S��m����J�$��Pcn?�^�<N'�R���]ܶs����|=�2��N&Z�pF�9�%�
y�>ǘ����z@M�~�^$��K=2�!�_�H�W/N2f=O�2lL��0��PF��iYX�c�Ov4�]M-�IP�rO��r�d�d~I�����S���D�J z�ӟ���y�A��S�r�\%νd�tt����.U�_��<���gF���:�r)�O��0;]T�9 �W(�T+���2���P�^����)�XlxVHYEB     400     150:pM��.����6vC�/ �^�z ���5s��z<U/Jo0	x_���b� �W��r���K#.�/�Kȉ�p���v7�n�O-ah#L�n�m����1u&�mK,��&X��Rr���Xc�DN�Y2A�K��\e�@���ۘ�'n��%ynD���tr۶�UL��!�x�mϑX�Y�W��ZE��iu)�t/c�j���+�0�ݭ�>�V��p�M�2�R��'b4x#���F����=.|2#��QUL,ޢV�=_@~�P��f�%�M�S9�a�'@0oJD����v�z@�*��i-�Z,���k"�p�0�����M��·�pՆ(Gū1)XXlxVHYEB     400     1b0��%Q!�}��{�cv\j�sLc��Z.�K�W��4�K
>[�͢�4����?e����5���>и��5޷�%���;2���:ix\_%��g�4�L,ML�`?`�/���Q!�8��Ln��s.a�
;�ud�Y������ʆÍ�ӻ,�f��\�
9'6��B��r���?f�z�Ѱ����Y$^_�2��s���(�|A@����i��R��)��,�͔�ϵ���Ys$�G�A��O�s8,|j6����wxC���p�^��2�K�7:�k�[��'V�Xp�+� ):��ےz�#��M���m!�!��;TC
T�x����E�G&P��̇
�r��=���~�i#]-������AMt��m���C� B��=�*���:z����
d%�n���~��A���s&o�Q-&ZL3mm���eUXlxVHYEB     400     100���G
{��q���c&�cʉ"��HU"��W|����L�R�A<��,�����g&���eU�@��3q�u�5i�$2�����'� �c���s�4&x��m��ZD��L�NSa�8�kCP�tװܓ$<�	�D��p�&S�`[��/��ݑG'%P��o�G��qӮ����q��6�F�k���{�XӜ�M��tw���zyE ����b��.��M�z\�6;=�?�Y����p�Fܑ4����*G�C���̊�XlxVHYEB     400     120ҦZ7�<[��p�z�,��&�*Kw�c���Ҥ���.)� !y�n�m��;�F%1]kG*kQQ#��WLo�)��ɉ8|d��ZO>�8&*| u��_�$c�)o5�M
�V��������ۢ)�<t��3�m��)�.8C���Z���j�#e=-�D��`G[[�p�q��O��
޼�+É���X�C!������.�`{R>�>�ng�(=(�`j���Јp���t���c"�I�G����k�;A�&d���p��fE�^xze�r35�����>��6���� �XlxVHYEB     400     160�%�İ*RiR�f�˟�j	hP�%<�î
i��Fz��nB��='���!��Z&%^��������zT�>�x�BgAɑ���ɵ)���C�R�(�6G�Y�TK;�'h�\�"��bT��IP�a8�.汻F��f�P���H���1čwb��:�8^{;����+��s�nyF�F�V��M���*�/ Mي�s�E�׫; �?�_��>NT�A~gz��qV�W=��%�����$�]��h��Qƭ�@�.����[��^����C><i=�Z�ݛgS��Y<�r:�Y�(��` #r�c��s���3QКN�8 *�R�?8k��!d�)�l�8V��Ι�NXlxVHYEB     400     110�T�M��SY�é���j�����l�0WrT���i�������36�l���cd�1e�wI����W���f��kh�����krEk�,���o��ʌ�X���9�9�d`��S7[��ZJa����Z���<^Wjo���p�-(O�����R8�Ȥj��,�U�K����8�o�w�Z߾e٩I���'�Wj�BS��^���"|j��v�퀠�5�N�$c���JO'�½dF:F�Ζ�i�|�[��H�n���㧺RXlxVHYEB     400     100�.�t�;��"i�O܅�<#�-�[
���Rl,��+t3i�*F��4Z��oQ�[��Rδ�.U�]��GK��8��h��fV螱.���|���,���ʐ򎌌��(�2�� ��:(�)�.���#a`�M~hy��K@05i
,gܧ=]m�x�o�CUr��ylR5<wo�xșJ�d���0�Ο����p���x�?���1��%]3�%/2�0�3bV�R+~7�^�HK�	�m؃�'O`��[f�xE��XlxVHYEB     400      d0���3��Ɯ�)�&���=��Q����4���(4c�����P����������l��P}�'hndou`�zqռ�*����u��/II	I4Ww���̑�k�Ы�B@q�ߞ���`�o�t�6��P�|���b��������w8��:~+di@C�G������8����T���xaf�������ik�~�����أ�ܾ&�XlxVHYEB     400      d0M3��||%%��H�P۝R��ܾ�|�z�;�q����s.#���<d�3��{�����B$r'n����iJ`N+҄�ݭ��`�B������c_���i��w?en��p,��'YG������k���ówlH��y��`��-�#VJ�K.�G���������3B�7��M��;Q���C���SC/��q��oJXlxVHYEB     400     130aҧ҉�\�'\�� Bl�d���t�V����{�J;����	���+�e���U����l+x��sFyC�ٶ6�$I����:�Ѭv��Y�E�*�Y�ң$�& q̸�{�[�Q�k�H��g���������W}�X��,�z����i�M���9l���CI���+D��h��E�I*f��5$���%�+Kk�ρ���%0�D\l��d�ڬ�y��<u�̅8S�L��y��?���o-�,Az��"����;9D��n���;|N�H�;[qv�@�>�L_�T�tLl^d����XlxVHYEB     400     150�T���������,�LʬFb��|�~�7��Tȃ�:;�;K����pg�Z�>5�+%����uZX�?���a1O�0Hu��B�iH���[�)�iiI�\@��3��R�eY�m�o=f��v�(7��wAh��z&�IKQAZï.ݔ�e��M��ܿ������k���;ĵ	�|0/�	��]�S��l@�>��-�]ㆤ-���\���e�Mᓢ���`�<���>�]�]�kl"�h���XŮ`�0_�~'}hYi�A}��JXO�ԝ�	P��y�b'����]�r)�1N�n5#a7��9�,u�/�-�i{n$��'6�:���v5�XlxVHYEB     400     170@{%��N5־ҳ�tI3�1ZG,�A՗jh ��m)�V�\�;Ϥ��=8ߵ�kP�]��Ő3�hܧ��_��$9��-�����ZV0q�����k�A�T-���h��5��#J���d�8|݁/�7f?*�t��j��Hqw�1�Q;�g����� 3��+?�_��(P�#
�V�iZ/l�$bN��pG�|c$������i�\<BJ%�o���Y1&O�0w�ܤ+a�3�C�;1��=���þf}�K�=Tk�ZC���RQ��3�p�ȿ�z�҈E6�����B'N��+ �[Q�(�C�~v��͵7��G���oe�Pטּg_Ld�t�Q����&h��ߒ;�N37�ٿ����dy����^��oXlxVHYEB     400     190 �������]a,�?a��<�Y��=�u=��k!XH����-ݜ�RHR�M��{ܫ��X��s�!����̔,�"5awg`	t���*��{�r��%�����Ό�~˲��<����Ѱ�8�L�b�|���?��-O9����P6����ڠ��3夼}F&��K5�f�%�\�9*�P�(V��xhw�Ռ��2�}��龕U��J)�ZuU�7�Ww0��\B�NL�(�,�F�����K���)��?ta{9=�J�{�+���h���/MJ�^�l�Ӗ����.Hn�Z�<���^K1({�-F�֧7�]g�}b����t��lI��0JV�Q��#�s��n��F�� l��|n�>�/v�O#���()|�sC��_8ĵ�
Q�}I����@�́XlxVHYEB     400     180��%ň�7�|�ޡ{8�q��4���+�4ō�T�B�*�����0 �tg��hR�7w�>���!%�w��Ϯ�C+�ő�}L62���8�=$��t��a�b�	�N��t�{3$iӸ�� &�Cȍ����LpR+��eMcy<=O�ǅ:/l��s��D��e ك��v��"ċ���$~ٟ���\8L �
�Ty��,���TK��:e�>�F�d+�#Zg�k��Ca��W��ļ�A�I�r������V�d�O�)�ۨ��r��n�5�$�zˆ9Ϙ̣���l�oG��>��$T�6���8V"8~ɿh$|�1�n��Ԏ?���X�us������Mߚp�I�_������rqVߔ�J���u�0D?�|�XlxVHYEB     400     140��s�o@�P�0t�!����t�K�l1�ީ�ɐBS����[�u+��w]*D֕*��@�&��&��c�N�ݾ��Y�8�Tb�a��,�A#���W�A��+�q���[�C��f�Ě�e2$&���֡q#5O� "4������iHD���r<�}z Pe^�9��j-$�tg�u�ȝ���b���]�i��G��)�+B�rY���n��/(�3�_����@�h���\㮀�6�#ٶ����ȝ�yOU4HxN�Q2kz�2�G�dI_��%'�(n��3�xH1��ů7�v��-
�Sm�U{CN]?XlxVHYEB     400     130[���(���V��ˑfڋD�Z���
FjnN�F�4����6��7.3�t��8K����_��7��Ԇ�s�cY�?��j���ɖ�nņv,j�OA�y㩠s nZ�[�Y1,E  d1gS�rs.KG$��_lP���o)J�Y��D�WO�H���u\���EH����yDi�9pKZ�����\��<�Ar��qb��yp=i[�V�p38/G��	�E(s��ri%���W]�RlS�kI��}���3�";n���`��:�-=}���O����.ג��sH�o便yS
�*�W�
XlxVHYEB     400     170e"<�����D�M���{k,G��|)���^�k*�����Kw�d��#u�K�b�?�Y�6�W4�~�|n㾎R�XDig�T�ӑM�A_jঁ×�)?��/�.>5�$ު�N[ϯ�hC�Ѧ���!F��{�nW;�0�MQg��P�w�_R�rhxb�e��_�����.iշb�֘V�D}���ߧ�ÿ��ю�� v ��	bC𶸝z0�T[�rbY�ƿ�V���;ymj�S:��_���#�1���{���z��ts�2�-٨}^R8�ũyr/�Su��E���9غ֒b�b��|�/�U����@�=Ʋf=Q-=Ua3����������6�w�)�c�l�5r]�Ţ�Lp2��XlxVHYEB     400     120vG�%$u�F��ՓP��H���
�r앾�Ěr�4&d6�,�<c%��誗����O8�B���3�H=!��FW<�([����Á0�I�K������Ҙܫ<`���ͩG����|�n�S�
"yR�+�o`��ĻX�(T�R���5h��D`��a��7$�]��jO��7X�E�ļ#uC[L
nAt�����'V���Wk ���iY�������0�qۡʹ�ZrFX�W��OUތ��cŸ�] �P1A���qZ�O��4+]�8־"l�H�XlxVHYEB     400     130�\��z`�i�����,@�me���Y�,2�Hc%/���r#����ii���ߛ��(EC�Y,Qig��J/��C�G8�u���Wm���+�����wf�-�VI�;�a��,�nC�׿S}>xv�jf�����-P�@�ѭ�_��g[�T��Q���\�K�����^��C1�(��6�����.UJ�W9T�;w�L��M��g7�?Z�O̲%���<��ϻ�=S�������~���Q q_��.��2tѵ��sK Y��a<A�X/ ���e񓯝�JE�7�K�����@��!�\�XlxVHYEB     400     140Ѱ�o-E���h)%~6H9+#��a?"�:�N�?p�
�ɕ-��	�x0u88��4ܿ����a��_�u+�ƥw���^���,5EPEk�q�f�������۟��e���}�ӣ�\�@���&���<���1��{[=�wrșȠ�x;=�ge�F��H���S6En�TP�C"k��f������8%���ĠWB�1'>ղ�ь�\��(��;��Z��M
h90�����ș�垻�U����'��OT	�y�����d��g�Y�-R'��x�vԂ��=���'��W��8j�������Ҙ+�L�5�8�	�^��h�XlxVHYEB     400     1a0;qd5N�v=s��O�-7@�r�H��V�h Qq�1ZlR���2gބ�U���M���T�1��4e�5���Gl��t�{���hM��5E�6��0n
ݯ��h�4JfH����P�afiD��ʉ�m%۝m}!_I��b��d���Ƿ�U���9������`�k����{�k3޺�'R��'�J�Yz�ȶ�|�Q�迻�K�]���o�vqgZ�x3R�Κ���l�E��pJuY��i�Rř��M������� kE���E�.O���b�E7h�R/f~A�§�8�����6Ҥ�Yb�&4Z��I�_�$���`T���Ŕ%j�������8�^bT�`��_�Xn9b��>�hgk���!��E��(��ֆ��($�y��󖚘�O�m�*�|q�j�XlxVHYEB     400     180u���87�X��Ue��I��q!�o�Ow�����ϥ��)����o�"��y��rPϚPe�j���)╭n���)��X���@Y���8�n4@��!�e� � �3C��APi�
�{;��� h�����;�Uc3�j�"K,�v/"�UQ a
c�oQ4�	C�vZ"f�l��	��Qaa���Q~���[�j{xiq�E~g��Y0�$�=�\��ɀ0��"I�2�2ٙB2u#a�2�;� ḫ��vC��2�����ϭ���Tv=W&7�mWO��nf�J+�x|<_E��s�X���� �1���+���c)x+�`L:?��,`����5�rp�%��K�uuN Sh���O�А:1DD�XlxVHYEB     400     170OMi=o������\c��o���� A8��@����0�H���vNp�,U<1��U�1�ԬCXD� ��o�e�ki�ŧA�7�(8�[��ƫn�����ju��J�5d���4��.�b��5�?�����"@��������L�������Եf�)��Y�-�Ws^Hy�����9���
���p]��o��r�CoUl��ͱm�>B!���"���!"2�o�5�3�^�X�U�Ƞ��v�|��h%��}�Jƒ�Wew=`$m���ڒqm��RC��2��V��'<+^!q���Ɉ���m�TN����$f��5��g��D�U�o��1�kZ���)��s�?)]rT̯�R�1(�	/
�Y`�XlxVHYEB     400     1e0�-�`�q���	ZA���1;�Y�Nh@���p�I���z-��*�1 ��+��J�?�t��o��O�~�8O:"���^Zmr22bϖc�]���(5���-�w<|�������ϐ��A�1 F���I@��"T}v#��tk��W#M����drY�n�<v>맾��{��3X��-�?5���=vR�c`]}ȋ]��J�9�a^)6u�`�r�A�5ѫUzǊ^5���t�o��5���!��8(�gf�X��e9�:��.��� !�0LƲ�kz���T�CC�ci
uR��k�X�lZb��S�i��/���.�����ƌ2��P��{�'B驪ހP�t�Z!�B�C����B�z��`���\�<�&[^l��Ӌ�ɺ���
81�o���ǝ��(������a2>�5��j74�̯/n{�fk�����ùEϔ	aMX����3��G�s'��OB	�-Ŋ*oG����.%ވ'��n�d�XlxVHYEB     400     1b0�@<yR>3!7��K�]�4�����ϗ0��7A/��������\'�4�`:�;�p6@RӛIp�|��ua���1�$��G���r�Lg1���X0�|Z�fYx�EQ+�4r� 1�r�}	$^��*qH�v{1ܢu�NQS��;�-Y����*�R�йS��i�=z٨�eu:��5�A�~y??Vn�y�2eAC��J�¢��F���f�P�ͤ�����b�,O�}~��.#�hxUw�*t���
~�~��84�X�ZP׶�â�e�3�׶� K��c�9W���r�=c�N��������@C˿�\���0v��@Xs�Ш��:s��XR>�%�v��� .?���x��4ij&��K��%��6��z��tF�m�(lUE>x"qf��s�h'N�o>{�*��ĝ^�c�%p|��&ށXlxVHYEB     400     160�{���|���b-4�g�������=���-K1Xو<�-��iz�m�����7�T�5����:����W��o/�Ŋ2��}W�Х
j�0_�����K�lL�&�a�VDHaZ7bR�٧�{�%��\ys��Y$l�G�T�{)�����-\u!w�� :�d%R���w��!#�9�z�ɶ����Ho��X����6�0FBx`f�����d����O�H	|v����8��l7g[�w�.$�sӥ�ZS��7yb�p��d�:�����$�I$�bp%Kɻ��9o�Ĥ����G�=bp����[�i�R�wryU�q%�4�^P��(-_�$kXlxVHYEB     400     150<�D�<�o
��1�����|@P���R���N̆�?��l���$M���UK�����Y�ΛF ֠vg,)�|xHy��w�43*�'���C���"�[A�_ռ�J$4鲚�3��
��@����nS��1�x��<��*�����:��g�#�[0�=��2��&�!_�PQ������0��m�H,bT�_߆ 7E���ń\&���㝫6����V���KB�K̫òK�H~� ȡ�o`�*wnL��to
H��l�B�
	E�oJF(Tu�i�-K�O����̃�ȅ���&�g�td^�TtW�_�R(W*�̴sQ^�֢XlxVHYEB     400     1a0��M|3n� �_��/h�$Ч.�%�PŃ��!�-j7"R��ҸoA�75zi��]^�^�wR6���-ix��$(e�߫�Dq7��s� B'�m����C�����[[X�WB�w����fm?��~-��$Xl!B�=f7���	�Aˋ����pR��� ��2�h�w��3;���-��3PF����'������#[yT�aV]@#��Z��xWց|�X���|�#�x��̄�`�t���5����c��|�֜��um���]��o�:C�w�U��1u��:� f���&������YѮh�lF����v:��ڏ�,�~w��o�W��g�[���K�EC��|xPk��u���A�=��:7�; r���ߐ;|�i�1��)��	w+t�XlxVHYEB     400     150���޷O���
��S��I=F�^#ޒ;��-��q�錶�[T�Ww&_9⠅�4mY�0sMQ،�8�t�uj{���2< l�Q�Ԕg��#\�$ql�KCN?5K-?ڧf%va_� ~!�U�YR�B}c�=6n�H�R������d�z#D�� u�Yt��U�I?C��̳�����[��H����~m���=qA�wc'�}�1_-���W�j�}�P�Z���i��2��Q2�̊���Qu�Bz�/�8Q��賞E�l/�*��xb��đ&�YU�#����g��L�H� R��R�Lق!P4���m�P&��:��:�eXlxVHYEB     400      e0|%��:Dn���������I�����.���KoXc��9���䝍�.����p�2�	>')/��bn����޺l_o�^���n��/4%
����F����/��R=���8�XD���P1����-(��}-��������@�C�p�8���v�����/�_T��x�Tj�0�Eӣ��[,P��Y�ј;Bx�Z����n�e�#�ęp'�}�ܴ���}XlxVHYEB     400      e01q���vI����]f�H�y#��$4r�c�ou��_��v2	�,���BbfSjg��:�r��$������xǹ�������sBl�?�+�VϿ��$�6/ns�j�I^�Lc=�$��	=��?�X6�eJk�R��}��)@�	�J{J�:�LP���L�
%
1eo����5|��mǔA�l�|�}K���ŧ�{��ô���݄�PU*(�2o��N_��tr-��xXlxVHYEB     400      f0��e�i�b��MP�!P�2	T!��J9HX�e��Cn��,�z��q��g���X�	��N1��������/|2v�{#�S�;?"(scn��m�NE��3���=_�	�)�#���yJj��wA��Ӑ���\�l����ŊfWX�{eB/�A9�$�I���O��5"�¢����S{�}�8c���`Ǜl��{Gh�G-��� f���!�-�&��&���iή���%�W���_��Ӳ>�5'�cXlxVHYEB     400      f0�":�߳k1���֩���e^엻�3�Y�������?�8Й�i��NK����k�*��ܺjd�+��v��\Cʔc���;�>��Oa�3{Pj�Bb-כf=+k���3��_R1�hL]Ͷ{)V�|l�2����0��9�6���k0� Wx���{[�Q�;B�u2����iL���vY��������-���r :�k~�W�o=��� H̠d_#��Lw̦A��$XlxVHYEB     400     110�9|�i�_ǋY���e�̍7��m�X��ޤ
(E���A��>{`�:^+�e���ANB�m�]�Z��܂61�CP��g���6�z��Á��T��tOh�(�M�����C  �Y�ƣ��Õhvd����П���0۱ծ����rSt���9�.qY�J�F�c� �&Z��.��辒Љr�	�~TB�pŌ~*��<	�LZ��,�p�鿚�1wx�&I'X�Xr��e]�	�-�ҵ��	��;_�4Ȅ>�f��$k�ͮ1X�Ժ�e�IXlxVHYEB     400     1b0�쌭Gtq�9J5o��BI���9f0�b��5Bu�<�tGzqR~tP�<��M�c��dq�w;��Z��PJj�RS.�hs�=kP�e>�5E�XW�Ϣ?���{_���} m�R8��}7ZM��yTd���9��M��	���ʦ�ݺ�e��N���6����F�x����~Q�~)�j��R5 N;'���2���nS#fC\	<��������l1ÜM��O,��)R��٩	f�8�y|���b<ak��^��Z�4� 8����9�&���x+�4mH�o�0s�� }�c\�#K��`�ix�fRm�-0z�=Tr�՟�e>��E��i��\��I Z�6�"^C54�di�;D$U�,���[�0N>���A~�T���ߜ��^��y��k���狸L��Dõ��T>A�_.ץ��)昃����WXlxVHYEB     400     140���}�H=$&��,�wA	�����e)BԈCN͒�Q���s�J��LԲ��p�����U�MI�,�5=����@g�,���~���1���3$ɼ��;�t�L뀌Ϡw�� ����փu�)a�� _@R+ȼ��'���Ҟȉ��L�����j���6�~�V�H�Jⓖ2�����
@'-�v�|�t�t�lYl�� ���e萕*EJ�6�b�2�t����.:pw=t�#':�%� k��>���Goh�Hڻ��ٛ��eH���+p��CH.zu$�x�a(�/�����F�=�aZ�Q��G�E�*�x��$XlxVHYEB     400     160'�Jǜܩ Y~aEatm	�5�!��?c�S�������B	>iv��R���)k��	�!���T���G���#�'�F8p�:A�1zm�����D͢'DJ6���l��DU��HK������5cMC�ҟ�J�i�y����5����qL��!]�O����|�3�c7�B>��T�M�`��͎�$e�9]��c�{ޣI��S2Y�M�8p.��� K�^Ȋ��W{3;è��A��0�/T ռ�x�&;fJ��G���Ǡ6���nV��F�貚f��B�5�3�/������Bu���Bە��1�A����J/��Fw��tU�� ��br�~w���Da,���tXlxVHYEB     400     140�n��9!b ���&HЉN�x:�s�M���g��Λ����ȲzM�]j���eec?K<��3�PҘ�G��n��P�VS	�Z�֕���gO�+���d|��j}��Ӭ~>F��=-�7ޘ�ŝ��X�5 qdEQ��1	v�n`uԀ�´�A�D )9_���A�r��	v"�1��s�&�9Nr����Q.X`3VI"�;��}/k�=k�����Oӥ���"8�Gb��|B��8��HѬ4h���8�{}H�P2r;�������8P@�8F5���v'N!n�)-��p��I�UA�*x�H�z\ȃ���:�L[->� *��\�XlxVHYEB     400     180���oPݟp<)�ڛ����D�Y����2(F�q�� ?�H�eK�"w̤��C���7��|�u�I*�r�c�4� m8�^"��O�a_�k|٠���#g�f����4/x�qW�N�ҕ�r2&`
Y��l��&q��OG`c�G������U��$yA����A�YF��`?*wA��v��o]�Ӗ�ѳ>]�/��B�0�t]�p���6����QN+l	�)��Mc����x��$t����ǂTՎ�o=��	V;ª4S�.���1Xn�F��j�D������`Ò� ���/�p3����{vgP6��>�a8`X,�r �t4��ߟ�x�L�
��8��б�e�w�d)w�7�Y[E�$��m�骐���
�XlxVHYEB     400     190��
��B��:��`ưNVH#��΁E�!���RL_�)
�P4��]��Qw�����&x$�E������l��@���M6�^<�ID����2���,�<QˊtG���K����G!)0���s�����r�׺���a��˽�P�?��U��j�Ii����%`,�czR�.�ힿ!+��
��j�g�y�IL�fuN�{+ci�$5[�:2c��4�F�r�d���#����̴��H�a��V��o���.;=�Y�X(A�p%#���7���������
v"7�P
="ߒ3�..}��ѐ{G�p4x[�*'��g�]&�yp-���'ǂ��B�*�!����r��q`����8�"�m�0◛��Wی���w<3Y(j��^]EC���47WXlxVHYEB     400     150��@p~��v�:����B�Ί]<��[垮�8}�ֈ^ziVI�"����� �.�{�w��#��мU�G�����G��#����]���clFw���rP��4L �"��4.�zo�<]k �����F<�|��|�*�ڸ*6��b?}U��|�����xK�ޥ+����V>�:Tc�}y� ���~����b�5\��E��,�`J"�Gf���$�C��\�ÆA�X�/Ԟ~��&��LHs4a�Z�<X�ZQ��V�Y����`�M�o���\�����T<��:KZ���rX��3y���L���BHi�J��;R�����.���G�ƁeXlxVHYEB     400     1a0���w��A����=����I�튧xu������2��C���P�L��b�1�P���杻�m���D�����R�ƲY޷�l���2~��9���6l�gxPR��5�A��a�O|2s3��bȿ>�̋�������P��M���h�m.׫��q !@-Nm���`�9p�;�W�0~q�iM*���|@��_��>q�k���Z��?ʙ����8[$�����}'3�V�����"M=���#.��N�%��S�1w[���fa¤���s^^�+�iE�U7�A�Ds�mJ'f ���ىH���~R�K�EV���~>2��c��B��h*cz�4��#�|E�?�!@���SS��,�0�m�B7X��~���fc?s"�1@����,���	ܶ�0{A_�º���:�S��1XlxVHYEB     400      f0�k9@��-eX���1���)׏�%�w�,!څ3�7dk�,���%�_����:��43C�_��;ٺ��F悈O04��4$��`Q�>��^�<��Jt���_B�	)��'�baU���V�B�ge/�+5x�MFVm��:�a~w�4���6a)��g���.�l���u�u���Ͳ��Y�E�����X�c����D7g�kx=�L���|����˯�_R�i7��`�^���"�$���XlxVHYEB     400     100���vKy��$@e<~�fRB�S�xX!��+��ߒ�9O9�3�{��~lO�CO�B �du�g$���Z�e$�����Ͳ!B��U������S�zح�~g�J���J ���|<B�	��S�r<dJ��b�V�%òg+rn>��~qrCތ�#28�LY7m�S��s�B�,��**;��k�9p�b\#���-������"�0��刁إ��0T���7��W�3 ��-�`#��P���/��
9��V2]XlxVHYEB     400      f0�#ߕP�*�4�4C���:8��?��|h\����T�A"^����Z.��1<ѭ��_e
�b��M�c�&��k�L�$}2?S��Ʉ�f���I\�d��f���ض.S~�yIl�?ld��!���[�2@�ZJ����L��
r����.�8��׏GS��/O� ��"˒̫(��5б"�|�AW�P]���(&�d��Q�$�9�+<��jH���0*�5o��:�7:�U~XlxVHYEB     400     120�;Vt�� �C�jI�֏8J�ܺ4A1�F��X�.����
f�n�U�VI����t&�����Z���q9��9q��
�쐀c��%��ܶ͞�ژ��� |p�N�� !54{�b#��G��&�j����p�=���X�C/���Ǹ�,�Wq�T��=(������!�n@p
}���&Ѐ��kO�ȷ�3#�7z��:	����S��X�f^���U��7���ç��*�mԏ�S���*��P�'�?Fn��qYmhˎs	*0H�DV�fd�x.�w���C�y�jr�XlxVHYEB     400      c0b��7�7���c���d,�����K� �?UD�%I6g0����^���}S���_��M�H�99�*��>S�U�#������;%o�I�LQ��m)�RS��
^�m!h�ي,y����W�#	�Ż�T�k��	��A���y��C�ѯI�U�GT�̂�T�+a#c����6��c�<E|��_���1"35XlxVHYEB     400     150��}{]N^0�:�p��rF5�<�m8�8%ѐ��{+f���xI->>�6M�Kخ��<�$�����Lg螘��&"��uvf�@0�3o�� �:p ��EC��]G����d����e��+�8�p�R1�'��Mh?�����(�NesZX���65D �RN�^����� P�t�kppk�FX�m��:���t��e����<;������SJ�g���t2�ۣ��J�����Ƨ{�Z�v���ų���D=B�
�ï��~+*��70�Gl\8�i-[*� �מ�:t�N����C�I�&>"�MC��O���eǰ��r!k�vXlxVHYEB     400     130���C�D5�^��r���j�����m8�9�oL�����O��n�π�I��}U���^H���DA"��<����hEMo�w\��2�c����Z��c�O�n{��G3��a���w��6 �'�5˙*��d���gC�F�;S���2��|Qn��njܴm��5NXMx��/�����`Z� ��+�*w�
M��F��)�U��$��w��PP/h7�`�\�&\3xy�H8��'�@�6�?kaD]BF���_���1�������)�mGx�`��4C0�Y�8��6�4I;ÿ<*o�U�� /XlxVHYEB     353     160ڬ�U\�����5bZ{VZs6�֩�;��gʢj�x���;n���.��P{g��U��k;�&3:�q�ޫ�Y<)���"�|�<�b�v����m�r+@���YPgxR�����u
�LL����i��r�A}��6�Z�/:W�/��+,�?�яaN{Л���Ux���2{X9��� � �;�c��Q�!U�9eu��8��^��EǪd���BdY�@���*j'��fd��p�������+dU�싯r%=�/J��x�UzTnZ$#���,���x]���UBCpՄdN����<��U{��m�1�%���n�a� ]U����F��Y&ZV��vw�C9�