`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45824)
`protect data_block
FBopDskpjdaV3reCBmCzAArFXR+j+9BRn0nimakY7nVFWWLDCZyQN8nxoCx8zyqWBb6YxZsrtp1Q
0F8opcBt2O//IRpP8zHxYRvr0gnymWHwtCQoxDF6ulwuqytavyUp/0iq59Zta3Hhg3x5ThIcPHMP
soehoVGMmMHWlW3etiDebPbH6tSL9Eb/4IvPQLIjybSkldmImD2untL1BOQrH0bHt4+XAbhJHqzC
duX4afyC54mFRWyRMDxcvyKLSlYOkIpWtXhGqD6DTCzzsKeqkzRApyFcOoqDO3fEiGUT6O7a2ucB
T22tYMjykbJPibwzbGyjkcNn0QeayEefpEWShIIczbm1GuIFzYk6wc1fml5hi942xSi9ILjyLsPB
M9IhbTQ0Ag/qCFRjsi9u1IY+H67lCjTnmoPjavj91kgOcqtrIwkXlGH9Y2bFpDGGbphDgFVN9gD6
YNhYNexiYpvJ6aF3+TJvTbjm6rpXBAZWvegGw+Rm3TBf4yvZsGfYZCT1bUKupz7lf93auHDAnHIs
vxA0bEmxQVQdEIwt2V+GH5FMgRN9/LMhP+qu6O1FeXdwDfQtJUzuHh/IqNGlnihdbswGXbte8r4z
THowJSOZqsMGN5e9XxWI4HlT7/kaXbqe1W1LzJ6gbqxSret6Z9FxMJMwCQoO2nTXvra6GLcicJIW
oKjFJl5d3Yp7QRsU1uAbvB9XRByyoQliIpixgtZ2AUdfygmMlzg3Xdn3790PnyHR5pQCKogxIE/E
gAiDwqJmo6aZoyEEZdljM/C7xq8oXxJYcyuWvlfSxX1FBjHRy84/TJjpFNgakNkw0YujdKWsKAXg
hsnakwGrbV2BAMGuRhvFYdXtu4D0CW4qOuIndrnOOdHOdFNyBFwcKvCRKjfbcyRFLP1xTAIiJpj7
QY6tXoMFu5MvWGqYQptzUfa9ikThExGstqBGqXFt1l9bUpzrhXdIm5SxeYCaEUOED4M0AmSZoOWX
BJ55QoW0wYWUYM8QWRE9Wlmgtb4L7rhF5nPx+JNZAtTdrzihagZxoGLmGTR9OzOK2kB+7Wsgtu4B
iBn4EStSN74aQYsrp8DNjDx0DKib4w9FYD1nTz1Oqtjr6ojLJIcLZibeDQBAyknYrQp7oZAw4MZl
d7/VGajmsbYF+SUiMuolQQzgnjvsq84iaWawEZvrj2VNYzXW4jCEWWQsrsID8gyEcuzFheA9oHzX
8SHX3chs8p1wFfyRenGdrRlCgPMBiY5SXEsK9DtorU+grz5wuZAbcphKO0hMXAEWncNpEpW611zR
9gUltudi6hL/5+WAL/zzauKIMuKlvmtUuMxl/esiigddlO12xfJ6ipqVBlgm4M+ScBHm5fQmsLHI
Gt0R/Z6A6cw+74uAADHmfNLAzSBiJPQ2gFXfLq1gsZV/2X6SNsdnj+zRl/t1xPm1mgg64ud6pQ8e
FKCSwtzyAnjuGBR8Y/irAzYsOwMQwHpJT6Dmwawv+L1Q9U8gBJ4YKrY0JfKdPa0VNlfpV+otHoqf
hAc2+MWlXPuKOrxbkNvB8gwQUEx8AnKLSd+kpD0GrSXgOcUROF7gsc5HB6hJQEKZp+4JY0xv8MIn
tD4979xPd4nwq/WONVWyUO0tAtpg5XM3kkhQ4Z9+V2A+u2J/olx82466wdF7Gc3UNmCVl2pooPmx
BfSC8RsIalps008MnXutr/TI7E5XeMqwXVKjgX0QwsXhWklJT8HUwX0KHTLUx39rImlKN/AV3BPC
/JxITC4ncDjxE5X0B9/v+8fgwgBM1m9ivn4EreIo+ZYZ2w5PljRetBTZBiyKFbSyJ0vS7y/Pi/7G
dLvj93d5UQI+LW4iPbEBm1XCxdIWuUo/fHPJacJBTZCvETs2o0OmzjodG0KGjxUbqOGNuePkYpJZ
5volcbsizO2W8fHXd8wiDG7eDLpYGIDwW06hBTN9SlCvyU8uv+scx7/eIR7g1Tz4HqgSsRefkz0m
GFv1tyA+2kC2XEDgXaVbOEfS6sl+T/oXx+UglhMqDh/kCfNTpFc1celaPZhRxc6EvEfkT+6EFU9/
NCpEHlEVVqRseHa+4PODtRTRSGQChXRDowS2QeUJ3iRZSDPgh5b8Kn+bK94RTwFKcVQsG7ZSE+iY
h1L9zFa1Ivp1olw3ZlIuGeBjEd0+cX5qqmofsyotgjNv7d9aCDihON+N29zgSNvFDOD5AGeAAuwd
UjcpMbOT6I7Qb8uKjwtAo4mtBUHm9M134ugVqFP2IHC/Ke/5Upm4yglwI8yaHcHMLGuWrV0yMgu0
qlcHSpWGJ/1jCLP2k8e2Z7FNaxoEQxwS0+AyCinJnWgE0LsSH2QSwurP01si1s8IVzIKhnqPzuga
yTJXrnGvWTOScymswUODaNxUaPVRvgcpPCCud5BdEqQ5ryRlK7UPDQFef7+BENxDjleRTdQqE3Ny
Yqc5YmHshmJNungvSyeXIZZTYJircZ3KgCwmCoXFzetH23qLvFcFWWLvzFmtURYzvXORaxTi7v3u
Hyw/YUGNyW7mo9yE1RrNgb8E18PENVTe1sbcLQyAdwDUlidc12zwf2pDl4+EJKQsW61TjQ5nV97P
HA18kIk4aqxghTR/JX0OeDUNQY+CkZ+HvV9+FLRYZDbyZA+lcbZYKQ9ejqdX8Q1eaRTdTeuZUS7Y
cwHV31/Hjd82tgGcCDm71g53ZOP7iGzNgVv8Ls8qgFvafk0krBfSAetNlEvu7gj0HRFdwX2wwBjz
q7PuG5qBPB9ghsq7fMi4HRfFP51BZC+C2hwgWJKWJswOc8aC4ng9QQ1ch/jyNl8tg7aRkvpUklkp
rOE6owCM3P532t9hHdw8LaIqvNJAQdg4kjZbnxR8NRhDGJ9I/WdrX7L0lFBn+BmkbsnUI9hyGXJd
fLPod0dq4kLwGCEonCFfMz48EwjkHO6a19vRsbxwLcwvPZKmTk/bs3Z9CBz/JsAVlzTStqXH48M3
YlLKj3XtAUznommMhwU5Qt7oaIcHsmvs7xlCu1e6ncz/M+zPr/JuOCx/VbV0+aB7s5+E/YeTTbp+
UWpWtBgKmXlyUX7aIhmpYlIsF11M+/HJITFJxnOVXNwXQML85MAy/iJwdzftFeSyBIpd2/6Ge4tY
B95HGoWlHotlYHvyuVJeLyiHI8WsEft4NWiU/IWlaL+ieABEyknXrcMmsN5D/eb2Sf3FzExf02dR
lOo5xaupsBccQSGB62zQhacGjHSKcPpZA+PrIZ3DwjhG4JESifrdQ+dpGxwNIaZ0fltZhxe2Spls
TDy5sFp1/a1PqjSPZ7mmLnbkZJou+VdTTRMEmcUYmMZYjg1qUykazlLrvGALm/RwlzdTMuJ46xvZ
u+iBFMYHPOoNK3/G3aAHyVi4EbRH3fiaNaO4TsXjimCKvwRz+qlZCxNMFCsNejh5ixplryG6Ix7x
2MbTPp0EFyhdBLOhZv4l9ZlJDMgT3BOHMedjPBPHfXAFcCq1ovvr+/luim0ganh7kwhrC0Yvl0za
dFOa+7H/O/zdlDqmZdTmvvrBnSgY90gqgrRzQjmp8/kWI6CBQ64GS5DBTX/65mIMiSL0UZ+erMOz
btCaE/CzUhKGf8VwPK6Z0CzHtwug1Sokp5zfU+htsfJf7yxSw0C8emzqgifp8rpYR352Qw36sb1G
75Gv1wqfrkf7WK3+GaQXa8GiQQGp5dM5AGa2SxBKTCtFUXmOdcfmjC1nLXeT05Ei6sBZJyJzjpDr
jwuxJvX/wDzdbx0GUwTjW50Q57tVxleCWMBjXYJbnmz5xtVPBI7RoMAK0zeq3mxh0GAzJVoc4zml
ZynHHbuwOiBGd1zdWa2M+0nQJcCbXy43gcULljqN4hd8gfbGjKM6SrnkLNINexWQiIwdkJQQAnzK
okhEFIqggxI8l5z3s3YssUyjzUDKi6jiYzlHVO90L+Y7QVe9Fn1hGxMK6go/DqcoB/c/G5+nmB/h
ZJU1bbxnYRubtp4pNTdWzfUCOfsmxB75y09hB6eHen3+DagqqinYMNGaY2DqSwYUORSBMu+57ElC
FQ/+ZVqYrkTDwfl9ynDWg6j/tpXa4estu62TVOd+h4/dRM+NEkgw8XRX6awmG7VNGbUyNk08dvKV
dKMTyAgx93jJKe5VtvTJjvr7PaoWINyBmTrZsOPAPnkwMQDB1tdTGnxG4zjXPD0BN9/p5hop2e1R
VvRVDwNzng+2QSVUCk5pJ0RsZWo9D8tyd38bw5UDVGexLi8qwWRTsisH6cDyLf5fyjlOaJ2j9P3W
LPJziLCfYVT67PvU6MGZ2q+VOMjSIUYTH1Bph/jBG5HQcC9ognbbJqAsa0up77iP1KskC+fZ4ziw
5qua85T13zUhy9xEgH0TnCzAGW7S/uQ90mQPaBAfkzrJjoOqBm8B8tmf9l7DJPak7M/9J/or6vIf
lj/xgbEMPshmdbCvAJt6F6qiLp2mccYtLBt8WjloGek5iuliV5IodzAC8LY4yIi4IQYL+MYirYTt
bluy7TEy6rNgzRLfHMI9EVUsxh4rby+HyYjqcDUGAcH+Ga/2hJfr0ao2XcXQ6JlBCC6qmOj+vy5Y
tl7l3qCK97txReU3nTwXT640SMno6+YKgs4b/QZx6Fscil2PDYQ01+ICxRSzNPQfVTCZvRQNsU0m
M94Ao84zwWQ+Rkr5E1eYruooXeGZEN3Wdt1mCTzpGKnH/dhXH1ORJ3bTPxzU6Lc0zw29CUvWplZK
MJ2PF/qmE8GVlTRdKzan7gkQvnqrvjIsVt+xFimGaH88tjv9u0+NUfeW5uG3LtpnYVN5cmHKn6dH
76NA6O81J2Mu7AdhyBnNXCEJ7qehD+AAZ7Ho1nPKTxHrXAfxGi7BAaVB+3ndTtrDm8UK3M0xvW13
PIEGIHiAQSBSXbnfDkl4ZT9uib/rz7qM//frpkdKQs8oQ+oWhqAf30MaPZXLOS/ViYWMdbuG06Sc
A0aqBcvNNNBviqsldWOQWptxO8CQlIOeVhockG0oQ7ZAPjjqrxhpO8PSjezMHJpu7iEuHfqGbpdm
QIFyeIFafU67cTkyKkUD9dH/hPd2WA6die40ZZc6/J7p5yuMXlgvAf7jSgxSIqCEkNaE5XqfcXpY
GF6u64S415dn153LbV37/z7JeuTOYOOcvSy+RdEO1HEPPd/WLOGweUMBXG4Nz+9wht2vaTUJSUER
PJshb0BDhJ26BLDBY3foFE/hGdvjWhOpYHjujf74UM37L/fNMV5HJ6zjruCUVMbDHpeX4EWGGgXU
OdmQj4gT5708SXyN+JRqbh6s3ajPTPdibhJOITxjFe9UMIS4iOuGIWzGSjfbpJD4Glk+AFKbm35C
GhX7pDsfJNbhDElnyNa88ssdB8MkuTzSxp49g477hbT+qfoBU31PjIepWcZG+geKylFkF3RljX/b
EjJ95GtYJhQeF5656lf/4w1iMFXqwxSAaqHFUHW2EkTC5smNNqv069wciCGwqPyTMgULqUkXoL1H
0Bv0R/4VM8t0j+dnHK0P6dhDcMfXxMXr3/YMcbNpsXaZJezWzS0BvITMsuq1SwcR5mcCwp9V89ZA
kX13N4kex22gpYFQ2bhgHmgU/XSIH3WULVE0TV5LbYcHUE0ZkeC32aTJEbe1hhO78ejq1RPxzbt7
q6nts+mPI81862pNEwIgVRXE5NhlFCFYGWX/yrEDt2+ebVC/Rmz1RB7lE8TqleB9ug0CGODU2Chr
M2feF9o3cbLOqp1WyS0QFGM3Ea8Xbj+XD4UWadvjPC55zUORHxehvk2JV43XAX2bUCxPEY4yr9tN
QGoYFhuUq9NpeUSnL2E+bmioMWGInZ/DMYzCJKFkzp0X9sS3nZcbbHg8FdkOK6LSvfDZLQCCQsyC
M4Eu7dLgxhpi+TGQJMpAOvuxhktPcBFi46UiQIOhGAcq/y31+sn2Vbqc1Vw8jqIRaVgV0DP8DLjy
8ckenQ0nGjblVJcddsW3ur7+mNYnrkHPHPvrhG4GQ8UxztXD7MvJM2cUybEeNb9ED1CCR+b+K+k0
+7gWGrO41+4x4tooszM9jXzlJAp2J7npaivHT78VrMG9JOvC+kH2HtcfHD+xHslhuScGYijQTcQK
6lHfanWoXgx0WH9xNUkBvhkYJdjTGSPXwaJOWtKCN8MkkK1j5wKINWErdVHal5Kz23vkgezL7m3e
aFXxzH0Ol5SRP3oalQWTMCBiMRIvigThFspzmAC3IdvtXmTxw4tCQphSVTI6thKSnuTV3dYKFAIZ
0paEwVra1RKiKJKqoSCcfBK6fvN6U88z4R0mWkur/C6yAYWTAJhnr7oHo5hsr+Txkp5ds+Ci3G7y
hutCXlDlopHwMOI0vP0R/gtVwZ0SZvWF4K9FUBeQ4I6wcnVSp+0s6vCVQnN7X00WyHgTuzFwqMAK
VI2cKqz0TKzXf4PFWWt2+f6Defnngasy+ULgME8vLG/CBsjBFd5olihP6dmwiMf+zTg86HBNeAby
K4ZbACideaLSQoLjZv/25SSVHIj96/4cM0m721WlpRDJFYwnykZg4eWMcPgRijE7PiI2nG7k6vPN
NRSsRew1EJpRHDMELx4UxQAl0v5aOvC6MuOq/N9CA7ZL/ZtcF2FQVe46Jcgx36t5H6MFSha3WHUX
/d5ZePjqi/raHSyIDGlgUoUr+BTn/y7MAeEVm7KI9uNDnflj8SFqas85+Dqg2jdLgNc98Z3Ms+S8
puwK/RIFW2uEDzcMhkIehmt/NA0zjWxXuOeqGCtD9FuA73gpRBStRnvEmmswCkOReGW/PN6MkQcR
tsHxtSe2vNYHZq0+wJhOZ1zpA7l7QRAN9MNaugf+FlPezwaZaLDjKtRsiRFTcTmtNGswk6Gz4qVE
JDe2igKCrFvCJ5RKqrLaBvrLLvNCiJWekRgRxYBigOGhznmO5WaH+Un+RGR1KCc0vMMz2SoF7HCi
/3e0N1gDiDYoBTv0BHZx4kP1W9O8e7HjYqd6aKP5T0WM2OMS7CPnXHagjBtA5YscBJa1EaivPtlo
fBJCTWpen3WkRScHYElHpuE6bIMAlIrQB149zbwNbfD0HvI3AhPyOx6sjIZMkJQOVPUT8v728gDj
/EBer0Km+CBrfEm+gQ8YQ90JKHiQoh9h5Og8rkaZySIAuS6QPfIRnjX1078t1pEXeGJ4k+LgAf2H
sFV3fA6hb7r9PVZnNn3oSh+PD4IX1esMTWGPV4RCboI0q7fHW4PkcXRJjrXInpBT/Qk2HmF9adMX
YbFdbBvLoLEQwHFXENuIDE3Da/mdoCw4EEW/FiR+sY+rqfIWme53asZHO7QUDq/+PqPoU2J3IvFM
HfKIeVcveOCRzKoptEMaNtR6WEow+UFMiTUErZRXPWxfAT4QYIrqZMwoFSFi0WGCASMQMROTxs/J
tWeWMrK6ZED3QDq3m91KVaztm2375JwtWlzwYVPF3gSYwkso22MbQxCC+FVLN8uKwhcH2ORzkXej
hUHp4byFJ5icpkcJwmo3DvTD4gvQ4vPgRjjR3cjErrCSmwDrGFsLIEKEKi06TP8w/QBjB8qaTDZw
LmpDYgCzpdZWED42gtpTFB7lP9dSzyY7JNc1I+WOqnRgKu4DMcpc2sFLcWeVwquiVSamu7EGjHlW
DjAH8WEBWXH6r+507cAAMsPtmhMuVqT8rdg7qKDlN1DKgERESSyRiA99vyEGByOVFuMBycSBLlDO
OeMFvuqrZiKEm3sj7IlLtDfalhVH/y1yMlO0MsQZxpD7vnrPQZPFrM/Ml45xwFQaES0Tuqvh9Fmg
oWxcZBaL9/IxCzwndikPPRKQZn2SdSQoYldvTU4XfrMTYXsoVqpGEw68W3FJu87VyLR2+n7K8fJC
VIXKAOmGhQccL8ICSXeTvaQEQ03Pqgr1l09BJw4GV3p5U4VEG0DVBTE2oioOHu/RA6yFY/3hYWId
PVrLdWh7iu0ybCJfZJ5h/IKmKb+PDNaLRRrZsK7AnFK3R5DwsPtMgabDKh2tccMsxsRWo8gogP2Z
NcESmRpLgTBCFbUosxjUv955dOkWwf11xvFwX8ZiU30EJfN1zGGLKcwQftvqp5MbX4FxfacBAECh
yXdT1RCevxAkEv7CzTHGNpSZ7yK7YThhHBDZIedirzbDgD8oGo2sUa88e4NCE22SdvOBFIY4SSSv
3pGzsPLwLn3q6+FQGoxSKwchmSVe7IegjIGS7FW127ig54X/9Nq0WCBO0OqQ7L1CLnvhHxXziDzB
B8EtiKZJVHJ38PE2L98u+jm2iisvxfl2YEwevPFzlrcuvRnFFKX6vbI8fUmcQcyavMmNMkDc5wFh
/pOhiNRFYaISnURsPWs4416zUEhY49ekBzuGcHG064gjRGgzKe5vleylCKGpnzsLnzgiEafN//SA
xs7eUOkRsfyFcsE7wXsoKDslJ+Qp1J/YTrmywQ2Bucdd2dWpllgcI6vp4vjqkH7O9kNv6JfD5ExT
N4y1VhiS1cGbZy6btv6JPqKYEQdkwI/6CoKT1M2Ewx0hBQ/y114AJW5eXR8KCHM0hzDR/AhWtP5e
XZHxulCf025F0dlr2uUSutW1HCBjMtDRGRZy72M2xRjuW5Ix+5PMgs+uBNim9LvqwTRJsdGX49Ur
lg4nlzmM77Alb7S3XnUsyeHfwlJ/bDOBvJ6aeOcAstAXF7m9FCnXC+7PZT3Xko7Z/eAwt9yVWgqX
l5dLQimM5XvKbffyYDtFIOh0tC/QJ47wJGxk4cbK0tw0mHuH6/XQQ77iYLvIusKucP63MeKg2Xpa
f7BYIdFYSK2Sy730bu3vlWxB0CAS64SILUEa+S6cVhDoqBulDgqQ6AV/ZL8krH4TkPpgpaLWn/ul
gjRzvGAkLnAXvPSzQA6fbrVe5ncKR6ukLNDPs/Aa+swwifJIzBMeu9wCVe9bbKJ6tpV3rSNhLPt3
bwh08wbyv6V45GXnhJ1D7fPRYqpQt83+IqO5SLZgUSNe0rMBybFH8Z5OTFM2ceZEDMZ//adALzTt
/IxlqKcecGQphPSCejBTUzCUlndCVR2uwFjUIMy3JnEEfj1m3x80dsXR2s0FPyNuDw568eazgZv4
dWTMiLOOCUmnIBgVJBuNOK59pPbrJJemu65AMTAoRh/VcGg3HwIboBgmf4bd34lyUdeT4njegD0l
0gLNZl/dtMCjRXa38ZBQTMpVk62qGYpuQEHpgOu3x+auU0xf5vvzK6UcVPYFiqQzplUlpUzj6I8Q
9KD4WFIB5SHeo12y4hf6bK1w2hi6PLgIybpq4gZI79AhGqetnIqJlxhWZXzSPKZs190eVMZ6ukHY
SHh1pfAKBj4xoOS5NY+fXitBwPZ3abM3hWYyeRzEu0xHRVJ3TZ/+lH6XtWLfyy0GnYyw4CWBUHqw
gGl29cnjQGZ4Z2qrmhKRyf42en6d8QvkcZzt9xDVN1TTTpxMZ1aSiTinF2BaDOuMhD28Krf391ew
XZupodi42NSDCrpKdwnkGCUrhIbCL8ToO9DbxlTdIgleUTxZ+QofWceFNnKXnGjUQYgNmK2YecfX
Mbb19dM7TSwFMu9YegwGyQYq69oxix7yjbbhITWt+ryod0keGJowgYg+GGu9yu1vhNqNacQXHWT+
DFHQV2yzhpzpJC0u2mLv/Pag+3la3qGUncoZ/qyKzfO30yW3aDsLFyWzqGc0wFEFppzB32tUqy+x
S2BEwVTmUmgbx0qHA3/utq2qF672LCT1Hoyq6TlNRR4J5go2dEzyFX37fWbU3Ct+DKd4SnByTG/m
vipE3ae98RyZ92/EudGGFmgfW7rVhrbAefraDqdCbuxS4/hIFDwYjr6lY97R/sJm/t6TOtAordFH
AyJXc+yWs2X/yHTojiId60ehLhyk6ssZripBCIb/Cyo6hPnTRIntsSTSvLB7+uaHLgksIDjm+WB+
LKBgk1JYbqX7wvtH731mSBX54FM8Y3WYADfnLMoSebwYtiPZau6zTlQxZvxwx+izPDlB/RLNtzxU
7qs9acLAA04iMOs3Xt/RWbgk2v0Ts1bERG8Gc4JyDQx3DTuKMUIaCD8PN9ytN7rGX/+U4aAcrqSN
d6rmO51Aalb2Q+VKpOAR7Pougbsl5UkXyoJq+ne3YiZzqqdSqvgd+k+pBFNuxGaYOjswpayLhfCX
erJDhNZIVPOO3BWd8mdOHjw5c+Yc6BGvnpnG5KF310hqeywJOyHqGGaPj8nWfaE2RREmBTc5n2rn
RqmXMNZeocQM4j/N/1QdXy+r/H5IG3zELZufHKgaB4i+phby/h8tjqbUgjpbXmjRLdvYzpK2Elba
GeYLes+hymM+DGqaWTqXb34lR9bGQbX/p0f7SEqRAfaTqTAgWx5b8rWE2a/nxoaqtWM9poW5mCF1
fFKTkXc0Brm5gus4AsZ8pL27NwV0k08MH3a/8xLDmq/0T+MQawEZo0gzASDs1smE2Te853BoxrJ6
XgXLo0ODczx7s6M+KlvhsE/yhFDtmHVDDMEwFTSPuQBK5vjn7qw2Vq0oSP3VeRNtG6GwD6TNgXf6
IVrczUWnEDKai+coZnrKQkq/tnimtXZRuY58XgPzbw8xTyLSHGn2ffiynxoJfzWrG25f8DW8/IfN
D5D6QUGDUazMv7a8yiUy4tGuFJ0aMEkWzmsin4iXz7Lr6Djebh1hnk0kkxkjAQgeAHF3JzS0ZnE3
nm0C62xftfiNzxStKCPVQYb+b2EHL8f9ld6EA+zX9uIGppIZnnBtjcCiS/2ZbZKLmTLnMBBdGqmz
PCWfN7y7BkPw27rQKeHbpSVoUYXuEyGqA0mKjko3WsRRaF7cbhEpfbiO6KpTu3grSPL/KvJjHZIb
0l33EKUGRNFBX+3SO9RvZuheR4AdLEiFZr2ZllFAPL5MD4igPlMxjkQ7+X8cZV9d99GKm3/kG3TP
88vew4fA8PFJQyFl9hYvNhfhMxhAcQ5zW1fqpJU/XwsTY4Uw+5tJCj7moLz6VewnKU+dSbJWPJ9O
IV1VFyx/36foFvJQ3nvITMVfJ8/kXkiwH8lfC+esah/ktp1IB51GEhcju6Ml47UWqAMazMzGnyRD
/fPV5AVwYPHvapwwWAtNF1E7A2MONb7+rsAOtt2HSPm6sjfC63Kyfg0kp+B4rviFDR5vQ+wfxkTA
H/5DXRnqk0k9URgxd5dV97LG6JnX5ZxMjaCnd7yay2x+INIbTNqFu2ckw4EO20y7+d7km9eCD/PP
BFBEQ/+n0tJNLAGtiMz9BduS57xE6yZC1t72+gIu8s52V8JUa71xW0ia5cz+ju9Bw9ScrXe9/S7x
F7AR4kdD8NkolCCYQd11CGnp264ZdwaiDPwzKTo8G0Bdxb4u+/7qsdwZeGbeNLT3YyqdHtneZ/9T
WF9/NIhpr3xwKpfr6AFRUKF5EbzVdSg33mNTUk5/2QNqajEzzHH/MlUpJ8Fi66Jrs8zTi5xNTF40
o+gKv+GcJIIxIeN+dQ5OHJGnKU+G0g0oHFWulS3ERY/ZqPhPuLYIhzZ4pIpomV/GoH8nEHuTFuMJ
O9plh3MW3FV7Q3vLlyDG6cgzDPgsQkJpDE8D813drujn30/zkFX4QTJgUQCWMT9NCf6Lle1q8G6G
TWOB9A/EOHfFvCF4qjmkp53YE6uRmrrXiCCeaz9K2X32ArLnI1i2ZHbjz+3CInlgjn5NnK/EOJ6f
XCDSTN3mhGzk6YdQoyj1cCHUUeGUny6gyrSpoZINVDmcxfGZGoTHrmRh/CmulKz/gMLAbSunXcve
0z3Atj2Mqj7HdHk6uSBrSjUs4JQqF++qLih5+0VmWrbBIGnlpJIll08baHJ/lJ9lbNwqSRueGeNg
YYsUiUHqGtvEoJ4QHLsSHbR3fBqSj2dA0s0IDTroR2RvaUaoGepJD8Wb3hI2Zlo/1VjQfT9njYIt
w/QJwTqe4SHwfVSJ/eDm7E9oDWrfb1AHVbcud/hZbk5T+julzpSv3f6pNQnZ7tJQSqZnoK3vp70V
mQZRWRDQnRZIzZwvIwdCYpphCg+CkxId1dWvD0tSYcKHtL4Iuu7BxqxB8CZ+HM4rukhs0MopNO2U
IHxKScFnrQKbNU/0l4vBgkZzcsWlm+Ja3t/+ATztra8IQhUp95OuPhFjR28OS+an6OR4jLMx7wUO
hzCySCzUOOmc1WbF3y7ySQB/fGYaENKKQGdQ+3g6RgNvdkap/5IGk/xZkPQwJh/4x5BIokBK1std
g4xwI4G/bUHu06Plt3fYCjLO/uduBDEkLnHkCgnQgOqrX3Flg3EtExDiXe2OM8RFcY9dwL3cJ+aR
PAbTPepunLGxWMcbzi0+mEkEKtUWbaNA5y8zXkTUbhhWKJQQ8VqIvJwkiRbDopmFEEG+eWM1CNOY
/IKV+dgx/EGGknUqfmnaBYyActV7N60XObVYmpahY0r7YyBYAgdf7GNIv4S18tljSFZDigYf0muc
CSev05QUDvWr4LX1s/Z+w/uOJ+TYAYiY6pZmBbEFBEgaLEKJ2zAg4ojoeJqNP6k5kkeyU5a5lKJp
Og8EueaIUicmq1nBwnLlUh85zYc7IoFMhMnZmVdqbcGWoICIg8fnbeM5GPSnF1MKaAPEFzwIyMow
LWhh1UA6keGt8wuRNakIyCyJ35fyG4R23kq/fUmFNvMuiKgA02Duq5d+U/q50JWC1A1ibm6fxbXL
XR05TGup9whaq5b91BDpipkdtcvIu7xjF5S6xWUmcTdkR43G10FxDYeMwfMHhEtLF6T7H8POJVdb
XsWClvALUsrYg5Hm2FMw27uF4HEqdNkhd9W9+wwcGEh+8mwCaqGMYs/tW3PAWZhWU4AQXL9LNrMJ
V0yuI9sXtHyZwlWaYbLwnAxs7ju8mpZhHSGNgwKcNsoBw20VrWL0KGDjTU+zOtDkeIqtxhRqyt5m
PKWC3swLf6Z79lHTgaKaOCQUTf3UNOx8uTjmGbzSQ+wYRLiBBOUgNS+3VZymAloGT8oFBsNzFUib
bdVZKC2WGBURGBSKnet+kwPD4icKeg3/MqN0RY9stbFtRvdkduaZiik0q70FkaJMnHcTWG6gs8kC
oKxdJ9PnAbzn4YwyLje/Gn3aFw2UtzFME3J54AuHfVNrwmuMmqbL+fZWauTgMuFZhjD8yTkkRLKI
uMtsjMzlxeVTlS+sTzTXO03dWXCtAVCOQdyVr1SOxb6iD7UR9t8i8BdgmwRAnIYxulqaRgG3aA8z
1GAAI+Y5xRTqqCqGlBSeWjOkEHdaFV1fhbwb1e+LzWXMWGedPA4ulgFoCmAWn0DT2K9+Kdabfb9X
h//3I+/QDCvW1yyRnZzZiBG2zZ7s3AzS/+SN4N5OtWOirSbd/vcmSsT14YIZbfOrQjXb3Esun3fD
7q3QDZ4RQGea4NvS2fx7fFtZ/DSgsn5FX5X6ggrmplj3Yra5eFoI5RXIDF2fS7EmX/gdZX7s5nmv
aWxZXPx0G5qL5JhHtPYB/j4MJnjWkeGJkZSE6idNiW4yxORaNo6H5Zgu0WhX0od7FTIZry4vTSx4
sX/RSa0OEbGeBTfffT2b8hJf8/jUks+soxDcKU/pnE132Tumq/OY83CB0rPwax15ae6/PGqb6Qjo
PTFFqoYIurmBZog9LYOpZgShTE/wGMxpywcz1SJDD71u+WqNPNwmc9ahGZI/2bw9IZY4Nv0OF007
BCTU1aVIKTZuuGablg/r7WsY/dp+2ZDiGDwN5plnKwsnuThEqjWKwP3v3k1ByjBHGdRTbfZJOw6x
kCcDhXScWaiTNcQGvfq3LOLsFERjV6pHeqXF8/XsRPoc0mu51Z4QwQfgl6d6SqfoZN3q9p4VSMjc
3B28uuuOKV9niEbnYnGXK6nMYe9K2tGy7p2aBypTiHO9m15D5dztv0DBJ8TVIKzSl+RnaCUUw6lO
JcSJ3wcXgDdkshcZRRoXk8wheWYK7WRaaVphivbBVZZkRI20n1DEIZh3gyZM4P6P/YYUZfLcKaOs
FwBuYM9vjg80FK+kkwOYPaHedwaNGBV8jUvvlOy3ayrTwIUB2PXCANX6HBf/sICxK4vqdjg+sUuc
cBLE2FLSyIkpyVQGoElPx9iAaJssHdz/r6nVAL8AlJtBeXJTnVOSIpYoZKogIjSGeVsV3qsdksDA
ecwZbWorr+ij/XHmCPiMPtJ9R3qgR3xJ7rHd1RzUZ1Dbd53kae9OqED0R4pJgAfYaQBSYBrFvzj5
PJxd33pYaEX3SD9C/qvkqMWaWE8ORXI71K14LYSw0dLJl4bs8KUzhFgILmHyawuf7lbH90M1Jzm4
KCkoWudfYCjLd22szZ/vR+2aQAVLo7WqLFK02NeGZnGLLGYsXGfnVoirm2J9JSt7WlYbx22Oh9hL
+nSOsC8vVTLXixMryIu391v/ufpy3qHXReu0zeNRKr9SBzSyQjiOfYp8FmljoTKhE8ZLFOv8cHjT
wbz2Rw1OiiCK1FbDdd+GWUvzb9ZU9MrVPJU5oL0m3Mbx3XcAENxsXFaLssRD/9MHvD7S1EFN08kz
vuQ2O/koEMIEVVcs8FQIvFugAN808nv/tBXkTkaxX0bHEMN8SiG+MDIUGeC3PUn5J6cb8xLiYqcm
H1dcYFzC7Mo81GZ+7OfaQjE7EoYctnaJ2kE6C0Bmz4Fgl52vRVtMaUlWsoY1p6FvQ2rPYPGD13y9
sVu389v4PTaTGnczpRjwqS07+UF5X09uwphIoaioOwX73lVwVoyucfyTTt6S8mj9NT28WxFxwfpa
QeevHvXIovXe+MhB3eyHt1324+GSGo/TsNmMd7vb4gsU7GIQcSuO4TusVvbE3JboqW4sSo2/g4DL
/mlLjO/CEmaLC0xawh/Ll3P+Efswse1PCSpuWxU8qIPMVhNk/rLM3qyQDoyAiF78i1KT6z2DIa0R
iezw1+WOOGY+0akoQkxilP3JQAqR7nLbyd4Ey/DMOkKCR1FHyXe1ow4z9xwbgrDuHfQqOb39qD0U
bBgoryuc2unhHU5ORwoVD/Wpkx7CH+94xB/FignMCvRZolpgxhRTqpw09YvjKyMmDvqvxVlgSXGg
wwP29zpptU7XBUZjNyGUcQyh160YklPGiB1W1vmYa9gSYgO6PtH06GNQm+wR+XLfBH2CtSMk3hU6
kaJtWnEmbXqBH2agxSVJX7Pc7Z359iw9tN6PZIMvVwpVHStsqZWjFxlF9F0E1fmOWuk6VijH9bPt
9zl/NZAoOkUR0pEz3v9Mlw6n384ZXZm3Nud+oez0ayPtemBdrPwW9psEMlRj7pMuE3L1+8K2YTwk
CkXIAHQWZATAeK1IDfbwoj/KNtxzQmOboKYSTAdfQih08vCJ/QKaEFLOaF30UdZPCsOo1NCTp24w
tVkujx7Bwve+oG85/IzYoHKX0rgAglyyfrY8Avmgsgz/E8nTqVSQLzCEm5SbLDv9+RdWapWfsxUU
8WAeUr9+xVpXin/XfYfKp2ZvtB6Gk8ds0ylUlOyTDN7kjIt0/47nXUR8jt9GIUhwFSggqXkr+KKD
SDOOUPrtzFDiF7usNY6wWsEzPCuDeQoCjRmTNC1vHf1RzRqUFpDu1Nc4WlfhDDLusizEW5WsLzCT
AEQ7ROXR8I0EE4TU6x7EYT32xUPl2GjSgj31QgGW0jZj3IB1qVqAGtDMhEQ93+YakCZt9HkVK2+d
XUcR/mdsROmZs7WJWolzw8xrNFvXYYwhdehptW3H/f+m/ZiI7/YswgdUCRdzHtOX6HmowgpWtdMk
Lqj22l2WpYzp0qWmdOLSfqqyNa+NtEV5LNoBpbxYPoKnkjNV4uBCrAeSA78wbJcB0JHxJ2p5eu8T
st+UfPa++kLBzfTN/phyL6tMpEmSSgMFNbo1fH19jc91ktLYLI3YDD3VEOQKf7ZarC6eQt71xbAW
l+wUixwYXN+/U0dZ20sym9jTrIBw/ceWuoy0XsdccNEhAt9KOn9TJlrdei2Ym9ddCO41mpPf+9r7
j+rqGDwXq8MV/Ut04qjgBaPcSZOLWFBMpGPUP2AZorvuo1Zpm2qNKQtZlry6SUJlIF5wMBAXQwq/
U6cz/S3Oxk28zEMrY3LhYl8YMXNzxmIPcFChAP4gGZrKeSdLOdcCSobgriGvBgLjdoxtDK3e/gS7
hoJ1JenmFdMRBEBgZzNdpQhgoWS1nYwqm+8SF1g9XJjbd4oXyo3Lg1E9xvunaHh1BTQlGUBRLiMY
taHmwjqC30mdAOrEYNntBXTLa4yza6qHV3UcFazwXAeArRGQ7SpovOq5dmKk65+OKNeA3Gp6fmNY
46nLhOasx/Qr8ClwT3atkBV5g2nnVvQTgk4uFvVMAKIlPgblMkL51j9YiCIk7gfkNtaVH+8QB/4+
UMFiyj75PZW/oRzENJl9LmqUD09a5rJ4CpB6pbMrdaY97JAGB83XgYt8dBp/jsOgLdI8l1+LRXJe
cyara+Z1g+VC7WCBFK4GOxorBmI4TstVJoSs0J+HFbamq8N+rTWfzoHHaC3y/vTJUeCo3iit0Ko7
V+m+1+2OeK87281vdSOy+3CZD25Nm79DO0w1YSyEKg/QXFNU7EicXPMZsnQoGUEGI8fspGNr8Y3O
a+r8877l5Wp3gt3aXfWXKcYG01yqzJ8vjxcQ09pNd8qORKzkbZZaizr3mnd3yudOFEPrA/TXIr+b
3XcT2sYVT/EIPQUHtPdOcYL1gGvirKWRWPl4FwmYmf9UdD60ad0Q36VX3WlDS+UV/q2q5iqps/zs
BMy38bQWRmo1D8gHH33iEFRU+qYpQiiG2cDlBZ5qFbU3MldSz+S3XKNo4h0Ro03jCc+3VnaTv1rg
3mCYuH54fOm9ncmjIGyfFCa98P3tFh9ZV9zFHZEF9NO64uqxpCdKBBqFGjqFZ6gelL1p5N7rDtgT
WtgV23i31Wwtb72hWLb0C/YO+9VQNGqFqZZYLQ1k3sWxGi9NVdnVgx8IjnmDP60qhrMnyrYPiyST
4pWnibT/t2oA302hd6qIJX/TJaKrVNTbe3mhtOlibeJf/3cnw+OMOic6rPWZligEdheiz2aVgF2a
dKsJ5Ovm80P8315XgbdwwEk34LosNPfKPNSXi0HiQIMJxcLgw2H29d7jNYY0JLLd8gfJxmwt+/e4
HvcqGhA8sQnlFiBNFnfPz0mIK033Or6bbkUlPiFhi8Z2fMlrnAC3mDu/3HxtNG6/IdeqTV6Fw73s
g8p3jtbSDta0LLFW5AYERucIGQJPdCbFa1vSaKgtcu0/DDjWiVyP06xPJ5uwhUKXoQGGVSj/Mi3v
OaU+tuBJQ72tezHMzwJdWpiyFrMtrCl4m8pTm4JGWeJoJd1mwZCarGfPPns16CHJ4NeMAfmdCk92
wLzjKhk3n6lWtO98u1IMtuPUUzmePmJdoOsksGugnW65CnJqhQyMU/QlRs8V08MVHE4XR3o8CP0+
5LfMikgsLEJRWU60T3kEvgK4gkVk4J6SbaO7Uki457XyU9b8abpbxWr3K0oJoc27g/RAn/Bkywrs
g99RRR5rvnJXW7K2mZfbnnKYxrQNtG4xSirfSPHA7zdq9gi4caDHprfr1SOukTIKHvgrjgvnvWhh
p1Q0dGMCOv8yEKxqMGQTDABGs9+37wOwU7pwegdv5Amby1ZEfIB5uiQMvWd63t0kuPZ/o9jLu8KZ
UwrMtS/blsVcl9vq6+yF/8fpYgH+UFbCuUvOJjV0mxJZ435wTQ0Je2Qxg07b1pyhkxOPvSvXX4He
Z1/8iPUQfzaazxtTYxsG3vVMIaStlZuKCkkLsWtFOObnZJdhYOIHtHr/T4b46SWDVkwQq5ngb5CJ
/J3fSqH/9HYwy2gtqT7YHRj7s0y0Sp7tp951wYBwTfB+YU/QxuwAYUER7BnAq9+yaTgOWqK4xxrH
5ZrgdWv3EzDJ3oMVSOghonE8c3Wqf0sq4t0RefXMhQUbhEqnJ5uMw5lYU58GhFcbXHYe98SLeQIU
oaXd7ZecOe4bcU3Lf6Vq01K1S2s9bC27dLPjUbVyue+oTEv/Fh68s5/a8t3Fm2lnnaCSweL+a8mm
kRLKJPVCOw+Qwi/53w990rQEnoslrqzFuRSXO00wIyliZsEBHVcLwD59TJWH3Vm7JXxRhx8oi1qg
t9snmK9Dx/4e9WE5GoNPQ7JArcIAduDbqXecPlHBPC7VPmocCLSGGszsGJtIaKCHKp8/wl4Bl9oV
DqQxWHNWzX4+KXIBMKC+KPpuRBYSgQDKWQFcTk1+VtNoATeKmcq4xaf/ZXtfQErpY1waCRMnJuTI
cbiXGrriD8jiItel7YKNZa2gQAbzT4k+kyQ0HA2nx5PdYLfHNUCVzPYfzsSRssi3P3neCtw0hURS
gjx131jQ/PGI9lRz43ppdTg9Pyqsdgg+EZmTQsAtxvHe8+20n1aIkUPy/ol8kT0JAyeYX1N2j9p7
OaM3N/NIMga1FJeBfboJfW5wrKRbKeCIDdWfS7KVynoX67OBQDXcTA1b4RWTVH+spR7eMf/nqmf1
ueyOjxJdR243qkLGtj2qJfPyDQPNOdixofJr/nwOnL9EjLB9SJzdD8EgEvunITaH2pleCdPswLgk
4ILIv9yDn7SYBjM95B3kuC1hUbt35Yr5j8yvbqhYyaCC8Tm7xR/FEZg0hymAiEnWrlJVk2SXqCuw
ijntTWfRAT5WbX+TUwGCUCrIfZec6rRLJbOW0ptnJrSXvjUv0fytRaCh9WKV2G/l0m0LbAMc0OvO
zpZKwru5SyMz+GnZWSdeMbpVReCcXE63vLc38I7vbj2WqL/dnLqxXeinyIEIpDcGGNmGepIpawM6
iA7f/pRDzwuw1+rtkW8Rr/UKywQnP4LaNwM2vaGlIlOllQLporifmFqAKa6nmyBn6sytyBGSNLi/
Qf1dl6aaxpTXD+HWP3r2n3O1S8KMnxoNv/KQVuweuBsnsGL7RlkZpuAUAPkLTuFGibTJORrz5jVU
iVi5I0y3b26vcS8MZ2C73jQ3L8mvN20Cb1l3TjmVkHhUhiw0VlK0Vg0n/sPZzzsxz3LmJ+AdGafp
Hv8v1SJ1E/iyKjitCsRWm5WeH9H4ih9KBEvDsDldPgAJIRH/hpf6PtKb0tPIVnLtZnzw9HyLNp3J
NH37YiT9LtPOs7n1jGVqSutmKHVB4TfwI+Xclx7bBOqVJzapDBC9oEG52FeDk+RCdcAyhAG70Hsp
sEZdtpVmmblp8s4nlmUkV+o4X7nAuXUXApuePVqMfOytQCGR00PI1eJ7h8n5PvRhvF1JaPyTL9/4
Gmgj8PFOOXjZRfnqJo4g6zGLYmSnjnAjgxeBsrcE2Er15ctCQ+++hnW7gNLQk3M2joaW1G8zCghC
7sXAY7b0Md6OAqblGYfuLiHVyhFU4AVHpDWkdRx6ZyRTcVIHjROsfHnijet5M4kj/yQDfkQRzBEz
Uj3xCTfJ4ytwRMNpNm7S5+mmLY995opGozlEDNuzIJ2D2W2tXQS5rsL1xzrNkdHUo2K/3jQW1zRa
A8AXqR0OAux2Zcz4tVP+KQlxkhMTNdye3wK2DJkCP4LxV0vGF6Gj2me/KtwNLHV0S8PKz7bgfmlK
YI5waGdlogQ7RFbi+HhBc0mvbcEz5ciBi7WmN85v8HkcjFpdqVuefxAzlWlgvNqyIKQiUcKP5P6J
mrQWB+UAaWPCgD2X6cO3waScE75LaUE0iwv209sDLzoFwIWqGieVXm9JMpbHKQuCsW2dJMXtWXU2
iLeFzjX0926rVNDPw/exZXiyOUTq4NHcQ0bsH5T7elb/ahpi1O3nYgrkKy7curSsnNBN9kM+pBD7
FJCurqSScocoKtNtm9GuYIb9t/S9FtBlYP5GUWW9VAPSnEfWXNJG+jgP57a9eiohpRfKOR/5TdcP
sQsK28oFmyMZ5tJChq9ZizFOiU2S37lLDWesV2fn7xjKtPAjnmURq6QE6yGUlbX7iRVP9O9eTpcq
bbFwKQL0Xn9nzlhtjI1/gepiKJaVv18WxhsCmIJLNZMWlSduIyvvckBHaqqEnt1e6Xf6yLAKQodg
KQdXCygPWAxnHKj/EsuiFHvsyxT5/GygYq2e1Jq9DMRkbDJ9YThrvynCC4frjSQu3R2upi+RLkLv
GvAEpiQ6PMhJoL9XM2WtTypmKbC5fsIVXee39niK0ZbxTHJ6HrIB44aLrKbbXntmdVBn1NA49abB
2mp+mXPGSbLMcCLvPg1QQckb7VxAZ+0gZRihcXKcNmby1SzA4K4olH4rnvTJXILU6AioNkFyK1lt
QOVvvbo4vwHDJvFO96yjNX6NBUGJpsw6kQg0pAmNWJI4LBlrTKKiY5PRFxexp7fsOMEKzov3MAs9
PYaoY65HSXViGc9XVZjTyonCNQ0WGnEx9OgZdN9k0csx2TTJYHkbgbEi05sjayL32WpY3PdYZzAJ
sKMj3FtSQCfYOKd+G5VK6nSWu5dDyVfwvwpVnjiQC0pLvFCibe/Ph8CHjud4MUPQMomo9/elFVas
GstNtPpEchiDx76dPlBtgp632rCZQ1ioJz3CmEgVDFSCvtt4xoaVU6TAGoD76euGEdwt4n594Lla
bEW7Wfiy002xodfz6RAbs39lrESCQZjCdh4kSm2s0KFuLoEqKx3B+0R/CACAPNjLPGanzNtf8rc/
uv0nx9D+PN9M4rvK/p3Lotxkus1wkfCiMTig9pCmxzj+n7tmFnUFwO/R5QbHtZ1CCKJvLD95qX8d
q14HAx9q1KPilpr6t0XNF1jRtrOKPVE/Xo6sOj1sMi/A/cUUiscMI76KGFTA0s+Sw+XEmjG3tLoZ
lKAcf2lMECH82yULs6wRJJ/UXf+zBHHLH7lMKuaslp8f03KZVXCKLfhUoGlEaMnsu6AHdi0rvHeZ
OcVayQdp+6440ZJmh6W9iG9pXrSfFP8NE23E3c39AEp8JsT9SA9ENwHN5k5nr/X5uNawEYdH8WO+
9u4PPPo1z/8VGCSce8Ka5ioUIyIZDZWi8RHHZdJKEBWHaMc6MPTYEZzyxb0VTLlXnxAXW+ib+WqY
lliYH84OtPZXfWZz7i71UsyKXSEdLCFEDjF2RZuekit2lzxgYPxSmkodVrFHE/4HBXuxNamaHpu+
ZjdsLEsGlPomFUKtE467BVQhasSXGXTHF066AHUdQzEqLDLexf3tPULJAY9RXOgeC/T6Ph1P1TJ1
DRk5CKqx65bcPMAvydOhksb5hkd/lYOIPNOJCqSPF8CZT+QugNLEH7Ht3K4vb9iDb8Y5Rul9MlJ3
W5R9cWewuHI6WWcPHv69cWGQHafuLNMP8wN1rZ1EpEX/nv7tXO6TPWSPEWDF4DmYViki1tNNpLpb
3AIkOtGb6OrbJJJgQzEJc5ANEKyzK5hxkjNOD0/cs+K4C097MvyGnRerf0a0Ss9C9JIsy5dzsx4W
4YqcCKr6cznyGPdHoPkvwI3G5d1ailJdz/Z4uIWKRvHgLGYuFP/iQH4NqJNLbCT7bSbaPp5EQ8GJ
NY5IMvhBVzNQSZ+B6MwzDEgyNNFByHi1uATEUb66Wa2kdvhEt9Me6gauWoXC900sf6rWWxjXo2cu
Z3vAb8HRbzvyPLAkyu2BuM+Josjn1PK4EoeWs6B0+F1j4JdsGlywoQzuY+2378StCEqI1yOluGYs
aUGwSTHHZQmbuDpzRkpqIfokPa6qs36U76WlbkbWoef0As+n8njefWYos9zg1YYMxUuoBmQaQV82
hZrBeMHMZkXb72AYlmYVU4Atf0IGtKpuf3VuPSRGdSYBahwRDaBi0TQ2+VQZqR79rIRPmvvXW/on
9X6I7l8RXhAhwRpeTuqR2ST768MpBD5qR7mbOwtjRZzJPbfB89kNZWh0dFFJmwHoYugOxhUw5Tpx
A4z5TvBAJCiyLe4cZSRemFnCox4+djMadzNChQn7b039jbm4QYjn3/p4pefMYIiHL6LERTZFN/l6
QWRfyXdc/LQ9iCY7nNdA+X7C5hNDLu+PYkgwp7TaJd+j3UEkQoE8rSD01/kdwWVT2z0yaAlPT1jL
xt47iLg68sOmaUSTyQ/jK0SyPqDTc0UQTqG2C4icd8g3iFki/QKAtGLvUrm+7xNFHdng99+tFHME
ZFuiDarbR3lz0PrBjjtKXYmY8VR9gm2j6vnw+sT1u+gb1hGxtm4ST6Jq6B6cfRb844kGifT80YKT
JBIB6IoscmlJhnuSV93HjF/v+9qEIEGuikEWej4Xo+02RySKpNiggkLAqqlodkGoJ2BYvWGwv3Oa
/45Z4slYSEOGDmDJpXo8Sy+o6wM3ksfhCHnFhgDcDWcz8Iz+Krmuse/h4qjyeSX/EaJBva6ayR4w
gDZ3vxc1Xj5ma0FXIjfVeM5+WpgreJ5tHiFLnJpTGN3yyrSZToisBYKiqaNzD3tc+X/7CUyAL4rU
EBuwKbpz64FnErwFK/kYHHPBIMb8iUnJvZ7OIuwhLl8Jkz7BynhmoCuT08Z8+5jA5Pfi4p8MLEoc
WStPZLNUmgT/HVwv3/FuOa/ucx341NKvyt6Fx+Um2kmRTrL6t7bLOqmdXPbiDTBDY5zNuz6Txa9/
ZgMTy/a2Lz+agWsNa1a1pMnKJfHIkVPei+GT1CGrrQBMkj/PX+8yLnAtyyGmlwiA8GEefyHSIpc1
HwmKlV9fVg2o2D+li9imSeG5YtNxCrTbKzwfUgWMSgkTqiUTyZVtm4sptFyvSVDVLE6lCzV8KH0V
vR3TH70Y+AFrCHzIuwQJVz9679IZb2Tht45mC5+UwYg1Qh6m8NzIWaGJ8Y4SZEzt5bo3kwYI+39o
+10kF2ugI/wGInbK7hxl5jn5oY25R2KrxhGMs27cEwqcs/vu/o7ryBgwgMkZHKNDZlls+gfBcse2
evf/z+KKyZhstWv6YvBEw+I6V7d7suzAfe/kWvKinz0eOZCcX/nMaxVJy4DO6O5JUSTwdAGBoW8A
7S6UsW5UmPtQhqLpF2OCVvqrZjYcF82pY7bvSe6nPjB44uFguPeoSA7pLvZQM1utgNqUzW2c8M2u
dX8TTScvbh6Asj5gkYh+ACffmAhM1JEiFOkC8B65MQmMZPa4g2ab9/q+sdP+oorFGGrwrYwEkFqA
Xy3Pkx6xzxh/PV8Cpp2ZL6Ym54KJF36Y2KFAemE2cvkg64KakiVTZ3BKYhzTNlpXPMSBAg5PVBDv
55ne//5MFpGXBkt6F4DrbEri9G5APVN25Db/EvfeUr6dzgtIrtmhafLGCCi3ZB3kBtEkBsLRJLLk
fECN0InBF0O24C0PKfb8WRx5ko0go4vprcBW95NPuaHv7JYYMgT0wxnDo2tfNEd7U017hiGQzOcs
wPb90SR1GMQaCyoEHy1ijZq1w4+uotajPusY2+qf96feeX2Dy056EsWsQYoaEJznL0HxwC0nQfNO
o8H5BB61yb0f6me8SMeoVEoJy23UfXRZKWNimhnhMDhOZtQnnVHNlx4ZNKDx6LU5KIdMg5D9GacZ
V+mouiIwdMDr1Uq10T/icBelUD8/RaSYn77tGZpSRsTzCNxaRiAJXbrwEXQeKvzg7d96TbqS+UIs
yXEkAmw/X1crXin7AZVV6V5bTuWrg1nrdXxdsq35wDQwRjbBZA6cicwJ+meFbXT1Sbopee5+1FW7
Cd5IONkChKxFLqNODcjEMzqBRZFtX9wbMLNCLHwVGg1tnhHk9XqpfblCPNs1jjs8DWnCVEr2Fjid
K+pZxiA+iFn3NCrRTEaIwQUefD+5O95Sz5TJQSRFcBNUje9UAMyA/RL3/qHisf5XRe6nv4cu48MN
Ovf1hEbksEWvltk/dnvS0WpLzsrLUAWmKJFjyd+8aLcMVGY24DekX/Sa4FHqKyne6bDBt3Ehzhr9
ukvTUhA0wwPe3EtNntd9FaWoXDIhIFcbm22IHyNW56scSyCXi4HayOYtUVGEiv5GpfyTfRVmbufA
D5O1hVO9LoJ45e7WLSHx2QQq1M/BP0aa+QNZWH88LRrUbvqj6UJGojpnYnSr32JJNql8/O/2EsN3
E4ONiotEINNd/Ph0pREkayGioo7EUc5V9M1Vg1K97qvWj6irrD4KvVgFEnDh1NsB2SwbxG5Pdn0U
z859Il5sTTQgZVAODzTZIn+GJfy7Febl1/ytp3B7unHZ/uUla55ZPlIq8b4QT8bYEDRhumNBstHx
AYxdArxfLsOpHNFLeiolcN6N1PENmaeSromQfl92ZH+sgkUM+nkhC4hJfJcPOBWFIF69HC4Z03Tl
1p/0xqEovs/OafplBkrxZLRsxh63qRX8zKmT/RoaIla8hUs5eax6dzu9bBeCr47WcGQqJ1RQWdfU
REgvHX1BueAjmc7pej3pODcrChXpkH+015einaW+hBhw0LmWDFOIbPlWWXcl453z4PZl9/7sDoa5
cOEsxjtaoKy2ET7Z/oeufaBjxY6iquE46+JGGn78396VIXmAdE9nQNjucF9OsnC/7ZRfWZueKvd5
TEyBnLrQK8zEfRwpQeA0m/4ae3JtKfCdNZebOqlKXsVUKagWfG24NSEFzB2oWAqWCx4OHtm4UNTS
/+vTDWf5eZA3zf+ap6ZaHnAY16tZ49v2SWR684Cll7peRs4DatNnKTm+vW5mKOFeh/8gH4QSNPJ6
aalf2guFalrPLDbj/w8U9wqszjBdQ7e9IPSCY+PKimpjfwLC0yl26wiWbVG9qhbXqABvA5R4gYVs
fmvJeOqEFXfyCXRwFAgwwknbe4NZHKumJAmu2F6XvBtD4qJ4wDkmJZhZsGcNnKGfUvi4mG5iQqhs
S2CQlpB+Y+tAytvHKAt7ztPDqpqVNnk6UMlQ3iMZmyqh7Xc3VS38lmVawe0XF1aypCGEM7LTdjig
W/O6bnNWIOhIQiYGTE8+fhlQhKjHXgNVCdycnX5CRmWl3ATkLRveiiqEZS4cy4HgeyEwNIjg8yyL
6BlnjrP143O7SIUTugk7C5Tq9IL/1bK3uNfB2jQQajmy3Tymo3CLYpYV5y0hyapSl6vvd6/Ws0Z+
ICmfipX9W9pSTi8Ey5creK0o13LFcCImG7b8zrIwzlsYZsLB7oJlz0kubfXzag/DYxOlTZAUeKDV
chJmpHnFhyO8ArOyOgTQspnH9fk/hldB+jVm/gdU0fHFijFwF9xwQqaREI9VCPBCwlIPPRX6ATU1
wNasNiqgvIIbap4a/C8nmtuzttUZooe9dwDOhPnbXg23W5Eu6yUYR1YQoPLnFvPZOFzMT5DS+lUY
Ya1KUeMaNdPDj/ikkS39IXFqZ3sxvfmbNGyb3TEBcENibDAOBFLch20TuDJvHpfK6CAjK67lCHM/
gQ0HJg15/il9TFcP3FSA98MWQEUeRrIcG81OKRAr8p/EmHWwpcF+h3TQ0xK+rxZ2dkasW3CtF1iY
9lWnXq0nEuNjgYOz/7JG5EFFyB2912EjXcppe8PB8vWuvCnocEho6TRwBza+9qZnxCihR7DMoA3a
TmOY2GzH8kjlZdLmuikBzUFQh7XjATFWsgShxXO0usyB73b/OwpLwKkzPnj7NHq56WEapMT4kdW3
ZgPt/W13jaVkYlGtcgZA22v27BYVXQ/ubCpb+fl9yMO85R2C0wTpnSfGx+y4zIxi8SBM4hQ4Borm
Tir2L2LD/dSG4KC2r5S3R6SqLHydeQiHK2rdydnK2FfMxSVgUf1UbSwQ6buYknjwZx709zUnx1P+
aFXVDTlydzkfRJhwnWLFJ4BEAaabWyS/RMK7kj+01AxykqEgX82+WOwrYreMnhBYyUSUIK1aAnsa
c34vA4bPYUm6ubXb/kQ6238cxnYTvgHjgC82ZwjqzmBekhVWMxHjHZ3hx0aGWzkuB07KeT+H3WAT
DBU3B51XkJ7iP0uTg/+aEIg2W+RoKj/1Gt/4UUuT35i9i9P8ByHBEDPEFybZ4NdkmELOFONpVuTg
YM/SvkEVfbSQPgqnXw9pCte8pB/zPPMlq8bXIOCR1lV4CQKme+KdqRKJ6aP8wudFjMSxJhrcEonq
DuIcXqGRXR0lrdxRHREQ+h/p0zVTIz66GLmqjeK+lgzp9AgsVpeuIcEjVRVenjMOtBgzSWjgU3in
jYSh04LEMlS7jzPP7BD6t6TyT6d4clug1QqVNJ4BXb5NUKpyAvSeltp39SAP7GRa4rfgNGlct8gv
TcVATLeOnrlOPJ0nYLyEW1C7RXH9aDojHIaPkeodGYAzZ35SDNAE6afEytnBEIdK+muyOQeUB+DK
9blNOWY6P6My/up0CSNa5SsagL/AAIZ4qzkqp/xebzqdDMZo9RPJg6TxIYLSB4EPV6uPG77efCKd
h9z2MO88XX1bS8a96UBGktERMYunCVlTsuk02gEszRFvZ7GqueRb4ktXDHYWdHjqxSbsfbTfh4vS
zRQ0tDuOx2SXXvzwl9QzjljVYjgZ0IYWb74owZSvhyyoySz/CJWo32CT6BqsZInCJJC0nvhLP/Ds
Sg2Brp9Uho6vPukqFZW1UhHVMNl3KUolnrtpDUSTP/0mcV6C7yFYxySWByi1GsRGS2y2C4fFI+ve
KKyiTOsKBaaIKTYmrGql55HEnpJ4ceEjFE6NAEFMzjE0BiAQf/FYcBTu+GEsAvPxUvMeIuPsSIGx
bRdXyWNCMBKMpvZCNn38dEBZAeBGhOPeB6OqG6QIZrwrmX2KvJpEC5Lj26bYTSaQJOEn5wy3WEly
V+P2ejyg+zktfcI1AqppFBZihmxaXvvrAU7rtufPIepSk6S7VxKPq7QOSBvKD2T2MOBZairaJ/eI
hEU+w+6nC5lHil8TxNooU+UxYNCjqH0k3OzW6koAbjCbMJAMw8/VkvgtgQyARVQiZPbM9dGxp+c7
OQZdk5yTGZpptpOjmL/QQg2JHnc5a5zdl6bAB4rponbijYGC4csiq5dhFXmGQAEuxVMaAd45nzji
ydnxAbAnEFa+U0sbPfmk4oK2u7b2Ooc18BGeaNpSlyM2PZQ9XfDR2++7jp8eUxb/FVmCSOoON6Xa
fYjf80mpiLsvytkjqkqPK8u0C26yoiAeLxCXsmnNKWer8ymonCx6BhDXK9TnFz4itNClSeao7c3l
Qv6gb05OY8KzCKD8NSXPUALqmHtY/28si9RQcKpYalHmVNVIsdFE+fe/M6gHyIvO3prGmBvy/bBP
e0D7ih8hMZ87o5kgb+1cCzj0Vt0p9R7t9eF+wMbDabW/DVEHPmlxSxdavgyF2YQnRc9Gs1kqMx3c
gW2Gir1DzG+zoXTzd3dCxde2mns/Ys0GfyZn//ho5NmaoY/sXu7VPgMnH4Q4nEbxDKWlha/P09v2
W5M1BHVgu+hJLOM8uDUwjLoMmRhq+okSoL+cK7HjVMWnUwuCOnEqjaxEn5zMnZlzaEOOpu3Hfgqu
GMetty/q+GBtXnkbquBBbB5PAXh2zSqTWcQgGE0UZ+Y/CB9Oyf7ZPOcKe3YXlhhcOZnIjdLbWmrp
gLfyjdZOZAwbuSMFww1MpaBd48OC+46xb9/Zt/PQq1at1hRt3xgucVhA8sM3p71ZMqooC4XbN7Av
Sp6+GLcPXA5k10LbVNWErN2/7SJSYsoPXf7GgheXIRq5H0WsActIVwIcOY9mCgkGnjL6wCihc2T5
susxfkn2yBvQ4bCws1fUPIHGKHArU3gVPbnr5a37z9xoj9X9j4sMnmmgzaWFuRSjdnawn3HHQ+pr
tpb9O5W6QVWCLR1Y1nPP6OjULnhC0wkA3ym9LxygPJXu13Iq+Uvbhv1rAiYIJ8qTAxhLJBBFFN+U
hrU0hhszoCtZ6g100F9lOgE+zuCzE9Yetc8WRs2kZXWhDnqyI5PCTBveGteUZuIa8S9bcAdI5PKd
3SDC0dyuHcTmac6oBbXC083A7lF1x1UcIPSGUX82EWwbvOIpKMEQhM8IsecRfQqcR/sT9e/g1ELz
jIOVya0JrzcVhE093IaLZ/ZCuDjYfaGiJPJSMbCyDfP7UptakSljVTUqXArdI8AMbk0lOhDd99Dt
0J8RRW5iFygt6cfZ9FrLvyreFZeKGdEAgBYVi6ws05OX9u+mV3m3FooHnkVn02j/7NvOiJyfUrXc
Vr6a539XI2wWl+kc6Jb15xEXKd0XK+W5rXpD3YT3waRFCS9dPy95n323XSxyFx4NP1wrFqBoweu1
IEUypy0uHCF/y/Ij5IMYGQWjck2mg/hkn0DBx6riqW3r+mB+CsfJJ5Ew/bMHHBsNw1fVkv2519Sp
IlciD3PeQ0ioeyHOjaQmaOGxPrx2dbvmsc74mltmTFj2QuAjHsaV2LNAF+RaQu592+nAa8pA5pSU
txhzeAVTbxPzH5TepDh2qZZ+Zbx5BRIgBwpAQ2S7MUBR2Uhq2LZXYIAeoHCjxZsFD39kMgjVLmbn
+1yTeXlQZSeoBwAU2BT8FI0wOoZ+mJGrbRiVRvsba6SfKlt0ohdQbf38Wa9qDDoW42FuRwjme2WG
83eF/TMOodG+GXkEqJFfLFOTjHhtXBLQIGX2oYnQNaeYhopyf5aWAecOszYisx+UxD4Lzl/qg6YZ
yaIxdyYMgVuBdQ8eJSXRNWTn+HCl5YE4veoVelIKDyzsvrrXo3GEJ7wrtnnK4bJvz0HLQzyr9ypK
e6mgygBRfGhlunbr5Vi18JI1zlyOJjxi56NOis7ooXqWwMKNuhPHwaGdsYli+LPJG6I68l4bsizp
JB4XoLabUQCI09zuw/IUO49DFfePJ3n7O95yo9syZy1ijd9gQlgIVpnQfRf1ZapPeasrf/O/KMgg
e5/85ZkJjdowVzRm1Hkk79T0W763JOQCtMc8gNMP+0oypZI+sD5UOQxJ9YN2emJcuRg/DNO0M1Nn
spzuYOaI0yT9CgTW+6vCfjDw4XXMAJVvG2TZ6Z1F5i6r4m6ItIJ83sDf8lmp8ijEv99Z7lh9Az1B
gfuZXlzwy//vQafuPz/dR8BZlZ7bG4FAitWrHOKzGMFM7R0kAwS6HESrL8hQNvcpfH02YdNdS1zo
snuFPnfGhGD15y27d9OAUDHe7Q5W7vZbRCBKMGkc7FupiS9ynmfWF2h47gz+LpSslDGLlx1podCM
Y58at/yxffqYf7Efq5e8LdAYLy8xqMxcKdLMaouSH1Gm15WyGLGZ8J/8kng8/hk+oGvmFnyaYB+7
CSkjlfcRISpe5bzNihrq2GHYsmJUh0OQfH5cVhO+y72rW83aW1//KOXvJR1nT8yvyJ7hK6azFsc5
acvCr1MjernH27EjM2C8NKEMhn+0/LVWH4D1mKd6pZW9pWLJ/1+R82tLzvUY/SNu/MqnAD74P3EF
j+e7c6iS3zeOGL8tm1m9JDwa9WuiIkkcwkyWNjsWqLFp07SZ0I96srBSodPvSRuWnMyxc0OiiyQm
QyoZMo41voX8QSbpx9fDbDkYScwCZZeYXMhNA29KudIiw3wa0l0W0doFqbwABmj016sKV+Zu7t50
U+cfmJ7AN6/MSzm5eZ5GaNSi2szC2zGZKQYOLhl+VYKKeB+NToQx07aQnpoFslDkTxOGPX3ER8oa
XWUu8QkKk8K2oiWaanc+WIL5E2wFnuJ74g8i/WhqFxGnkJfM6Zub2fc8tp61bFyTl6GYMm2eKFpE
+rGwlGvaRpeQbwkt8lsg/wf/1ee4bqHt6YFLMuDh+narUTkHRMTBCFVwA2sy5co/H93/oBPDb1EH
IOOmZ1ZGeG37oGluCk11HFxKy4f24/rnsoAfT4R9jiECIJaYNruCFSQpbRxx8dKFpwViNN4ZM9DN
xQT8BNrvDd1Ki2Z6w0d0nUxfrFFvXZ8SMtP3njikDIOA4u0aL1cjdIQb2FAmp2behg3WMgHkKIze
KblGW7AWA8Rc3ct9xu5y0RhxJo4E9jag7GdyYAU0VeB+MJ4LyOQVngAKjB0xevK5qhSQxrCPLrqb
guOyAy7bkY0vHEgmJRxnh2qPg2tjQ2B81a/MW25xHgZ4Y+B6Zz+DBJNWri4BmHm3DqdTbxekKNhj
zlkWcmQi4sTm+zuARQjNqcRWD6T1Pd32JcVgyPxW6iJfdzi0rYJht85wbQkj6V6jAFMllb4Tp34k
8LUjM+AMCKIUYoNjx8uC+5QJ/I/+XpZkh4RxhcCOIrUDn++wb8Qd73dM33bxb/v6PbAGWfA1gnRq
ycumZz7xzNk+b47713vj/bePR9UFtjalXfFCBpnrwefTdlOIOWqhLFsClNA3iVDAD3X4H9QQAhHL
Km4jd994eaO55tjEHKaL0Ex7PtG62YihH0iIRGGVd6HDa4jDGtIjgAPg//JyXap9vKu4Fv7yTW9W
Am4EYSJxjd9bpOBOFhRdHuu84fMDY5KvTnKlSrW6TJTj/xwF3NRdy6867TmmRjU0bsQY+xq55M/U
TdZhfVWTOAonBnXS4uUH3wRjsxbixRpd0jMStNWwc8vu+cnAvohspGDOwf+cuvdmuaAYyhbiOh7p
jkBC88sY89pxOZ0Of1XXhTeKwHKp23xkcnYgRzbp8BsRfDFv0z5uKW1/cwwPlGwGQh/2kOyZyC22
KvH3VWcWdoYv6/BP19IhXX2U825fTBhm0tXnGbKkUqg+vl6/+orhU9Y6W9b2NWJuN4Dc8jlLvXSZ
rZ3V/aWEsjaPrCFqzF3QjAVyMx4GmBpMEWS1g5NOuRFlAX+DnYgLCqGTI12d4qFvmWxK7mUIulHE
xhpvI9aSBpxaD3E2cSLF85nrljLxBBTA/loTr6xFyLZ8Z305dO1gZCEdPF12ixnA9FuEaF9jClrP
u9fhK9xaxXgONH0yoxx/PjfNpMzQ+MxbcOBhlCSZNiKPIGHVFf1VMexqwKYeShpGY4mU8jvgloRQ
HKn8r/4eZIGXanHPQdLBdYNFXppd2vEjcrLZ3QTAKJEPtQl82oIBYzJXWkoufyMF0POoWzRmtar6
sQ41vV4U/jwQkNpQV+D2FwwZ+XN9nbTCriKmfRvBpREzpagaPJyXPeo7WVRj4Re9DvttElQ8Xo8v
mWsYkUFFHjej5QwyEW0dainC+toiODjMsVLB/OWJ7V9QzO/3zVYTh3QrBW5yOwvfqCXgSg7XwLkc
5+4uex7OByxjDv66AUxAscXQbERE30l31JeX+D99MtqiOKvVMQYJFKE5BukzmRmsSGDBYKZfFWPu
x3LZ8rU9FKNLzOBQdn0aP1P33ZlogTZpXqRHp3CSUhpzWVkuePg2O3iSkMaLrDSVdMAQprkE0MFf
Jc6q3dkhD2IQEOBP0xZOfO5uUwAnvk6H0ckkKIK4zrjrh8nL1+tiT8r/Qe941YpdeBxsz63KE/7h
tC4jWsvocz2xA2vZA1ZubMima9ZL6cmk0ZByD5jqt9qo521T66xXDPCSqHbTi2pZcKKABPQ0ok4n
sBG29Bi9Rn5HBLEn/dIAVKj630aKdiuhtyCzGJhJdpQlOEKZDA2uro3drGdOl7GaWejtY0l5vlFU
CavbyEiC0w+K0uaOt+0Pgx8bU2rZ44//m5pdRkJT+yTqoZZeFk+DOVvtZmUaMMT81GCt26AfgfFg
xms1TDe4H6lbQEnurbMbTGcU8e1HPXJhkpzXVPBdToSEfUoTSAdWFpH6Bz11PLrv0Lln/ZFNyfxU
DrzhyS4NT6ZhGxNpHrdsG6iBZKWnAZMpHln6IzF6V/4CIGX1nxM6pR28bFJGa7fMoOYX7Og3OUdt
mv5glNQPCfnq/fRAsqN/kA1iLLo/+uttTO5+68IwZJdUWDkw59jVik21aZgUFmdfKHkDf6k45DUQ
0ReCCqs+ty6WSJw0qMIEBkPQFgGNAQQ7mgjZJH72+YMfzsn9Ebtui5zjONys2LXhLvdMUknj2Mzw
CnWo16yV1TKoPiIriNiqi9va2B/yX4EDu8gnZLgLVNJOoLDhhvWt1FF2SciySUOLeGn7Drj+pa3K
51UNHlKv1/9ob53CBZmspz+SJrsCMN/Cvb03dCi3crNqWGYvvLuH5nBxTDJUHa8Vj1kJUs/wMaW6
QzWCgMahjAhY7bPUGZ1WH+Cwo9fs5Zsl+IkPd4WupzNyO1cqF/ta/Ge+l2pXC7k+cQZCl4yNXqP4
RtrCJi1YJ52DqqOz4L1uLLiRMNEVQlfKX+JzOkKkifMEqKUmmcPRnZBib1rha0ZZ+hAkFZQ/mGRo
AGmehp0p02/BR7W4A1O7dlKVP94rRB3urWK58rR9ojhuopneQwKrOvOdcYSNRtW14QZAPFZOu9sD
83LFIyvSyrjo6kHjh/2QL0K1PIFnfrofTwYOrNiXsKmXl4cjtj7RwD3r+ySJopZQk9ITjvC/sm9z
9+1eL0fvDSQsiwAWu/evsOcydF09NEK7oS9ftPd2bRTunHYF+ihFmf4qNpBxVi8caUmHi7TfSCCu
sCLllEyffYWDm6p81s4XsIBdqErzJnMsdUtvJOSuBqZpiVbpnf1vdkcZv+naYQvUOjQ7qxhV0+h6
teGHnO0tTo14k+NcIcc2atKtDqG+C7xu3O6xc/lo3py6FweG3Pe/rxd7ADpx5QUGdl3xR111z/YT
rCArRBI/GVSF0qTLCHfiAbwFkqiXoLHSQnt5Zhe8j2zaHrwgDJ0h76RP2dBp7o0T/xwsmxsQItg5
UK3NB5ypJfz0IiQ6rp28y3WdIy1Ko5a4+10/8Ov+TZw90ZVymjKWuf8OpdtiybldFMgpZpGfUAxD
h0TG1y+VYCpRPgNCH+ugUDh5bdDFAP8AsPu8exaqpVoWW9wCv++fqpHKf+FdlDpPrMYp9HDpFi0n
1ZTxLyVAevM+e8OnmaT8aDIt/2A+q2nqva5KBkxVt750g74c9+4gAidhltzibNARWe38MpU8UDYy
7eCN8/4NjgK7emqFt1ivqw6VRgo3Apnk0IGaemQHK305seJ+bMUAqBOY2Bb1K0rW6dQenTkpujF8
h5QejvC8sgvs+PZkyd+O58BCI0Vn7wWFxOqe26aZGAY9bIQs7D14kyNQZlyK7tOT6cqq/f8vgJkG
6Yfxc9+Fat5yyby9pG2nuugQ9pjYrQhVcKzIWISnvDDERBcopV4YQqxXa2X2i1KJ0jmRqowuf22q
ZEMfbBSG6fx0MLcBVekPyE2wmoqWvlDXYyrvRrQgj6eDzOyCIH79cmryQ5jaK0p08AEykbCM2Ww6
Hk0f+i6MlMs635WxGv3tC2F8Nt0LxxOxDRWRZ4KYDX/RVoj2kI4ymUhNcdfrt5WwfFjGlZSBg9dv
z1CQVUI4spuZ6xkpFgnGGUiHOtSnCpnJ4CcJmLxCbsz2ib3deCWc0w4W+PMgFO4Srz/89T8XG1ae
RbwCJURA0VocW3oYbLkkJBmMhrPPvxQLOjAJ7iHyWtkz/K8Van6Zz5AVYLPTM93rWXxZuidyIUPH
sREJu6a9UonnP0TmldY3XqrJs93EmyO//d0eDtibu3O7ZE60ziCXDqOnm2ngw89L/TZl+ynY3bSW
ESJkeFiO2vsY7SSy1qUpZaeQf8eESx6GejvDMiYYFweDouAsjO3ZSyrRHpvTrHeF4fugZVHZ1nM7
tnZsS5ptVOqNg7ihW0I2uhtcW+m7rmy/RzE17bNETPZF7hsXyY7mtrCvfc6iYCw99hkQS8CMC+m4
fCW2mTRe0e/N6pDffC76stVLGwrvJsKmXjgvcm3Qx6gi0tlvjLD1OVxZZcWwIgaqQggGZgj2WxNs
YCEyLBUS/9Pw1wwTBkoZX6hY15BQZqcNuuhKPb2rWO5dZ0gZFB0pYZ+20BKFjeGRf3IxeyM+mLMZ
AWuERHnM15n54wJhtaXPKBhjj2wx8XHrqLqDEsV6JslFVL+pzkYnN/COuwkHC9rm05NWM7N+oWpX
q2BgMHy4IaazjJLfWOPBQuoiWL89ZP+01+ctSG7yn7xRrkKwlKudhLJoIJ2PiEf9MPx5SriU0+0Y
UQ+H6lUjNcRfSR7N9SFDcj7ZWFeD5ToNLSKhChuZQDtTD8kLmONl22SQkcMdj3rwZR4pUruvHwdt
H1GScMzmYspkZnj4tRWVk8JvjqrsTbvM4+ByDNVHhZS8CksKqGzXCusiN9osXrpEISfFADwzRWaI
ucEcs+EvPHWPho3IL00s1hyErT5iVM5H1/MPmvYoyp0vZagpmHsANeLssHH2UxIAbA3EJ3fKeKUt
VemKyPzpjV+/25ulqrvphd7kxpdfXXJr0nm/ABS5HUHMXRZAfPYAQ6rUC8OcqfCevA1KsttxL3ln
i4MhLR5vM1lNrvRodj2P4k1w9aeqmYYfkKuI85AbgyPDUftPioHcd5ra48BSTHGRPK8DUkbXvsx0
FxwZQohgMmc+p7eVrHeXyWzgQiQVjYryt5OchFGcsoHWr0SZ9Yh+rW4+bkwgoGnSekbmOMvmf92W
D1bdH/2gr5Qz7EuEavqVieVMkYVHu3Cy0RTHqv63+LQo9Di3gDVZuFXXGdEPgpDlX8QrV0EyDNUO
eSBNsF4jJ7xcPfgD5TAjfmkZ1x0xI/CXp8z8zEaGsClAKqHhSo3O+92plzzunZu8J//eU3a9rioX
9/yzzClfXB/4ORQ+dpQf2eGWaG95b5C7PDLO2C76khGy70xQRh1SOhZhRJK1F0cCfnG7GqnxrO9a
1tz3RyNnETHdq7xPaw6VoHaNzbjkiQAp/U10oi9riKx+j1Z4E9Akx9nsT+cmfC871Z9XPKT7d1ws
SFwXV8EckrMqxQmHtZMZmyBSRclro0oi6v4jmFwTxR120GwfaMJFH390/19BhprCfEZKI/cbnnKK
rlnGSrxDMssO5zo/vZPvmFQTMJEnHGYcIqaDhzjSYBZjxiIWUalb6avln/0XFSNwcBRzLVKydhMF
h/ungNTW7nU2NknP3FE6zDthIJn8hCYLpCC49G1mKqRyKdac6Qj2M1J5Jf6kgh7hOweqHhPFDwZy
aXGwdyUARlTIyLWAhWogf3/c4tLgWjoKQvZeQpPXzc96SYZtVA2NTKBZqKSfBLAZzj2oPIwf30Rn
xp45mATFduJ1JSIUZnLT8eCJb3OB9kLjfND/yTbTnfR4Y0WU09VXEZoTCRmJRGybUHlXovewDmRx
CU6ys91iWKWhMZbVgYza9rwjaRYONU85uvZgAay0L1y8e3YmUSqpilyh3CVAECmIbQ7l+qkCx8vG
z31SIorVMerThp6VkGQr3QUOnZMb8shTPQn5mpDmaUoUGxyBPN3Xx2aBOxcB9C7EYOQZCRcz6Byh
sUQoJeZYJZQO4kT0crxAPJxGEDd45yB8nXaItjFM2BM+QPWgP+O4GVeZubSyMaDNPMeLCC7IBXdi
NVa8novh7knVKy3bM3FJwGJFxby6XF9bL0gaMHc+FAiH2tnfi2IcNlVCU0LI9+e6k/+STuBfc5o+
e14WzzZQUN9/WJ38eG+S6LRlEYwRUEKHdRcbbh/7rychnI4Migd3Q2HpA99z1vhxSP049596Gk5N
s1l4S5wNu/q9cv7UjiQoRI9IcLxTKPFpkDLrMcIWWbHcLCWLpuz5D3YYtRGyTOPJRA1ccA98ljiD
0syzdUqBWnu9AsaaPGv4SooOjgmcLj40THF2WLqYiRKkOUWB5hOPQWcYQBFSYOmwQ6a2aOz7oKhq
1+ZMKO//31Q6IoxkrC16uTkjCi1e7fVPLJkvhCvG3teIVigLDy0GLgPBN4pGLVFVQhZC9msYUkhd
BiRZvdrfu3qNbhmuMMHFAvU9BY6Rag7eKw9/H6gR3Egr+DGRQ77nM0OVq+61V+JKEDLNcbbzGR++
m3Xr6QF+IL1CsV7JPHajgQGft1a3tv9dQ/thggleP+8C5e+gaExYXEYpjFA4ZMQdvZM/tmIe60CN
EvvpHJTziw+AkJ00aA21LPfD5YzUSxn24MaWqiYyUUk5oaUBShTvhsJSaSFeMwMew94G3C/8L3vI
doXHqPZzwPvrmfTV5YwynJSJyExZlmsmAQP5vzPvyxnpbWvhkJgS0dW0ucvBk3XlRaGYXYNraDNu
+Y6tseq13vTvAs3Mf/e1WB+jIvit3h7m2F8HvKkkhy1Rfmgb82ZXX2E5ySmx9XM+Xj3W4n0iBfCA
GjKTQvDT+BciO5WD023T1Bk8SrC3kG5wrkOPyxQQgCjEQkUzZ759Gl8hI/FjtbQ9nzlaY6bK6Zsi
/liA2uHvXtSOtvl2/V3M+LByvzipbtNJRrOiVzKLsX72tadIwzFXSBV15jY7o6Sy46pqsxGuLLAD
7QhFGpz0oSXUFyuTGFD1aUnQG27iRN38kYZUPBlrVFMjK+4GoV+wH+mDM8WKVtE2JZsQqi5zcTUo
YbYaayuViABsyDPUbA9w+CNqC9FkWPvIN4FJc3dWxVFRlLr9Bh5MizroOOxUMbl1xz5T4I0pgsru
3K+Ynzrw3xjIwerbehCzJTw1mdBhf4h0k3zwT67Kj/z8vO0vReq6YNpbmw/fsGbtZbzSbEM/ef3P
z909czHhebkSGznfdhNVySQOEvsgmTmqmzNZ1ziLZJtlSJjTqI8Nmy8e/HmYTEinqell1Siwchzu
ZcDu4bgO5Q7TxYwtM2Hl98IsNukW4dzO7dxHZYS2qamWIZqeWZc+chEqqpLWl1GIxY9w8S8PrXmG
Pif5MMiGs2u8ktYod1MqRmyQhKwp7xp0jcYw0latI+yZmeYhe8GI6jjIHAxo53c26aex4HWmw+wQ
0vqLD8A26aXC5qjDtuQROnlaV5QrPedLdnM27OziJpgWbgSabu0xqR+/nZePQkC8QnL3LumAbzto
9efJ466o3rXw6/VTjWgOE84R5xCuPgBQuAssJHPNVZjGlK6hFD+Lds/YU14OZdEpv8t91azv6MS2
3eVnwspvLF5Uqj8nieoDo58vPsrDqz3rOKltUbQ07C6bpvmAuZTodPjfp8ar2togVA1JlGYyDbDJ
J0DlDg3zR3yPMhy5zpLVK/f3bpXD3zDjmILF9cSb2qEXCd9cKTcan3aiLU7GlGgrcyRT/PJdIZPO
mdqUylmxuocJyEgZCQQJi65l3UValzZCh9p44k31+z8Q6a4cY8O8FrYdimBelLIldL9spP3Yki2Y
Z7ZfalTDTH3wQxYI+d0tiXMIXSD6vtm0ahGvW8VXE0WENzXiT79zngzCc+9aGs+lAyiGkmcnsm55
IwhD+enuIgwDkqqNyuyb27TDADmIQycQDu9KYtZTjDES0uw55b9saE2iYPBLxn7gw9OTk+ISDnVw
AwfvPHSifu4RQ+U02FfkUIoeKMZGXEJUqfAv0KEu0jvNQdZnLML5E7kWMLzSMgZK0cGouB1gkW8t
l1nGI3AKefMZ7w9zdnTAWFT0bcoOBjiXFlPA2l+I7W/Up4tHg/Y+hyQjwOxZ7dhkFM9F0xOpr1Ou
RJy0lh8xLDAbXCYPueISFgoAL//qkzGa9g5rzX3w/NtHbO3EE9rZ6/ii26tIv9e3sN+Qwi0vvtpT
yIFc6Rp/ujP6X4+1TB7l2udvImuoeAtvX5iMLOtR1oeZ6zDr5xscfNJvBzsJd0I7MaahMTuH2ZuM
+nB0LY2QW7J9sqLsF7NIDVhAPgjtprd6GnwXThDcJ3PSC7Ar1etbxAWC6oNKXdPv0EyTCU71BbG9
D2BGL0hKP5aMqzh7E1KwtLzo62VTF+P/Ntbs8Wi/MnoCRD6uasRbWti8hp8F98LOnYobIxWFst9f
JhouMTr1CUdaPNNerBk+DNHmqz2bWVFWK2nqqW9bkqUUOl6uGpEVhF/GxEFNPOJn3J7ak3o09Org
/leSVrWVusiPTSW4iL4RWC/TB9MW9VTzjRMZItV7LhWe1yNkyJYqhil5lwQyQPUzzdWygl+ePMU9
KTVl5oeSzNPR/oiP1/LUn/yNMQ5QoDa2T2gc695pE6RVNp+bcLVM4gs1ZBRgroFWOBXW552M/Jj1
yS2ROfFm82iMe6n0VrmNYpwZifQR2DVfGIyXpZB83UI1VMUPfdtgVPgon2QC7pIFpnWH/1IRHQkV
oVK2B3tU8eufl/xjnHou7PSpgadlXczfnuHiCkfS1jtcNsA+e32sPcPsbhLuciBKMLgOFBN/Xf90
wP+DAM3ED9GIgxZKz/svKqT1DPe93dZtRam+8vYUvu/rcG7XAdBkssWanMGC0k3gpc54B9cvH2Dy
P9bdZhR7DlOClwZXWsshfrtLLskxEltLBg/MtD9qUxPEnMvYDD8vmaBnmWu+/gS2EcoFnnDVNvtR
QwyqzuTIUvGY2veYJ6tdl9IUkLS9IPAjsj9Ii6SwtwxhbzBAXBqgI68XV51IGQRwZoAjAp7OPeuv
8ekcd0jntw5STzIuZrhdTHG19RfQbTnQvf3cbLdNHrquhTOtUswda1eVQgjwv+paeaKRnlpMOHlk
5uoGdhpmZIGaXQm5NCmI8A4QO8o9RyBm40zFf0mmz52YQRdFAqi4KnmWqFCCMyW07iwZK1JPWE7Z
l06BIRdFEfpm8aF/YoZDycSjRBMcKaC15xe/fgnxBtfReIS62TMlzpt3c4WbDOcV/aLJeQ95CiCe
K5wpJ5L0xQnhzB+VcAkg77BsZBVi08+GHYWCyK39Lm6FOStVGj6Fggi8nB4ZdrXbStL7mAhBUM/M
9DDvkdWiYgObgRaMtzVBetMBJzcYrG6yADaeEZM8XllXr07ng3lxKtFeihPQBDUa9rNFOubg7jiZ
btR3SJ2ufEbv/Z/WP/dFuHTv+U4E0ipjj3KxpJsVDiPZM/6m9R628M2/FFe5LNfD5sB1P0y0Z3v9
d5l9H7kblSUa8fSp0jOgiXSxtncGCNAvdaiDhBqcVb/LcX6Yj2GxdBf3wH8sJGI2iIQflOZDHkVq
DpHippmDVNOhcDvYnZADZ+36L1XSG7tkTOaOF99mv5AHwKJNSShbwAiWwGnjLYOAC/2JBds1zEPo
gamwlNVM+ijTtwEpF9lDfNAO7ZQAdlav/d/SsP7v0dnAtr+TZO0CZyxqU0CclANj9vtXGv/Nnkj/
m0uSygFDyqsG7p7LGouW1Wi2hxwZXB7wjrG5im4fRfobW9iXHaXeton8aObIDPejAYwaJSKRWEyT
+rlYWQdpg/G2/+AZvuiPlztK8C0x8nrxj26VPndoL+zRwecincnjQngo4HZOld1XxIJfwAjwNIT8
ulkcNLpjGm5/J4ATSFAAtk01PIJF3lLsJOpYYl3FL+KntubfmROHydMVvrIFCFMpL25Y6ScK+HLV
fSMBxTyf603wM2OpJsZi6qqALjQD//GQt9ZG8NVDwafKI9XH77DO8JaPM9WUrSMR7z3lpaWO4y3s
ZsIL+XHsiVzdQKgafcxzA86QK9zu/y6VzF7DdWl/fyJ0hAMXsUENC+mgjAt3QQAjV4G0KElBDfQL
lKT8EbUE7wFBBdJWTqhhe1RrJkEORJQcOecHZE5CVXGr2bicc822ohB4QPDFtwgfSLR0gEGcmKCX
DAH45EgGsgw8T8VFM2XCAqXNf8myM9rofnaiwrHwEt8kJkATHTMK79gPO6n9X2KfZCcAlsYLuA5W
1QTcCbUvJJAC+T1h6Fu/Jz08e/13UbQHufEU/fPwxf6Vk3yfzZw0oc7j683/LU+bSCriYbyR3Cwz
ldurz09vF9QkEKA6v0Gch7YMVa6IIEpfjlnRSFLHYO1lNfuL1sjbernWUOAbA0T68hfCPhMYSWVK
uhNDmtQy279OUDmhHA4z4YIJUwzhI6u3h6ooCy4VTlnDB78Y/N6/ztekBO444eBSvPVQg8XlCS7K
LdgEHjs/gE7UcJOvGNkh7X4z8LO/2EKbgPsvLuQX+it2uyqCDDzhn3NTFSByuKsSgt0FJiRJs4Zz
5IM1wrbpA5geKjHTJ5F9lOutwLysfOtgPndqJKnSXW3uWy3Fjj1wQbAsSpxPOU/tFF2ShXG6PYEa
gjfPwl45VA1rVAmuhEpzUNxLUBVR4hu2+YXouXm2+7d0XISxaKugIJiCY7Nx4LW/jGymh8PGciXl
KHtZCfNHLMXSqhSzjATPkfLw6ONAmYGgU1cehvneMWHk4IAmYuASPYk9wD3UuNIS2jfFRb7J0Jaf
KZ7hO5FPVKiRKK/cpdN9/ev4AY8EWBfAlqGUl2yDDQzCvMF0zA2wLc8Vq9zuow7Ggkmo/82X+4NQ
EnZ9bEMW6XrscvJ3IBhJRGKzvLWdqyacSn7P/SQpzy46VDpax/f9xZZahqVzxLDHI+CshFoZYOvY
3rwLA5z218mWPxX34wRSvUiGBvHCHnc6qMCrssPttd0nbn4LlzlzuqI6bxAerb8kSVSphWeWD+X2
WJUQDSH2okUlE3SYqHEhz6wkMdzfvdH1IEKcGVAvB3TzuP/UAF5Ydv6yI41olL/NRrYZd7wfRTBe
wNBRyboKEY34FTP7JqBYbyYhtgQRoMh7c59r41VhPUpp56GTjM51sHCLG37OOuynUC64A84E01ni
3+j4gzlw6lxk2KrW3/Lx3B5xzBhjRKEuLNkoQ3G4NZG+sfjt7Dt9Z8YdgpoJ1csJelpBI4sPfTVS
kuOVWY2dewQbk28PUQQ+f3OVBoMKuLRE/xHg1o/FCTmvVMM5R55CVxVbE0I961wOyYtd0clpDqjr
WuQJgRLqLsOEIBgZY6XYRFYw8embzerH+396ZzhDUWYxNMcMqWjReaYTmtoUoS1YGyclg6A776YB
ogLEYM6wfvjLRNVAwNoTO2Pt/xKFObALB8nCNthww3zIwSJClNjl6jvEn9Wq2xr/uJf+VBQUB3T1
UGO/cKAvTpmdBaGGJiUHOj5RHOU1xs4vL+7CINg/SayFFaoaRVEa89oMu6lMplQy+usli6jU1yho
mgOUza/NLHoZ4kDZk3dQ3QSa2zvdyha4PJ4Glwk6TfMrq99orb9P7Qaa18EVMydZ59i/gAlQQr/W
GWuLoeSik1Kaj5FonCAOlPwAt14oztMLZ1huw25f6sqipgo9/zR+cI4/Dr/VWtPtA3wxJd2WbYwg
DD43WXb+eMRT1oTcCpSTIaGHm7YkIgp+76bvQjXh6aQlI0ded2FyrMlo7O+nkrDWMj3wKfzRGptb
VbUHOsYzgcjXKV1H9UFkk621xHsSc7RUlXcZ9yEdVbwjaZxPpDTKTBmS8WkM+sNcRP9tkDI8yd1u
2cCMZ09ZU7/nnR1ZyPYDMN5J3TfkZcLX94ylw7gmucWXASTXudZl/7zEyYtAjS4dGwY24e+yE+1b
CEBzj1OhWD1PKUy/T13CuGcMCrHOxL+Z5MJhp1IXOMPorgfRfojTFXfcA5dqk5LxWOz+0LOwARnP
VDEJg20Xe1taqtaBGofheZlG3X967JPhFa7rnuShA0oGikbYFNFizpBbMxV0Us+U6Ph2Mf7z7UMK
yX3kq0XjaP0QHgVqcSlX5l5ahG2LYgtez+RiL4iRCcrwrzGgKyv7IbsMX+tfPHqPZUYvTpa0LSeZ
jK5gyJoQRKTFyzn0J0rNmnTtK8+7DxW+hCn3kqgRXpfxuRwBpWdVRBwqEJ3HHDeDmEa5s4h7hhrD
mdKX0T3X4IAgQQoidpNLEF1MJbjSDha7/9b9QEKbwHXidoOUvCcCmjWKbIQnMijby0rnYZ6a8QYw
GGTpVKK4jeeEt48AnHPXyRPzLaUV8U9xFlXWLElux7XAoWMxTo9SAZ9w0HiNy7ls4UMo/PRRoAgB
1rSSi/OrA9FjcKIbbdpR3AajviSmrsWs3H1c7mM5yka8NQ7SEfyQIm9cP1+O6WQEBV7N9xm7EGv1
pokKAehS/clcgOSZOAVTQYWaWoR6o+OrgIioIPD9JtQorgtbltuZ52bY23CQHcqASfv8uSOJCFKl
t+KfRvyY8Kl0M1VbaShBJQtcS0kBrMFARp8KCRXwL9/wHVIEo9fzA4/+UvwYuY/iHat66R6tfocY
YVzDPVAt7DpNROsOYOkJtdgSzd6AL5W2duf/WU5VfzWM63s4sy3TygGq0Z8cU1aVaVEivnfjLRbv
+pD6w2yylxIKXNz+1BcwbH13fjVr+eEUQpMBj78e3nWyqWtI6SIm6UmXlR9jX0VrF0spKw28oZdk
44F6hSbKk3wCHgZz646gfpbrn77z5YnOXKMVi8tbGuS6XcCDmxSfp97Av/3jm29XhngatkL/TFZa
01zW9kEccNmAX2Tbk1tBNflda6ifAx662AJ5BIv9yfPTsAsyQ11jGgYMnxSmJU+CiONVzA4fBqwD
vIbuQ1UN2Hmnrz4r2ZtLCbdZaB355t0RjJPoUWW2hHatJBlhEAL1Oz0xIYTPjwzb2+h917utkG9Q
O3IFDWI2tRlaW+CxRxFivJRs8Caxe+jXsjNJ6SoIn1dz45Oed2ZZPlmrJ/WCCsntmEN0+QCdHhum
lrrWhIDECOD9BkKZWmRLGs4Bm8U8m2AIw4qd+M+v/oZeVOIYcR+99LiOP908rEyy7pWHwX2pinDP
rGIbqUA85Kt9/qBUZ2EGgxG35vjNzwx4aOACiov83kCWAlP6At6YTXamHIDs6t7wL05aduycODwL
yF8pmXGaGwbvse0hWetPMkyl49Q8hOBw4FO+/AfM+QyNjsYWtkqTvoVg4QvGKmkEIYep+l08En5Y
4VJMxQ8bNokmRMOexJrpsuxrlVJkKJ7wWmWxHOQwdjERJmD49kBYdLcxKAVVWyca279jvj8MA5rh
VrGSBiWT3nrjjuctKPPN7F0uRclcrij4QIu5T/8bUQqXLgyiz6wGP4yvcPXf9Vzq7XLeT+/6NsSx
d4lLLibHYnEm0GBo4yyBohy/CGDMvuLFtVXMCGSH5D0rZVfl1q9EwMNg3RtpxEteqoNA/ISQ3rT8
lMcXj3enzaqCrS3oDvy1ATeMSKX15J+7Z6hSfKQb5vTTtIe9bMOp5SEBSznWZyQcXwDhBPlvM+Jo
HNQZEmIg0hgcXljc3iXyQjjPh4fnX7MAuA90umQO14mBK3+G0f9rI975qHUeRGdLH8VnZlbdzwCE
bFVWoUYzYrhuVG1F0997l1w0K7bgZBpNU+ftBfvFKdT+jybG2g5cc8dw22weDJ1GMhIxLQokA+H9
MnK5wrMu0zBmawZ9JqJmkdrvjBk25WTQPs3atbq0+ZJED7KQP/xMsUM8pf5XzD3gNQU/wV56beab
CLZUmy+WXHqKSwm2LnmHeZWBIxvJJ0BFV7/6J8jvgEczLdkUCk6QERTTGqM9spr+kQWUE7KwYIJ5
RDdB/DmiG33BIDb5FdPHdsYiAvmuip+bpoD8+/M/ZGtoZBrh//MWW1lSsU+Xfc5Uj/JBAGGvYL5M
ddbw3/MSIXOcUdYd1Xp03nSWzDiAPZu1Hg2ixH7rx3XeR3qqsCSAVeSGT3WV1gp9Y7VQCLEi26pg
/ArVus0W2qyxfEMfHaJrvsyXBY8rnrh29L5iFphWm2uTDSPgBlLqcPGRv9T/TXeyK5RYMTqmpVYL
CTLISDZwzZICTHQGnxsZ+Vo68vrNiZ6/4TMcnd0rT2FcxjTyVOIySEI7Bjd65LptwHDYxKwTXI8c
KksTMq7UqN5vR4bqSbw3d8jOw6of3w6GoTHWd7sOKsuqeJmgHEwsK7wjPQxawB0g1IurEWhnfup6
64w3MMati6s5qWIbKLHBE3ZgdIH/CZtqQdHL3IXaPxrhQVQVXKPIfAomavKTomrN9eFNPSvEcY/e
dKy9TVfFgAqhFgVjlqGo1Rk1wmNy+k1bh0Gf1GUbxnG3+hxHbJ1zZidpbKy4wf9WtqtD5oW2WIHv
ReU6AsohKka+iH+SJFsHlMaFMsmdqJWLAYXjcvOuN8TY6MwqS9758oVKgc1fIeorEfexJkLqahCz
/y3uoAPqwnPWnNN34SwBvvHnuaxJ7ZQRPyvCLy73lbJC0ES+UEKyaBs4dWDuzQUiq2DnTWCpc9YU
U86B8TNNNf/NnznjmG4wGMOZdvMzolYQSYTtgZIpJ0htuzWU9KOJrkGtTgpAN2toiU8lFLxP8QHo
RHkSLawfTOz8Xcq2EZFmhEdmyUAfqoEo62Vua7TXveasxdwWy/0p2g4l5UzIykTEkvU3pzKmT7jd
l2oE1HwzL5019ABR520WjOgYHydXFodZfN2PT5FdnWB1jboviIUoHOz4cqp2ksWldEPx2vqFijlx
RIvMtWk6FJD/N/Bt5CbfJwk+Atxs/emMJdDcN7g7ZpVCoj6mpnxuOxgyK1L7qkXnJGk5mbwVTPqI
9xWSuyruhB9fkTpSkctHVPKGQdTFtdZjz2ZXU+6cLnc3pSl8M67qpo9cWE5hMUOwZneK3ygoAfXY
jllJprRt3JNVXSuhS8pUnRRmnVUkxVmOCiqqbQXe0Kny6Kn2tjsyR7Vk5C9GNlWSyUWxdVV1C+lJ
NY6RF51mEEbM4ZINbsdz/SLnPRo6mBnfToDb86a6So9iZW51VnsC4E4x+ujOFiFPfegkqDk6Ngqx
8Sd48/oPHjPjehL+NQG0uy0/5UDt1bqWpnMtm1x0eVbDA9DZkIlg9b0g+7r5fEwQE80rWjTc0NgG
xPIoqAEWDzpJ00p2ioaHZ+xlz6a6OrCodWnWc+m5GFLgwYhPd5eRnWMZE0ptc7p6nr/8k1fia23p
0CMGV+ElBWA+484fjiJlUL90QNJdtFZxB0NInx7ds1VJFquv79YklIwvlDAMEksWC7jY8QtuyAri
Kbs+qGd4xEWCMGcrUMAXRCL4NMkNs3LGcqQvx+2hlEUnVECkir+IIL23ieHrgvfFHLU1oxZS70YQ
dBf6eXQ53OX6LtzzB11alUUcaK/SdSHJrqNBhV01C/ryIdVDBfd+7bDDSpNW0kLH+1zlvJsogSXF
qEguVDRYZ2/hxxOm+XK8yF4hShV1X04ATyvpxletxi+c+FziWOkmWSakxS5pEJ1BOMeAvsfxwE6D
1Nf9s1VNIO9QvmlqNVH8stecuBk4kGcxpQ1coEuT22WBDvXRzpWjPq/aSf6kEIO8JQ7fWNoCnVin
+Uyg3YkiKs4SYYSa/bF3U3HT97UUEIeftfmpCcRaiUzZoImitCDbJpb1OwxipgDFMpKS8J0ovswF
h8xJL2Ki5nVhgKDu+zeqDKKQZFm/jqMPNqsQen4aqJUZ+Ki3mdHz2M9yD/CiiUwXXcWbZM+4fGr9
gDpiMIoyPZDndLntcAqIe3nYkJ4HxSrV5+L057dqjbk84uMwKYdPSCAeKLyV28xS7U9lz8Glm4KA
TQqPOWiPLf0fO3uFXzWRGfr4quA3VDEVmkpPUfxDf8exxvn+TJXjD5/VG72qmlZRu/RqbjZl2mmP
V2+HWr+ZA3oeVmMTpBkWjKriWQtM5+hWYJq6RpRp/TbfuTiiEZoMzL5xkkjJVJ0FSW/SANrT0jw8
muCj26FnvIWynUlsWLIq0L1JGD1p99FkFhzGu17Fgu4Fb/kPUv5NL5N4sHUshacRcw8FOOII4ndo
gSqkO65UL3wilE8yZYnMxP0i+WQiVptQeomFPcs1O0PRY9uzvbamWimqDryUKhEOLNU4AEHllIyL
BTXWTY1D7d2m5CFJTpeGa0+QT4vESBdwzpMrdbFGUfpMbRoR4rxFwOmhDb1y94jrJgX/g+ICLwWu
Wg5/QvZWJDwmQKBmAWHqa5UD+K8NU+fg3kLAtbxJQhehkwDHBZkx/s5M595mvH3LmIxZMuE26XnZ
vp976ABWKnLmjOSGuM8Ld/1J0xP937ubSPRQP5Wg87FxhPPnkK9h4s/4YhCBHKhEXZEkCFcLUsoY
+31cRdLrsj1RFydlSmTm0dtNKPeAhfdNuuGRNZ+PHRDHUNWorZXpHLBK85Up2ysSVTAqjNqlZV5w
+8vafeUtP8X2dSKSVBOiC5JLHW6D1uoNJtNTTkn7cGD86zoKeaLlqS8dRLKQvc1MYEf457eMNWdg
ndb+Vc3IJxust6DMJhtT2nDH74hkyGl4WAqnCL5IMDsonVSzKsU8l+hhlR2gu2t+YhBwbRTdcU+V
wiGcro8+yCT44cdmnF0UuT8w0/2/owzc/z47mzAogG1oSSgdjfdWroRUi+QdIqlIY4azjgIxi6WI
l1wbOIzzNDw+kA//enO2kkLE6FJ1tt+7Q57nMilIVZobfrP9eHaqXyK028xWKj5yVc/YunCD9eC2
3DuhMecB8byHwbkJeCHl6n9tjPvsISdRYST/LlW9S9GuOCWo5xlAcZzhi/ZAHEGughxZHzgDsc+F
Yb2CZiG4wYYKfqgfn85VT6Ks7dJ4lhUKis7QjOybkFEb7rvMgBBXJ4ocJHjcu8ZNmNjA1bK0jI45
rcnWxJYBkD4F5ZI7xVJagh1eoBDouCC3GRA+Ro/JHksQ4CY0CPyAX8dupUxeMVFEdiLYFQeQGrfZ
+SQaTdgalDAEnDkMaUj5QPQqp7iqtTYKyFBWCkS8bBrcqHwrXpARtSa6GPNASt44iP7aLjLVXYjF
vRdrA49h+EGgjP37vf0KAkWh2WEnCLYYjyzsv68dCHyWcX3/udtpMBUSd0MbOZ5I1wYdizrZVtKQ
o692AIswuVU+2fqZ6x7UwQtculFHZ1j4BpdReZuips5PYEIsKaBNvSIU4BbTAoUDp+1/OQHv5ITk
s18ZYXB1kk1wU4b+SeHd6u1hX6vLwWPaYA8gnoDJXTPNde9p4289aPbj7dRFT1n4ffJOvbEgHQV0
kltA0+GeiRij/6jOQS+k0vs9Y1q/s5oog9ezluvSw4n6Qg+wMxoJlrQKWLWt5tqqUOOwn5QgKcaj
r2xV/l1q9435Ec2wwyJRSjLmWD8OpOJEEQsUQn37rTpLzsdD7ZbDU5oWSHYQrTAsuK14qSc98I+w
ZZk5AWxj8OMesYwyUx2rA6eE0UZ35X2vuTzni6LYzFnkzn2OObL3034qYq45e2BjsEkos1GVdn6N
72MOpbKiQszJavhbn65SHhimSEkJRPqRNbZrYTNBmliCWaQEIcxUn1aMPjrnYIZlX3Pp1/Y0KzDw
urR6fjHKYgdR08oTwPZgUd/2b5NANznex4wVT2FEM5jr+qwE94+0rZFBZ3KzGk7hU25Mw2AfsA5g
ehCP2wkqzUMIuVWzqQBBrt+jNBYiJPd87hs2oB0TD4PHubFUgq3cK531XGnHVEvFa3PbEH5H3MBA
RYbw7D50VYMD4pY+t+UYkf2Sh5e8SxOgZeHZGmDDaL423EUdP76Y7beS6KgD+ZbnmESM8RmPHX4l
zB1AWZEJQhAujj52qbHvR1Sbb5P0KdmlgJbGJK/fhXBPHN0J2AxBb5SKnDXwV7bDFsn6FBKErr2f
kwY4HXORN5N0gUO94Tletrkq7KHLSuagvFfAyx8z5o0pTbj1AYXrL4AKWG6EqEB3Ol/sK0Jb0XUF
9T4he9JMALKvsx4UuBL4diqjhi4FOj+rYrFF55joVYnD7X9hNaLhj3iXjrHdK/dBscm57vEyjE75
oXGU7YBpCd6AP7G2dyGb7nMDdhSDlQ3tiszbU3db75v17dSdvEiMYaaosvNdkqYvci1/wTG5Nou7
pOrQ6+arMVOhhQzC9jsgZy724DVSKxvL4BLvpNaTDYrjlMys+4jkCsleioOxjQQzhizLkJJCP+Ea
b2zfZnhFisP7vIfOu+DHHxxgkOIeesUmwSWCGj8xNiAx39ejw/D/shHPvcY7bFYBkIInOM5RH2RB
GGsSAam8IwYgFOfzpG8AWzLfVWVHKIIZjjoT/PqA5vzn0qmYBW+o6Cawt/WpUVViqe4e7EZ0NHWH
TFmJcVqg0AlJxnUoqDOXTyMkch0CN80t36GWLBfL+luKfaA/MnyqAQ6fI05DM9lElVOgEtrjbN41
JlrLHPLrpLe0qta+Iq4sxlNlTTRrWDsVX5gYZ/odG+oPUkbPs/U/3hXIErke/EpM04bC8bX8CBN/
ZoyXGmxrAhNIWP2VHpAyu7DiQ00uC4E3hHWwxwpJArnxuSGlCYvYdMqPKVv+7+vi3r8SPjM5i5dy
MShBJRCK+xONXrQIjcYIaZ2FCisUqVGpea9uXR0SOaiVJwT7HrsRhV9oLuTfJHPtSBA8+hqNRXzg
Kn/UvUMBiRR0XMvuJa1+uKlCxpUQIW3VHTm6jVO9WM8k2DK0GrkVJCWEzBt52MedSeQDZVIN7/FT
+aZvou+fo34nrgWE4+OMG+SO17Heb9aD2t60oKspG/slPypfzI/wUhz+MedywWz0vYTOC8NUJaJl
Z81nj1cD6IpKBo/qVlxKF+TeRbArvlIfpVzm/j0iLejRRMSCbC/vFYGsdRWivbvd3V1Zi4lQ98fv
GJfRODOwnucJwzYP9B/OEdChMJJyiqMiLPqAReqz5OFUcQZLkURzB05bFu9slZQpLywc+CPJ6dyh
AA66WCr2u0dRqq9b4YV+1kuqsGqe6cEfWtErms2s19Z8TXbRvueEaTng9KE0LrvN9GXbCtlwfRt1
lItGf0Mh78fyZWVs3ll69QP1Ijx5m3JlEo/tSZjuccE5gzJsyGa8mHMa/afms5zFDBTq+Fi/LQzS
3uMwWI3OhX3nsMaHrPj/KlUUhEY9+Z3e+L7DWHZvXVAX0COMCz6S1VWPh9MZ74eXgw/2Agfihtcg
1xvMI7wpxvfSqCdSpWPy2mtedmGoc//87AdKBcG3rzmMDJeR+6PdJKq5hEkKajn67b6fq8rmeQ5S
cmT3dWswvj5ZCmidgbXJ7BbtqizUqL+HEs0Hgkw4JmTQDDiEVNBIkuq84Ou8VREhg0luWZMRpioK
HxSKSg2YdCSf+3D3Eiiv7Ch3omnX6Pbdllw5CZ81sjRpM6VFzku7Xlg0twsoDSSSGnp0bF1uvudo
gjmr4908ZI5r6EgGd2tKvL8pRvDQQP6RTta+corAKwZR4gx1IT4HyD5vPv1U6y8TBFPEau75UaSQ
Oe+TXU42CuOPt1UX8Bg35dpuojs3XYXm5v+AdWpyYw2hIqbiTJ4sEPIKo3AWwaWpDSNcNFLgFdkG
k0xWGYhy9AvGRHJctWdriUnwjbsZbY9HjKuSWXwEfVJR97vy4Dhsln840C5QQJ66983+hnv3xpIo
5v8AOe+sGe5Qsv2y4ldajKD6z1uf8j+yS0G8hyRRBpayrRMdhTWzv811X0A5Cy1IYD+VwlrmYDkk
c43p+tTHWIxggeI7rOOiAJ0rjwA6jx1TKNjHMQ/fIft0QzM4vKUKI2aj/ODSXwTRuvdnGTFFfIAT
VH280YAk/Q9QTkWaGSAoemy7Ex2uwfrJfJKZHoh9FNNUWFUvbcYZv2Q9AhyTwkwAEZEi7DA8uaLr
itbsIDDsNmW0LZ/VaFXdSqsfCzwWsr8oReOBdDUAh+VGgSI/pyG/lBnc1YbLzfXQ/ZCnoIK1y+6m
u23pAQtRB2qdc8h/PIJ/Q7m4o844dCq6y7ViQ1+F4a4hxqbvBT4cNHhM1mHj/UTrjQJJZfZOYiD0
8cnIRRAUWLk49bVgR0cI8Y8bXKlk5ckw6zvr3ff6n2gh2LabXUHD9Z88sYlJNrAijdM2O0Es3hW8
KffUxqJyn5LlzN+XOppAbshsNzQCKPKR///vJTYxb5hA6rutC2TFG/kHSxZrqipUWY2fNHsmnQS0
kDjBcWkvh36XWKgSwTBQ8d9KejibZqBxLIkIcl2ea3kPszFaROTTS4k04d3EqiAZf4/k8yxqTR4F
qEih04tgbbzu9KIYf/JcPNtg3BeyCVJ5qKuC6QP+GICuiL8RovuRgWd41FLIfBhjyEkI7qktsmiQ
mb/tzBe+mwa/WqLz5FJ1O7mNqIao8tK7drAsOSjMHveCxfQFR7ppUMa10jo8yoRVMmolO6Qc+cU7
TVgEKheQYJkruLmdg1aQGviCp/+lRz0IV/XAwJD5GZUZbl9x7LFSyC5jHqlYrpxVj/cM+a72MXw5
FEkfmnEeiT17ltOzL0tr8zr5000xFHBHCkJR1E+PHl/iQQW/WaF39GfeKNlFDGu7rxtNUfFrWESV
Eyl7sAEpoi9QRsDa3nkhOiQGfgGRQCbTU9DgHE9I8hoj/5kM1i17xK4CLGTXZBtrCMmzgimwrwdX
16hJPdK7JQ84Jl6lgfBxuc1/Z/fZaKRu16aiOYsYJ+ZB9fNN9YrPv0Mm1yhtwmBZbntXflNaTvWt
YeVshh5gWF/3zkcMjtKUvV1JgTcAOc7JOQAtFxJgNqTHWiSWIrh9ZSfAUWcLIGM8tpUFQyeq0zxp
V2d4VhEq+kRhaIh89v13Nx3IZQJT8W+BxSEiceyR/lfGXdaFTc6za/7x0QqxCXxqgN1jcTQ5uQj7
QpZTU4Zz0uHNJMpUzUjuwxOGf6mHu9o+Jk0Q+TMC7hF/db24XlRILNAOopNHdIPoAdSPBzdaFzEt
kyFgkIkTOz+oaOzh/LT27Qiy2LFJM2omJJBYGYxQaI92ue/pdkp1d9adVNAyFAsYJrpyIsKJleYk
48GV0brpRkFl9kQPaz1Z6xMY43jEgqzAQUlUX8oYv++NCiTplbAGjWGI7fFx6nAPOYYQPXkyF9X3
WxCamISXQK8pnpughOf2cbJDZhlTBuHlF5baP2UDako3UcUDWDHIYZieesrjc1NVQMYQpoQeTRPE
845RaUs1ZFQh9tgU8faAKrL6DLJns3ycNSvkDdQz/OSUG68i0Ol3kQnLguDsjzTHC9vUIR9eev76
NUPRTfEDvpQEv5sfn/kysHKd5YAvy+ZaJdD06zIv6YTISMWMwAc8ZbZV8EI5TIumWq6z1toEQ2qQ
dWVgYa0zGzCykBseibFSgXj0fjVfoUmFLpZ73sxPxJcL7LqBKMMrIiAfrpEsGlWW5OAG84LPcdxr
efOsh+6p37hVM/wndAfd6fFMRfKd8tobPPdJuf4dy+NDCOCbewZECrdjm6JBkXhM65PIKNore/pM
7Jh2USeaY4ASBv3DaXFhTc3FwpphrU3KAztxhm/YtEGF091FZrP9Fgn4iwA5YrEiX/s3rBCIVPbP
2b1vftvs5OVFByaiDw6HEGMKeffScCN9PN3eg8eoFNmSCG/Y5Ve4aKKcZupi3hC7izf0qK+gjeC3
e3WueF+Ntl283W+rMr6fh6EsAhc07S+a7PPPNFewck9g7E/BI2C69IS50SK4BPnaZvZ/vyUkLMxv
l3DpvyfEUkPPTrvytisGVD+THLryrTR1Y1SUDIZ50vZMNfY+2rc7JLZ/rUkssIgtqgOR70PQ/QsA
DOCQMHqv6UGNvp3hca0ihElTYBKavGXtHh+x8kPYEuwPa4OFW+2hJkNUFochiR9J29avqa6V5YAg
caH7YnHk5IEvEn42SdU7tmZAxF9DkESbRUN6RRIHaVCZ3g+3SVeprA1fJoTWUAWZkUq+o8t7kKKy
dnR/0c4X3aT/tGf6FdJu8ghxmtMmSKGK2HosFFB3c0GFgZD9RfrZKGFz8h5VKt4KQw3zgRvQwa2W
cB14QWGm7dzLmjFCtBlNTczkP9UfyoezI1jdWKkCTRHtXAjR9pXgIt6u4QkjsMB/bfj1aBcDzDd8
eWGI/BQNrp9o5m1P2qADFdoBwuLANDzcfFzb86nFAM4n/GL6QcEoxYYjJgAeYSG9yvcZaKnS59An
IIDFY2duaHzgD5RDskdYo+YzqNsDlY4qITjOszCGRssigcL5F2lDl5Izl6Wdjjr3aepjJ0YdKjbC
3kAtbAShJxIENuonz2+jh+qM8ICl/nRwrJum2aF4VKrKU1oYryrsuXKLetwar3LpOCV5Nkp/v2E7
78VTkYXT5IhqDG3wBxV8fS22pyFkjUYIbOufRQ0JljsF/3fjTR2XHb00BF19qQ1rvAQ5cMd5rCTV
MbeaStnd2Udbsu4+BE5I3vgzo3/JXaTFBYuQOfVfoqxXb7Z1I0hn0POQb2rTBG3L353WFYofx9nP
AUCx+Xbv8Nu6S8RcDB78ZTKZYFCPc4bRJW42dU4JNNlMIQJM7Tri4z74KIije56CALI/NLorZo5k
QB796GhObzMYw8VkCHdtRGAC2znFjDcpHZAMnhqz4NTamBcPrWkhm05rKxzgAj3cjV1QTjyqlhlh
HfzVUTfMkSFSjpZpi0T82M86X3Lyg7n7087eJbKV25G3aOX8b1fJi+RqeY5bI9I34Fy/gbMVnDRk
AP+kb8h1lwdkzqezjVAOw+lqKuhN6AdkoM0PUlBGcZnqwY7VGjOk96viKTXj/bDxhNEBhHXjiGHj
HovFstZzVDJA4VIbjbI91FY/jnwxO+tK6t61rF5gNbAxhhKEkovRGvGJKhqQg6CVT591K6ejOtla
5yfJw4TNuwy0sw8lgT06uvnndN7C6qDSEAxKpbjB8JzOr5eeIfTuCaptf+xkKEtXZwzLErCF4O9L
3RLoGD/E+oKTFg0Rk5ySt3KwIirydt4Dj0b+LyLiCXDzv2DO2XxRP6Qls1so7kNdXA6a+6u/Tan4
J1Fa6ceCB05DN4U9Au798buwM2eeZAyl5Ai7UmMRFh1YD/D+1eks9V5f6Op6bQ4ktsHtChjh2rF5
ilTep/PU/dMMkbDovMHf3JQn5TNM/PBpLt6YKDtcuae8sX6/673dS4AHv0C2TesJWuREaUW+Lldb
Gsy5J468QUr4bdCoMGcf/F5ZWv81AVEVm698Y4v4q5FgjjHXLA2ImcIhj8mdoW/a8IILw6Ru3l0D
7JOQHzupRflVTrlGnVYBKEflilbx7S3T7t+AgK5g9c6nLXi0V0VI5Tt3QZaxK9rBigqv/W3CyHCy
4rsZK8KwsexAVIs7sMj8l71DSJWgOqTDjP6tX4GtnBo6jj88VDPj2ENkopY8jtPnrZMYZ4598nOM
z2/nGSF4r+cBixlKCzvUCVqQ87KY0ogj+iGQOb8DlBV86YxYJH7py9wP9+5smezX3P0SsNobmpW/
hcIpQAXUNkqwSVDliPPeQ3lNjfhAMR/DnDhpqT9aMtAzLuDSA3+sj6blXRMvssz2JHB8Zvn3VcZB
t8rzLWkxToIjd7pAiVs2m/UGMZte2vM/vNubia9/j9trAyo8tDJ847eToKJ8HnvMKExN91tN12+i
vVrljjxTk3yyHGJm8EXhVjz9rTZJojUq/BkoOfrK/eNRQrtJidES/bg3x88s19vYSnLhlXsI9B6/
GB3fs3J6Ys/UHI3eTIfpBghBgCkBhPWCInufiqgEvT3NI2+0W//XBbJcGh/DOyU7oUQAnvLQCoho
v+WJsFMKMJzJ8CGxRM54vnrFFue99stZwjZnJUVhJW+eVg3lCCexWexmBdcApDfB/jNWaEXM1EUF
P8fNfwFeZPDZjFoPPctXhejn2UHmvUDe8ZlQTHuo115Q8svrjGn0IKdAMYY55PaLtKPURoxeYrmf
F+UQNCeeMjJzLarUDjFICP+fLm6RF9gmhuU/jOkuOGZekNgb9ZiIAIw7/nDvWQALcawGc/57ubqV
Lv64MQLKr3Yk4beHl26vqVPq3ToyD5Mz0jGeEbqr6cUkT7jKlyAcZ82TlUqV/91YKbu8ZlIV7Rcm
cjasKaCdhJ19Cm2GaaK5U91PxKSju+v96XTlU0HiZPZbCHC5FTfvCT/102jA+mWEx2O4C5O+Eu7O
yU5D7aHotzC4tpKLCJN/xAZJf3se0CJWNQRWAOEkRgZ6MXVtBrlFTr1nyKDJvI1vtiNqtg8zjA+T
EyW5yCBeNdpYLZBTa5QEPatl2VY1Eqj5OU+L3DcGnou4Wles97YR4/6/yymtvzMCWo9FfNDht2Mp
trzqXg7TgzkwEQJNpOaqwGdWCGdDeMBiJYvsahBPw+pFTBp/yV7glWcvdqLs8Ggb1liPJfkB/vsZ
/MHWlVfEQudfHkGVcqlEM3+Tv/PczrKWU+7UhtlCU0FhU6lcqoQ22Eg73d4jklnnE3kJNfJcgoUq
wASMncP0quxujT+7ILtC9VN/I6CkjNV/n5LBLIrIOanEGXPoVrgt3fLUyDG1ipkq0vvMGLp+87qA
m1t1rIM7UrMLHO3rfyRJ0eJyfNQZj31ZOLEiHkDjIodBsFxgwU5WHNLUCBdE6yDHhaNQZhCm8MoJ
dUfJr7mKw9u5EU9eIMGWh2LS63GMij6EDTD1W1TtZrwfkhDMAUMVjuBi3Ui2Ht6OJv2L2j1CpcgT
YOA8zfJb7MwXkkLXXqmtatwV1LnmQf2WCF1M56z4CXsavsmlNPdXbHLKjIn3PsFb9MOl6jLNthG4
VUn7YFnbyUD0b5tXnRxVu0YcHW+gI7cVIdwwBG4a823Y0to462Z8zbYWumdmJRsFOlkSBie4WXTb
4rjkI0Pe05oTKcU+rkJrEykQJK3bLMq42sL2kG0pSmZEynCZSRKRkHUIPrDfXx3om6LFMaK6ggyg
K1o5+kYEmRrBm0wAv8g7zvI2zCi+EMeO4aTYWGDvC1fLj+8/HrMjaUmINcJNulaI0SFxFL3m2sqT
LSxenrQ1WUwGgEiKtOSVc2kWKhJl66s6WYjrbGLnUtGSfQXovYuJHEqOX5BddGkCPPqnWPDbRKnz
9zS6qeymVKxNwG5EwyDv92SmrDhMviZrGnfFLYoQj9+67aijIzjZGLVAFDzg7e2nLsTj9HeLa4Vc
E1uaadUX1CRrDK0/J+01WvRzKr0E1YpW5Kdnfon0uz4QRKceVLAluWJ3ehAskKSb097WsbD45j3c
ZtU1uZFu/jASsgljIpxbmpTT/A5yTvreZ3vwssPKlyrVlAFpuv/UMCgk3Ro28QP0I61i+wcApzyZ
09n7ia+VS9Z4ZpAxCWTv46ocB65OjtzQDIc84LPMmLlkyUfEWSsGACE4uZf0KXHUzChFZBgYM0jL
jWOlUZ0zCKipiUuKUS/IFKB5y1iTu2/vQR1N394OJ550WmFsg/AbXpToT6yUyQqXA+8NNm6vwFYR
5Ae9db5nyvJokT7tBpVuxwKl38IQctbJrGg5LAWrq7H+aoiOxdepaQquw2/ppJE3SFXSOwZOXcCc
K1o6+JAMVsVklEMxM6yArhI6kI9TcP5UVt1Iz+z2fS81ApVUU+iMo+jlYmafw83eb5/FXqsK1KYL
t4KLMfSlloewjLBRygG76vbcku8g0sWIykmMz6dQXfbgIwJH8DGdMy8xiOznGDPpZt53QAmg3pQE
AZyf9FAerncBFZwbhsLCkyqqoPQWRmc7CNI4Wc8c1TEygPlVWMwm8qzGSzDjQ12XzmjV+6fRgcLb
GtLJcAxFi2V6AX55MFbl8S5rFGA2Wic5uHh8LufB5MZsovsX0FRV2NDqCwSfwQ4jv0QQKgE28Kvj
VbTLnsGw9cTUdfkiOOK7mVFkB/LhnQrsnvA4MG3S0JVKjbh8WIttx61S25FDCMkG5i7W7SEIhlB1
GPXBmtcx9f4rnP+zHz62eL/VMdk2HXnwZT3MwlGWef4Vcnx0kLHvbralky8AsynoC+bYuwtAh4HJ
aj6dEzQbWsBolG0h4nFUlIy6pxBQP9dKwjDj0amydwY5y52iRJbXT5iXzTOYbDK18Fw00I9U/57B
TO3FWHC0yqL8/ZffbDc2QGrZUrRmDFH1SfzHVf0Od1/jm2y2OycapvoqtugEK4p+7KNeTKVOQlvn
GWxQO1RvopMFertZi9Yveku3oxxSgC2lb7DBt2gFgEYggOmRFH76q2ogxHFgRHrrr94xb2X3iihl
U9x9jibzHm0/70GMUZ9PmJ4KbcKVpatPB0X4PYg0OLKCum5lZ8JhkczH0EBeb1QC04W3zKB4wqbj
IGqA+BeC3rTOKGdaqxqCsNwSlWGk0dsGArIau7xjtxHXmC9jUdLnQhYeZ5qchYIfmmT+oG4FuuOB
+Es8EOc+NdbntdE2ENYwKN/dgKhTENXGFA2MftBtpn+ERH1yozIncsSYtlyuXNfxhmImhql4VR5F
VPln43ggsOUQjmjSJRVNqewd5RSjT6aUsAb+EXW7GIOVXvkH1f+UjaMc4cdOCYa2focr6WzvItfK
wmvoXVaWPFTJcDBiZk/+WDk8/IyqQ2oyIbJnfAPnHRmZtTpujKCswTvY07LAEt0myZ5cQT1aCiuL
kpglOAIJKQEPUoPFIl0CUziJYkBWbCxJ2pSxLzTRozcxhL3B4O2TvtbLvGv1AdGW1TKjvHL+4jNb
IdjAunzSsl3BPEao3G8qrk4MnRs1WyT1mxFvtJWw7A2bOVZ2UESr3+BJ9ismiiyAub1L0nHbcfSy
KMrVKErDPVgt6W7fV4GubNFmxgjGjzUeh3eY62UONL8ZJ8O6QrHEu1CIEHV+7pn5flLU9degU1fJ
6XpcYSVq4eQV0pyNZDf78i6D3Gp26p1ouorhBBNLGVo1xyuSUrJ8LI09jdemLnusxuocYsB8ebfZ
DjFbFZjjf9pPJ4MQOP/x/SdlLHZv7qJK6nSk/uZTvDAsT8e/wDKa+XsYiWn9S/IEr+f+sE0uCYDw
fDXkYjld7873dohMk97hZ79qJTXmN9SrMpXbDnofLeMpKym2Ct4kWUknXgfK+aDhX5XHpyqolgK0
+ntckUv4YobDbljLC8xcrChD0dw836ky3HB0AnFBCeMRoagbBjWpvncLq1Hwbq2BJp4O0LNAjzZn
s7VjSPL7wf1gem5eNWFL8ovyOK1jC8dJaN6Kd6lhR7n5GRUm0AOdRzaoFVs+8HnTZMaRYlMMZMK2
uJg30yej18QbYItYxHJ6MOSAdndkl1vxSTXdUQ3R+HrPXKPxRkDufxlgLNVB83MpQXPecC4iXMZd
DYxtjTdAL2MdK0JF3hdRCUyMlzhGQm6ScbxwiBGlYH07q52u4BpngdadkcCx5TEHZer9cbJsfD/7
XygVA2b3DfSrpzIUuFckDf8Fm8QETCw4EzhdiBjH5GqfkSbSM1G2X+PUb5HlKqNp4G1edqo7Btvp
f6q4iFUXvljcaYhcVXVgoRBEaoqR+8WTEM6pBlkY2ayakXhM0reKUlHOFHFxXkPAmBrCKmw0Jq6O
FlHsiqIXzaX/IBC9Ur62bzo31//5m5eqis4miG8oiFqEAWL3V4sTNXB71EsCQEHGai3KaIjWwBHW
42DahFIwJwSD9A4ZCbMzlqeSAxX7ABLgTwdWxbBh1G7OHf25UDxWQN3P7Ttn4h6qbwC3roLSXdrk
C7DFfpq+ng812f8N1QjGr0tJEOmcAy3B5kGBGsxuWjMD/EFqO8blt4hYDKVnM/hioB+QIxvTOLUW
gwUE/GUwjm5rHwnsINwMJejGXkFjSz6bbWr0nH25ERHHDsn/VzK0ahXbh4edaYVa/62Y/7q9eBW7
01adlfc3Be7lbaa0V1aSqAoVYJT3VwS+mGSEvDgmbrOlyx265+pJDfDBwj9xxHmuAHMgyRUOJ/7l
mOyud4JVhUoEl1ybPiL7gpp5xNKpAdN4yGWNtG0T3WY8uIz6jB1Y6tUTWpeTzUvK9s1Mj+XHH7U2
UNv8dls/i6srp8TUzBXOIRD946ZvxjXlXigS/OQCZ5q3cIAs2/7m/oHQpnS7Zjj8FIsbEvzcGpv1
jjpP42jmN+rvYAOjAwcEUgEZIxbh7CKjQiSrPBu2FzkQ9kJIZh6rRIxpSXIKL3Qd2wo5EKtQvvFN
vEyRl316Bz58RwsnrUhMLwk5s1kfZgCLoOAV/lTQVdbPWghVmEXtIVT30Dwqgza0r1ghFb8Yd9Zn
HW0R0LGtLk+r8rwoKW9SfGZXEglhu5q/QV0C+fD+rkXaWnBvjsJDkDvrFuI+cY4lt3mNm0krQL1q
Npup5rA/UG5nz2hz+6R/Jg5B8JiHmC12VL4sPWy8DSXU5o4bg/3RCwzAVihEsLQPT5iDudIfDaBw
0aN/FLpSL58/aVAkHjIqj64cfOFXIrIQZaGLKNv13tazqF+1XlUL5gA1/QDeAcMTXS8iWZ8qwSWP
8rpQwDheTA2qzeQjI2v7vCN5yJi+I6z3mqYmzxfAmIdMwMq+R4BWzeBIHVInDWPR4oORUoSFk+WL
xVdskvRnuXqlFyodrZ4TmEbrHdybA5Wmnwf/UrFjHnJjs0n3pL9VzEewJA1+L9LPexijGBooG7oM
4wt1dAx01BxoPasl8BOLOJVT8FKwF26filt/869zMI0laDXLj65Q5uhuvc2TjXwMJcDWMIHVv/29
0tpjbSf3wT0VmGly4JK1GbOFHpRIVSQXZn4VWxtK6UYJfKLqXw+WAHJoTLC3+tuu037zvZhe4WdM
nrw35dV/PPjfWub30BEdlW9zb7grvxVDg2sQ/zNZCdWkZ8M5u48mPItDgW2FN2qra2fTe3T8b3fZ
QtBw+3NNvToFrEeFqu+/GKDpcnmSApGFJ8WeCeWtiKFPfYR9jAfMqW1pdb6YApBUBhWkxGLdICr/
1MCP6np7pGF4+2yHKCfnG5mmm+SJ3dy1kIPDBeTU5iHcicGDDaCcfpbJRz2ZvYnRFGyjkcKBY1Fo
FGEhQHcv8KCjGoeWKcEoT2PIETSgWZz0H7J5lnamyEjbAZRdpzYF6nAkRocGJrtQ47f4N0alaeX8
Pb8HrAU8hXbKdlD6IkYEy9LvpVcxtvh6tUwpJp/S+lMgezwAHOLRL+bSMQOMlERKg65tRwe5Q4es
fw9AhLO3pTqOA6C6r4IQ+i7iJXiZbL3/xPYgQ0dryr1bTzQtm2Y2WqXF6sfk5p7Skc3il0A08vbq
ACk4XQ272gUe2uzOjHw0FhxgeuNETeN97kNW/edXkBd8RQzJlPQAGLWcVGqAblGvRHPLs3N8T6GL
1Zf+MxmIMHIitzODKliXRlF+Tfrrrl98UgAWQi8t6XCiXyXNiA4aGrnZIO4fuGN56eSuXbeG4zgf
IEhFaPkB9jbgkaCeNIldBmPlaxPrygEerXZ/RI5Z4UKpIiw1Lc5KDPMwsM0etGEAlTb5I7TkVtxd
QNqmlwrdAau3lt2ZjVrd8kT3BfM1wiJqXOpnwhJTiUnWdCXWgsEvKkt2NR4ewe3vdMd6xmi4Ubvu
KGy3yUj8jFuKPSbEsnS5XnPkEfOhbGzHoHSZ6EGT4264DLMkUnosQTiK1rk9N5S52vOrkPzRl1tE
WPVV0DsJL5yV/0RMhZ6jT3tG1YeBrIQm6PPTOmKAtJ9ZtRJ192wwAgjjZAhSTOTcqL6smp0/z3W6
lWrdtNtL4tER8+UtKK3Bz/Gonb93Z5qhRaP8zYo13fQnPJoDWir28KT81GC+24gMuNDSSY6dz2hK
YeNwoK+larjRujyZ6A7QfBeBR/7Cb3PhOhK+3HJTruUXgKkKyF2pPyBzdX+Ipxu8h1pxiLX+lQsM
n1ET3+TyHdIrx3EVbv+aQChrHRZuOdcTAXn4gORLzt4ns+/3XkrZD+67dgm/uHdejct6JsBKc36v
700pj557bLdcZtNOcLZWhrqk2eQOCfe3woIvrrmQj8JA/uRTKV5jaixD12h0vYSwepQUpuT5QdsY
WzBnDUR8yRGOilP4jKJSkyukT5qKrjoQBEhfGU7PjXnX3AKzuc5s3k0ZDqa7/yK46yCFIYiiIsgH
KJWYxeX9zSx7+D3qf8wXOfOsMMLnGbJgxLEBAajB4v4ZsSsHWm1EthbZisP7StypyczoqSeuG+r/
BickPSFqRCdWzvPlOhyKbu5zN+bjWS/nnfbDh1ALkX2t0OHXf26Xu5fSnE+4tJ6SaYGoi2kteoOt
2PlD7a/ZsLSwBUUNy8SxFXkjBoIQ+mgR14L/vMb9xeEiY2Zok6IjVk6gyyEpBXPRAK7UD02v9Bl8
7Y54xExBSfWJeGgmg5K0xOE9hYCejLc6h7e95Me9KLmgnBfmKOt5Tquh+uBVtEqiwU/PH+8aPWtv
+h6r0NOq5Mi8slQaMSXZIA8Zpps2jhT8S8uxG2Z0iU4Mt60w1h1sDtvYKH/bcuXjINbzGEi5WD7I
NHzzzUdcF6DJoPS7ZxqeyqI+vWP3Vj3g+G1O3C9lvUztR4JJsQiJT6RcwsvfQCOR2hijZQ4F7WbD
ICJtOBh85PVa46v+fRlr7TWIalDQl6y6+HAwtN26eCv4bBT8j65APOdhKsDgld8fbUwqRFRrnNEl
KhYe9XY7m8/th0IYuFJlDCCBj7pmA+eDeP8PNWGwHv45VCtp0hPdjJ254nnpZleG0zlyfn9MtgF2
clievfZR333WxFzHH0xdvhZx/K8IlTfoEnauM0BHYlrllQvZLKm2FB1honSlAmQd1eQOg+AbsteG
IbECN5RLj/WaY4EeE1Pg3UOSptXYXfPjLoty6gy4MXygxOvIIyhtUO7AtJTntT48iY/gJvRvCNeD
vobBkQaWRK18lRI07PLSiF10r5l1eM7rAyQSYh4+ncpkLdSMjtQjks3wXLJ56nwdJugdnK9TzywL
c3dJCs9K3JWAP3OJiC2M4XBZHRRzOoKUdYWQEsaBc1Rp/7TLOD9SZNvOkqol9lQKtERiW4aQ8y+e
bzkJD9n5LdDoqreYxycZ/q4DZ9L3gVXqgLLL+xDH2CqtshUkTai0rHO8jDQzcwQM1QDebPZB88Ms
l8Nr3MT3NaQEosgrGncLQawXuyOmHcJtRvEIM9TP6FKFAEnaSd9+/OOPQUdzKywwqlB8cvTMH0Mw
TsxTTr07zIkfyknayLYNNLlg+2QHRiF2mHuqzAS4AODGpocimEOe/OhT9XHzkuK++maMhWjFeCXQ
TKM+5ihyczb4EsTXDvtzf5LYzuQNkAoga7lN/9j5kBuGjXtqPeDDZ9zc8OqJzFcxL1kUcrmiVW5G
cBXqYTvpNhpQ1fQwCWFTvhP5PUPFq8Egzj/3+xmhqnRUrhenQL0R4rp0H4FIRfNkFUbgnmUF1wmE
q0YM7p/tRF2jRaVJ9ZcBh8P8thbXwtD6djMACJclv9pTx1HUL/Pu3la5sP7TXFPb/JGWQv7UP/7m
bB6wlkhG01pDVzQY+U/pfmZoQxhc+bhTrnXnOIkEPiWaGrj24R+O0J9JPNk0dvayjNzW2SH02i87
wXuRz2otgCcxw/c9r+tZ0EHd074Vo4oPUG9JfCoMbwr3rU1kJqWcYs9sgmuNX2CajYDLOxG4Hm7/
/kQ44Me0FZj4Y3UcNkBKVM6DZTN8egr30MvlWr8A6Wm7ENrfK2r4fuoi9AKK/t7nBPEsDOfSV0tE
Rhw5r2B8K+BGZzKkGL5khLYhL+8jfQy+d76/25LZyrP1P34wb7TXSET2yhrY6el4w3dHmJW4hLyP
hFTBxRhZnOECo7UN3+CU+cDIaNA1f1V0UIapqVB25S6yBfbo86miQFJUtOWlLpSDIfuVVXnhP8ms
U9Unegi5Acn4Dv359L9zbryGgpmG4hPH7B8NWqFyen83NqUY6aE/5GHpHyQgpKf9Lpbn6qtfWDOi
eKVsIjD+Trzjo4RFl8p5sGgyvvVbFwCeupsqttN/yTFB3AfKZYOG73IlubS6Kaq/Hk8ZHcbcA6E8
Eg748TrZhb8CEo1FtMzVvdL2c7fCIDLvP+HlDS3rZd29Wc1S5b3UCIIvF2AOcL8iKOYx0JPMj6Y+
a4XlZ/sJNpTL10AHA6s35nwbgqPHTHKARcidmn1lxSExuwgdfGSiZBjYRMzfnzRLvGitqVglc7tN
AId4hUOVzgLq9Z1/9E/ptrlFKxKJPDuy+f5FKc1CeBSF2y3Gb2rvGsLOjNouBNS523OupoE=
`protect end_protected
