`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69072)
`protect data_block
6+eMG2D627Vbx8Pu7wCt2HAsXijREaEJN0w5Q+SahYSJB3/J2eRh4QzlII3TVy0MFHRSl/C0dVBC
hKbzut0H/klgy2uiBwQI7D7A8mP9RdL/YXepobZp0mQZlGU8hhqcvU+ZiOKaUYsrs78/qfvbnSTi
Hb74622H7DMPzkiiUnUJAy5FMQFX/qGIzHjCs1Q3NsTqYEm5GWHHzAEaAWfS9MHDRGkwvJdY3PXI
cHO/mqUhWp84riBDhapeFF8aUJeB/9Zj4vq3WS2whLematlXOX4XBbpvjVYAKaj2W1Pyzc375Jks
yubC5IgmHDrNO1g8LjzccEZJFS/QzHp98j0TCUOFeGMbIALxMP3Ei1pPw1jCeFDQSEKLgh92XIcO
X4EJEobi5iHVIt6Sm3RI/PxazOP2SHJJCdPqj9UzzSrgH0FK1fkEgYa+KND1jdvZ7WiDOksZh3D7
wtT2WpZQeh6LPO+ElTtaV0qHbv1vbflScd2L6lJmoPzhAM5a6I/H1zKZhyRrfK/XJosoFhJIvvtY
vE+6atHo9cLgrP5iZJ838B6UOE50bU0vxkof+wbxpSNHdoIXQ0PxDxc2nC5RKaF4yZ+QQa9ZHe4I
Ak3aAmxwIB1lc2Wcpz0HC3Uw1+h0YUtzmeQANjxjjM7C+fKTag/ewBGJZoaAay/WaKBLqDsEH9yo
pdUQgQOAZ4zLjvu656r+1ZdvasrguMxCZxzMwJYHb+EpJn2dyS+ei6EpH4n5L/5O/kZEsey1slVf
kUXPUgbV1CzPqLFvT1ha5yrIESS2TKtyhtFfqSmdlmanBKmcKnssmzDoeWkieMlXHZIQTmFt3bad
S1VMohFHeKmvMop1X2Q0gh7aqvOODbj+KzrJHorcBZrQoa3Z0zH1vOy1HwQXxrVfbOGjvy1CJ25n
axIkgqeEZvArdBW/cxP7igq6YC0E0P7F4hkYFPetok/+PD8uOaCbZubq4/WJNlOZcCUCHrT3pUTx
92jMpRvRs1bHCUuAk5L3FhGYpDdRFIKbFs5SerRmyBbF7bc1MWh3Siph0OTcAtHx9LoMLA8UzBYP
gOdQqu4RNwKC3UUw7OZFy4RuI8L5G8OxtVBWrk+4tJ7ziGCcotRSHZyoOEouh8ZR0WPoqldzySK0
aDlwwgd1VVoeZQjtxG3rLHIkONeWhFrl7PoAE0cwV4jPK1rygnYJs9f7CGa2tp1zIl5Tuz0a6i/D
mWDmzc6UY/8RzlTCPLVHGUtVxAUd+1VdCVKFNHrVaC3uaubAoovv4m9PxmjehE+QsVkq3C6i0fJn
y+Kv/Y+sNrp5x1IUPsS7baGcytoI9ZPT+8z2GRJA5lzFFePN3UlIJFwD8qQvoBBnjZXpNTAihc5G
0NrZ5O3vIrGOyBQPkXjYPX0Gdi9hq+1RztOJKIyXh6V1ve8CWiyMu+R2IH/AsDrFzCH09HqxUdyC
HqET46AcE/caKJJqcYfJNYGFAzpv+HqaUQUDvYihEDkpl66i33XAy8ShGpB+IBuUah55kSGISUzd
aPDGBBTvIIgKZcAMjNcsuGi7R9pYlKrTfu448v/NosESoAtCn4oT08KMOZ8A+w2WjWznYVtboYTa
LhUiBSDsmuQVWNvB7RW3wgu0pOSyNWMnA5qfLpOJe3hO7L/I68MaU4Dz96whsAiglLJf6RslVbSg
R83pZn9v/StqnPpnh0aeEr9JieZ41TNr2mtognY6Er0szt50URlnNis5N5O4Ahx93aKu9tXA13hf
i0+Tzk2mUtdBLbg8lKYzjEcKtA4tGEyO71zxPfMKjc8Td7SVow/QtLwU3vv+bSh+FD6rq628F0Eg
Xy9jRCsVVRWozkj3I1bn66Qmd9PzQt3ZKbbLocC7FAcmXczFSbHfNQ9SZ73wL6spCFjsT1wO5JKo
ajy1IHx6O71R+L7/bgHO4p/5RRu+DufeTLaGE/sJFvkZ7ejVuRvlVRqRX5juMoFqDcKbkKHVDOP+
gr62PB2PL/eVJzs95xbp7YwLVUJcJG21YOsDjbf6zsGQAWA1gG1n15kz1izOHO1yIz5lz5I/Wye2
olLort+Z3oORMM7vsF7HtNfhQwflY577ORW5qEWrbPWl5wZdpPyXiz47ZeOs3OgadybjqZWFVcSm
77UUDgWAaQ2YaV+9pIkOs8v7U8R2vA50gNW2xLOLMjZJgvmpaNliQmqtbLsVPcE614V4pfatQfLV
exherXlWI3Qodb/C8xBO92rB/QAPIyLTOCbzFKVaDihP8Z5qBUu7s5Y6MHwOQMGNRQ4/AynCnNsw
vVbt7M6p4tdyX1XdV/dZksbT8MKhABgwlVZtcvVdOzLvDieFl8xdegT1Kruck4FV2nOjMAplGPZM
jmzffzdI6mrT/Br3C5JErbOxeKBtrxv7eIGGXxFacH0CqBNyZgCJwEAXcMElsZWHeHDOfHb6gSJ/
HKGpxRc79vi6RZ+kVOeI0ruBfFek5Hvzg5X8ueRKtq8Yc83qzZd0jPF+ilGWkmPOpK0Z7T4FXm5R
xDvVe8MK8UTduhr7DXSZ1yY/8HJZvS7KhVaEQK0NDRQdYlz8UVSBkQStSGLEdEOW4vu+tfhiEnrX
GzvhK/HS8BvC8D44x6HuIVEyY8kuZdSFd0CSZjLUDRtmqsyUryvbYE4poY7OsFGwi/zCiPLWTYgo
x4hJIsbR/SBGEm8haG05H3k8Nz+0mP0f/nrXtaQB0yxkqv7vI9KsjeZ2yKdi2aUGhzgN09BTmmf2
BzFn3IjmZNqBvEmCtXYAILJckFkGqlxqfSBCx1fxoAD0fXZpJqQzlHGgHr7p5983BOq31+wyxLIp
GWggg+bIkdxfMIEqP7r6z/gu/pweRYT4ArMVD900xW/jk+23TAt0AdlwhAQmTrOYRX8fJsp8gkZU
Mz+bugyqw7HD4HyoyKyHHWPt4wzLY+Svr8Zk3mOy/KnX/U0CG9zmxCLrZDcAwFYfrEVIASFGfV5d
5OoCFP+ARVqZg4OTXlay439zcvRIWvOuX0Y9RaIavnRDaY9x+QmUJrK1Nh595u7nc18qIqVerPde
/5ZSDzl8zbxuDHcc97J0GuiP7GXQB/xFIzA0e/1yFeIzbX1kSNWrJNjI1WB9BPUqCwNY8i93C467
31mUOQ0SkVb6/1i3Z3r9DvMtgI3qFcOzpKkkdjBp+FA6+ypCDN6kz9YHc6i94kwuuUwnkxlVt+5A
d9iL/M3vLrXS8kqH4cyPjbTGGiDMgUQ3GnRQ6J3Y+Hh1+KWHALtOqWOeF8W21g9sBAkPU/oVgqfn
58QuO2KlUVvHMGgY6bF+NWJbxyfLwvRxFV7lzAbKsr/buZrALNbUHZvddQDFROfeSxZRykfQE+Bf
QFlEyF6fqD8uf722v+w3nB8VPrjVehhL+1WqX2cBto/BaEUXQdFsp1FSnwW9SArKxXKPrzr47+Pc
hEXC2V0PQW671/piFs8isvBlzW+wGpKVIAiaQKggE85W4hgTkOk9iu9Ln6nC2eQYYKMRopnP1I1i
tqARAAKWHZvrIYIBC7UYJOUpim0WTqApussk2mWN6NpF6pxVLRmLzfTFcmdUUpRNmEphLslbuLA7
MMkBgGv3jTDNWuVLfH7JOFzaiupyEufCfhnGcde8daEN0k9D1tYZH6ZJXQUXObgz/G9mCQVTELsE
+q9Yk440SwXyoMoUwSzDRulMRBf5zwiVrS0gSDlbgSHKud/F8X+GG3PVxInrraoCi2v73a+u1ksy
ZluZzqVtXA25EaxJMs5PcLvSlV61JkrIekJmr9HnI7ERkw43f6RxnF9iiqXZCAfVhQIWISkK5za6
24Fzduu+/oPklWQ9LZwfw53/4eR/Veol6YR6dsGbmjChTb5Yjc6F76cs1Mcr1QlHh98PsM0k9IOc
iq5G/5vwMhZjvoEAGVgPw1RcQcK+DoQm9keubJGzU7Kkpzw9/7N1srFryLno3+VdDYQEPqKfla8C
dCoyUzZvdqGHOOcuu4nCa0oaaT6QQpgAEg0aZPV3baYNGjXJdw3+2FKP6gJv7FmPEEtsQ6cfCwww
0IsmU/IvtIQpvx0GPYPBLbNR9KMkmWbKa3vNS8zSWmnQgO1bMU+tuNbYduGZq1/W0ormVLOJ3izN
GiYxjvAfGzP6HMZt7ZAgfq9J+MjzT4vSuM7j7lW3KT4HcC44KUb/RFO7V0JoGfI7RZCUFILcqRcy
+Qf4J8zHY0VSmOEm0AONgfhuaop8ujklEY6AdTSjKIFdtgXiDTWeHlELLkrwoAU52SoPPJ1C1e09
QPjNZAS3JxrdhIfWMgyOuZRS/P6Cj8pQAjrHLRHHixUjk664Hzn/N80jXan0LmC1aRFMLmqFAZM8
y91X3V/J4cEJIxCgKmNt231bLMSZoRK4ZzQ9b4Wv7jKW2wcaKFyEGHWiN92XD8zcTK06dgc1uP9r
/4wu4pad7bIQOp24GbFfFRMNa4VytGPWsKoEQcyGIiWPLDBQE/yYovFl97u2/R6vUXvjP4j/CGTj
LvR8Rl38rtzbsKHste7w+SD7YhQ4ueuSLwNjSqYyUrOkkD41JMTljPAkAzwvSh+CCsZlm7nutF2j
PE+fhMKfOLSX50yFjMm/J5Iyt5wauqTmgiLUxA2k8cej5G+xMZrila5yzKAwgufySPZ1SW49SSZF
J7KE7+i9HqCR6azTCuWkAcICekvUgy+Pu95Y/uD+6iyZVbZezU9jIeWa89utLOJvDBTzw+4e4oc/
9FzASp/o4gNgKv0J9TFW+jkjG6HuVXmyoqL3TZ5Bar9kMPnU0smX+TbxCBvV5yDAME83qz5cEYFW
C31pRehz9p4tamt/rNTcneR9MDDRPPWFFjHN4pQAnQ1hJxqaJ/SStLqhxbimGTitIV35lJhZGnfJ
Bp2GERsNqNMn/EYJ3bnGDXHfOASJ4kDZxEPDzsCxKf6FzIC+E8NGU2DAYPzh+f+eRPdF6qZxqrlh
pU/8PpTNw/30BfJGP6mn0htgfhgp3lKOZDSlludRKfCQIgZiFGjmW452PN5sjsd3R//YqAicJCEU
Htrb2c1+GnYP4R9Y9uN20xvFF1mfs720tJZmPWMzl+/2cmw8OjtmMnrF98c8QuobSAU3zouj83TF
hWCZw2XsWnfsKD9OfghqS/Bk4yaiGu98984ZicmpDuVk5kraRQN+clbyqe+qUfQ7IXotVCpKUm44
KCh5gAkcgmNKtCZo4EWyMw3WqkzOaC9p0pIZ/nlUGYgycn8cCfPtvyjwBj3iV9urwNMVVF1I8iiH
RIm7GaGJ50rRmT4hGq/gjQe9QKZynR9R4070Q0nhCtVPRotnwEP9bLDyR+YS9DpCoim5lCSEAzoV
/Gpv6Oqr2LBR0IemYHN358eH7KQb+H/QHOyjOhBT7k0YfYiiUOGgTx620Ta7kYOC9ck0gcXJz5L7
eqeU8Gjd6KdxlKzMoU9vvQAjlrcX1kXep5pLR0LeEUf8xOCACMDcPrFDld0EDeA9D+OzNgAiD7zD
l74UHVNRQg8CAM+QX31GBaKaorPRlseb55xzZVrGZ3Agl8hmdLV0YvZJTxQHTCZmAOETNm8hva7d
eADiJRC87PBJ6zSURsUhi+GtG50FPIOnLvyYs3LUtmH05O+Cco0Xw87dPm1MGUJ7dXmgLjG6JL+v
LE3hnQBrttDdD3I4pLOFWhKEZaVp09HWtFyYuiFQ08Q9msi4pSo6PXRhcp96lVHBdNr2iVxLQbSM
r0aXHib4SCnGGw/W/VLytxnqMGQ+n6voD09FmYNqErFFWMWhSfUXEpuQJTBggHGP3Tn+GbSmXPhf
pQtD703GX3Sso3dzMddT+XrjxdSpyZThZSUnSycnHhLxWo2ZpJdRXx7hpWSfg/fyewOzOCyC3aWv
RwbA2Pukr85NDlPb9h9UuoXqch39gITFikkVhD+OrsbVswrxMQLTNcMD0pXFVY3wv9l0yjTEO+6X
2pu2ZZgCOeUe/803HFblya53LrmonqOBFYQlE+nF8wU+zFexbmBUJxPGl7E2Cq50PNC0ybDNSMS0
RtwQyecZQkczLOaiJEjkiC4YW4595+RjrTPaXg+QqzLyPIi0ySii9mbXJq3yvZYQ+8lCLUb9MItE
7dxKQiYq/rKf8eUzLTGp2fpJkV4+vodAifQKFqI+B7bCPnyCPtGe6ARw3gAKL7jgDZMh46kEjY3p
9RfReU0zTNEJCVbArhBbWsNzwFOw2+CyRMg46zYP9cECTcQ/MlbefROhQzOHYUZhbZz+T9hpb6ep
Y0pfBqABIu+nBeswItmoIg8cbQA5/lK1ak00LcH3FlUkDx4bY2Z2RnkQvVryJnO2vPmyhIprB9Qj
DgPqX8v5XXe8EO24n4ggkz5Y/8kwsV0V46pt8tIuy7eHwT5n3hQzIM2O9nhwIrHpdJPUOEBPkkim
joN2h5d3mJVN426X+PGlsZcQKZO9HcMkRae14eB/TQsogJntHy2hziyHLzKtPfOsJUBatlRBRTFO
mQ52yOYfVE9Xz7BEH7zWS1eGECCsWJ6bT0ZOuic7aau4O1B9GS9sfTH398pfLeCd+G7Ld50LPJRi
BxngrVv9IPEZ7uZsIEu56KSV5NBZGk97dmHQKd6ZQEZQF/iMdrTCNc455CDSYMoTUHbubwrPuPEo
6AeZuzPtGszp0PhuRUW+9mp+4AAQt6P4kFEC/rpo/Elxbbgpx1vg9HDJ2PZYyc/EAQ1h4kUL9ECA
Y4PsHeGOJBYcZJ2sd26IToUw+B5/b16JIf3tPommI9wU+k8YEGlqqlB/xz1LDMrtKjegGdgJ+5nR
MUn2L8tztcTM5N2/FRPBl+PeIrMFm0f4Z/ViYFg+rxwYSt+JQtxnKBtzLh7HfSFxlY7hhIHIlxe6
7Prs22oxqGdFinpXeGy2fgX1gIWDADWawV6CWR35IT6ePTGMFHJIfSzfB7nu/X4g8yXVXM8Zw6fm
oHXUDsJ17YgFn/JJZLfIhViWlz0/RZGPIS5v0RBlq9UvbiRO9DRER02vCOXEmficNrvs0YhvmZG8
8M1dMEaHNw328Sl8Gict+Rzcv+bt6qPqxD72/ZnanQqmPMugy84IUx/PfY8Vs1bMIiwZl77xFGe3
dUKn1DOIT9nKPlT291n89DM9utvLk3Cm8Nhi7kJcdmgnHyH/uZ7oK+Lhln0ZXH50Fa2cnKGjtNkE
R85ngDtzMX0ZMiNBTiZDxIl9OVuNHVZI+osdi6+VBicm7+E8+Kw33CEJ3eYXdwP6vnS6M6E+SXXf
w9KLS8JtkYxSN/piXpFkOa73HeXX3gYHXlPfhHBqpA7OxkVUeLijcVxTTJQbMrP48RT6XacUKzCf
uUt53Dd4BSpndd+pvxxB9xZOKxbnNOyzaF1Tren+oHGmkaR66ay2Y3eDxHSa0sIYhbnkyURlLJrZ
2phCfwMBwJKJ9Z+224nOpzmrHUp6Um3/9VichnLhq8CF4c4LPt/sH27sDPcS7XgL+JLUJW8E4J7f
8L26NlDB8RZ3Ywk9df8slSJ2yeFQ+ZTmYrB2UvB00OHQWsYDMDMIWmDDH5SsIJ0Mt743WtU7tfYx
xsd7gnkpv2fM/l1hIsUck1Rl1+1oMACVipUuz4pn8h3IQH04TO+rzkdLvYwgBEBAAFBBPQDkFwdD
3G5gjIwsao/bFG8ogjJHUSp88qrTAM83ZCAY66sNv4DwaaV9w+qabmNctI479pdlx3CYX7E02AXg
k69TsEtqOgp6dqVdXChtTMEnnkntKwVUovk00zshunscV7qz1FIZ182OtcSkwBEWAGfMFmSkaQp/
Wp45jfSP+Xyq/N2vggGTpQzb26EVUt4p69qR1ezP1SPwm1wNGZwc5MPJ7qdL3f72FuwfWD9fke5R
KF4ginnJA63ahG0I6AMZKgCW7l0c26g6UE1T3NZPM+IHYt7dVmxN1MGmMuZelm8HHHaqZSah9jN5
mga3f8xhB0t0+ojRqQhfL5c2oYjD8S/n8cSaUbW8c77BWBH1Xb+dXniH/ukzgjP6lgGXXtAA4Stz
IgpYyZI8i8AwGOR2lm6HXcS18op12tPzbN+7+zBFVPHVa7qZoEiLtbQonLz5bhIrvia+2EIGvyEA
Tn87gl1dE/PllCCbjw/8ZpAffhdzUHmTfnwMs9ZaJmFnUy4hIPeUlbGYnPDl2n6aniglC+1k1E/T
xJaiRpzbt7+CsjRMzoJeTt+qYUArnkKHYlULUfqU1TcxfUEPL9OWMf4K9NyQAMYQN7SXnCIEAEse
gKODbMMyw82U60gbjgOPpHgHide2RqvDQT/8Y7HxcsPi0h1d+bRptrJrILvF26nmSdwOySEWdYBC
VopcfqxDBvt+EMfwGp2RGWD6iAxl8DBJPyoVQev1uAk/xycy8pZfxTS1wjGQ1oWnLRHqhGljFJ63
uE+ruY3ZU/4FT3zQJB+3JPWBcYZfAVozlUbhxqP0RMbOvHvGYxx33Sa4Synq0hDmEN9uIECUVG2z
ucjVF/c3R8m17x8LF1tCrCuqBnHsUx2gjZDwEf4d6FlH/h2UkPn1oad1ciBHFtpKOy0WONmU4KJo
u4ty7bA9wLibw4R/6VrnsXS1y+kMQyXoDEUKVmJaoUgg9RxyglGytcvWfRLwDypvv4ebTgAUhxsj
GXp6fY6tkT3cD2hNxlLJccxgL73EIrfItdeCk7FIdWDJAJFLE3DcbD+cChvX0plwxCE6Oj3LF+Is
CeaUqTvQ4d3jkX8fOnemwBYhvpluewc0hnjcxaw0H9/tVawPzM8+Kb4sEyXWGKlKzNLeL69ngeTL
pwEm6qvWT6TQ2wVKnchN76WAw+TwWTYxbHH80qBF2MbCvaVQyVwiWfgGnliv3+mxbYHpeDS6Vaxq
b5N25EC+r8//2Zs/9rz8pdDZnWumLt2pCmHLISfKWZWw3GO7YgfeDW+xb04+owDuwM/JnhDllMUE
QgjMsxFufJORvv/I7eCuOg37XydBRy0Vn/MSz0YF8U5Qqpwic2nrFwDk2BmsWK/HKC+bepOn30e8
fY+X7ee1KmByBc8sk8QitUmIgaGX44mXKwhhc3dRiqpHZCbnsQ6ylsyzg9GUn8MqvbTB6sndKB+x
WsYUC4aR1dc+UsC0hcu6ZiFtY3TWCGFn7OKoMvJdm0Xo+VGFlkL/zbRWn8FJ0c+AZiidD9vq7REA
ldMe2UPqBqijU7zDlWVInRN1nV8HizpIYWvfQxOaTXyshrEBKzcUcVuEpLJixO7MLEu3cz0LAUHb
QwAmsTUVhtr56p/DZ5y8pJ4+fvWucaOh2gERzsNQc/AjxkdPIChZV5ptpRHmAkPdu6eFXDL55w0/
J5zEfdvYw59/ZZGUR9nJ4a3mTvlqSIxW/alAeLKuaMa2nElep9DHLOeOVMoFC9A/yYAFDYx64R9X
O9KdJL26QW+mgC2t0qHokoNn5QdRYZ+i27AWcT7p4eHrUpt9U8YKxNtCMEVW+Md6ZDCPKIuaL3II
PEet6Psm6bSfUjTA6Bl77vbSxD1hg7logns6anz50LEsJ0vZuJTWBwGceXYG/GEIjjZL1Y3NhLJP
hUq/TDoEsyDrb1DoezJJZdESf7fW28ted8pbcNms2JThS4BbXnBA6b+pScObbEEFfS5drNuAt/Rp
2SxhcUQ0G5djsN+oHFAHvY7oxpesz8kxjEWr0uvHsVEzCWv0FBJYsVj6aYnV6RD359xFURJWCdxf
8/qdKJSeG+2ofupZdy7wVEEsNVrk6EHGZVWZl5DllSlLZsPtyWJ3T4ntJCi3NXzKC5TuBnrcw7wy
6MIEYpcgWSdIz6ICcOol99zxZN2rGeku0K2L24GUKfk/7rbhulRofGIHb13Vcv1bWxNtKf0eo9QL
0k6+0JZlibbfd8zIRztnA6uLRH6Q05GcnkUG6pbWXVhWA6aav8u8f9NKWDc35DkHhCyCGAhk/tXT
HHc8ok/vfiEpnR5hH6v5QcdaAKpx4RQLfvCmAbtHE8AIF2jxsba1Eds1OrSWNL6T+SU4C/uFxidz
LY0VJE0lbiPIfNeIc8X1k8EaKb1qc5yTaq4OZIEhSfMEWVc8cZMoRvNYRqq6UIncruiOWHdiTuLk
Y6I5CH+lqmNihiRLhmxDtVJhHh7uqHsy0qh28OTVNzQZP8t+lKeW7UzSp9+Kfag7PR2LtWcnC8RR
Qk+EbAvWhGRRC6WwxeXapqWlrCAEepE9lfQkrnNCok9oxTjsp4pICkzZQdlU457jJb1nmYuD+GLC
ZsbKIm56JjV755lKaWILV3TnweURD3u6YoLAet84BAbCc6WFDVzqTH2gLGUKJUoGf83ckHR8nf8u
A1ApslLygqQShWEUbXrX2KBDxi7pS6hmxQAZ5zSwASyw0YC3HIu6X35VcTIEhLmR2B4ryZUCHt2a
GA4yJmMKaaArPM0x4HR5utVnZAH7fTHvbWN5Qd4i/Z3p5V+zPkkku7NfQZ8zlbUA1OdTlJ5ghuuH
PwAbRCc/Y7U1VdrlepexY1jt0RA1he+TD1uk5q5zPmE69k/sr7e2D+u5bgmcDcwoghebeFbU1df4
23oIOj2OAjtJHVH9JIQOHaEZMdlJon/H/Cca/NUtn23d92Q3MXWe7/9FuOz/HJj4vj8b9HLCFL7i
Bu35CaytWfZxFmSFTF8+aVPiEuRPJSXav8ZDtkPSE9WxmteQiy9YlGgqMHeyafTYagOdGagu6jL5
umxNOq/O5NPTwTPHz9A6jPEfPjl/jV1ItZfR7G0jY/KqCBOlIhd5DKq8ZVPNOBZaBOlh6vJYrSr0
OEQPLxd3jKsmSKUdCeKL0gkwRj3wGQVlzMkC/ZV2YKDOhHIuHazbN3epD9L5wGuRrxVCzCiguIP/
UUS5wyOgouQat3Z1hsHpnM69FACBYRQsqBGY1Qr/Gk6KlT/gEzJwfKK5NIwx5Oanh2sCYbc4OAsR
l+k1EpowVmsseFmhjUijEQD2YtGtfq9fb5oqyCif/kDBu2YARBem7Hd4UIss9HpasdhBB9ZQ43JF
6VMbQz2YP5hZ4Nb9F/qMeh7oOcGFun7QgdtlrxaDf/lJM2RBbPwJE0qfF9dElt3QpwIIEOHpzEA/
je9vt0pZWLxLhvIAV2t0ghaFKSCzDLRMixGr0jJyb16nYpR2JR3TeKZ/iDnDwClnF8j00zxTiI5B
ylNYzxF18TrsGDb9KfrAsMpXP6Zgf0oqKpw9AOqFlpLz+1L8vODcS7IGcu//KcaULlsGGvGYre4t
jJij0l5bEFcJvBDYNsUYh5moseoTNQQYrplJ8YOwmOIENB7f+JRRJXHmk1DLPYYe2jEXnP3Noc36
UYMC1PlPuQFBNm0Pz7+W8OOJppzJMBExATosSk517y1ootjdrjFvHPCAEs8s+Op5397pUgR93xS1
v9y0ewIBd9p3pxRzzIqcXowTJcgGN+1rJwlG1AZwXqbpaKAml33217MaFzBdjy9YK/9q7mLvGR6e
7cAYQ9wIgFp1mn8NyxNf8YGAutY2sz8dCFtZln9gI0dtBGOAtcrNSiPPw6fVnN+BsoJ/5dhfW+vs
6l1GQPK3GYYAJ1aXwyQIn+bfHqQNWbtx+1WCRDdKDvZ10Wg/faD+pnZGEZAb3+OAUZ+wXvfOWBGB
b5a5v1WIu/G7pT/VG7hzaz5y1hOfFWQjC0uu/Eylk+xN95l/Zpz0FzD1+4zCNbY++cSwiFyvhu/v
UDS9W+k/EmhmN15hZtTucUE96VrYwlFuQg6iCWBXNWrjQS5hzt9BpGXSMFcrKF8XXH0Exov4hLbg
sEs4/KRI9rC4q36D+Uru6A3hFyrOkSa03cMu4MRDaacC75VogDbfs3U887v6QAhE4ESIRsiEBIwH
do0HAP8YROd7ywyKpNvE4Ibt7eXr3bCIkK0JvZ1tdSWpbGbMCOLihE8n6zEZylX369zoVXJYCpie
X7IgSuQmYbZm2pgKFpUFXCJkKpJckTMoEZntxADH3huvD8vMidIfdpn9lMl6Zm5fl2/CzhTKXEtl
l5UrPuimLeCPPrwHT7E+WkJTwW0wf600rMYbjjNoXu9PXujOOXaelo2fCnZaNw/1ihD4N7EF5KrQ
UZPIJFjKTW95zSlZARsW2YHnbNmvkFBahBCNydjrnlmRPRd8KD6140ccn0kVsyJNU//hSAfu0VmQ
nkY2+ywpb9rWspv6uaiYqetykbCnqj32g3qnQlHn3CUjoG+LjPZe1Xh+lJk1DVJpoTHtg8Lf8JxA
i9hwZjzin18Ofj4ntgQxk+Z8ohaK9GZj3LwzM9n02iGp7aHLeqIlmnYZJYzGhwWfydd2SAXBrQ8F
dIyYUR991UX8gcggXoLbURniHKQOA3/MZr6OyyUJMhS7a10t0scv77vdXoGgxvAafE0SnuDW32Wb
y9b3pSlvcsSIJqV2K//OeKVaa8M7ljCvxY2HA+0Az7ICaF7ntIHpwgkYZmjl5bEA3acgVJM/p+q4
q7xLGJPvsWL0/veb81KeCxWMNeXtXitZZQQbsBCDtjSorWJgmQLzZTDRi6WL8oh5jNFsX3wm797S
45McAhmTy73XrQ+Crl6sDSHGK0oaY8LVny23z4xkBhlReuHF1JCuUqQqOL0YidFgO+TecbNq2uy3
ILSMQJbo3GIYJtRzY38R0/ClGPY6KHd6SQ7EkGtw0FGy0cCQoDoO9kYtRKWSLgDDrx+IibYqq5K0
tDQTb2T6IU8YrLuUYd3TUIWR+QyYGIfgdGzVjptalHO+4AxQ/5yw7ELZrF1ZlTYbshCSyYnx/YVi
+MCyPq6JbUVS4TVe60rv3ycxzATp9RtCg6umlizEI7saII+1keKhh0WIOXC3BvcytxT1aXf5eofR
0okpCGmLnnyVM6ZOj4ZVehKK/eI7TymXt900J8+vP06ZPrD5M9qhZoM586btNkwAroVH5mUTaAKK
nJ6+AkA+pMH6pYAb80kXJB8BpCOXyYJcCp6Ov7iT00JpHThANFn3zYSJbPHDHYGdIwfWqvKbrQEH
ow936B1omTLP9cN/F0F7A+eyNmTYyi/nqo2DGX+wraT7zsZWO75GaOvGMPhSIrbZ6pxbGoXDfPfu
3wwcmz3nQxrJu18neNfDf9Ri3sy3a1ff7/FxY8AaR5aWE8oXgSyrnYgCfLVYe0WnHnwH6kNq5fg6
bSjAg8lGXBKI7WtX+ntd+YF93WleSmaBLAL8ygeyXPKftI3GKndI/wi+qL87wOBlGSN9srTkiKxF
RnnQvZHvAkY6Rx1qytwRoBCM926EEui3UsKpcJzf5WalMWPgSYG81B5fHN3o9SlJCjtGD6SxfedE
e+L4Q6/qpunYrjWAX8tkzfcI0C9s/25vX6TvzO9IQ4yeHa/CJoALtG04I0T3qhP2mETN3zCnpPpP
QkeRjhxx859oSK8EvWMBtH+4hjNwuge6J1yla7pvbceIb6bGdOL1pgNg0H9avK+FtPfHLCUMvpiC
oIbehV3HpKbV4TLbzlSYDVGTh96ya2IwhH4fDwS8MEghJNmSMkWhPXDE459snOXOizASmcF4fL8i
tZJi/zE8L93nYVFGfrwJ2xs4hqosEJkPqbUvLLslPJW49eL+/asDROZIfRISSjBH/3Nxa2Sl6Wmt
Zo1++ppw5g7x3t8fhGHJdj6uQWWpuI5DyC4DbKfZxSV3V5Z+TSOjhDT1uF7JsT3VvbGUhBPkQ+ER
RW9iEW2lldhDGqoqkOoalQcyIgqQMbTWHRNI50cikeQ23+9d5g776Qr4gr3qeVKvUEh8EWoTGUFY
ljmOuLx+rrhzxOaB5U28bp5oLmv3c/VeR3Svk7jp5lH6r35dKJysxV2lfWnz1BLy8Wor/1zn1b/D
k7DzG+b87ENA53fiYEhfm8COimr2BbFglxURrwdWLojEKqjh2ayn6uw7IPhfsmgIK47o3IZUA9mo
6GjboLy00SXx1R73EZI+sPDaXhzjSkfClCOXJrOPGpovIHpsTB7BQHx7BK9i+HXBIoSMXaawZ1/c
LIY4EwFYlmdFRrxwlh/D05r9oWoK8X66qpeWfbmxQlj/iidsF0PLqBocejk9GqoKCPqTJEBiavs0
lKjdq4OvhxDbzDhT0Q3rRVTyjQa9gMepAVXZun6Kxk8GLhTkW0oNShLoaqeXjw9weCNetEs3MXTq
DxstME2DAopiM+vJRZ2+caJ7Ld+8RJuQEI04Hm9N510kMa1DBzT820ksAx+XbPzEXdDVfJwe3Sy3
AMpnJO/f0QVo2LXlPXf1Yfp1fbkZ4Ewws3JHGhb0+4Ae8OvVOg0nuepI3f2xeyX+iuMzpjqi4kIq
EN9szX4uv9lVHjgMotxbOW5R/87FfqA+QcOcd6gKPZhui0c9yvbG3EMEzsnW+W0QB67MjmuUSIsS
/rjzaev/QjPiDyq78Nya2NHbGCdwOibddILXC/UvBFh9cqEExtRbWzAgv2FEYs3HK7uxny2m6dBQ
K16faHGCqbB2WeY1cHaAdbpSCoBcTodiztYrvl2dFnedso1bG2+onLfqg0ohlpK5hLPCAv3Q9JRK
64E/tm+s88DeReH1NTZFvtsS/IronccAMM5/UPN6hJnapASYuSyZ8h277v0yx8NkFVBP/fRCc0uo
uSOPN4GVIR+FyN6UprGyug9sYdAiyzYMnAU+cjnPFDnHu98Rt/DGrR9f8DTN4Dd6hTK/EivJ72zT
lsNgRXFAIVNYmJH6ZLuFZ4HY6vY2MZFzGQTgeUA/tqZf8xTt/Mi/N6/gttbaDIhi0IZos56KbFKB
5ZVbmztbmbWdwKgw7Xj33spUp89E+xfEjH9W9hOo0ltJuj6r6bsSYSWCKslMwa2+Qgf9q9hAbxig
AM7aMI+NONYsD+CbBm41Q1phHfCBob0zN9+RaWy8GkV5+DnxuiNVVy1lCIvbomED2ghICHU6s3zT
JHg7cHG+PXgD1zsfZ2th0OevV2HO7ln7jw+lmUp5QSzKLfEPx/G5Zlwt6DNFpFAXi0U1lBn1wyXp
ia2dG8CcS8ZUSSBRtgFhFZwJk3ekVHJSu63J+zgSKmyxZZlJG/VeoexSdd+NvEd/gUdZ4lSaQLX0
zIPvR+fYZnF4WwM2PP8JNEUZkeLtz6h0fDPWQAIIPp1qU71bTuOmci8GPHZbqHMAa7gTYGIj3pr6
6W+cZ8prdpZixtHuJbZDgNiUcwSNCxMctqkQNEvRN63lOpZ6EPbomc10v0Wxd+DxaIbE3ryiMz6M
pqAuZrCS/8x8RZkOY3rezMUNijNkPxhDacHtxsyvGc6nTWqqSjyZrycUTMVFxIK/GgytRVYqDI+y
UFMz/AUX3lU4h6fLBfgZr93uojn8y206pNtiLPxlBNqOobGt/P17XX8kM+QfLMTfv3+HnK5sxqVT
pjNHalqA1AgRA/hZfY71RW5Uzp9WPpbjhzcOTkldOOJe/NB1vs3IgF/VOLepI6H5DlmmIx5RuJGM
+2Yhd9A6jhtq5AFMOVTDglMYERVCjKQfX2f5M6I6DPZqFZGg0ct8qGC227QBSI7XfASI6Z8T8x1Q
MukjxF/qeMyev1IbJxOOaYgWjwML/UlspP+s2QyrQ9wz1G9jzo747JsoVKscW//I7Dwc7uGkxj3b
75PDiNeZLyXRofzPzRxYWF+6sVezqU5aLcQuYpNOrQCETkdm+t6ZtzfZgl/yAtXlFH1ZZwtHHtiZ
L5TYAOx62FRW7vOenfXqSzxL9GEI6ODcfeR+JwrcbSD/aCztchJLnlK2Ok74UzIPXNvBknhJChko
ekPNBbRg+wyEkpyaywj+0CREwFYl8Gt1pqnYjvLTacpsd++6OSm/4BMn2AXFlvbD6daLr9wJJSo/
oi5DyJykZCI7poganTxvqgxdA0BiwaJNuqiztX+5myAXeGEEDmfxQY4lbS5ensKqPOT+VIpSk5wv
ckDvcGAdTKAqLEzyfkFpxDLlPPteiwpIoE5cK8ISW1WDzqAo7Mudeyl3+4d9cFGUSZETcdcAmw7+
HIY+YgmGS33V379fTQXxHg/ZGUJZDR2QWGh4BoXg+eI9pZqyH4fvhEGmFrnFE1Ahe/Wx7HAWC9yi
Rtn6QmMVonthgMzUW4Y7I9PETMdZeqpcxDCOqrtdXjh8gmbms5BcnPFhH191uZZ9MMQ4hNRQVr+u
rOtdiPPkRh9BCg+oCHUq8gs+VrcHKXWxykvAJ5DWZXrY9TDM4c+I5dP2QXko9tX3NeyH3Lh3nM9e
fRbbpIH+oJDzdfEs7s9bqeMhen6CljD/KGzQvmVTixe7objkxuQf8v/rzwiPcJS+aqPvklMO1kSO
LsLTM8MarzMHPqk/2cHYNCw4zKZitfE0tDG0d+qGPqXy7SsHUbCnbVFjXcXpm1Ts5zn0vzNc1qGO
yKtMkYTbPPAifMn/FVvNYCSrebi8o539okEOvT/+3f2VIC8SCQ4NnTlvXSwanyKV59W/Pb3EdJIw
NoxVa9j82QPlJuAvmxpO5E3uQTqML9bBknuEaajhPvbCAQD0SL8nmvGi3BPkzI7nlTwOcLEf7lWP
fs9bJg1/sk7ebueo2Y+1ySynN26nZVNa89/4hfRHt5PhxSUpWwA9BEGAuQ9twvonGBNL0YC6JbcP
jRPTaOKCkIeOr8PK+ZdKS4MRp0DXnlbC63icqZS56A1jLq/tN5BwblND74qJcohL7hbf+z+1balj
ZIe05/s5V65PlbCBnQnrjTgq+qig4CHht7XPFWBtEpyjcQGlHMOArfZtjQAJ6ZRz38qvJw673wvM
dJNlTCXOfv4CaM7OUEa5iPP+XZVbsYtalKM+dSayxJ00cVYE4AJJbyOl2B5cgLj+ot87fbIXsyPn
0huxp9Z4DF6IdJe2c4fgfHY9lrIHxp3KVPIzO0byV255KbjTtW1yIwCjI8eIoqPvLkwRRWT5A8qD
ESs8DqWKHLzwHIqsCpi2YeU8P9DfeqjaxEgc1zAVSLuDnau4rNrjawh0XqJzRD4ywRmA6rby29mL
v0EWfRhoirxRSbXgUh7imdSb92hKeuYY7ejlrY/CQWK8Tu9ULZo4kYwqLNpQcKMNOmuZXIl9RfbM
O6gDSI+PwxelKEEGT4LAr29doElELLuTaoSJIwgAEwG2Pdlf06yqiR9PN6JSRSmItdavFEYRNHiK
1b5qZTZ510VhdQwLBeonTlrOMBeCrmbjZZ7sYW95KTJduwLFgp4gPoE07Agm+WSHSUuSK3vIzrR2
5d+/w7Wbpt9I+zBBUDxL/+33Ayj362LA8yzzdkIuKhD03QpGkuyJNM7iYdosu3DexBL2JzhBYByE
+55Se+QBjIZAqkpIzj6GKTt1by72ckWl+P2GFLGSxz8Vmc6FyPTJdP5O4+G8mapOd+pcBPPBz2D/
WmupY2ub7U9bT3R7dm4tqts9fuz4Btsd6SDWlXCNZiewlnB2oML3OEGWAJYr+Ls28pwin+q8Pwvu
dx2bauepJHMRRsw/OuqWYbAB/g1ce4lE/tYA/NvLIuUUgarwAc7N2riYFXGFEsS7Dq9fGD7m4f9d
3mstmPGJiMCo1Fz4hWMck8nq0or9aRpge9IpHm+r/woDcaBVHgHcDm+LLlSrpuHOuaMlLc/2ZgWm
3pUNh1D5453fH2zCDKXmOUib5FZcuR5e3dA6hlNocQ2Cnt8sURjMHeC8OEWfwPlt+LVjgJdhUMrc
xuyoes7cpomRYJzdMNLW1xgb+CbONSAsncdaILZ9kqT2dizm8MXVBEtJwUaw7sF7g8STL945xl6e
X0nCnq/YV7mEqy1WK9UQnwjb0MI3c4QR6Z1CmRG/5XnOt1lr6fpwBkSqcjsBUfvPGOjoRSy86B2+
vNTwsHg11BNSPKkLgOoh8dsuE/LwWHHRxWfuhf+W80LaWy7mQX0CRohOmeZ6TbRbF/fi9YVAfLPs
qEWAU9UDB2c7PFkw5p07a5D+ErLS3KVWW27UakmjIL9tWVZD+s4jG2qNFIOyQcF4rRpaVmZkNQhh
T1FtVz1az28XPPwkoUxblo0tUusRn5pmd4yD1VrAwKvlFoLRz+AVPepY+NvkJoB+x6FOves0Y5F6
1sTVZOfnKH1dniLHExDlnos54Df2ya/9F5rOQKQE3foj+BS0DdDS0x4hZSIZQwODysQ2puGOUjM0
LqxEcykdZYwu/Ym8IMn3E5N5oq5Zmw80b9m4mCpkAR9AKMv5KqeTNgXGQU+hE+NEsfZi2TA4tjzM
7z58+KKh844V91jpfiWk8qj1qhEBIMFXiZilN+JTQjLMO7Wkbq1ib8dfi061tCT7WmruDdsQFUdC
G4t0FmCzXvodxqAWlG1uQIdrGBY0H0IdZ5FSgWs3y/iuyzLeAfzfZ73HJZRiSgj/TqsIU3S3/yhI
fR/zEsZ2jIJnJ00ANotyhsjZuUCXdvnuqNkYIWloDckc/0/IesW9cahipXbBvbQ4mIkA/V7GbIJK
/n4RlbNI/9ve6cHhSi9l3N4TfX2Nd1H/GXFxiYWTcLxHEdE1r5clwa4Zvs7wRhqBcMDQ65uLvcuT
cR6eDugrHifjt+zjT6Kb30BlrNYcNc2jOgKMPZuxynaNx0v4KWQC1aP55vdolx3UKqOVSlRzunuo
uxRTqcuT21exhWnkiTO2Fdkg5Gw43TIT82FHPqLm9g+6XNN5lOxq0NdEVxYeRwPMbq1QOcfLeTm3
6J9LkqRbNdo64fvNh5JQ1bjqGxhLggs7OD8aHdjDbs5YFjizV3yQeIVs5EkVhXqcKAsrGkuNkRym
2rLreQQPmsbkOQkylPH5P3g6WqcDhsahec9MQS5+uZByevI1VPXS8uDJi7MFNUSDQHKtBbsmjAXI
o7Htkd8BiSdC9L0ExK/D1mNnXDaBj3lMkfj711cQcFWVfCEsgyXMHk0u1fjpHUo5Oi5rrGzwee+G
1maUAy3umPNAhVz+zgp6Ry14thQayI/q9Erwoa+jipIcq92yjWjprc70JS6btjt5ghR04bIOxY7x
wcOjI88mT2gDgi0n0cOaFup44jRRIRiWTpLzpFwwzQ6Oh0ACw3gOIUlqT2kpq4pw52Sh1GleEqng
8bwR0eeLogCzp4ilOPQ6/CZ/57bR6kW9vWCe1IJWBwboXC6JmYsV6YVoNkAYaTwPyErM/UFat3JB
cVq9NpDOsZwOpc8ajkr4R8L9PQ0ZaMQDrUB70yKiAFpTCcaecNVKvq1rbhfoFrmZ5Q0NX2f4SWIT
tPgzcRZhffktx92Y3G8UqF697KqJZycANV0M78CH8gRwvACr4mQ0Zua9Agvjf9f83w2rN8yZEDeT
mk1lLz4wOQEsBW3lIftzy311KfGBuP4ZGSp8rnv3+CC53d9ed7xin//FhgMQoFvC8NCtdm/5K2JV
o+Mf1Od0Wtm9Tqx8aHMray6SuLiK2zsudyadv4L8yZu2ZOMbX/9FQEscS96L/IsQ83sCXYTX0yOM
M0Qmic64FIXHO2VJ/TwU6DPHDoJCRfymX6oTyKhQCnV28McadHW0pAJUQ7bSBR8yAHdHzMcqtZFw
B3NVv/ovob36JGKeXQHmIEcANu5gKF44XsftYZ5SRPfGpVpnU6mUOPVxu2hQ59aTsLpC44RDRHpp
4tn0FDpYfRWnMJIWg/UHXyDFKecw4c7Q+opt6ZqNZ8vQhufIkJTZaxVwxFX3DgdHb1ahTp/chfb2
idBZKIpOXWLbyiR4qV4lQqBj9GCFHPtZclA+d/2E53UQkq5RbyUQ5+awyGtghbVJJxR1GpE2JJxk
gZ4sUUObT8AaBCYLXW2Qc0Z0Gs3wGV9ubKKwwoLc/m2hb18J4UQGtmaAGVWCYnZQ9oitQL/T22aG
h25LelelGlBmZ3dcL8rRKZwIgpLBGNkVIqXH33irjMoLl1NBX+h2wUbpt2Y3mxD0VkbS7R67JZKv
eZFfGje0THdB+NIJrZzfO5Ud980g6jrJ42CQvcBIv1VaHykvJJWHvev0swyW9v91SxfSjqvF7Rs3
tilAS3y6UELuYTG0SLuuGCq0AJyMXFkmoT9AzrY+cciNEjNuHJSIlS+DHVY66OyJCTI2RYrRg1nb
6uBWn9oozFQV1UuTPNA96w7U/Mr68V0mM7NV5AiSKx87bXx/sI3nUURlJTOeVPyNPXCqIBm/Tz+g
bzOm4MDJ9+N9gmA1265oqhOZbfnDWz6cJXS2Qt3eZ2LTB2E/9/p6PelHcKZHTJntSbAuHVw7EKdc
ol5/gApHRRmNUCYAnjM7yNzFB3pXV7XZOhVzyPTw1m+AwrEin3ltgoJNEfUgqiXGqBTQmSqPKmKA
wzLZdACTlMcpHxgpOB+5JLaXVEZpf7iXd+bhwqQr7VWRblvVOkuky9AsBsOQjfNUDWpePT8ZnioI
HWVEGfgGYryxiV6e24D7o8PsCr4PAbHVp2c6BmhmRmpG96DqDp3qYFIXTUj6cmnPtgONyEFd8qv/
tdkkbFY2d0KiQZGFLGeoY+3A8DDsEZbzlc5Adf081UNgcbXpeeCkG0nnP0Yu81qFzna8tCup9Fad
5SjcTS4abwIIqLgyoZF1iEhjtB2r1cYq3G9nMC5/baQaGkkcaNJr2TKppbb7k8FDGWjD5zGoUh3n
PKaHPHevU88moxUEF0nbPXVb3YBiQbURXjoyYADeoP4wDt+K2NZDBfUMOdVGHIuUk2yQ6GGOdKAO
CCTDbNhVZMcI+kSykIyp7R+ym1bmWrFA2IMwRQm7vNrFw6C0uT/TGceXHALT/P/nklk6Fmf+m8I8
mbuVq67rZ+/pzdQA5p87yCl/Z6/S9fPyKjPm3anRO8Dvxrx0rQBK1fbVTnVFVg/rBi30UmY92avW
/fcGdH7KjvCKwYxcVLkqjeFsvzfvyx0XSoRfxaO/vLOL407EwHBW2gs8F9eeP3rq30t3HuWrypJf
/mX60wk8hEmrBiRSIqSCg//jNCMlJMx7QHmJbA/GJV1PHJulaPsQLhNLZYUi9O14uyo8nnbbV3CA
MFHmr0E+cgPhWwXJeZlCmHLCacNeFZhBXdSrB3BvXZfYAHCHnQuX4L/dxcEbnXtXQjTDgIUJ5/3J
PRgc3HlKbKL9CrKht7bNE8Z93Tn5ie7lt9uOjSRUcZwS6iBInrWdmx80WpEOE7ogH/9u4hXk/+/s
orOr5529TNDRS7YeS5SU6GaIBTNMapycpyJwdGF0Vi6oylQM0CvXvuxJ0deHFibM83JgnTCJbahT
SOSR7YukNQRSkWIBHGyOAu0IIF+UcCNRNpluXT1mOy5REJoxqUYOc6WPnZe/K3vr8ANSqGR4Bq6c
D0TM6pw9rb+WhDq899xD5ehsZDr623lattk67zoUr4JkdU4YpXRgCe0wbUckhuk7/CJ9Q9MQ0k1O
eIuDdd4wIpnJpK8DYqy2ws9qRCt7341WZEpqNQVvB58Zd6lnBum7GT/aPLuX6W4U3sE/y7nFlG6C
DtaOxR7r/2OL7oediEqaRSHXs+Neco7DszORHGFapzIbNXceZgg86eDNidV9LqxGfLELJ5H850OK
r7DSpXGx7WtaMgnqqIzM19Jtk6jRWiq+IWfnYfEasfK1YDMzBC4QymW5nKviDSogLEn9+i/Z+uq+
ss2h108QEvXdlwLQgTa3fVAs9OEuwxGjrOgeDh2nnCtayr67bU6V8fDSEzNRVJJrYMy+UFVSMemM
wWUnvdjNQKIJ7j8nKRrD7XCBuVtwhndtZwcNssoC3l6nxyDNkRe5I/EWv3Wr7jpxPdhkluWYoBia
Hdeeqggz3IRJy9+I57iXb9smARqLp//xtL3IBba6hesN3/n5apVO+CR4UBm0SI/t28Cl0UbHVbvt
j7KgMq9/Kxq2Sd8RpzCMSy2fq5qGDMnsfu4fslr91GD3U/XvKz/gJoFKMrKEVy2ve3vbotYJLTx6
1wiXvyt2p8fgSU2865Twp/qMzmA44S2jG3JCB42NFSFnYnaFjXO9kLXeTOLgzMtO50SXNGKea1zC
WeDG77Jqawgc1hw3SD7+grYu5uvKWv79F4+qau/OsQ22/z4nR9WGXfsv5aOU7KaOsFi0jtMN7frk
KHaFa/Dgh1RiDwSEBCt2s9XZEXxbpv8sIeXu3PAWMqR/PZ1H9vVXdVcLdr5DA9R+dehssdQwl9dO
5zTTOnjEWfX0eIN0y816PDTAPQmnuHv3CxVXGbxLHvKlwI9irulFnotGVgeTg8ihJPeyayVzRTy1
af9Rijl/AA1rfysJyVo9oJVeTKrYprHze+sgzuVhEBx5VIymPXCtorlWKDuNdw5OWOGigCEJKql2
QX+hmmj8F07btVUq4A0FSoS39Zc0rxy3NuwtaODLqMgJETuOeXlRcdVSBRJy7WW4NYx/CKWJ/Y62
6rbf+mWrJ97iB7hLfTsRWFycjP+T0T3poID0dRKh86E/f+mwEXglRv6BFT+YU7ruC+sQrA3URvrX
QoU+QR2gdBa4aqdNCDAaRbztMYBxmWYnvoIWe3BbLfyI5lfTcP1a0zftc0Wt11bEPdIyg6mUUmgA
oJY0mATK+d4tWd1+wOEeMZh7GWconcJp3iM2S06gpw3yo1TP0wS5eBbIfWxx+6qXpHfyGOITdO0H
4EVzxpZPURMVX2JqUG5wghFTvFEnIVXdSx/msedOF17TCfPch6mRmc/T0Zs9eKgKPeTfJ5oulrbR
siW3by5xP0I531odnNtdfv37fZEcK1PymKg6A4NFLowH0STqNsPCIN5FNmfN+RNkKHjQHipDiGVm
1equlOJO44z99O4CU8U7/QqUZetC4Dl8oEmR/zCp6Yljdr7K5u9ETucuCezwIW/Aqv+uoRrul9qI
Ad2ro5JL/Fups+tIySJ2a/4R9bsaTC05PmaexGIu2Kj2TyRl6fVXlVRdbfsP6Hf1mHLmpqN5otLe
7PlrfIJtxaZt4+rnVhaGFsKcyvP3iUTx+Q899xjmc6yTa1ym0W7/9YSMmre/7rMHRKidXYiYQ/pP
HXUw/IukvsMYAFF2fiScbEHjBb2k2r5ib5T2sdKDnPm9NJZIdgbjri89TfnKByjh/j0URk/rU2Q1
Ak1HuyHK2W+P8MSGN8YojmMG04+vG1p61obBHsHJqeDnQy81S9/ZS5bevLlKCQn7TuuXxI6SwIoQ
bOmJ5TuZe+I3vvd2dkQB3M5DmRELcsTrm+RqqzZEi6zMo5ZqKLv4ZBmSSruFNekAW49yC6qwJIWm
SpFlqMyfWJ9Qf1BF9KzoT5oGyQs2GqrKGuSV6Wz6f5yeyhFABHFfLBZCvT7+j4KSnOpmApMZGSVD
KnSENNyWkrCNsBocBdwSrB2FwhNYH7IJIXVnevdtaf9HnGoh9a/996JOa37Hf+QahcBIvGK9c4G+
c8M6ZapKRybGb/++V4hrqoDICM4a2+EiwfHXfYaQ/4JQG0VA0ph+L80KDNhIwKQ8hvtKsSLPztuL
HOB+sejnOB0Vh1NVqgSlkObAVDcS2PELRrhn24OzPMMnzHF2H+miswtTuarkDel265t1N3NuMST2
fdC8fs/CHFmW0sopVPkmbTTE0gV+wIISxCcdB2snb/VB3YcIkQ7ZavXichSy/7Z/1iDk4p6kAH/i
6mw/ooWzPHu9aJfDqigdd90zkujvxFrdqd+cv0eZZa+7EaG5ZHBXdDBLIDYMxeokhcIcnT65PCJS
WcSfqHjniZtCgC1Uy448pa9mxz84vgg6UfjkKGqMbfq4/2NhHrdG1KNy8Jsp4A+NVP95S8hXxdHg
6l4tT+N7EY7ozn3DOKHzw6DGIhdVvfoU08/VIUeaVi4HD0OVb87JL3KW5HnSiUDhRxcxhDm1PjMt
hECS3y+w5+NekmHjK2UenFYhUBzlhSAhFw5RgqM0j4hsx14+WM6jCHgFwSyrFYq/WK9fKVr40qgD
r6bNkYpvBrcVAF+C3unQK2tOVrdlLxRXICZ724yinOOZcB9NDlLRafWquKcWW/xpsxV5IG6Tudxr
djCo34xnq+hnjnv6VBCTgHqL0hXd1bx02HXg5JVDCmlG1lfwH4Aa4DeiKysrDp+mkaOJzuDhEi0P
l7o4sxbRjTYWBaugqLQ1McUOGipFQmXovi4eVX/jyRTZa9Mosrfpesrha6pdbyIRXXBl2GPAGAxC
WHM1HnEUVe4h+FvN75AlZDaw8aGKjF3GdJbGG3qWvgG4qs9BG9woQpSUsEtYBsmnDzSH9HlsuUo6
aZOOPICGr23FL3f3fv4BomQLGqSbze8GYAUewUG3SugCFiBjNVKNK8/TX7oXqzU6RqPf50T5d7qk
2BNTgAKHd7b/UvdekkM5Wo7z/so6SP7+jdIQ+PZAmuGkUtgujEtTuFcZzdvSO9v/HrEzQn07WY99
oed1Xl6UJnaIt1yI2Aq98vq1Q4OoCNrjIKo6UwObXppLC3bZSTbi31isxjmPIMrF7KysdHit1s+U
dPPSfycNdPRCv52/KZbUw4cyeq0syfIjUDjw3utWEkUsuIHC4AUh1m6mEivxIg4p0rma8JBkCgoV
ZT2XX5HbFyuOO+LRmsPL6JY4BafFvi+4DkO4IA9RTy+1QXveNPynvCl8gH4NKd/td2E4sK2zpLls
pr+X2AmFanH0D8NVSpl4rlV38sFyQBKEFpR5uiSDCUEBop2fSjYjkqBhGNLFOYICUVBtmR0eQ12n
Ju1giBaKd2ZPrf0Cd+q0KwyE/rjBquQ83AHjcV8FHKu8TEjMBpi2NNK9FCUMwqu+4UqUON0nCOVP
aiZ9ZMDUrA2CZ8uCCtRMM2gUgosvEoAtoehX6FFA9dEHvfZb3K1+puhVmADt6O9oIw5q8/5qfRU0
yUe1lCGmHROvPzkIUx7hf2VLnizavOclnPJwDdgO3tS4R1LnT/vh+ASF94rGA2OKEL6INnjwbwmn
LPS4tvbYcEx2Wqxsc1LlNGpeUDrJTQQ7kEwbY0G8CBuL6jjlf2jDLYmeosxxG47D7iAzh1F9OK/5
lK71fuCSo0ID1vWMmxvS6pmGdMkxk8q981wznKjxQJznoo9xlbI+CrciUY09nEsciiBz+Goomo2X
7vrw1ljR8a/p/ld2RGEt6ccNdZvZLTV98w+oLKZ3s9YPP3zKXzKGlEqxChaE1X7q2LWKivLXR7W8
QeM5wjLxE076t84BFRvS45m1zPxPrHLvOsgR3bGMK79RusHvlJASBPspbbm/dmNwwBZj88en86h9
WiUYsYapoyOpVkDMJkpgMWr2Z5dAs6SXZObDJ2zxhSeIEd0cCet12u56tIID1pEeM/IrNo+8YJJG
avKoLlbUkXfoMnkDkXZVkCyLIy2X3KufkoD2YXrj/PXaP/G8uZU20wlJM5TzBKRtoU79sNH5jWn0
ZBrDbwoOgY9KSFeM2maEEtfL+v3aiLwOizEPKHxeHaj1eiHEWzTWdQA77oSHdXdQDEk0jiVMbvn4
5m+4ssEidL2mHaMIlUgdUHI1BPuQuDeufnCK3UOiaJ7x8QvDNK22Xkd5Xz7WRiXYmk2SVO4Xe091
ZdanWXR1+0zemTIBTogq01AC+xtqy9z9F0Tsu0ANNHOsARysJPDIhoPVmS7OWMtUhU4lCwwZvPbF
94McP+YmeuGyf0orRYorgCY3uVGcLAvogaf0WarIr9RdfEU6DsHXEUyPvrGRB0xPLoTYJy0r7Imn
zIRxBLvWObqQAGZjnK/PczMS1pKEG1LO05XcQOtLpIhXa1UclyxOxveGmCYfxblMNcy1ARh1bR4K
J/Zjay7K2P1KVdcSQ0LSupXo80r513P3Sk15jUnKiV7F1DLdR2gBnQmak0zlJ36PBBrM5J+RRvgL
JGUG87s/GFnL/adpX2UW7JaxilAn2tQAu3PiSIjhcqxyP5tuEzkjTUl2RIjHFtV7r73erOFUURh1
7fkQpod8eyHx59DL8AEMKpkPRuklCcLN1lsbHQOlxgK0yxIEQPn990RLmxmedLaB+hrrb45awN2H
VnfnqBeQOU74OXnE6P+2L6E0lhh7oOBMrbITxUV6C2jTv/oigvXqjkfcZZI8/LLqqfUPZBOU7Of0
YWZtbNKFzRGIgxqFU+iEMPg4NUZvkXgLXNntxvSLQuvKT2AunUwf1dBq0y2Htp5neSD+2imL5Czr
5bM5+H3yl5M8ZI9oUeVASVcfQCJzp+4hYAYSnodhhWbRLhGrkV0KRI7s/9S+JFe4I+A1WSruSJS5
RGfP9z+Cg+KzfTf6SaRvQp/IsD6Cz2wcFAc7aWslu7qVR45vy8n/e/HAx9WYB1jxWABFHTbNIAP/
TZZH06OW2u7Br0sQmxrXB4V2UZHLZUSleR+u1D/kM9qwdjkNg/KjLDyV2/Lp5wMfJ2EzZJmELxdy
lDC54vKzIdD74eQkiHzVtzPa219oYIdyfOgVGaNAdWSdjoCn3gLHFb8K1ytBmN/RvZ8bUR6oCs1J
6KbftSKwz9KeX10QU4JEYuohhAWRiwbBwjCsoF9arqH7Qm6Ho11RHtjIDmC+TcpMes/NXsNCTOqK
VhW+BcDOBoTouh0Dzl6a6NebQIirRp6x2kFaoooJUDcBYXNg4szR2+HhfSwI2M343oukOSbaK28T
saNtxXoGpwj4uBbFo82nb1xKqCOyhastLHGFyJtC6b5baxZ5196VdtVl1BgNB+XpJmAh+KsYZyDU
Irq/a6Ncq6ElSWX/2fU5rgNf+Q0aLmL90dF/DBObsxq7pP9HqcY95b3/UgolmVkL2EavnROyvtTR
mjokNzh9IxkZqh23eruD+8069hocyXJMW2/Ygzp7x/qiRQ9dHKUhqP+H6CfNxr2innNVoTL7Id+G
NXuO75U1kjLlNZVJbmPWpuxs1y8WO4ttKNt03q9rqmZMLLc/CEL0A52lJa6uHbqKCjSlVypkOMe4
5A2S8sMIYVt7qQ57gsTsw6hJ2Z6TUD3pioAiNmf5kbNIkXOv+unH+zPNmvvnbMhXdbT8QpyGiqPL
TV2i9edIcQOWL+UHKtbrYTVGDwpBtOf3vr/10bDlwkvCy2PLLURVjSf50wQ0WDbzrWCxCvmF6SIQ
fpHZ4g+4yzOu8F3+356c2VgT5xBO6dE/BKhC2daznuPPTgBGLdA+wq99w94vPIe5I2b46o7SZG8P
aWmWXwtSzP3V21qAshL0yYWIBMFJG4d5lQ+383yU8LJy7MrTAkeLcYGKd9czH4S1aDj5/s5GP66V
5ea+W95L9ApcJyBuctWzODcjBqXVhziSTk5GewlCe+N8O4XnHxW0N0ZxkCltpAlpyj+6TuHo81Ix
H2NhN1K+phsCHTyi01Fkii7q6vy8EjxDCb0FXix1ClNWJu4EtZbquH3Snh6paDXN4rgQCE4AalWh
DhaHepOudPUDQtmyePHR8vUEyZcq9NdY8mJ0JaGT8n4hl3SZ/yAub/0dB0onDawj72wHQBbwhevV
/ETdxr/M//cHuuLHw9muHFxzVRfIs94r4C9b1k/4//YRU9aHhhm68GAdfHO6Q+FoReKUiL0EljQj
vuM0xT7QQVkI+ka7eMsE3n4LMDjGbWaqco15y/j+nc5w0ZtTrsBJMDewTN/ymWDx37BbuHsM6kUU
DPZ/J5943GLt03pnHYATobfDWNgfFvDojMTz+xaFoLdJiLZwNuL+pIkDjBPcIZg/0Pbazn/T8cRC
xfNsiFIxwywV7MY03A1SfRwmF0L276u01L2YqX4yGElYLD4cxUTluOpJ4t7x1/pTvJHelXJsvaX8
pUmNHHtqVlan5ODn0nF3YsJV+HCFmabDkKWyMdD4sAW+g9KMIiMgoeM+ThNaBsa5gxjm3UwO17dU
XgToeFq4+v2pxSzbIAb2G/zsbCp0UoJ3m5EJhr3tWsNn42XvAnE4OxqVxkJnhvAL7J/z9A9Jpj30
BeVHBI4/AF3uHgzoa5tP46XaeA6ZiP5g/q9729NqwQ3K7EER7MUO5rWPhKpzjOr9yguO4Cxf1BbB
qsbF+xTiONfwXcgW4XhH4WEW+vns3A6V0c77KMEe3u5naKWTyuxPh2WWiDMd9bHWXVQgGVcgOpWS
IAg1x4ewz3nh+Ulf32WHuWUSw1G5LTxXtlEo1ZVNRKDE+VmDdBT8dLSce1ulPpKHTb3Sp0SEoaOT
Y0bMD3rLucPyYLp4r7sEgt3rAUT/+hLuH37yddVHVC0LGNlbuooLT1MXxdXTnGE8IWayTgVufNUm
BEVbkHhI12jzq85nZFsJP/M0otksuwn1PhAl8vTXBhCJF0H68hhi0Czj4DrrDSzvaFzfflGzEBCs
lZYqykRcbZMBDXwnbsp9Cml4c8/i2fOWGTuJsS+kSL3lHgzq6gdUH+L3NPxDqpCA+sQMbo7uL62J
+dSseAciXvIGKArXmumRNOthWHVqRVJN37WfQIxCQDAXikM1iZO7qQ6g0A5uOgzIcQGvR1MEzlfI
lVkZXDouOmG2/4ii3s1UCC8yiU2nU/YKamAc+UUjuDpv084qvO4SvTuOktY43unzJjpB/KovzeHp
3WrS+Ip/h1zN43ZA1kmJL46zr3idqz7KGUYl+Rt+ZliMaDkQxBKAPA6Wl9rEI+y0qSh586qKrzEw
pc0Md6C0Ut7gpxi+sZ1BcskgVLns4wJ6voghipELgogrFul8xSv6rAwZ8o5oJJwXaGj8nPvZreXF
+Xfhdt+qT2yr+HnBZmNOsisKfGpF+EIb74HcRKY2iEfqFpUg8BaLn+iIIjp4EL4D9bCHGHbKTiY+
GhosLkgs5luxfSck+jhxEvKicBWtukWGUMQCb4rI0Pk8fm2AO9oQBkUCOvfqA3FELVgU8cyQAIAB
J3AfKx3retOY4Y/dDx0qwYqh5QiHI+lOaO41qLuoC6ikBjqa/QUfcT4EWy0PWbIoWlNDK30QzMTi
i30sDOLa1iofYJnXaZMBZlRf5extl2R1GonWH43nKUuNUeaYx+5BQLjc6KTaLm6hLI7qyPSByOWG
w854Hmi9MdRU8mH9v38wTmu9nFGyn8k+ndloCf7cLj1i0YM4OPsjh3mT665JWJRor2WFTDJSiRz1
68aePTGSzhR+2E+z/nb7Ubwpl4mYOpxRk6BDvmbg9GfsuCIn3qcU0jtV7rUKgDiWDUwUfWp7irP/
mNdMGUEe+M4R86rXcX5NIScaxsoJ8lBiS2ml3znKcZu3EAAtKH361zinb3HWXIN2QnaT+G3doDlU
OBpggF2Hwok7/Fq16A0DfGAY7g0sjSCN49ogEw541vSk3HsmCe4uhBt1UOE+GPKzQK0Fn84JhFSI
Gr0j04tUlBzjyUKYUhd+mmOjjKLBRWZ44zl1ZaNynUQbPYYpM7vGc8pnbQ8QVC2Mh/ewPNI4ev9J
qIYflqHgQ3wsnly3RzLDpDFlae0KGqX35LgBZ/BP/gdp1qS4Ba5tuBNlw/jsn8htVIEfTtv6vgsM
36dUsWsCAa/WHnsyvqMnNrmktX2bv/GYxM5IrRS7eWnWxvK523QF57S/5RKU5yEqn72bWmuB8Wpw
FXoLIcjPcVG1+nhGeLwGrkj3S/XP6l8r6xsT3fhUGFrfIFWVO74G4UANci/NrU5QVLog27tKZ83Y
h0XL3aejitzFCsXaNpGMxwaS8Mq0oQrZrpaBJqv8LXCi2tsbCR0UisASjHFBHqAKI0OsjzJ25Pdj
Dr8Zk05MW20mHsez/Ke05cwBSDLJzOn19lfH1CZGrf/9wu2EaVHHgRf28tFmeavJT4Bh71EihBgI
KKSoaXCqlUwWruBnUlB4bbXVtIvPZkQ48gqTQ3KSEkJAq6Iv1eiDGzCn89eq1XbHN+pOXSNPytg4
5WhmKHIRVpGMfKmUpfQVw+zSw+t4MhcxPIlaXEUb26hbitpV6j9gehzhJFlA2U666k04AB4ENzvS
OtCz8tXxmIb1eDFrtr8xzq3aTOBoD/ahLRs8T0y7E7whPepIDfAss8cixDYmL93cJ57vILRSFajA
aSt9dYFh/2vM4Rd0scgXN+Mu69P9tupAfW9HPbdAAbvnOOaBfS/VajEzHupZhAxQKaqztlxeYulz
jEjcyC8SMrIYfashLPXw79WeB8/Sr1ZkEln4P9tH3luZr59toKu6N4On1IBekBztv/Mm9qeL0fle
Ms9uC5/Fo7VEkkYVCN+RsbIMByrR1iy/+gRsgy6V1dWOtMSS/OpySYtGRKwrj6HUSsU8zHJjCIOM
iOvjttn0cqXj/WpqDEx/04jJzXY+r1Qb5K3JLLqbZrlYciSCy8fkhS0TowC6MjnWn34ghjC8EOiq
sIblbNWzq9Kl5fw/B2/Uyixi9T5IwfI9+wyRVbMjmb7bltA3F28sR7DzORs2PWTtNam97Xbz76Ze
C9PxhpmCzSnlsGDFDwo7PuDEtwlzeQYAgdwjBFqXlTqh5pP2Ok1TlheUaVmpm+L8qa6USI/zyY03
sezBbhilAAtGSv6yKdcLvyKpnbdSR50UwyMRXwf23L7ePGDZonlPsm6piy3RLSe+WF4sJwzFAoMx
yaUCupsHqZ3U5V15aOaW7LlZa86hTcpMKBOnJo2nMmc82/Ev7XoXVWIDbqGV6Y9goqkTAX4YVBCF
wgDqJ6GOxlIvE0yuBUgOk34XVAsHdgbbvfv1tlMKwD4aPHFRiDOXAC8NlbgJx6aevm1U23yAWlGP
DD3d1VgEAXl/ifA6HBXJ9o4yB6MM+zEscxLEb0cHChvnRJ36WVMb3rAldt9Rh3NW+ILRS8rGtQqH
WQvv+yG21MiwCSf3xXiNo3CpyV3jxhyQz1n7Bp7Y0CeT3jrF6Kv/6zdVCS7eog1EJMNlr1mJApkX
afv+Cc45xOOd7PETYfHPXTaJmFBPoUCH2XnYMKqezqZbyVEDyEN4NZ0dApxUaePJ+YMCrXO7t3mE
PqePUVWkQeMUiflmnG2Ge5d6PihWK90BsbZci1MCPn7V+AB59p4WuGUebSma0FDsrziLX61JfDog
sybmww/2+5ljy9HQSZVTLPHxqJI3fKKC8Ly0Fif0evnl7WA1X4rw7RAxvnkLGGuhlTWfnHuIKE8x
8JtnXG8APCIrmJUVgHy+L3gVFa31YNPQEObh5LeO3bTdIyG1IdWD51UKod492ZsA+zMYLNDVHx+b
Xpyt5Hdw61S+tHO0WyRvWVBrRKBLHMqYjr2BBtwYm7PIMpq55poGzzywFF6mIzcV8jDDUYvA9fEb
2KUinyhbNxwi4F9zkNE1HPOuwExGOGsGrhVAVd1cEKXFAy7fEZEfgn+oMMxjOAbW5HkEOKDS868D
ljQ5tqdNXW6n0lTzyHZvCNJJjDv8URI3d/wrK1MNqPGg2PjVakaDeMJOY97ZKi5WQFVCglY7TIZl
r2GlK8ebAxAddN5eSlzf6F/ANZA9RMgqWjNSI36RW2kdUPe2OuXdaikx6+GmYC3QBVgD3cjdMMDZ
gFeq207KxsBIib8ot3GXaOMXqKGmfFPSeClUm9E9tRLttkSnJozJN+ImleHULvMSQeDx85nt4p9D
n1qTYXE+IxYiPdACSqtnpGda7Ad3GMxOSoo46j/Pku+J+nN36HxCP3YCczc1Bqujp7a9gEAc1cVZ
RBls0bvz1XRM7hhQ5JF/ORZHqVLHPnNFrRhVdEYfcYFrgcaGwbY9xJcrRFCwPwRrmu/0ISvYng1Z
kg39svh1/nzRyl/weOsKkJ3XKgrWjjKYYsVAJvGoldD3byT/2J+oOi9v/hUDQJcPC6K4YMjnI0Ax
irTeZJzYUHo0ToXzF1xWyK62Kou9KJyRm/NnC7vQw87/SwWbxRGZyPRxB2CumcqEOi+OurauI9DF
xDwrb/MSaFFN0C4SEk92D7XfLj6VS7axkxswRhrzgRE5yCWh4C3yNxxOc30YJVuJ0VE3s22s1AE9
GpRZlTaDcZXQOIxf8WSJBPhNqSS+ruLzTDSmP9to7KECdsp+m8F7JOwvUkwP+hDhLr/g9dtzJip8
zfo8bY16pt1CRDgBUMZE1EDuZp9eOmP8UfeBeixTbtHE0aHqbIhSCbsHn7mpFtCd/CjlOv0GyBVV
+bUHO9vVcvnUMuexfZgvSOQf0Wo2TQedkX241H2k2DDWWGyAzeXi1qLw9aCxMXutm4cOsTYCvlWt
MPqE6kNAzvAIuoHZZgLeLm/9Zdgrkh1FEr782Z+zhYrljwXQZt2Grj88rTArE1KRNo3rUUJ+Ztap
0fYq3qPHcDQP0lZPH3WJPBjOOAB02oBep2wPVXb4M6zDBtPJGp3YS/xLfJevgTJQIX3bueKIojZB
N8vEGW43a1u3rriG00VUZEuCSNqfz7bQvdwbi7iRiJCzvMsjm9OhDMRD0NrGBA0kb13L7zhElRW6
oLrhTUE0KaKKezhGsXwUxF80BR/37EgB1vl2kl1/QqoehHwtUMrGzz+/d3Qt4/LT1naDIUNZbr66
FOqtTjEQyWxzfJAnAJx+tGUuvLYpXIHOoccuJ3bN178o+zuy6d2sfxPRL3mjwbSHhQHqzl5LtQPX
RTkoHZg4YgwcGcWq0Uhb+JK+2Ldp5FFIqXIX8Fo9TGxu6Jv5WiNhLAwRfw3+OBUGMvjl84Cx7P4B
EHSMx2USuRQn9HtNuy7CFZd/T4lbX5r1L/3w4hRub2lD/0XHovRpB+ytq4CipLrG6w4kq7jBDmjo
8SCsdbIvImiNPVw0+ptLKwcgkBsSNBSXGt3A2+emcV7t1FQMHgMkIS7VFbOx6VAqLQtwQk7OMha6
iFKuqI4Rw04nf87m5/YeixJMW1cW1Ay1XK8mjXC0uBXL+uDROPWXlFhJ3VI2wHP2wY6uICnVu/4s
221fc+vM4W6XNCYRPjdcgpNjiAC+/hIX2sW1nSQ/KKlVG7LNkPSeWF7SuotEU4xE/yt5AKL3p7Ld
Lxcs3FWlxAX4GM+zQ7fhL1J3wTE6ROUIzIulk46OcOVtWsj6Vw7CjGJbT7f6YzHn34HGBl/o3p1w
63UOEof0rfvG/PZFPVi5zZnwwaSfc9iAl7uQQha32IsmahS6fgjDaDdKNZAGQdC/2reyE11h8UlV
T5R5YSaSAEX1XMMg36LwY1XF5NmU0ACPP50q79o/GYzv99rnWq89hzHLGCF9PV3vEgzmcFoHRcps
lHVUig6mW2jE0aA3ALRQeYKDJ6J5ErVP9djO5e/29CKpgIs9KZUavxbWcSUCEUfam2ee3OARcoNN
TXn6zBaL2q8TORWfc1kJWgS/6sIMSkCP64c8JlYi3Au3WMEOi68SNkODreNs9U5ZAtSG0pz5ETdk
gpucOH/XlIgjzltOlp5NLREEBITtFL6qBGiXe6IY8DTmssLFcJp1ZOD3JHGbTBLhWuhHIha4HkRn
hSnpHEMDrH6cvqeH4CWnt9izQe5bCAtrPBetrMiaHgwBg+x2CGzCWZVdI2tZUbjjeuXtlcU5LP4T
GaCBELG7keopK0M8NEE/nU9Ios0zOkEp5bbWe7byCzjvx9xkgX9TrdbX+JvoiTYdkjfehf2bKcEa
CXntB2QXiFTLH9MUsVxD88pbgPGEuA5h1YGoREbyM1M9cidkN73VS8ETxsK64Vi9jytYRN00pWT4
TNU4GxwjFJQ7RonqyDcGNKP2APoxjjN3MW9kgUOh5xYI49vLQx+Yiv99fUXynvjKjOF53Gq+OP7Z
sgO87GnJNUsnKZEU9/H4hKJ79TTAcrTmYfO9O2h5d4DipeS9UfryzUi2/fLNW3ic4Yg85yGNjvK9
nxGpYV/XkTriFepNE239aASRzHlktvpkrA/LfDBhzWCPg1MgMeN9YXsbEhCguKYUPYlHffI16Ln7
rRhi4uS0iHjlY51R9NC+oQHcp5RD/QWkApYy8czzvTxy3HvsTR0vekiFW7XW5kJH06Jr8AK3qdEo
rKjES8FJBYX2pnLCG3whiuLHx8ean9bUNQ4g0efjqAQzZemsA5hm+rR34ClyPoxnEH4JT7g2xZbe
Z9WzPeXF3N7BurU7e0/7VILsxR3Rf0dB7nFoAiXU5OxptyNy1LwfoqPVJ3dI/dONn1XyDqE0UC90
kgyTYIiLML3Gk89S318HPIXz/tiTA1q27hLx26NyGf3Rn16NJtAN1POyToNzEPBO6skKnypWjfSH
79Ak90luSd0si0s3poYAi1AkfdgRcI4bcDDc3tBWc+Uk1tIwcP2qEuzIDJsp7+pkPFW9fY3fZOE+
F7jyECLVo9vCTz4RFaS5s7qFqZaAgBuqtfN9Itz09qf+fkUJLjAIZX7Tc0FGY6VHGcFxT0N9dUGY
2H8WjuT/vJSbNVIPEatJW/EIFAI8qBg+kMlQIRTBILGbNnb7HYoCsEBvzPNawfhU9s9TBrevlM8Y
KbpbqpBuzPcaYFZW0dLBvtbb6/639qKWMyHRGQhpT18Oz8XT8+rHh9ACrbdSjAlTPooNV1EhJA3a
Gg3t1NF8y9X5L+FN7Uy46IAurMfjhwJoNdFtJ1lc3iux7Y58pyi6Ec0/qEaFT0Y5gT0Jzg6tzsjV
2m2NAHliLBEmQ52JiR4oqwgjefBP1ht7b0FPyqakY56bXW3l/kkDAd8mCEh79koEbV/zK4re+YQQ
cZ6WhiDtAA6tCyHftMvYRXQEhrMQmplWY1RNLJp0qkeuvUbDRAtfXDe615L4W8gxrnxdnYEA7vOS
Eh3sM8Bhsp2UoSDWect5JpUzb4C6Fvcd8tMgOz+pFkwVx0vYr6Fh7Fa4uUHghgryYTdd7mSFOgS+
s7XB4JKTsYNpoteBy86s66KgrYH6iXdOGnw8NfckHdO4gWyyB681WgMD5rDGUARYQooCKCrrl8DF
fQtF69frZfeZsjG88uBLMAw2B9ijh/aunQPRpxDBFnn12mCjmhvoZgmuacQkYSq4kp8dsxKZM+S+
Tl55bANwf7xIGbb0Yia8jgFJ6AF7hRS9AbygCHShw+hmIYqP5mLDtcYnCwR+W/nqCzlJB9Sdh1J0
9YrMzc1fohi2c7T3nqv5b6oYfTMR3u3n2bu6+d2SwdhpOF1nAW/qGr20gOGNHA+JRwfj85RgTYtw
Ffm+6qPIPY+I7D5i++Hhtbha3HYEgeGPo4BauPNiS6TyKgqL92/YGD389+bopcDPKGt5IHpdOpjJ
ovJ2JbeZeFR4iWRVhs6NyLTBmfdL1/fkUkYRx8hRviQIHI1p2FBoi48YNTffoq42CTibNLCzIBsN
NKzZBVY5p4b4uaa8hK034JaddXzbSWbl6QRzLKpaL9ckdMHk7MA8B++lpJqNPNT+RLiITvbWUo9B
OCOosKpVl7ZWjdQZc1GK6R55dqzxffrRokGmsZH+6VLd6oivc4gqR7Bf0HlrZOYWEUPvQOrBSlxT
31BH2IWZ8eNfp70QUJNQ77IwlHAZTAfRP8J2uuPe+IoN2jgkl5rDi0aN5KdH3J+YCz5GzCo3CxWi
lJTRrddw/FV6x2EzMIUJT+NqM4my6gx9vn1za4IMwHZpd5ZHTr1gCjXhOizdH2WvuAiKvlZOQI3B
IuSaQrsrrZyMMderZcsLqTUJgvgGaK58CfaSqHvATl/zS5fhoY4nSpwjlq8IRU67LKedEgyaLSuO
5eruVHvLCUoBibH4uaPsxDCYg7Ye7mVHCEcoJkEx7LvC6jmTPM0ofZ8wQGLu1J7xrRCllUdmJl8g
LbfpHZj5QSor1kjVDArWdRFpcsvlJnu+ukOWaqQTa8T/ZJOsq1KsIqbeQIIN1q35Z7LLnXfYmxZF
HMW0B+X3w+yDtwB9PP+rinNecZ9f5ViYTZEmOzZ3St6IvYIYdZeqjNrOIgSmw4WAc2OeAK9WuCjI
xLhMCJKUINkR+XPHhc0vLREe0DcE6iKvqMa11ObBzPziz3isfXh5Q4V2/qqzGoObpYtjGWAJh/3y
q/9AbF/j6gxMjPqz7Fbp6f1X7eL1K30qVm2X/AElI+xV1mhKDwlUkMl7jjJuHnZTBcMvmxRh8O4T
tZgoHJyZ2mKa7AkH4ECSuMQ/0qw2+29uxQpm0jHHgrSoau5SKwoe7oxzfbe0T3pXUJfRpt/Lrhof
l4DRTQFXeU8sybQ3gWzjHfnlG+cyUvDn0fJ7Nbwyg3YaUIO4YANtY0bEOEri+l2AZSRm4R5Iuz14
oQOHj0k3M/GkH4qwhPsiPvEHkagm4Dzdm6S1jqcqpd0KDwhKL4S7C0NlGEserk4RFdxeJmKJgHZM
KA1H5v+5nsqO1BNljpfk/pp0SqEc9eARPXhUpU6zn1h44Wp9qok3RynGd1OAcqDKr5vOJFpkqg3G
r9xCJWw3Rzs2ClPEnHTBVOt+NYGjRjG390hSc+ST6iLTiatm0EDIKRxLd8EMyfCm1qEqhUyHFdBc
/WhKOiIIFYYKmgoJXGEYPK8LgWvG8wJQVK1euVz49/sQze1pMRxnkBNQ+tuTQr34C1bMi4IDFNTs
hJJdRb0Trn4pHBr17IG2A4TBA/TckG+0i+0uIZhRABgjf6WAjlEHdu1fpoeHMgKGpbD3qE7YjQE3
l6D9OHCwR4lroMW5FKpj9D/OBQK9T0PsmIxYDxW3Di4hYc3ZLrAOln4fRrKbDVGtk7HxlDEjqGqW
oSSN2JxhALhl8NNz4YuglJZpOXNQkdXMm3GxEiZksGdiiLUGAGY2PDFqE89Evtgafcrhg3OJv0rh
XDSTcFbdFJ4f1ITD9yYDnvRgal3QYdT0ZX6OoeIf/+re7wp9ouOdB/hx+8H/L5QNG228G+7Y7AiD
6hFf4/dNxnSDP27AxyWcBS4D9hWaxb8N+bleowb3FHztgTl6Z9sK3g11RAQwKbLQIfWUgbPRFIDr
qhx2hMqr2SxEA6ku0m4SvYS6v9bkym7sSh0p0IG62DLIvVP60v5JNndODbfEfTc8WGPci/Sbchv4
BMUJXjxkwmhkO+H//wAjjD6RJ03xz6ybF2ZRHqbPYrRLrOCngy4IoELBdQ1W2qRf2MqU8Tz/RmaN
qFC7h4Np2+D4BsUsjr1VDf6gYSZBYKXJV+YIodiEYeOobP+s7V9LtBhvSS8cC7w7NE37RDUDvBAI
vswSXsySWkvSDAko9bOQ6dMZNL3Ttn8buyC7lCYCAFXdAGzhCgG9T/0WqkXBMDiM3kWSIC0xGtXx
t8JXrOkXbP4HNKT435z6YX2dIK65DmOJ86tAVzVNQ0TbfFESxZKo8c0Uc6tsNT+06dahJwdtvlYI
1uPMyRPkT/i9pNqm7cvjpX1NhdUhu1zRKb/dD61F+bRvK07ejHOkep2WECQbn6zuE5L+2VWwyaht
a0xiWsGIC85YLBm5Vz9mUPB1W7yAFyZtZDR5VmX9/6C/q2nA3XqVv01RlNKSG4NEbMTO0ht6xz2v
YszXMOYUiCHTLdtGo+PC0z8v/L9pupMV5qnUETsWHtQaJIkkUalqbqZHQ0QdnTTLJJRdggu8x6y8
bqhd+pCJoiBKTvDv1LdsmX9estBaKkONC2Qnh21NdyhR4H6vxojgwDqMaRb3aX3qKCsd4LwEI00w
c+PCOnfhCXrf3PND0nIym3/viti6m+HaScOCq0q/XuyRY3jso8nFbKqQ9IYvahv/3MYocnHm7iOU
XjbvJkf1OYub9prz5ZenrvSI9yHv3L1JZbQnZzkXFsa1pE7l/uvxHH1VC3SXY6BI2J1i501cGSzO
SAFjL+4D7pgNRp1Ua6uynFLfd7O856oQ2cbr+X0505giWmpBII8/qA+op7SFXPBW04pYTs6QzVKq
j8BJqulBPb/D9PlDZaTGDb1qsqAA538/Pvi3tlo7faAz54rycUl67JxUG1D/bML3gUmI1EzehIbI
qyfXPJwyO9DQwIbztcpjUib76umvyz1du+9lt1NG+yftHZPhOqLeDk+DtYBJWnSWR+xf6e4a/MId
DqjTQBhXNG4MIdwZOJAoD4ydj2MoTy0cVdrNmqDegScaQauuYOD0kQEdeX6ZCdTazZsknmHnQSCK
sd8Mxryr6qi5YpF/0Rbo5utLjf6UW1rsxHnL69jafP3z8u+e/hwqPZvqEW1MYN28FM3eC/wsC5p1
W2YKMjM98MBinXiKMMfGXwiS1lXMsFiGf3CTD/JCo8wHp80VH/PL7b/awKhHsJRjXyqtZ3ZRT5XV
dMpN8B9CBifA8VPR4Ebkcx1ZJZa/elibrh9RL4XB8aCFitM0PdIqDaS2NUkPUxRbUhzF5XqprTPr
A2ycqYnMz/EbtO5Uoj0CgcH85f6Dwqh4xumJSZ9keuSPUz8Nxq06QU75cQox9DNyVZfwnLX/4J7h
JN8XfQNtpf9v92NUcm4WJd90BE0BqEJJpxHpI6IEifa1DrTXqEh8lwtRUO8UpB6+OlcYE7k6hG65
uRzjmLznrvjQS/Lq31Y9ig+Oq2AJv0dZbfkxzyA848ydzB1LrFZKa8t0knL/92840xsHZS2tm1ix
02NxCU8aKGdLsAPUT9iM3g8poa6rP9gJ2A74T0NLQxJDx4v+bgtEBHNj/2bfwzBSyWO+rW4Agkx8
Ykmt6P8pTrZ/RvDFHKIxiBvfpMmeWOoIea+aK4MAeblNYHVFE2SKAHFUBSq+FnTouuSBN0r3jzk+
s08haZRX94dfpQGmQnRtbwSSAg4iybI0/lU+kJgktScWQv4cQuBAzjmVLzmp2v05FJkILVYesc+/
c2wDm4q38YRJofG3tOU4UeypZo7ocoIF2ygr7ESjAS/eF4ws2rHKacQoHUmcn0l1ZxQpxdR3TsZd
ZnVv756sSRCmyWM95bsPbX5qpdk7JTuimoWN+lC/yNnvetS3yCWgSAanA/COtYoF+WucaPw0YEGO
bYVlN7tzeFInqRljRzMLCtCmOCWnLH/5hXqo020fiWX6L7FudaZC22SKcphTGU39yrzcydaq1rUz
zMwl90KBMgE/bEhThjVYbuBGb4lSZbz36it31REc/zH8eaaOozc6hJuqpDUqeuHmpn/UPzFEQfYh
eLTHX8MI93gQcRiM2hIyopzawoDinq0jQf7IY6joXwoyHpU2apgxuWjTCOqdXBXVJSFPrr5mCvDL
9LIiUf+I9lNoRzEOxtYTaXNvpwD29gReTcxajsfDZnG7Xw1p9HL5Wl5imGzswidyyLK/XOrVbKwY
/JxsHID0iYd2Vej5MEBnxaQoTkl0Mp9DxoMm8ZWiC0wdhLuSNVquHFViM99BfNFb615YtlXwcvL4
+TJTpHS9aCtHZMf3waEhaqjo5fGPMlKvA18TsnVEIg3vwtQB7Hm+hl6U/d0EQoi1Guue5UtFSVQc
JkrzfjfSh7yoI8rmTZAJAZEgeBbex7Ec08AMrRZ2QvHXDv9eYVkWwnooB7/cxjPDxYyTbZvcsZ3D
0vWk6qUGnPBeRSBxmKLOqer5ZnkOawg0hSn7ZkQse//LGhWVKLE5JfwQxa282cJqntI0KgDuFwdE
U9B1PWEC/iAwlIIoNsOl76m29gzXu2dNAi+VDbqX9P+EMHfnirKYjGVqKZ8FyOMNLYXLRf1ifK7Z
W9QRt+JTCvm8nctBaiRhCEvsao4lEcscUXgNLJ9x0TYJVbVXsk/LMiNGSv0M/tNcv1SmQeHs5JbG
lD+KnzsHlVCMT4yWc+j8PI60IN0c9DCjEcCblFGroGt5OpWhy/Q/Pi/3V/r3op6zWTLSAOAE06WE
afhH9pNRHfSTONWafI5l62KjH1PorEJG2EIg43aKtRbnc7Nx5JOgUkYcpS0PWvt0p8PP/T1YnPS/
XAWvdaHzHT/ZVgGMyht4xK37Wk2cqv0HAg+bY/XZLP+g3pZ/HpBixVd/HgjY6ktTAq2OoutgHIQI
DL1cAFW/zuZhSKgbHjTSOHGXBMwd1tSOGQ0oARyUoBuJn9sBwm9xRXGqdPPElxN2BZADnAAl6/IT
KLSljRZD+bCeWOCBZb+kyZdiZM0GdUFgQLXj+lBHrC9b9VGcrYJiuIxILaO6sTxLVIFVbyhq3v4L
/PFELamqs7dFIyNKMWKZ/l3zzuFJNcsTojkxI0rtInZqZF1NEyFVu5+R+JNPkVvsYvxFYWJcvnxo
oe6wvFoJ0VXMnfBq247g5oeJOWMYLvWEbIuIqqpZyV9ygLg+btvMu72f2lGBnYXnFxXFIiE3YAzT
cjH1bQNcVHCk3amCnoAlq7EkT/qP6gW83xnrTPK5jtS/XuxCmjvgPbT1HXJhDvIAVJ1kArZnkgK7
WoO01uw5PXZXPZ1YSojwTL/7RZXXkVugsoOkjkn9ORXPSklFRI9sXKuJzCZ7e2vqqL8xvgFlm7nr
R3nU8ta7b1cln5pHqb81Rz3MEWM58gVMhhlmqkmuRYN4TVRB9jfVmIqXaDSYPNO7O7p0epqSXa5N
vgXVpRb+LzvkX7RWpKZD1PotkC+LdkjjiNiIaBdzKyysWF5zrZkKl6eS3d7hHDhcGoNGUj7D0zhO
8SDQMQ/gegsf7saRv4CE4giKla4NcMZ+sIXhcGKlSoR7FpdM8Z1eH2b0j3g7BOd416KvwEfTKPy5
3vL1e9z+WHN3vHmsZLhF0/e2mHwVeEyhQQWLyhD12ymaMYsijGvyptffuw3qCVA1NQaZ3rjwvmva
2lPHXpeSRa0NYQ3iFau8RV2h8v3R2zMZIWbj01HV1MfOASUieEoHthv0K0/7c/w2vHVRHKMIgOke
1/VePs436wbaYD+0KgtY8x5WoFaJao1oivpD7KFjivw1LlL1HSUZjfBDl6EvnIIJXTklkeEudad/
CJdW9eWwsk9DpC9gtU6g/86d2bwnDltp+aJdtNe0bVoSc4mmc22BnoOsTMp78xQNQFgBosBG9t6J
JcTy3S3O8uwjaXZpx7mbqnqrZQHStD4WKWoymJuYoUH8Fd7gq7GEdgtgihYsJyq5QkKjvXbb86lE
VUgVvNCJJ0IjNwh2gNgz3i8qMBBrh9a3GTzAFNEKpME2Ml9/E5R+zvHV5EsNDro7kIPX7z5nlkwG
fx0RAN957zxYX9Zeg5ZuX7EkmscTPdMckSMsl/flN1fSLPIHkkt7Re7RH2cjFXu+MqcGuO61gXs4
wOBXKAY9hSXuzoVc16oz7xtYzQAdkcirZD3CMSNK+PnbUp+XMlHlSzfiKrQN0BfHqXo/0XiI81XR
Lv+gm7KOfS6igrHE+I9TC/P/EeVC5DazlsnCke1hkrh7Fc8jkMkgxivknqJZ4dQ6ri5dYzMjCdlH
ZlBwzL5qyYgxBVk013tES0bFIm5F4mDMpCe+zEWVOzaOV/cLOgtsku7XJWn0ErLmrN+gv1eqYsTW
+CIpOXepVZVFDpy+i46uT5RUWv7aN/XvWskBdqzq4F6dm9RZ/MdQNW7XrSQjHmmjWcyAzhqh1FPf
6iUvPGj+BecBnkRzBT4ClliczlL1cc8VC+yKxIavSO/G/Oc3NaAt6HIVQQuN/rdO0vkshvfXGAEL
p5cKCTE7xBzmS8Qib2o6eiYVGtKobVd0n5h3iDkbZQ4WgFG7e5AfdEJ0dnXXD79qU87Kx1MVPTVn
6OtFLPBfVzc6yUExX+Hw8XAh2d65KQS226ew0U3vLi3bbBMZujYAlLecGCWbBDvQortQ0WYKGKF/
3OtIVqS4TdGTH3d47N/bv5yG+G/EhHUslUJ+qe7W1MaL6kbNbPXxSs5wD1Dd2P8d1y3iaVl6GbzV
bKAB+bmolu0nZm6Nmt/KHiO6Dem/VFFEGeAgk+LcM55BKREcKm33yd9NqL+gxhkt4myimm5jiAab
3YuabS93JcaJ7RtkPJnRZEgzPh/M/7ELF5TJn0D6mp0v95D3Gy+C/7qvudodgbRjeNYnkd1veMFQ
ESF9DANWYpO2OC2a4VnvZKOZ29o7ejWFdlnmv8B/mNntm30aDw+xWw4KDLn9CvCg9ugtw5MFanjR
tqUKpQICVnVHpsXYsnCw91CTEl5/ju0MKgOasz97oy2FnH46p1jDlGXNInXWm5pkCPHHAZBFqKd/
my7aPC5q8hFEWMLETvtiK6uTLEKSJcelOd/jvFPA71n7fWMI+Wgw7TA2ZSJSlO4F4sOzK5tjXZgA
PyTeBO9+FjkYTHUQ+PFu+SswJlXwCGR/21lBmbTDOXe2ixdFIUkCGoJVD5dDq/GwfEQ54gAcjN6x
i4UwagRffIuNdbwiCkuJ2GXHG+qT8cU2BjF96kjxlWYtKSzZvO3A049wWC3TMBGg3yjlug6/Abe7
NwWcFYLrlzzu7uJhGoYh0U7vqO9Hodgv2Ny+hcSWdcrztovbi0+lvJwCopcyPIQObXAXBnBkGpJM
32FW52HEM9BhC5TqcNNCp3hprPMGQNtanws4hqjAPeUCrMX6d8idWaQTGydZU1frn/xe3NgyhMMt
L/e2F0HyIzahBuSh1nAafsxlNHrCE11R7lFCnIIxGUWa6dGuR+EnEbOQ0vpDCeaQsyc4zOCvjIuN
qw+Ayys5wfpwaoKGbU1wp9ql4uR/2x1ZY4byWDGZ3yaG+PhFkFvp9fHpoWSLE8CmCNaZPpvIGWPE
6yX7+A+UtD8htMQ9sMSXLLzoP5Mkz8eMIhHmM7cdApFFf3YDH3FlzjkoM981ABnHRYiddH5sQNp/
XAuzXBzAs4I58BYM9yFBLxpDwnQu1+3Dh7Yhh/lqRCsjURIwjmqPVUQuXdgNWEfYJcCSBcGjTXp2
mxpXygRwp9VWu6XkHmjUhTBdBI44wfgGgSop20MJmkoq3We+rO97SKVMcjQ0wnNzmQI1YRhue8Wj
QRa25aaSAwG3sCk9pJVUqrPrZUHsTwA+Drp8y6AckIGXUP2PKRy9mATby0eTSwjkm/au1VXujaBn
1DNC0vn2sjwZJohJj+TNxvU6bveQcmSR6qpdGzi2S6jS2/keY05h3Dk4jqxCRRSmLT4ljBnURXbA
UNNiieswManSghom3vgVRbqu1/RCqR2ccX5ajZgSNpaoO+aoGvZb53Lpkb0yOsgAoHeKMVEBKLnk
eQsx9U7DAFPm578vkHv8sz3+nJ99BncIgqVtOP6/m1xKRqs4IE/exqtTCuBYMEm5xB3OqCQSD4wK
Pv0KINJ062A5q9UTgYfqdHyGAHDr+lf5nG+Ngw6jOmB26qLrBRsWUmVtnh6nso733iDTDcgL6Wg/
vNGx1wn0OXBtb66ggD5K/hz6TovyNNT8T+AYjhYHVl/qmkRFAWgFyDy4JyWtzXfwWTvxvp6dd5OI
AP/FyfvOYzSmoTL1k9GIVLvQm2UXGwlQZ6IScBK7BLN+aeIHafQ4A+zwxikb/otxmNCqoZR90l7U
egW5BMpFu9eaSEwQAzwObJEf52MXZ++VeeYeY51ctJREnGcB9jln4HgHfIn+8YvFjQSdMVnkxSfo
T01QvAmVTbDe2iR703WPttkL+NIVe5f50ct0HDC6yUSMC/t/fCVIfYqWwu3lOFM72LoWb7FAJFvc
V+Ecr1ILYlwlRxVkQEqPmTvw6/U8CLirKr/tGcLUXVCauaZuz7lU3+u2eemNA8DFdOghvpXwaWYs
ixjsB1yd5QfJimcJgXPEcSogH2A+jXUyVjMtxuqnDLzfQCm6rAiG9wBm+Q8up4bcPqvFvb/YziLZ
0XdqpLljvU4kHdqGnb3fPs1/LQZigBOadfRNknL9uLaSXrjFTHGoKpq7BewGbVynQ5io/xuBpdtw
fHUeLjGnCZLJBAcVPyFRqM990fSZv4Wvhup/aHjV5SnYHElO0r/3bTOO6hjVWyu9Obh+gcBUU28R
8t6efCDsdRjD9NI/ySx/EqbViF/FSy4Xej2TqDPZSwzNL1BbMsJGJL00X4ruKMvbNQFLVhgMdWAa
+MKqnyL+ZkepY8fC46e4mAbZPQI5gjYPXxz27+Ot+aMJZaGJSF8t7MBknK1ogK32RJsWZfkqwaWJ
v/9iqZo1NE8b+ISrTxckg0PeOlaJOYrvL0ZnUqhhEwJ+8MgFH25E4JnNenSu8M1KjjTqrFyVcESM
Ryap3gGCbalcgYx0IhLeIOuOODWbz6pEdgnKYhLIT72BNNb64d5U/3EjrtFYAlGep/ilHho4tILV
5c6H6QTHz+5utIbDKaG40XFI1//Bis+mhTM1VBwHjz0SPXsFircLbp6+wS3oosshBuS1RFocYY6z
dbqUALYjTOetSQrM90ikrBgsM2Hmvwfpz3P644DrEIvO5EgooT0N0dOQEGWGeJavC3JkpKNRjs1Q
TVQ+WDNkuzQv090SS3ye4HqD2EOjDLMThZ4TgoUkqkjZTyBnW+pdEw7y2dWMe7xpYjHqS8lVUp2z
Ev1sRsHLeFK20xcfmO2maSmBVFG1ingXqRv0m6ORYCo3VSZxWJ6MyAXB5SD/oAup7HloM579RVrH
hazvVE2F/eg++RQy8LMooG1/H5vwPu6VRF2fna/aaeEuUexfy8h5pqzvjqcphCoZJAr+8TnHuZrt
t1Y011tx5wU7ph45siqqTekq7Nl0lb+t2ixT3Xljt2lCQDNMhKd80yXkTkXwE8HWZ/9uhwrYnQD8
zA+zQJ2DGz1IOgehHw+R7aCcMUNEu9aGkTQNbICDg3/vzmSFsbO9k/z8xQROZNRj68K3cv4okxXh
KySTFZoscmuRlaWj99QzaCSTRpkpATKl4BUqmi6EHJVSNPgkK/XI5bI4oFKBolKlI8fekR4QD1JE
zw1a4cX4EBCba6U/YjSgKMVyZ11BUPe8rkM9cb3JGVa3QRaFwEojrDWndfNxAhhtA0Vko/40gAWq
kYR1Mh3Wg6F+iVFHPjUTb9ZhOzFmTAdZ2ucIAf2KXt9RKAsZBTEejAx8QdIJ4nd1IiyK0leGslu8
Vcl3mx7trUPOpPzMIuWIy3nOgykI/HznmS27TVQNsi2tg3WKVa4W7+zDBBa6jW7IkATIHkZR/rR2
ldGcAsXKtv1UFfVLDEM/mvxRU7Py+ul9sxbnPPKaVD0xdIT3Wlly/SO7jgj6MYoUoUKv431wl9aV
ql+19kN2mNaA6Tx7EPEBTz+lg4ruDHW4claSatwnrECBr0sT0LD11f+dW0mkg1E3Xs1OEMvvAvPI
5QWTdp3+J6TGGivUoE30nQ6xp/TDr4Xpb2MVjzsCuFe3xyX4tAfGrBXgPu+gCm8IQ8XS4FWgspcZ
+fC+yJ0b2hydry8nnO3ZWrlweDsjfqGcsbKLuLoruxgf7UqoyyWIMNk01IIjhz+OCRReoNJ2CBCV
H6uLs5s5hLtk8q7crQRCPWnnPyo6RLa5YXswZmlLCIPjTnkC5kYFVv9DU6vWG0Io/8qvPQscCFSv
3MvANinVdEy7eUF0OtfntLTysqTpyBAJL8QuKPg/Jo9ZaeWF0H8yGUjj4BqdNKTQhGXGisxCcqIO
96K2IgQ8jEIRp/R/rcOpIQ96hhbYluorTkV1YzmzJvZMzayKmoLndFd9vicluEIYavqpjJbPke4v
wXwzqICmWL1sVit583ylRq+g89jvEkuDbRr6Y5SMftAD249Q+0l16VVTeNteKfKiHrkk8okWOFAX
3fHhuBs96hC04yK2HUYSnTgCatdLIiC8rSb6m4YW7D1lYcha7OzOEM2t8DtOl8qMr7CM87iTseDE
Dokidm3+A+/A8kUINaW/ASrquWp2v0uH5wznaiBStT1YSIYrXJ+rXUlD2GC0ppgEHUTjCZ2zxd6Q
VAXKGNvAYpAmoBTlG9OO2Cxutn8MfINvVoOxc0kQZ9GYVwCfztHzy0RbwPR6O23os6zQplN5+QtA
RtwQHZnISwKEPjCOcKI5nbXgSmX+db18MjasrnRD0nRdO7uDh4A9g6qUvbJXzpO2X2Re1XAlI81P
1KcmOz27fCfnyHnJcCrJraxYRIkhnroEKa8ljzd6+FWzLJz5MeVmVM7ylgAPecccRPrGZI0TkEAv
DS+N9c9cdj89qFZpem1apfE1b2zJALLrI1yEVXrA5JOSD1EEZxv9CvsmAflNkXJOR4QATBiYPY6n
Ar+/Scy4OBBRq2aDpWTfMXO7D6iuteJbaKm6zRU/30Rg4k32UMgAm8EQ1P0Fnz33eXWNTMoedraa
MoD7XOl6c6X/vlscYVkNsZ34eJBpH8WSeaNYNJZFS9B1WITIi3oPg9811exyeWUhebJk24B+e8HC
ytXGuxIw47A93RR6vGYsXEfuKCcl8DnYU30R7gbazGrwZjyChUKF6JbAt1Y28Tj/mwzpgqr8PdrB
as3+rFZDvriKG2obACeW6VLKbYE0xcKffn9ypqRyZk8NyEeDUPUx6rXhXr8kKg9Rkw3fk9+FnYGL
txKTHI1BN/EoxxfpXMZvsvRH2C/YGdm7KXnvWeHvGYJXirQGkrXD2g6IzACAcaruTaYzYtBow7fx
EKGGaT9i6etNEDcQGRfH4J+miYTAAnasHsoddTHD8awIhbuC8IP9hyCvV8jRMQJdXADRxWC8xK5W
O4EGVKykzTNPqsdr4N+pyMzWAdKIfB8TCVs9fiq6sXJZSFU74419/E13/oBhN1LEPtAM9L0z7GCV
Inyk5Efe+y1Iv6PiQnDZPHu8jBwFu2CWzy+qY7Mc7DXNE6tw4BbK77O9Oa6XNvLotkkpCeldu0tr
I/gRfT5ERaASEI1fAe2OUjLbxWgcrUTu/MHrUNejWpKLtHtjZtn/ekY9EQaTRmOp8xYLJKvm0dMh
HMkD1nzHkNiP4trW26FCyAv+sx3R8ZlAqZEQdqzDHAkGfimHYcyiRoaJGiYzxvni6tnkcjBw1OfP
VXjq4jpAZQZ3zpINGLZEzKNTKRd+J11wD+Yf210qSUQFRrkxPQr5pQMYuHbMUy7P+BrmxWRpA1mJ
FXXbDQRPR0o68LS5CqMkusTNCUD0YpYvTpoY+mWWL+VZecdI4zV9+u7+HhOt+LsZXcRzwUj33G7I
LEdI+6wq5r5var0Nmsymq+juMEGuosmZMf5IF0HnjCBPQCkyu+t7DETMeMoglRfIUkTt2KMpOhjW
ZgFa+pmQQSviKhhX8ewoHCnI9KAQqoxP8/2BnpisACuO9JMSR5kF7KKsL4rXQSmphD4mXq2/36ol
VwPgb6F6ngqQ1r5gEYuS4YOuUx3gD2U3Xwh383plDPp8//gDmMA9MgN0HhM/g1enrFN62LGXzVIR
GUsRoaGeV+y34gfNFKpfv0xDFZ6tJnhS45FtleOMRH+zvbsBkV7jTZwTwOFKDnSJckUKO/LX7tIe
J/REXeRD7nZ2Y7pOAazE++fri2WnVsuZQo5/oFNwqxkaA5AhJTpC95RD4U4AeEUyvIFEcVLgLEOo
Qk8bol4hUqs93dVidntSnGV9BQF5uz37yArLii6afFxR0VmsHoXvfcWVcwv8dkod0IoujyO+O97e
zSFD9xc2tlprKPIB1qXzIfrA8rGV25d/STW5B/RBjBLub8h0HxXCGTlo1MdGNTunsvLp82Fzhh7h
d1MIzWWUIWgVvkbDatUWF2BmHfL2gQFQeVbyYucvC3DHdyjFLzSx4s+dTh/2SpR/9rdvCz1I6eCP
sZ3CqoWjqzqsMflIYpno+vKsLcRbsNmGAJ3zV3yIMOKW7quJZ6Qrpd34gm/GnPAGvFwf6yW1XjXk
VvHp7P5aqkU2h2/mfdL4efpgpmr0RPwpGozJKOl2kvOY0deWqjBbmVlUNRyzMbjVQzggbCy0Thri
0Rzuc6sd7rV9X+giOlYqojYNC8B7u62FBuBwaDiOOvqEFYkRzQMO2A2leuFEojInhefVanyU0zt6
qW/Qr2mAchYGXac3G22w3Ges8TN0YYy/aI6xxuiEe5cH86HxfdsVmu/Vyanrd0i9ELiwL+HmbHww
YkJ65spCSbxfNeyR34NP6/dVEj/+y9jVYYb3dKoP4gJUOq5TgvgUA1ukuByhs5Hsz3eJp1Of3J0b
2Vr3PRSEhPClAkiIs4ewGll1daIaVqQJmy5U0rhR4b7Ab8RF+NPeNbscJx5sNpF8ZJjYywGYfMhP
7H++RvJ+2+a06bTiUVgpX117Jdh8wDoSj/Cjpk0r9ZiUrVCyqJXE9R9UQpko8TNkqaLALpqSXeEN
F0sp63OIhkGXi0a8IX0r0CX5EWNNBtRErQuEmmOZU9fr0CAq6XJckFHcW1S4DmlN5dgwi0A9Uv9U
BuTsJLy6fnVB0JlwUAZiqU5jCURlbhbjfxxc5pQn2N/yiux5GPDIstI3mDw1OSXjYPOn4eZGaGqL
CJosdqK7iPiZcIOXj+M+sQKpsKt02kkBSZLR42LNE7K5NygeWzvgJ6h3+RpFo+j7V78BU9lRKhCk
HzEQ+06XvN2/YCUrgR0NrVa5BYLRLXRZlA8v+jE2yDJV7XRswdtatmxMTqW+0IumW/n7mLUQevp3
OlrIs2l3nDDa6smaDTBrKqUySAC0ThZXrdT5rK5U4rK6QNelCYH1gOcBSbOQLV6u8HgEVetxxkFt
Xf4u2Hkci9kOkz51vAT/fEGoLzTk148fDF/184ADHzG28xs+xXPEZbfTu5l3nOFdO7pX/qaHg3Z3
ZmfCUYN7RCtX78qifsOq8oUkdvUsADhGN7krvvrJ2ao92Kr3hE/eZUrXp+baHcYKjTh0ONg0DpJ3
zwNtzv1BKNrFGRwfAxCIJtQRnAw/lJSSRcT1u3BlU/gFjWM5zBCly5BwP1Hdtrbb3hBFjPDo8J0Y
noyK690/ns+RTo/yncTlGVAGYJzYhdrCxPlpnp3/x69RYGsR8B08C0rgHQg8FoJsghoDJsJWMZwl
l8cHbUp0VReUQaBZDlG1K7/QYVURESdqD/Slnz2RfxsoVnUmFD6PkBj232KKvwgWFbE/mYZ0OrKG
KM7VNWsYWbcQlcWotoDfFuypCkEbw9aDr1yx/pephZclOZjslpnPphK5oR0yprR1rNGwpwRFkd0k
AKX1r0hvnrRzO922gwQN6Z5jo3C8WOqNvcaMCQ3p0i6IwtEjZ/9ygrYxSe3p7XRYB8ZTDr25cCrt
ESSTk8maBWGiPTzIowt3eFH4AtOSUPVdvvfs9Hnw6O9Tolgh3XpmTYl/A6/UrKRZLQT1pvsaummd
/SxfCvHHvSA0iBatJDIUdOkc/PpAJKXkjPPCsWKbZJC5p/k4lIZve4/66pgqbuV16s2QKAaF8MM7
dXvK2cts1grJ9KA5vttws1Wh4bWAQj4q5TyxOCLhfpTORbWcO7GTNHS43LU2s85t0mrOdrOSzGTu
JNx9fRzYXv9tZB7sFLl/eXQCMj0XcqzoLgj082HPlPz0GdD1voyxRY0rnCEhbiiaPoXTWBvEhrcs
PMQULHCWRCPn4WCBITYxRPYmfk9IzwLt1Hqdw8GOxvtEnuBTYMXkbSOjaZA+eIE/saiypbQ+3JSp
d3byg0thvohhNUDKWYanvBagoR/L9x84ob4ayg/r6TZja7RcPVNaZxi+BCl6W+1FK9kK7ZVvB+17
g+IuFrjc0UIaXULsenu38gn+QPZod2lOmuWcBzs7LT0mAyCu6mmefSfpBZwUEkf77mTx0zGQWJ0+
galU03HXefK62Q0/V+cTsojAA0eWbAm00LJCTVvEMPR3deKc5S+wDBQirVnjTHnu629uOvSntkMZ
1nGCTm8TY6ND4QGU9vzePTVLluNjrpe8wvsJkee6OrdABjjDOB9uOvlj1rj+M1oChu9rvLq+qKPS
gwZspARldPFxcgKtvY5FwirX6S1rwroberDDwD36JMnTeJ5qOcKsQJ48F3ml+rEBqRF3SCCRDfUy
dY6eAzS8W+RfWbigyAi0xJUqWcX++KuwP9m8ccOj+cjvs6Ln9pmkBL4zWEJ4X/MzCsu+509m9hcu
Gm1sukMkSnooYGEc0Mxp6k5rZ0NZR0hQcM+U4hszP50ZFOEgx5/7ExVKU3bc/a6a7Hd526z5eWfT
ReeEsp5bg7SSTzVLHXcgLaWEFkiIED3WK56fhUVURjLemH4Q65jDL9vMzLGb9msRKKN7Ww+/o+C4
SgqacfvQADFji8N+IM8nO05+U23BPOXT4DMHcWsyoAcCyQ8Qv6nGzzXXZkYQcpnjxI4sVa/Y8sC1
pwhlNa9UHlqMaEot3u+5kDwabZAVi2s4IEALxulOGjENRDDMmYP1WIHN3W7qD8kw95do7d4p3FKy
WJ46+sXK2JLn7yWLKWG2MeBx3497bD8z/ITnIaZLuyoGKKALHCzHgdhVYd7O5X3cUwccW0q+LXtB
IkQkoJuJMSxmSV66/zQxKz4RdwB/nIXevbAHF4BgvGvX9mCTiS90jGdQ9eewEy1oXXbauc0lLf3J
L68GQSeLH19Dn7xJZAoWuwa5eRMgDZU4TJ7JF4WZJPPRt+940Q3eW2r7ixY/nUMAWNqyokrW1HCk
V8ruJV6PHJCemyb2rPZUB6DAdpK6LBahVSEHUYJFNiKaAOrDKPmxDGGqTZ+JZJc1NOxcJ0Z6GpHO
KsQzzpmoYHlSzuFhxMa04sVs0QRFVwb/f8E3Z7VAHfPetnQvjX6noq6BDNcmZYxHlXV5gVMUwOsP
lrgvWrYKUUyXmvV6KJMixNBnrxLwuETWcF6N6bNRW8umM2fX62z9/a4HST7kjsnAqu7ikDIMlNmR
/mrLo3O1TfQ0oeuYmU4ZtnvxbuhTuy+aC64rkWQekoNLIwCuWU3DoplXNUAwiuEtvsEWDpMW7ftA
6n4gySVOuvQI7j+xMIu0uFixAupwyGS1JdW9e+IahEP1y+Rv6yBqV1e6/KCMuhR6Xret93llf0vd
2rEbt4F/WGAUH9H2ZHYnfK9cR/S9DNRDAVca5U/zAa4xU5O9nrtng0s+97LSlbm/EqvLvwcmAGfb
cs35h9nupL1wQnoZzAYPlOYWqrKjXPUrtj7sD4pBahpTBl6j30RxXpn7oizOsw6GuQm11+Df2BRs
3AvhofwFSc0uWmhULWlsEz8U3ccMmDkN9l0BPPskE9n0tVZ2y7XTti1Q+HrAQQaK4ydi/4N50DJF
6hHo1RR0RmBJP1QxtNwpogIKL3ZjY3/CtKbcgVDvNRRCCFUKpJd5aRw02lLswjvZazxFD7LEFmDD
Gb0MNS8imaGxVaz/ORyQqa8y2bhxIl8xZyMeHZzShoGor0mAKUjdrygAvXV7Y3UmUaCBvXyIMOs9
C63B80fLc5+urkxa/Uz6cPGWoKCgPvzLTug8eVR74B8S+5JyObrXJF8Ayy3zU81p7wVrTLIR53ex
9bTGNJBhAF+1HZsZqnTcM7BCs+9JrbuOBpxAqgmNmplvjr7hbx53I/sb5qhz2KkqgOheMB9Zse1t
qxcnlJLsL3ICYJPGvUAuBvo5xwswsjqoOnIiuCbBxspKymbwe3SCqV6vc28DrixfaT62VbtlGiCT
3B0ysH3g30u6FRS+wtgjBU62VkQkyOTg/XALR1uOhUyMeERow1KnfK5SF2Qe5hRpfvfRqL4ZkD8/
FEavJfpuuf8I5oCgiMmmr9kwyUxtrCswVov3XkR5Lc4XyGKBLJJ5upz/Jy5EnrpWhYvuCjAekwyC
5Lr29lYf5qtvpVw2uqitouMEJ9FgQmA/suPLGCthxGaq+k7jhgfXk1DGvgQfSvRl5rnOEGZSPFp7
Kc+zGHE2nNqkhfwP6X8eBWm7lBmJuNBjUtNRz51mDs01A9duBzRttCn35f36ri4U+/6WnxbKc7HY
DK5c0sSfOuAXvOzDzEZHW47eLXoDVqXOqDsfZKYy7/2yh3ZQCvkhiUg7/IRhkEWfhDRXdEhA6oRy
/KEdWPfo8j5CGQkwaOCo26wXGJaYdEP9S1wxW+MpKRHrt6ToHU3Z4Sz6ejStMWxxF1I+z6b2lMaS
AY0LbELbmH89//xx4bhPaCMvEVI2MWZOSQIUWM9Am4PqNYBhw9GRrDmltve8fwV5tMsUmoW9pkyB
11XGtyFOUS+zamX+kNfSlCb8Pu/ehcTD3eDD2L2L9U74lARX0yaQkY1rVAvfhZUHCocnd+JTOCAv
mF3wHeyY5GX4yySErPT8byL5b5gAUldKll2GOPv96lkFQ+0M59AxX+lXb4oBfkWbNwhxQXLqyGWL
24SFa1z3Niuy0+T1ZBJNehulKAJhdz20ABfu3Ph9jY8Hmh1d+bxTXMVoMhDx2p0kFsYzzIy5zJLV
18mreJj1ilUKcFgVnC7qZSXpWaMLoem+67sdUfVpIM+S/wUj5EQjf+KFOOrfujJWPx+Kmy1eUQai
qtDvFKKL8qFDs5d++U+hOdxc9y+FuX5xj29IKQ6dQWSVzZzwr+YLT8hbmq7cf0pMODa8nSH9DE4K
ZFFM0CM3jIsWvheQAqR+lcP0AUU7i1wtUR+hA11Xc9t4GbBjUw2Sga7n6RdodJOjIvxdUAMWGPPs
ZSsqKX18damyhBo9SmmhjPSjk5w5R0Wl93HugGds/8lGcNXrbMDhxAd/zPri9AY9OdFIheg6qTDX
Z1Qgygj74PnfPcImeBhzd9V1y8e0E3UioKTL+ebHzyofrU3+/aQpbGjy86sbYlHTO3Zxj6Yu2eTi
V1FvwVmStapg0s2+0FXNwJV2nX2LmhP/r/rmZE2sqwXLf3wKA1b/ONjdJqTDvlirUkfrp9aqLywm
Ad+qBu+5SD0sSAGI07dbY/5m19fvPj797k0yjovgboOEF/UbMOAhK3rExb1WBfqCwkowEaFvRs27
T0aPoDvPWURq+u4DL2C7XXWjzwetpY6j0n/aFvB2OhMXl26fi9ZnCj8mU31Jew5GoW64EABejHjM
bXLonadAScS0YqaGhMPNFVlbCXKu5i+Tco4Sn4uzSp5tZNkLTxbE+Nf4jXrs+l2vmlaw0ePnla9d
qVCww9xaN5abqolkDW8g0/ckVHhbaNSq5UmAzRPqW6HeGkB0Xt+IcJ8Zgjsi0QIyC3T4FXjNyAXO
YBTAqBDy2HimPx552VcuG9THCnI8rqrCk4NPJ/Wr68nzmYQrBtzpILgnrFNqNI+X/WCpS1I6ALAo
Nl5sCKBqoCRCfaP9PP1l36/FBw8foSfpNVAD+Nze8lquJ6fo89iaDYDAYwuLbIKHwy6wAXQHndGN
ttzAmcbuIiKhrz4/Y66quEKlcRegslFIFBNaHBPzc4hCjp3GnbCIIcCcRQc4XmBMsacoUsOoVcp5
ANx1s69XwQadG3yZdypAL5mhL+TC3W7t77eh8UqV5a18h8DTCiYJXJg6sQ3ytuGQaFb/OtlFu/AW
QbkvsdO1ZYjhpI/lYau93HX5wt3+KnVHpuIGJis3KLcKehlK+p4hKrvG5Jk9vBJl6F5R6DNSrmay
TlTQj6ROLBvZji1UNhMWF+7eqvki8Uwl8CsgRDg1MdZtQ8xMK9iwCzAm4yckcOlz9Qdju/VZeK4Y
8ScN62Ue7bDVs1l1bQ0aSuSn2AL2xftDdN24sib+LG2WxzYfpVWRqpNjvJNxy4S8sZx5EeQg4NV1
8T4DbcryyY8RvLsLqNWHC8PdC/JOC585H1yhPC6Wz8F8jL3PjUH5Z9vBisC933OiGfaflB/HAsup
XgDHZSTjKv0EngUNMrqKMkx+KXoRrkYOcmExughbraTwS+s9FAsWCUBmrLz810AEtvTJchp8v6tL
wEZGLmCPSdN1QFY951yESfLN6ewN4AvcQU7XDsdSGrxlKSUodNnAHQ99P4LZWpbtqS6vbf64VsmM
SQs0ihYQAcGYopMVPrfN5z+paQ5+kQY6Zi3My+6yj4IY86g+1yTOn3mB1ncWusOJKImroWEqkZL8
PBDG0ju4tQFmTEULxB5LR433XD4sWn2lBuyiuJiZtLCVM5wLFyqXdWagj5nlT6uFNoE6+WbxXts6
u0xbA9+PsmD+a/PLe0ePRm+wWxcmDjlzNw+byyjJapMPp0fYFWtCkEH1kl9PszY8PiQHFwJUcUmZ
IyQznQ5mB3HwuPLG8KSJCO9xZDn689Jo+r+hBVhwMuCJdpR9+qZHCi8jn1l+lQKC7goKvOcApEw3
esRExwB52tN7JKlxGwlwugbYwKGgZGszYgCyit9jBxgXaf/0sK9RMw9lBTgPP8J0+Nwj81OBL89W
DVcHv/knsJf8kFXl/OyRmKcHL83tS7SSvlhsLfMd7FKHv0K3ANxM5PvvBicaqGFknZACteG5dFiP
dYuFLgrym05BOMggKeStm4OZydp+01DHFt9Bg13e43ldUmEa3/UzJTJ61rGd41MfKyWwzuDBGM4l
i89MMp0FloJH4OOFcMyXwbGJXX9v5LFfFLCSmwbaq8Lbr2q+iB63E05XDT39ypOq/vzq5Eejhoww
hh23mLSmT/gjHXt6aN26dc1gFdf5DgQmlyOItQVK4jkxMdyzZjw9cDzkZbDGICfYPB+Qdkz4H2Ei
V3tlDvEHYFvx4lN8kHireRvLhc4bUZr0tbENXTnos/EsPDR/0Q3jPjAxzoYkei2GdhKhL5r9RHob
/QhK7fY+OGRLEDQtB5yHg2Ynf/amE0pUHcEBfck6qeg+CKFGoxM7wPWSDmRR5PGxjffc7p7DQB4z
wASQJt6RN141KAs41wHSZqvvHQJNV79mjaAxs/A+Zh+j2vwu0LyoCFhZIsZ/Y3kJ8YLkT2JMsOTJ
1Dk9gsgmtL+akqOGDp2oVRC6uflUxMpoMMBY0WLEP5W/Mqv5Ceh+cbZ692khfn2zvO6rZwo+0EHb
5FOAJpUiBXM+Z+HQ1O9w3gqhtu/Xn8c8A18fbua4SFVLAtBC5hvybssmSOoeyUSP02Rh2ZGMgPC8
PNSESTFOAM3lCdM/v8JN3w74ryvdTPtWVoWW5JIC4QnwXG9ophK8SH3fRcrDkZlpn4mAToZhFc7f
5YWAIj/nyYZZb/M5qDaUjBGJ3APgfXOSODwjMRxR9WF1Cxev96PX3GLx4a24pkaT+rMR8c19HVfP
bROPcT1V8yVK+1a2VhmJ/m//BoNAUqivHUhBWqXAWlnghbc498N+pCLLi/ya195ndxPxOZxxFzSQ
yXVIgXsJZ9sflsE3zsVXrV0cix/GXBuVxU4w53hjDVu7KAtGEkoBfH/8B7tFlsnvao1t1WWvZyoq
xiyr7vhC0dSEHd0Zc5Ubh/NkCbh6ehxUx7ZAh+OFhLwh3+OmtOXgdVx5N2UXwmcn/b7FV9+916Sv
QVkW2S/qV5pJAF3jzKeQufPkLwfXf4DOHgAlY6hqigpN9jq5sY6JVqwj2HzMqWOA+NAzBpO81Nx/
IBlxDeeRaXkkxyQudBYk6S7EFo25QZ7bR/o6wTVD1tBZvx+0m8587vBq5rduJ++IzKLE9zyu4Wvd
vdJnsMxA1rrwaqTu3DaOAQhWBq2pR6/PPptR1onPAhFp36ANF5+2y81M0CGunq4h02ZjyrALo34U
NKiSLH1HCbgx/4/PL0rsyh9aqcXRaqc1thy7Y85pdb53el0EdzWrwjpi427Z5BuW5NET7w/NDB17
SwjghG8O7U/1gemDnZ/gbqSq+HmM5MIREjQpdXI4xKncTdiVzcW8GKQM5QSDRPJpn12Nb/klCp3N
TIjW+62s//xjUK/JP3+7d0v7KaMAAVZ+IMz4jiNE4bAk2zR9J0o4et2+KiaD/pI5/md3tnNnxfYJ
9ZsH63oCuaTy2UYk+mVQpdI4ys3R3zXpF9HI479AKuEJyaATf/D1HcOzxcqeeSNkdriuOhd42epo
D4WL7pAt7VwSpAagdJmgkSu7hLDwHjguWcp2aB7dX4q0QWmav6jo92OXXTWDSVzUl4Q++KA5IodU
Go2LrXIF9L0cBr/u+GnVy/vwo0s7Cq361Kw8NzmW0bPc/BAYrbUQfgOTmBArS/7vQtlTruXydzu9
Xq6GGEMzSvheSdoxw4DiwlFMxDK0RiCTVOkTlxtrFvC7T9l7jaPI0eg//4CyshyHvRnmTbpR+5OI
D5F8i/Uz4JAfgKuY6rvpVf3ODkoYBeKnbNoRIzNpSlDa5VWidJu+u+JOmfy8zdtwpxSaplg3e50q
DMIGGJxrYptZV6/EFhdmpYTc+Q0hWUExMg8+joaBWrIerKKW0ZWh+ESLOxwq/VEJcJAGEG3S6nxX
zdK9x/TeohJbNzPQEJFWRa/ZcVb7FeDH0fbGnCQqgCoX1fLWeDmJKAX/Rwofzfo4IM5bQ5BEDwpa
YUi/dHz+Wvqb8WxTi+Ljd28PKsWO0NR5eiIlOoNF+ZMwlNap4D1d5a/IszT/Qt4wjOiKgU+Iv/jG
oFZ9vLQ4+ZvfJS8rEZqCH7nUSpNZ0SwbEOi9LFEQ8/dnnDDpUlP5+vnqR/0zyd8Y+g0klStY27hL
GJWslXcnG7wbGEoJ20T+P6ojuXYob9LZlXsOvP2hGI8EaC7SqUnhTgQL6GER5JmN4DNU/krNisMT
vcT1tDezrwhdYcFMRFciv+AQ74Omdhb29wUNTQJZ1odXyHVm3/ya/hIZfiTsHQScZYVnuCApQEQc
OjOSz6qBQBySnL7GjO34XsHbcWkuvGLZ1gCm6+aEzdEA4gQL+AyzQSl1+GukI+0IPGMvtXR3go3R
8XKYDxHz8wKWp6I78Q7c33IKfBx2ybaX6eJwJcyYPZ0hf4cvo+Ro4Jm7cZQA7RHDQfAmyHOsYEjc
ZyAmYkmla5Se4CspYPiJw/hjektdyqyVjZPeftPfipIxgR0jhQDvzQK4VqYbg1w1JtwXLI/ShsKt
/ulCSymu5/3+Z7FQQO9FVi2u8emEJ/mAIm7/CrfS0pDG1gba5Yg9N4h2OiUQXT6JWnCjXxR/odmj
izbtK4WbPYrg8ZRFI9PM2lvrzIGf10wKOTwgV9drQgHaN0+4fpXE+HLRmWdY1LnPXVgYhPx5a78H
tBdi+NtlhOrRdPwut2j6fExtjIFeiEVRx3C1Phm/n3zyTmS/h0PnPq0mEN+DjTbe8IySos4vBMlb
wrTi45E40vchjUggOihtbUGpuoVF8wRBnshVODElBE7Vwq/C/R0eRM1dg/n1rg/YQzBFdsMjgG/S
xPEk+QiVXv17weeCEsvTT57alK5BgjclKrsd/cG3UCKeFQmhQQuhwqx/SVF82PV0nwWIhaLCbwuR
rkhpBFKFZyX0mSeXP6xmgRiOTzM1uZmy8ygyZV1dob9NbO5hwFfjgwfxwwLytIP9YKdmvYlQhsMm
dwzUx8x6Yft/XZaC0MzBRo7pm03jxtMYuxq39ZtJegIuZ7A4sV/GIu2/DK+1vTiQCTIKq8bAJNlO
EAd2J0MbOAEKwn/H0pDH0NIOt6cSlW3jEINoGxO7k7fL/MtQBAFO8Lv0iSP9DNeBjBfgLs4IgfVC
7TtPXZNUnipbVwlkRsN+N5Y1B8ikmnpaRiJ7sylRpMskvCB6EpbFRMCmyxR2cAZt/j8PBmcF3mPx
mm/9s4ftrGs8Lp5CAH+CmUobVHAcjrDUIZJGV7zfOSwlIsu5hXe/clo0pGRVITjVuv8YV0tvAbDd
v/6RgdVum/sZZuqTw8A9I8QAM6v5b/DhhNZlykektHin/MKHMNh/7DubrbUyQqoRjIo8pSBuJKV6
8BmlSrstEpl2NUv2eBoZ2Z3KpQt5BGekr9UscjFvJp+26+muXfFR7dpONpb9AIizQcGYu28EVRph
I+vlWizNK53PH6Ei0PQ82vLQNq2tB/tGnNRRU2ytMVyZtr6jZxC+vw0FClWdW2BLTZ9kw7W1JsUy
+nR1ziieNTW/3tW+mXIxA71G8kXZ7Nb9zBjf5XNfe1XP/cja0/H5eJr0eb7rVpVxMT2XxfdxmCH9
F1pWMd5X6b/aHQleJAK/9Gla7OGFnHshAXFHaxa7zyrNwMGofAnYakjk1+HEFVdww2Cx31kTKzTH
3sQYgn2Q7Vis907uCe405yh5WJDmYFfoT0I1+9nuFqdvve0Iwu2hGWR/B/ULOJTcnT5LR8GeH9BR
4zZpk05FORoSccZ68/bSMu4rvGHZJ/pFcoA3ac0Puu0LI7xBB1aq8KvuSHkkt7N4UhGt5flaQuUw
SxjlpXtftmEq7ly5/La4drteYpYMhr3uWSXhehgOWcUiNqWrhyE5ecFhGhOX3eCTaSIQO6fXGcyX
KWQca8L0frBijjDd3WFh6WEYY55pzuTz3mI+yisqn7s5WuHLcAQ2wn4Jvhfr2ARQ34BYugqoRJvT
9juM/Ifmy+JyHyJC7F7J64XIP+gBvZko3pudGPNmYN++CEB3f+EqLz28pGd7NiSA6vi5PTA+eOy2
IN8cR1dhlbpCmXYtXZtkI+8z9M3zSxDqI7ZTvJeodMrECGnQKbHp84nJGV9zQx1QFmx6FvhgTgtE
Ok3c/UvfxuXVESu3waCh+vxD1m77F63can9keaip1RplEPAjKYRf10zpfUVklUCHY/jjy+RA9GG4
Us2FxiwYUHbTX7CGP/2cfmzzvDzYVOMgu/uNWo6Du5GaB13rUXd0VG7KBTww7lXeFQTHJo0+HPmi
UsPBvTFjA/ErfL0af9UBI4efINIwu+UjI3NKi4H+Mf7mNbizZF56sgV38EVZTUDOp67VdnB2CoyE
fBVhggtUqI9oVwbFSVcaW5wD4lkwH0PMfwtyY9WC6g8VfsuNkQ/NRhzTfSlW94hjnevq1KAv1fDs
b+FQDE43VJSxc+iUOwLG6Vl8y4VKIImlYDv4p6pQxp0wFaftdiIeI+nS5ElgDPt427KE58nyhhpP
W1uk1fgbKsQYiuWS3+dPNJgDi7QsDj1GQT27LahBoOoFK73cMsyyKENpn6tc6QI1opHQhldnEtmX
O0tBCEK4nsqwG+43QUx0pVUSn5rmv4QFUYoYn3xgLVDMNDFLYqI7FgT2TbYx7P22bHRosLOyPwcW
moxpWf8jyzHcUvzGEFsI48pcLgcCYOCA1/+s2CwJS9fvznoSlnwHxJkjOflTt+5DlBQDUKwnbAWH
pHxM761iUUkqifWxKzhy0rZPducY+IaKJDNWtPlDfvWeRxmRUMp2vS2McQ5Pb/oQgvlBoDLfSBxC
fyHlxfb3youe71/PrmX8GPzHl9jfCw5NSlVxog1DdahHCfKIodNZDETWsCnGh8VgB4B+QtAQzFWV
s43yqybs7ka7uTnZ36dUDVRqQl2i6dTxjCVYl355CiFkEMHP98YDmyv0zUcXTrGzxnv/a+J8hFPy
LcIHYKulg10huGzfUkebsy27wD7mkjPUrCk+2s9ViOkQnaNuUpZPMn66g+FBiGq5aa4c4ODSx6xj
SWI0pnVl+ukOBkjC/x4LVpkECVON2tCTPcbxVpABi4lfswkw81NmWyHrFG6KuMIRWcMP5fwO6ufM
l7l2oG0tp5MWOKfF7Y33iagNyEAu1IJAJqviJ47JqLUIhkmQ7W6rOcDrsOSB9hp7EmJTnn4J2vbd
Js8PJy0JZbD8yd5myYLaCt1PY+r1jehbJBVTVk7Ekql+cPw9vFKgdI9JXWiWgPiuZVdQkAhrdJYh
CASxom19P1Hdp6S/GSLexHq88cHa+jjHD05kxerR3+xiCrEIdgkeAJzC/v8hCnE7jVFWez2AFbZr
nXnOxPhU+lT760UejSav/Klqr2p7fkwybv9PGFdnnLc6uY1Km0f8bhspylg/4sBqDIBZFvkENkQf
QQsXBWWptRBxIyB1AzPUQqsjZaWf+UZ4YmUMNXTT+q9Gyi3FyyKl9enY37tSbua0UWcg2VDBg1zb
zgXhUGPrEneBbcwzcbgPvQ58IXp3y9NAciXE/0/GuUMhDF296bqi4AJhA1td/jbjU+6vZgCPyeDx
xDZsXndYr9KLRW67GuYb5ruU13xUP3kA/0brUH/E4qyVcSOKv5rrxlJC8o2slkFdtWaR7IF5LIJs
4kCvFHx1zJPSb8KmwSuwhsVct1gpVs0y8Z3hB5k5xAiowXh6qjDs0Ynnr9I25QA9SyjNXbw637Pr
komRM6A/39VWhn1DCB1ccFxXmnHiqbDmEh+5tiSYdgCwTvjsPr4sf2gdynczA6e232FhGmyvQFsa
6STPZahUX3+sVN2kAP4PHe7pH7MVZqBEaEuZDmMKOOZASiQk+8HTbz5V6WoZPVe1LTyoOn1lAim9
ssDOS6FgDl0+RjCXY6aH1kar/yyI8n6FG977tKDBYWlRZzQp6oGDahOAYydwwVVEvHbsMZ16BwoB
0hbgtabyINr9hC1nssP6skOFrtXfFyuDwJELXSXWrHeNgZU4XGHOT+5+NkDps7b3RGiw4+j60Y6I
s5PRlIororn2WcZjFjg9gpY8ouWI9hRkB+NCVUPNGryePrY+jJVcFISwwkYG4hP98N/1DChGa2l9
nxAoUdRz5cvwuaY+Bb8KxOsXkPG/NaprrlLSKER+wOPEpJY2Q07XbSntO8lRZLdbOEcmHvQGZG2a
fWZrfePbOe45P28UV8KUnti3PNvYwCsKVuu/rannnNWJzqwHhKa1M3UE+aK2eJJcRirTmEON8NCd
rcHOJoUyYnOSO+HHsV0qlP19jZmL38iv8HG/8bTRjudNfh+V1cBSV/gYWH2cNKzFCwinPCsuvr1O
LwcOYcxJJUwIH/Q1RwpHUfh1jXN6uNLiuex1sAJiZxnKeXua1Q8UJlYFdzg0O9Uy0p4Sac+zDzhz
8Py48QimGowlA4tb2bspSahIqUD1yElYYEf6oLNSv4Ce6SKyy2x4D2225IWYc/yvGjzNkv5s6C6q
ZrQH4/pU/HvNUGK4IwtAh2EEIP70U81cypVdFfHTJ2hHyaLN2x4sa/LE1dp+2LmKlM73eq7iR47m
TvawWH721/XD6vqpsBauQJ7KqjOrFDj1s+Zw7Yb1wk1vjwP4aGZkEqrhfTJ9jCw86/sXFxmJZEgl
YThIwKKekhBh/YVbsVVDAHVl7v+Uvl9J9Sd5Avk0eiA8EF6yb+aXeZ9mUGSh19yk/ziQPVqRe4Tt
+2b2zFM/EBgp2TLi5MkW9ZvDK0XV1W8ergC+2yXWBgKdEPWKP6eeW7EnIO6nyaNbaCniODk6h0m+
cT/ra0N5CraI11Mc1oiDwiDJ1KeKJ72JQvtJhB4Vu3xE7Wc4tnpWw3EbZrwXmvcl9pOgX0VrJPZX
/dxQh8p1gDWVRurBKo0n1K5ZN7AouBQyeLkxFXPTsioUqOlruPLl29dXRLKYQN8M6/V8QM50tTXJ
vjsf2ygNpjDVXo3+0rp5GGkIaU907T9HDzoAiHvLt0CjHAj4BKJtRCTuOH3caQ1szEzuhNboLYjG
tXTVI9a8QhcPOru4Et9OTNroJLaQXuZdQeX5inyhqEoKWRkSRI5q2Wm1p3RSoPTaKSPENeYNKjCU
giR9UABs1iN+0WJCB0fevvt3I9G2pBGpzeP5o1QoxoYETFDUIVDrpe7nOJySLxdR33t5ZHGeQJUZ
9miI4xT/osNmHoTBTKPTtCNGSFm5Nizpcm/J15Udbo/KIL2NIQc8wlY+ubzP6D4HGxZHdl1CsbUO
5e+6r0qACy7yQo8wUcLFmRdMXNi2zxsd3VkrdfHuG5+DUBt6HJsbKDWwNGIMfi8hMHGWCA44WOV3
s913tsHVAC1Tdop0qK4t2ILvF7/1eKSxS4DR01KqptMqsufemY6FXY9qaeQ7ue9XWQCFyPplGTpg
bRWKxB9eVIRFZSBtg9ynoZcrZEtcPz8M/pp5doxrPLReKhceoDPQc0KsW3sbSXlb4hsWDUu+WoSp
K49Li0rLnjVWN/L2MYDgZqIlznORgwktwrOomgsz7lfhSTbuWuQ3142da92ifciotzHW7BrSytbD
S5XYc9Sk5fk1bPRit+vPpmcGMD3lIHnBPkUOcVBtdp8l+2Ak6CQhIqFV5+prnyqDA1iEJlDuXK1z
wR5p170w0ODt84TerYQ2Z03bAAj/aaJf8OfHin75nAnLpVrI17A77baVZbzRj7AOtgtyRUSQHFk+
TBeFXxRXrwyXsCbSHiJBlsipngkjgqSbKMaKleuhS9fB8cW0tAC7xqaYS5VrupXxiCxyr39F/NUQ
W6nZ6jI+miYhzuvWhFiumuu99SlmI15OPOowTLZxGIWAGbGVbfreLUnAErbFA6zsuOxuW6JKvC5e
t706cmEIdfjSZ6FC5JaFmyJn7FeKXAdkR+qY1TuIQWVGMSAqpftnqE1g1MyI0D+9JNq8yjoPKXmm
PjYWPh+zd/Mf0UUCmEnwd2FMb8ckWj6KNJrD3V56E9/yiOSXGn6eAKqbUEDUXXHm0eA3ORn667Sy
saatk6ZH37iqI+lUBV+FZvFrt05Z07IQAotph2cMpPe0F96duVEHfEbrAWtBUwnFxB0QL1W1aoc8
NWqWvwX/JGtrWwUSKoXTrrLOufNuPGf7YfDzKSUNZf2UxO9pvvrb/m6wAdpLunnkbiqAztiyxh2Y
QuAzg6j/YHsia7evRWgarmFAZXHT27aKVl6EvHxEznDK0jXykUfrm1j3hbB5Rs6/E/UZawhL0vyM
31pQMkGop8Acm03if84AMNBbUYzBO6tox81hTFB02Lak7WVtSA+YIKB3LK3IfTzRdkYzFEarNq0F
1tAGAa7wlhznq1eOXsO1ZBB+zvXgxgpRHtYL2rFWbHvCcnIRCdffqvCwX4nVSqZalMXAdRULaUu6
qm6X8qOfsHDoaVGrTd/oHLidV7wl3TheNBAWc8/J++Mj+EsYcaF9r9BIauOvY2ylNsco/+IYnVtI
uloXCjo0XwvaLWLb8+C0xA79hKfhZNQ5EykAJ1Inidq370JkEhgmUwHrV8tzPUge5VlvkAgZ/sgJ
D8fPzuQ2bEMJ9SK210ioD11f4UKl3QnwBMKKu5m8tQcdc5B19QqLjQTPaYKQPhRMlf5cqzqw1OuB
aCGJvNPuqSuRt+ss0YLEscARmapyiw77/d3KjzNkbJDNVddJPDm5wh+0fLY10xkBNhDkOZokCoBf
Og3SJnb81jdCtC+QtbsmVLcg8sF6sK+N9vI4M5RwdsLPRtjaXQ1qC8xGF8D41VcCXO2MYPCC81UK
cVjqzTvBOqKmVP9KDqtG2wxl1t7ovaUC/dxETnaGcEzHK1YlJtdbuUvZAaHZBKvKlqNIfMqg+YUP
xuytjJ73D1rxs/0WZnErMvzCQqi/FDq0MZiYI6GrJZqr2jPJAFcBFdEJtLhzIYbQ73YLuoql5y1i
/ogUh3D2YuThTJIFEzOMjIMV1m0t0j9v8nk6jDMEYjeii1IVPWFqFGtqf/qOViiB2MEONa5fvo5C
NKos8DwDjZsHYbfvsy9p+IiAejyStnM2eWI04pDBqPHfo2ZkaP4/QUiihwS5APwJi85EjpEWJsto
X32s9GXws+/9qXliw2g+kcNdKOI3mDS9TlzpeIqDD7FpbtibPW46XJ6YoV8LckHtU5YNchfFcWZq
NhOghKzOAJEpCv8m3SYivAlsPqPFMnTE7dD0xzl1FChRVr2cGVVwYNYS09qtzPA9WnGsMJm89hZ3
nQJPmeulA3uzY8pv4X5983GOka6AXzPTFF1ZpqlhTGRrSy4CqviKWYy6v5dKqbPYg4u6BaxqpFwX
8W2w76Yi9FuRgZ0cf8+ZQKTn2EL/0/uXVRY42fR5N6RQf1NDBBivgL28oB83TtXHzEpOGN+u71DQ
yapFi6eB+W35bn4D76sSqBiuHiOZL/2Sffc+421P8YF2V/d0x7HIIT7lDgN9M1wsYA73ATrJHcej
o1qFg61Zx/Ub8RCMXQ7YZkQd+qZvtnxoe4CcXvYjXUw6umbsDNNhoMf6e6HiZheQb8vusW3vwVYQ
h+EeyeQlWnoa7MytAYTyZR9C7qN7VzDoBAw10fgmJCo31g7Yd9/BBoRPJCHObr0EbIRIHbF6aSGq
eiNlo0Ogc4cUJrQ7l3EUeBujojB0Ng8h9GpymWixCbX4QsXZW80IBT1XcG4FYXcTb0I1SqgUcAbD
ynNftoXjqq+d/apzDoryN1GcORpkbzfCywt03NZnjCt2KxomnTlmH+3KHUACoGi5/Rd8wChF02b4
nkLj6x/5cFYH5qzSZcbnsSZZdBiqKYsniFAnRGEU/ADdl3lqwRKtkGkZxenFVukMbeC6w7a/12H5
xt/tvSyql5LRjxlc3zER7F2vmF1sKto44u16P8Gig3Tj5fQUAeUsklGPMa18sCNv8PqUA6jigzWQ
NY4XPWeXk32EZADcu105gu139r9EmbFEJfBLqguyD8hp7iGTwhIhDw6fd75/rBYtP8iQefujaaIX
mjUCZ1xwzl2ehb0Cy+ETAe1kksj4x+IAwI1TKjAAEa15feYPzd/1Ouvjg29UrNMUnji02QlPPvKo
OUl5hG75vQVvxwfOyHaOIiQFEsLhUrmH7yHDVWHM7nJDlEI9zQ/kkE2/r6vm/kYV6LLE7CaOo1FC
gbw9NE8O46jI/8fBIzXOnNspFCGZtfgvWWQoyGuJ3eh4Dq0+8HnPOEBoyIeIEiGRh8BjQE9OlvLH
4aqr9OKCHZKzrIV9TcEE6quQqvRj1M4fJEqpeEI30GizfWMJRVF0ZdoSbs3JGtmNYKyMInwOPeIl
gkvKNq2emwzQwo1m+fx95zwyvS0ONLW4B49MeJc+hqxWG1Puu9/31/Djqc7jj/ksjW52v+aXFIuL
uFOxXfrVH7I7hL0YbZw3MTQJ1LALK5V4EUni0YdGVtuDjXA2EGQxsM2TlnTb2qKUquDhRnmqG+xm
8fig5wLevIvSJ3OPv2ICa6rorhc/Yoa7rQWOaj9FSpjBwZL23mtfhbTFxOqx/T/C8fYyK1M4FlXs
v6qw+ZQX7nGRkX6RilMllrpbvWDVjNmlXRRFFirp1rqJp+1/bvUlXG7SJAU3YtBMSGSJe4lIJJjF
4vuMMANc9qb6IRlvKNN1LRl8v23VBuqkmC3mBQyUvF4rs3Fbi46VHUSAI/eX7yF6nnruBBaEoED0
C6jMJSze2UeR8LX6guk5QupwnN7DXo0rGyNbLbPECD7FYSpt2FhQ7S7noe7ZE6n1poPMOAloCyhJ
4FW+Y5XASEYzd3lIsNYq2D5m2e77rq6+adotDnZXzkY/g3cVhSPWggJHMK4bSJRU/UwhQsPwYH+V
+sKfXfAYMQT3J/gyBItY+lxl80euHAng2cq8FwAfOX39bZ+iSnliwTUq5bNzM4uiir4xG5zmVOM4
e4IhgXe61BBtrpShStYk9ZEQBBODJOqRpgMCTHwnXlSXmWraWZGtrvgAVd0Bc7w7KZAzcdRvdXlm
RAMhxuLi/Xw4sysde9d7EszISsAIO3u8YLwaWKBoCuxKSpp/Vl7ZRB4AO3VHtDV2gKUsnrxGvNsK
oiJD6TMdOYrIUBKm/CV5KoaTd1hnw2O6XKl5Ofl4NuS9BZGGjfW7Bu3gRtNOYQUabokYF+5mV/u4
/MEtHARzf2OS9xJ9eaDLMGH7iTdyHZO6xZPncW7bmt2nxFZOx3Isc/w2uutkAG4yqCFgQjENveqO
aIVrmhW9mEuebFp4SWueY8y0aPKyeO6dkZIe2GlwU0wXJaTNOxQ2lZTsJ//o3N64yb8RZdnchrNv
F32a936aZHY2M+Aa6SLrcr1aW0FCyitf2+QAjWR6YH7tgmDtABpN2sLRqKAClwhXgu0Yyohop90d
JHHJw5Oxq4kkAYE9f5XBv13h1T9KTr6xTY9dK/NDHbEqiO44Z7qzVdyP2E7O044M582G5kKCoNLt
aIwWh03U+MCbNsD/ImwIjJgOim+ikXPTKZUzlLdKc+PaJw68Lt5jxpcB4xAsLzfror893enpAiC6
EWIzx3L6WaTyzf+uqZyfQKDvNQowXVe71GPB4rTEkOVx8kErVWHj3RDkv+p4z+wgkQYfc2C0zkQw
1QlT8wAftQytA//Oo6XNaiXWITmCywSfhHY79ipo24bmm03+xPYuylFvi9T+P750j6l5DL1g232v
FDkEqTsfIRedFP6o2FBYMih/hT7giliO38M9tsV6bKRs0WsXtbmZ05jlYfb9FhYi9MyKDkOJzJPc
B56tt5JgS+8tsCE3hv1NWQZ6Og7qnQlBaqC9W2/SZkgfCOPaQjBYKu4DfvsO3Yiy+WEJ0jg49PCV
RZiMiuoXJnqFFcoxCW4teIJWmQAyroEOp8SnZRPUESgaFcSPnTQnQrxijUMcMV5QVtD28Nh5C3T1
DPkVP7QddTZ2Nj5s9RZYYgl9G5gelnwHxUN9d6+gViyQxWJw/LqHaLuNaLm0jw3szwfNAznJZmt5
mkHvWW56zHeCO7eaxXfwg7mNfHzXwVfNMWI5OoHB1O1NMwDNJ1f10ma6b7zaCO4pHzURDaudIogx
qS9gG60cnczJrxAoBET7r3sExHyUUEvz+9qwVyWsJN1/gyhSW//8hwVJfKjIe1CJmUzZCqnkxU5y
I+pS1HkaYCkfIdfpHSzI8eEIhKGjeAnfr7oPBxGc8boGVd2xLfULJYekW7/yMR4XdilXg+oQc5ZI
uIf+tk94uTdo155P/pQbcdqypME4Zyk6xa7q72K43yRAQDc5pjybGrGz/f9lfAihVcvcXSL8yb2E
b77zbWIDcP8iBI1P+8pSQoK2Zs56yE5FTR5w0BXzs8HSHKmHTi/M/bEpQ5TX8H+CacvAuM84+kax
XQAV8R443M//e42kZEEt50QWBBl3CY+jHsEQhdmz2QNlBmsAP86FTKPvYgoN50ROfX9iR8nQ727n
fCWxque2HKMbIaFe/gaBGeOs/3kk+L/U8DztFR7cJoOtNaxQspA+S6J+G8zMm4Ivvpdje+KrCrzm
rs3Y3bEx/4EYys2jhJ8iaX7km3+VrWW/xjj/76Rq43pMotJ0wk1QIDR/uLYHGC/XJgPWbuiJUIhS
JTE4xPVQZj0lmpz4r9O7Ku8aZ58KsBMC6+vMr0V88kxo8g6mSf2kpk5ZO4UHLJk2REKAv3N5/wVr
YNDDZVyloBSsqeHg1Gw+c4QI/pZACMldpmoCozcbAV2O2KR8xDwTnf3zVeYBPE9nZ1xc4fHC9ukb
gblSGUMLDxrpYYZx6GuAQGDdFQ9ge4o9mLnUAYIRHJOgp95YvFr+gRXvk+TWle9nHpcLsJ4Ag1x+
7TY7IRx/uBTXcZPyo6err03eie22CMfb9VSQtaXZ0Z3KOYmrYsX2AehjWcc88zRx6dhxl7iNlVi9
y4//sveWaID1pe6uXIzTbdN2nYSjMRO5MyxcTyYxY1NcaFt3mIGohh1lcQw451PGDGjF7zXhCmJj
+yygzLRdygeVo7goSi2S/X1B1JoaNGTbbO1msd0ANUiGMfOgXPa5MENoxB0sFwITI+c0oTNJ3ojB
kDOtHfKXR6sc8Qk/HjCTTvQUd4gYF1y5y64LING08OMgQlhZj3+MGj6X1/cH+LVfMVSD/IGfWbB6
u97LJIuHAoYcs01fIqzWqZ3LQYevaTCpEzxqaksOJpDwDCWS0DO2shUv57BlC3YrOPbzbztEOAFE
39cCniw/HH+C7EcO+yHXhuJW6sdFriBljtM4QYPh/33pBjFsn9YAuJbIqJt1cet8p7L9wNXWEm+5
GHq7pHgfdkp4S3JpozEY5f0QmrOnSfnKlAqk/uDVFaELLf0DEFLi04TbsBZlnu2o9cJiechxdq4a
HijUj7EbYKpISKq5xpd7OqblAs3xdrpUUhXCBz3InS7yy0NG17lNxnlwLXjzphG2m4ZC2oCSuM7+
RYwVyxH1lq8x9VdR+9+C/5l7r1U8ItUmkDKSp2s8/eL/KQhNpxwOHapP37wFxcF/sefeF12rljAW
GQ4jnbTkgudPaj0udg/Pq0xRpzaPJ58Z+1yrZPfmilvzek+w/4fJmQ4NKIrHPTGBGDkfHjHLFm9d
h82v6ZiSOP3Tt1E3uPiU1wGwI6bGFaUwGLdH3cLQ1qpf59m6JHlQmq36kYZ0Pl82KxYfrtdYjAG0
N1/Nni4YzW5+HebD7jHRqIfNiPTIH7HT4MMAqm08W2K9hwizeFwrjxOltqWOKZmcijQ762cwxf8W
hR+EHkgSAbkBIkw5Zpupni6SQuCHjeOVhnDRY1KXGJHk7wMmAwHzd6ex3GuUVsBIqZ3IwQ0ehzq0
dr76BDHpoJUbyGT6/lySSlOoS/cyizuL5360WIO5PYQnnT4gmws95+XK0qPvRQoky7G8WesF465M
LQrAnSI1NkHO8g4R9/htSkXbw1lnlGN4D1DlRSqqPPjPJByXbT5KRMWore3dP+WnYrj4fAQ1xt5g
YMA6M1+t4K7LFn572yEGB/1f1KFVUDw6a77ISxzlg3c0zq36icgW/EoPGjTu5I6RK+3xyXP7p+M0
LDRnk/x09Ba3Udelwt9TkofSS83AW34422Ou2k1ydO5fk4FUgLJtpw9aB2jrNOjqM9is8mqMc6jk
BF/zfhOY7jDeUN8liPNZ3hxDfXGWO6uJuE09h+hH0C1MRRlPZbIPYIqsvGXRMw6mWJFrfr172++T
XwBvFJz2CTIaPXLlcirmZFU/+cjijiT7Zw/PZ53vvxyqpHwT5DbfTaef9S578IcfWrHltGYoD9ux
feycFU+aAJL4cpCPUm634ieh1Cw+67FUZwYeU7qctTkP8cskqNZQ/vNK+bhncIe/3Nhk4UiXn5Mp
QsozyZRWpaNmZA+QICZ2Ns7vko/M3FgDbpLR88JsjmbiPQ9PSVG+DHsNlRhZVkly7/cJhUR5c9sl
FsFU9t41aiObLiCcyb2cIMChYse/NBHWCnm+nSaJaBi31gqJ4EVEFZgcjhUQirjBCTzjrgFdwSPE
gPphxLblz2Zg8atF9T5GQ8GYAR3chZswTFIeOS4VpYlDk/BvcJrXasac1a0B13e+WlS7TPTDC1QI
rWTTahsSrqWf54oxM6/lZ0yLY9mIrayACqv9IpESTnV3V9FdxJQev/P1JALxCFogmQhgbwwLjqru
sH1XhAmNxKsMwfPCRnBE5kWVbT7ssEb668VqiKE+G4KksRsT3abaKrraVvOzWSuynIUnSRih/CNR
N2aOjKI+kyquKRJZdgNHj0dR/wGhoDtAWqT1YO6dQgkPmddap57oQ2QNUGjKlgsEGzIYyvI0cR+y
D4KAs74eQuCtNXSWFGwcP4vIdqpOSXgkQJNGVRYkt1CmqYBoprl+J2ryqh4F/dgfSpEVWXtS8yyz
k6JAHYnI6Y8uInBD2gt9QJBfAEjGDvBAXC2cn6ZzT7hHeHlVdpG0DxUKJdL1i9E0lc4/vet961gz
HSNaWbMwojg34niQlQTz97JnNcTlBYvf+Ncln/6yPBvs4LaNkdM4p77b5M+6KorQPdFchGa6tjz7
WvRkssUv7NIDhy7N8ti6OaLFw1S3zs+lW1clf2TqC6qUQMyMLwx7RacjtgNdDvuZwfy4UJUyC/++
36pcvXoVlZSDAJvMGLMEgUGA+cssAd29e9IJOItS3S5hea+93NUAF3BaiBDQwgOyygGOgNOoHPvK
tzMoHoqNgXtl7Jk4amCtsZsa5fm09QUiPpWp0PwZbAj5JV1/hy3uux16UyKO5tJQDMDgVBn6h4W+
MkKRJwxxd+bFp8HBMcO53NnuU41YQxXOFAXEu3VVk0MiMVvY8CC2whOeS119Drsano91ygIoe7t7
IYw5QhWOum9JmjVC+VHxKpfe6s1TQ66WiNIzwAvHUTFvjMkV63RIYWzrygAd/y/rgnt+cB20E/L4
qxKpr4f/S+tjnonboatWb5SnkzVXjfjQqWFwzgfuP9YghqUpdE3bjTO6gs23fGsbeGPRcjQHiZ2B
VMlgt5nw2Vw8Q2EJF+hreNkmz55tyg6bmjYERTF4X4Hlto6XRO2pWsCSQG3GhEwM6zFDMCj2PhNw
Z3xkFcuWMC0IR0MVHmI6BRWZvLJY761nBwrWpSOLok3/zEMujIyBcnC4/fZ8TP3Thlf8nqzcHxfh
AMYHqM630H5yUqpEEVOW0F+RhQfx9Oy6WTnuw0wTta6DTCpawvPslbZf7mB74SwsxmJTHAqvRwLe
GpEvkYHVQo0miRl0YtSth3EyP7uf9JVAPHGgeveNkjarIcqI9yKhOjVNPo0hgYr60W5BfgVZfncx
nwY+xFOaz9mMI7Gdr2bsNKPCde4yxzXfZsC5WwQmvREnqQIifsvOkPqiFT1SNjrS41djcw8j0xfa
nJwCJYM8QhqKj5C8OLkh6Ex6udPe9BDH03MVizYE7a8SL3NkT8KYNsIjMr0DSiB2R12dFy6+w56C
upN6onYKQdh+ZuOmiRCgN+eAghk41WdgOsbCChZfSixM76Cnw/DTZeEeMiAbJbXhQAcvU2kSg8At
BGZaMHJQU7/wBoqpx2P++03eth11AhKzLiNlgeD2iWPnTj68d6n7iRK64LkPX1+aOa2wwMO/2fix
C/hKZgohflhDMIzEmLBpsRbG6WIlEU3BcrB4gCCFl+El8Xf8ZWmCQ7o4YHVYPOZTg1n4vrKEADrk
F4n4CV54KQVA+SN79hzXEW0+F90ISGxtRCms9zH0P4vAS7el1oXeo/V0xOYQq5DDiRHcIBkIKM4c
8Zoi4MVZX2EBmq6C8UAwX6vPsGUvjS7TzbbLFrEuFUqOEPVvBAfr/yOkQhTbjXAMtJj7HQshh979
BqckAD8We+GoyjohlzFUJ+1OP8cIq1jODgwGRQAnEPnupfhgaR0FXIwhVbVhbp3/AaJq33CR6mcM
NYrMYKLPuhi6nlOCu4qoWuGI6mE1JsHrshTxXxpbnNjnFhAXPLRAMGE3KLuACzm1dFftk14mtfRv
lLNzSfRIRxThwWEZ0vzkGgCTV0pfAFgLxoIqiAnBRf2r45mVnmj/6WPGR7mOCzl5oywTQkvWRbDn
f/XNkfyu4lfhSOjI1fi5YxULO0j+BCx1Fp/tQKjzst+HcClPB6DwAYoDwnLSIZ9kIJzq9AeXZg+H
LQhRuJi0diMRVP/ZkiUctA8zH5O8mFHZnWtQiDGaAOXAasCom2l1F3PjlU4sctY72eGhFaoPWi3+
nJHt6+SCzmRIHZZtr42QIpOjFv0RYTWbq9W5YhyyULT5QVz1Bzc9iW5JrNRSfKxveehtbHLEw0/Z
c86v+ImErsxFOUYAQFtfv/N5/JUa4cE7wwYlZAPZg0RiNKN7swF/FkGtbl/myx3a9V55xWrJX7ot
m4FKb0JNmK0wMdSpQ8/9YZppR3k6O4woofjpdX3HitHr9Uhy7XK4paOZeMV7rfTqhcpL/qEEMHU1
QAOLPFESwAtu9hHH4UlwtMUSw7tu/4JU/0ixPg6GPT1ELhMl4hKv55LQRdxp3MTU+lrWatFDoy+N
N34xcLrCQpr9chKikWiMV91vXN20g5ZDRi5yiO9YJa7Z9QUOZtgI3ZuCoVv0QQZtoG4A8fDkD1Mw
G4zLbXkhUHzqszbw+loCvrpXl4o8CbI86DlRY25Ak78iJGZXX7fSS7tpB99uBPBmP5VyeuV5S4oC
sR7s4WgMOkauC6DUR4FyuEW5Wk2LuzupYdp5sqTSn6DGOpAU9klHmb7LtwCXG7ozneflwN1lT4Zx
AY5+ajIX9UZR6D3taLvFBpML9S0Nkc9elIYjZE2ROOD8W4/5aTTrCyAnHA6j7cXqjLn76jPNcwFT
x7AUQ6tKG1Pyb19QTHeXoSzH6Axee0FgHaf2X7Ob26RzQtxI6Up//9qb99bFRXtff/iTPO8dtHIq
3AluhKAq3dXG+g32hfRIV5do5YEFkn+YVIoXqS7Ac/cEthJesTItbZUzOWqUYF2RRd1U99BnZ7Fl
XDMcoIlAe/s7kV8Akcu92KrMqzMopI0zRebDqK5/DA7+3ebAU+ZDO+WSOpq0N53yHEWzHgTG51qW
mktIJMDIMdXbUJX28TO/X1NDhRFhG2Uw/SJ9LrT9HMFGlvYMw11L0qIdbTbhfMuUSA+ippZDg0GE
UC4J3GtfGVfcHPZLIvw6xKOJ2GKNVzJ/GVNSKFVansGMZSq8RPwS7qFW0DZCz/TJQ924Ic1qlFsA
0wVR7LgfTZnHNpJqvH6yKHDBD8J1/90SNJwKagCwdEp7nivUQTCFvD6illR2dLdQkU9pjkEhDusA
FUxxxUPrNHsTTgJhY4B6Kdyk3MuS2AR3vQpONHAePNbShyNy8pI1XYa22SJDN7Jmc3ij8cgehPm0
QrqQNtWYRwbKVyb/oCBKv2vrif+vMo7fhOvruBfzKdHd9KGkG/5V6gZB34X4q7UGrLGRTyXmgXi5
86Uffpyk0CpHVxSMfUmBew7vtqrCFaSuFEITHCldfj6G5PK+lNPAGQP+JlV3UzF73B9/qfPf7Fva
oLjVCfZhXGEUb9Kj8YV+cH5HXD4drP/e2LSgLOFI11SSrOKBcc+Of7CNMjUWWfGPn5oyOjt9uwZj
9Zx5QKd0s6qN4PoZ6zGWSV5FxwW4pBIpzYpVuoLXVRvxkBff/QXKsVbTNhUSRUzTrHsufXqDksPX
UDanvCP86QIfFbPpCRUGyOvtQxut2b6CIRl3uVKqF16i54jhkl0lRj6htDv0pYaIHmHpIE9eXrBG
Iw6oNv2/DWsD+lhHjbYg8REJjRz0uiUk54dgXF4B4cGceMu4R02SkD7mCaC+MTXljyE6CvCrgQPz
Vuyiv8TOJS3ujYR6gGLqRm1EYUAEXRBKL0blsugwr9AdrJKp2QNgg/WAWp7nfOoiVFLWGGEnYAqX
hgCezEfXDjK83/whmLeEHGyyNere/aOIGxnJrJT7GqVZfkhn9Mx/RHxoa9j5TI9mOS+VbEiO6k3/
/+R2DZFRqUZEAaDzgF8LhfFYoUKIdXQonlX/df23x8YCQolFBxhNBJ5iDU45To10MkoRTBEHmN8B
NxpGISETLByDA696s3BJX/cXYMU2KpmN7phGx4gzPg+9STRLKntyuUnf0mC91oOlrdJYFZa69LnD
GJ9A2LF8pjNW69kkMncg4r5qlPsyWi2/WfdY4I4AFUqsn+18v8wnrzP+/FkPZdO5QPwwJ18kNJ8b
NajZlLwEz2aQWyXp0wZoyPyiTuvKH35taUmlHeVjEtbX19JFkMh31X6QIQ738hHl4uu2W2m7xrpM
wdqA2EFndv1hLWlZD9AvBN2HabZAxOWbZsvJb/vHx0p6PUsjjHd87QfHLGP7v1ch5GxHcDx3timg
up1KQ2wexd0mZGAMO5ackdQutYuHG1HIl3tZCQvAn3wgD2o3uI1Vo2T+HnIFZdVNSOZ8jjSphOcm
5tylhssAZ62xAEA5luyfMn0CzdG7E7Rb1HatEe/jNrepRLwF1+7xOT4vNCkqagLim4DS2Dlh4m93
Koih9Qoer8mVfpkx5N30hfw6m37nn1s5NoK3oxpO818r2AogJjEOECNTiCnhvk9UmPoT9MJ8shdO
2UJmaCyTDiTIMK8LLKGkMZdWyI+jspcWJBZXEAJ3l45AVqF4IIkPSTIWBoKHuKdBe2g8OyGvjUmL
hy+4MF2uRU0d/lnnYcCcnxopCnk4bpnZZjalcVGaQxIsOw7+Ut2ypdVjkN1g6wlqxA45rMPiQdko
eU90kHx9A70bH1wR+GIK376Q5L4qhuR3AIdXRwW5byhVlRrwR8lstSMER6R0aCcLPxymHhTTbJIv
YckhPP1d9toBZYnvEXoqiJb+s2ErhIQPWotszvPeT5MzR9mUN/eGhN4ewdwCHsVh3zeBDZ52zaGg
UiJa93mpuD9XmnaRV9CH0YyrFOeN4/YqpcsD5aafWpapEz1hQWb1x7qDzVM+Hp01U3Fia1mhYQSv
2uJMcZ54G4jvBUNWQb7gyzsWRw+GLlOyv92aHHZaTDf+NMI7u2WK+VA00wd56kQrpWohMaqOS73D
X0BO+UgrFqqaA/+DfaQvNMT/5vIGdkPlPMT8hrDNKYDvSeEjbnCWeGw3PeV06sZms1gjNkG3VxDh
0pm5OQ157tBGikApCJJj09kHS+w98a0LvAY6g2zpCA1IQmIHqeNPYoGPKGQqcvm5p6c8oTrihp+X
MLL3+/ZYdGyb0nZdOWGzp65QHPnLxsNkTbnLoYOL1crYdEoseJASIeuvpb0XjOASunlJSZoAeWJr
NIh2Qr7u0v9dOPGx1xnvPRMVl4YCfeoj+0Utgbkj26GvNtXVDJyP26zPdSjU/NrI+VHAWDKDhcrM
PpuLpP0RhbBk862ifttAuZP8js4lc8WvabksA3MZomkD8RITQp7wslgKpRv+aFl4Rlxz7GphBLrQ
+gjC4NV/lc6Du2nyejK9jwkfjvJyzIoO86QfQ1/nCmQ0e55klRT3MgN3fgvAeq14zmkJw0skj6wO
4RXLa8ZLdvh7xAovJVgukOkcwdU5/pr4gpqWQECRe8r7ua40MsrDCawo1QkaCTnyd+y+MemLeNeH
BWJbkCTRem0CjoWWDcZGMC8ue4iORXYhvWu7f8UjZGm/wQ6broTJc1iqizhkhSp0X/ARJwuicroH
X7d6ojPd73Baxb6yvLLE4FU0/b344gB33iIZ5ypBkH8FAtYahajK7ZTuRLlp3oJ69qKpKC3IQinW
upIZPgrBGg+PS5M5qqWzV9MwKxvlsm2gieIQCBLy+pEoi1FVZMhs8pBIBEN0xYdDBugT01g5eXDk
uJ/XeiDlSKR0byQZtxvrOrfb7MBtus778jEPRSaiDAGUYxl0U/dk0D2qNh2w4lsOcN03xQDBelbP
zif+QeSB2PVUaAf9EdrtA3Xp52z03xUfhA2Tb3yHp9jgT3sfKb0XU4HnplfpcErqr5X63djtRDCE
XqTq+r5FkI4W8HH6dBGWs/KxtW8H5/6o+bkt7MUH5br3JGEUG7AH3pgLOKdlXTYUCQkk1pc0uKMR
ggK0VNa/laxE5Jo1EBrmv1fQmmb9mv2hAZavbaMaQ049nBXUB3OB00SLe5OZz0FlNzSc4BH14hYF
kwzoBpS7A0oUOLMFQgipq+4/EM0Rd3ZXxlTXdHCJ/ev+RStjUpOVxzaRjCc+SbWw8U4/SYWDjDfu
NQQouZ3wQ1EUsWd/z3lrw5tXoGCbqfQClI4ux48algAvPqZWZ39OxuywGK1hfax0CXYjZ+rD0P0w
DG8Vej5FNSJaOiPVl3KYmrFcj1YZFKxeOmXD3bK2EZMGhbYDlksqk4ROc7arqPYFb+O4sGwVen0m
SXdI/tkZNQimbuka3b7SBn6Uk6If1b9b5gwT7PKD/lvSz21eQ9EB+xtsZGJenabndJ/aAqRQ5Riv
XOASC+tL+WhNmky3yux6TmMWJ7N5Uu4hTPOVZCPOArUxepwRX/L8vZpX496GtUnLeeSv/cAnXOuD
rVZ9N0yi2KEpSCe45Hv9ATxBKtLi0pAl6bl3OdBS5Mfuo+gGUFFlmXRYj/Kc3nShnYiETira2HZR
+ObOmh/+eIuOSUU3beD2QuQm2+SQiLi2GVjsW82VFGGFfjTKSe0wsnKis6EwKrKel5wO8l2BODbF
M3gu/4coyFt1GgUee6F+F7TWOAFc65wSUwvEs0mJ6SwVzMq9NXSzEPDy33lJi0AsYviPZ8dvCWPr
5vW5rVHtPA4s+5fe2QNJBw70bJYGUSNhaFKAkHLMIGjYLS5xCBO2sgMBzNbX1UPIZCn5RtpUmDzI
L0onvj04njlNCaswwP422rTMpe4VaSdWkRBUh2eSZyxOwQFJGaFqTjWYVKb3bdV5LmzGCQblx1cn
q1Wcii+VbTZo80c3wksROnQUhiRiqDVxnaccrRAMFCv1lNn/PgymEQEdgI3WsjinR6JGG5wjR14B
4OM3C9pw7LzbEVrIyJpvugvk78l+SVVmyRRM/5jm09r3tS3Xw6hA66MfPXj36N7+oYtN5U2qKAIE
9g2WXVnvLgNfGB2Z66mr+AAJyJr2Gnms3ch4rT311wJUYWLi5kPQR0Gycam9N5NKQRYw4xLcAkHP
vP19uAIt3o9ZF3WCCkfwld5LBaKb7V+Jsmwkj18ezG7S8tbhwC1oLxHKUbRJ+2yCbR2/bOx6+fxe
ycVk+1TfBiCsWgDp5aC23alQFLscRHzOWPjt6TR/3QE0/d+If+Ph4oLAJKvm4oVpKjIHeU4Bh9tz
1CJhmiFWBDmIuEEhalkGGDLyGORcsfVUVLmhHKj8sX/MqsQKTet7aiHpdFiINK1Dj+TE0fphgmqn
2NgdK9XMRTtuHXiEQRKKfowVLH0825lg6esn4J2h6U/qGcUiY1qI+LWuPGFxHrKlFMWkGEvm/Avx
ciQRLrHjNg91yhaJYmMzSleWmB3JFBcVqwuIROG0RDCqJ8XAhTNZhhXhYmZVZwZEuasIVmWYMOD6
vhBTCxDVPfjcEvlAP3rvfkllBRtWFRhVlx00CiyrA8PYL1uDenzPxFgdEnEhbdIJa6L2VIxXg3wj
NtnBVjWzInxixlEfmXXdSFkgmR6M7mBCwokN/OSnxiVrc3L4Yb1XBiuC76kyvmLHWxs2mRmtLmQX
MAXxxmFLLfyRHxOczN3egf1bZZ731vng/aLRqBbiFAZknBnlQNnKSuK8CDBjyz4GUoPQyWwvTsdC
3hmPBIDKCZBLNpAoCg+y2eq/YmSn/dhFY4N+eIX7obZ/kQ8PzkVPHQJYJFZYLVfN1okWDSb5o9f6
nXwgXucMBdy73vPBu8J/CYl8IBe4Be0rSpRuyUaf+zsNuz2UNkvBX2t0oavxRGPc+I7kUNL6FmC2
yE5IGsYgMoKq65lNBTYDpTxGIevFc2QGZNnnCzWzKsoAo1U8dNzeslX8k+NRjpBewZg/fJnQzi8n
PqSnGn+i/IP8pl33hi5cBjkDl40OibYHosYCucJtKChUTD4oYFzavIIkKN7O3U18l/ivDK4YxumG
qeRpTDZO6NYQOUby03MEsO/gQxgLU0sH58WtD0t6VrCn+eqMN45cYRPSt1xwpzVxjGhaltPOpjD8
M0N6SI89JZiF1LMtw0b1OdHHCq5wgtsRIgZ2T3EV8tM7xdxDWpvzAtHEwDfoGDB5n4TD1Bjo9B0x
8Io+Ma4NMlZvXcwJKPlnoMn2BH3T0k5jwv2k61cWUX0+J9esXv6I0WG1O7AsdnlhHxtYEEPirEIg
YC42+mJQ6j3/t1lE0V3JOdkWOxZdHnxHBPxJQpi7ZRLz3zmGpTAPciiNxVZhA6tlqzaqsDZz5y6n
yCo4UoBcrAfEej21smzdG3pfryjA1SdvfFsqk5oZH9nU92eDfbaHcUL+sbEU4iBY3izagB02GD1L
zKdpIObOn4bBUJcFBWHSAEa6ho9Ea1ie80F5+smojHekaXBcVOx+IcWTQM4uqRIm8vTGaSHNRMjE
wdA+Ljp97bv8PkaX3oSVQriWxX8ZEelwvmlbV2J3xAcd7HHXDFOWJWFYDDdzHzOezuzSepHNK9Ax
r8cSZV0rMsDj3jLy2eP0GEuqwrEbnEJUIht+iJybcnN7j8M5Uu1e4l3xlsnsQ/AGui6dUm4VXkx6
RbWrRjjgjWX62oRToCajkcLHQrOc96ISrsOPEsuaO4p47gqzHbd/eqJbrgCVlXYlQacbWgb2ksFz
9LvJjKuoq9uYefMKyaD/NcJoJ6KREDFRvDIL6UuoSWWfAuEixP+0rjNOhVxxQvjkJOKhQhJMHo89
B/jBkrtofmq3iQebKGKcXg6GfIwJY+kMh2NBgMp4Wdb1uYTT9GKh+0osRKX3CK/MM/+8O1c+8nya
mgU53cPSNJGYPrxNV5A9CGDDwslSqDKolf4cN2QXyxsdVl4PcwIz3kJ+o8OeI5zg4sOzyzARz/ZF
X/2rh6qzPvhe2bQ21JGgi9AoFtZRx9gJMXSBGhJwbdXtAH4/LeDeRkeK58NEbtq0AXKWr0P0lTCR
Iys4BlN5RZFDhnl6O/ygYJq3tsGwO/v8JNLLAKofKwZ4vv7CjUfa3mzyhkdk5KQnNOCAZ4yJVJGk
VBy1GwEqQt104diID+R8EEjSpvgw0qfFcib/JBlOR1auPHHWO4rbtwPt+/0qPPgHYo4RTQOlATy0
x2a8iIQw+S2LZGHAZ5YpXXWMAOo416FNYkIvxr9vRE/HUxfhPqOTdy4A0TSbpHqlwI4rBm6qtfZb
XTYQIPOdYiGR1SkX7JS8hJMDuoaijUwCbnlX/k9nfMhLggYblILp7oXWSW5bO2FMnFjK1wbVggmo
J1uNncH7Szhj0R4JU9/WlpmU2oVZhZGHWaA/HG30J7rzoOCW7mGYEl0dg05zH5UfJ0Ysi9df/Gkt
6gXrtCAE5c99bD8KNRSZ0vVw4eatS2X2NJKpgKW1Z0ScB4lry2a48Zi4IwTD2TVHQ77hDh6JMwTb
a7NBsM95GhGfhA+Xj+PYZigrq9jSDvtHN4qPXJ/poRm3JwkUz9tqXmaqxXUImmoPZ2f0l/XHJVtE
lpL+SL81EXwzYcA1WIQN94K66GRwS7nqcjL6Ek76T3FK06SO6P0OlUtC/syM0n0Vfyxbfi033KUM
rL322FTbIkR7XbDchzXSyRZ6jj5dNkGYIxZ/INzefi/bebdGMSDZ2w1IRrg7OWIGy0g/BJVFuu7Q
1G9XvbFr/ho9EIG2LRUdHs3tPk8sglfurt5HarHTqs3UFFbiReqkPJBsjTN8wqAA3/9hbujbBMbE
oVjtDKkBeyQWTk55da6dNF5V/1eu/SgjYQtDWYyDh0WVfzO20ef/Do4apRw5PggJYGQSbV9yJFmM
ZfE8Bk+cOw7onN7eC4WAldHPCGOC6Z56VU03NLvXTtSmtJrHxnowJ9v9xDX+CRzoDTj5nGPHqZfb
NK+Dli1BO1VFQp86bG21Ve5Ww6AlllGYd61ZS6NXW2o6APMga/d+OroFTrSILtyVyNh+QTEFUxKS
O1jUkeCfH9IIcacvhuqszlf2pmaIj1TkQkEVWmcLvoUN5MZKjfaTmFg9lltAdHpml4ecyRL3KCfS
AyMdAIPD3a8LUgRM5gq4K6/8ThnSMgtfDmb8ASoNLcS67RuHeAkignmW6cNhEW1UmUwV8VRUHcVR
xbPom4Ph8kxs9BVADXvOWT7cRs56+eTF9IBrWZharoJ2vxIbkpcDfs/izisSuBoaffqE1QxvtwEF
VrB9TfkC9I7g+1BY+pFbsUkDFhL2F87cW/NXMcBB/oQy06h7sfhgXF7EBkEEdKxxDbiXzG5WisWz
ffzJJMSPce0iAUlWh2/GJKSUf6xSSQRsYVQVPC6sC/eTWB/5FxAWAQ3NT1vT184fE/N+6K6e/U39
0RcUG19WAhyrHTVmgE5yi5yFACgi6uRpQzRl7NENkNl5ogQXkAKQypu4WOMaUgtps+8s4/oxr6sd
uLkOn2vMqhtsmXjmFQTlBf+8cI+QH6KQ8jL8C08Pja3z1d2lfsCIRUHKBL3pikTas7axUMN4pX0w
qNyooBPnibmuwtSDW/hK2bwiK4MiuvRU4YA8WhnwOHZxUckvM0wgmcOEYNhxCp0Zl3Wkhsvd0XQK
lL15GxVyYMJZUDq7EwHK5xClzNML6bLVxC93IHHxp71bUxxQjOXEGL7Yt4BSTyF7z5quJlQLm1Nu
1wlewwgFbHo2aoDdd9JfiB0K3HZgKvd7HtLAmoY7egCUWnPmsTvEpKUzfzio7wHHBsKPNUTbStWI
ienWmF6zzwGIICw99M7ntEKjEjSrBe688FCMiPgh47Ly8Kef4c8eZqEWYwrlrUwbgvD7fITTlxHF
I1gpOwr0ZM1B95PC4xoweFzTQXC7f7vRYlRr9QWPFeycnkozPybNN8biLS42AudyULYVEDH1Hwwi
8ySWXjlY3B0f91fmIUEBpUIJBsLNjWyunl3dC/kWsdJiP3ubaG2VCW+BO3Q9TyY+zuZtYicGXW/J
zvTLngz38vpNw4M2KNmtfdR3iiciwFRk9UBykpVZMsZACfY9lSkN/DJQgR1B+CVNKUOqvWaVpFaF
4iia+sW3H4IS6KGF1p7uwT/PAVy8fjG0Mz2fBORqHDKbNZyZDAVb2rVbNihKcyGIA0FZ7M12cAyi
iVWsAhT+ExHlD+BDxNCy4VpBBgoxPG3d9xMrjMyw1L6Ile8x0yquDoJxk+s2pXZU2WNbsiTxN3UQ
mQuEJFnguF20INdi1I7P2g+Kt8xWNta2jzdoDzuzEvfed4XUuqnoqdlKcO6z4sBqHpXqC7+9Bi9/
OiEc28cXbmbDKaSvUc5/hX5v6YiKRvDEg3nDgTtgrYQ3RkADG50kZPB1oZBSqKtmIY546I9peY1/
Kz//gEKlbRyyKOfp56k7X+V1KSATFz86CJaZbFKIN4yiU92ZKGOEGfJgWxqG+fFg9G4M+71cokPP
KMawGH3YSxSVYWEqxNkffJAxQs+DHiXovABK4tXTywIf/8MzJbTseljNHZbw/td2Pja9CmMNVF3J
pr8ghfl4BsiaCNUbRX2OJrB54j7B+r2PnHEWszskvWVAXIWKXAkWBzH0xOKS6E04kzgpeabHReHm
ZCTKjJgsQye/t6wZreiMpvIRUBrke0esopJpOqrx1xnIwndLHV7wgml2cU5ifzltKIXnEGLj02sI
eF//8ioL0eKDqAkFHvTakS+cNEFsxZqB1C23aIohN5VnUu8QiZgy9NJk9yki3yEXf58NbLJNjLTI
laJm7iDyB0SUm5RwvpdVzPtP1mSXliDNxE9f+F5KcWEmlQD73Fnxw6a6WMQqZtmQtNbOvNDaUn6n
Dzpr306PhRFXmlbbxXM2Df9T5eX/sRpQ3hdylEkR3Jn0AtybhoIsO4JCKmDi4MVsE/v1OnCAyJRP
qyhtoa/KIRDgBfx5vnu4sUo+WqTscCPfmlUunfubDraVLrgDczeKt8v1IvszYMsVgzBid86WXC2B
8zwK6Tik091UyoRQX4KmvGhycMUtdP4jIBrcYqyYNhkYAbK87CP282m/2r8HsefZDLhigNszxYV9
IXgiXCIMwfizIrxvVsOkkPQWQg+YeuA/MYNWDN4iDlImNVloQT/AU9zQCI5HKl46MpRzDkGT2EBs
YP1msJUeRrM3+ov/+FfD6E9bSAQllq8OdHUjgMO/OD4EVRPv4/zlvNljygb8vMAWkmOdItBh+i/P
XzvToaaCnteGQX9BxxKY9m8uE6CbHEHECmXo/FyDK64kE92pY4mk18lHHEpi74nDWXG6A7kir0KC
fLHExe4pdT/345wmtbTjyt2xWxrpCOttOWp1zqCpGO1Xq5ddW1z2SN1yBDqTU1KsA0BqTuLNWWOU
4lCrYRudn7qZL5zdVYJ6A7QFKOfvORwdIxL2T9NQ68VlTzkVMj2rmbVUZcNAm80oynYP1EAurBPr
3bMjkymXz1igH3xjNRr6b4dqiprpge2NPshlOBiFWNgFa+zEGewAVzecrhmhcIzcgmVghpzTnU3b
OPXkDPYm/RqAhLT1X9abS+pe5J03RUtOOkvQe4QBl1m4F62/nKBbdxpsIM80iRL1TfsomRM+N2A/
rmvd/KdoJ/17ybmJEODAtZRcgjlq5hN5IyPzl24aqnK2o+2etavccilYe0mYzgiMOiF4BC2Yn8uC
mJ9fZH7CKWRDlO1b+pZtnAkKaC4mVy/ZcUsIdZETr1lDN5t8o1Sygb4bEMd++3P8sgTUqqXREMcD
hGIJtvibht/UEHYTAFaGLJXynvzDdXkpP+ctOHCZzROYpPMHbpJXl3wkyIIuCV4GFD7sagbGdIgC
l1KaHdjzC6uMnFQXdXjBAaK4Gt7PjPmfty5G0gYJcdh5qlLHE8q1W4P2/7tAhC9DTiiAwG9EGZ2O
HQ14oGEfob1TaEOTPZy27MvsvmrS79Qy0L6K/sSerb5PRPPH4R1XojPpKnkmX3JfbOodjJE3Qlm3
RFrCzDg6FRsnrRkBHF++L/SIgCpNHaDXIFzZV0oHpuYXU/w5IxQjs339wvrzwq9AF2O5esVAXMU1
TcpJH3AW3zTaHgi+Qu8Fi4faoSgas6YdhmxTy3rftdIXV63PzCUgIgOp3PYoLnpN082LMhVJtCG1
wcH1TW8bs/mFfhkFZdhYPzJ3pBNBETy1qKr6cS+4449OTudJhbijhSHjcELaGnH+JzkCZ0LSXLoE
rlYW7rqdCkfPBKWadclQPtX3/qYgrgXA3KiysjeKvAR3yNjfAOkglz1qhUnCco4fCUlzd+xfvlKv
LdPvK/3A0ueY2saN3PB7/AfludfAvsiqEk41YbVmU43OOPOzpDn8huxYDjaxc6ztKQnP8cGPkZuy
KAIN1X0qHBNjQ7yG/9lbVlGjNbpATCkEHxtF7eD2x3fFsFm60NZ4abth4vCKe20LKe2UONAwcOvU
QwgmB2LlDOxmpOwf1jBbjY+25jgj3MEEesuwu5jazkqQgv1Hdroh2D81wdEt7sWWR0iRnp0oOq8p
HeszC6gRUI6OB5xM2uBwC4HKuWGePLQQTTLqHd3wfn5hZJ1Q7v+oxBKI1CK+CGHkiRMOY2e01auF
xAlUGX0q9Xx6oHW8Ua8rgNRkT1JOHu0/+Uby1+NDGrnX+GgTlvNXqP+1l2cvxV8bxLXHQMvKy6ru
txlWBEfJxIBEQLnLAh9MlDAYF+O/1I+mYyJ7P89QBODmoafDbV+vrMC/b3CSr4wmrt1Fi9nQPCtd
yJrndW1Vw/qmtpRp3tttlT7SU9fcYaSTcCgHLHu/E1dkC+WtlefJnorT0hhGvs4uWBZKS3B8Gcy2
3TnzacbKDT5/I2uzrPpNiziXp1VqfSPwqeGV/vDhx8r5QWnlGV9fxQuC0tEZeYdOAvdzS02sgLlm
+2nXMpzr/OGmp5ipryWYgxZpH+pPC7n+D3AhcboEZeZkUTl2rYrvFUn/BYUNiASE9VroCvtE6t/0
MBAI32p1aLjAOMs44pGWU2U5loDHdECLbgXuaqW99Iwen/8BXdD68Mj66TlJTjpGiEBsjSkLHyi8
3rBqTxKkCoqqOF/nFs3aAN8t3dMUKUQcWFEL+eTOOHzAREDCcY/dwTciY0DvmgwOXsVyH+guLu6m
tqLkZO4Am2hBzaj8LX9I2UgnsCdfRkfILG8pPu2/EAEV9cfBynYAAYd7IuAkkA+Yon32pbvgWGEa
5UAfnHJZwQpv6mt4BTkKpOPZpeyu5ji3UZnn0BJ1EjlNpmIphnzMU6ehPDpKgMizRljf9HVb8A86
K8VG4NQc1dAEmJd1FjKzRN4UWGAL+5WZIf0I50tpnamtEtd5JeAfXtLEwcTkZvD+AH9u+qKmjwNL
br39hCxIDhMxM6QWVZudo5+/2mDmbjcikaDiai9eNZ3UUqJBHJeFVtFJ18Ks+PvJxudcE9htj5Pv
sJf/VG8PargrbzW2UZ1G/gnHTjEsbl8V05kLSuY1vENYz100NtsoAncWPDSyn3QJww34e8Xvp/SR
oTN4zytYh12Tf/msOdo7jQs0eA9AoO+MzrhmimQkUxFDnlXMtp2GA9Dc7BuoF7ukr+O5LYlzDolR
oNvxkXYJS8srTAuNWvBKy88+P1TC3VnIRL9geUcuw29yXL69uqhBcj3qX1iy5itSa8QihgQ6w4Je
YXEwdJ0bRX2qwgYHjOcsPPCiwoFm6vIpKV7I06FWl8REZ9QiPRKsef8IoJWMM9rclfUi6k8dFJap
owpxUuNVea9n6pvABpy60lvLvBNvpQiKX3LWWJBf2DZAQa0y1fLGjcdtKmlZZPUh9gVv4gXheYax
9OWBtncXdVXIjtakd8g4J90R4dlBQrk+EYZrKDbW05P0Ua0kjpyDdNZwy8i6sq9zC0TyAcLQ+XnB
FvgStNz5dVbvueAvZCqWgua6m/UoMLLS19kRWRku6x1qrSGtsYjjJK4ji4nRzhFncl4162CN+k+y
yAjN5/fw4lqV8KZopZ2f+cyjciY2KGBCI50lt4cE+HaZUXJmVod40B8JLhuQxybeD4Tv4yREmGRD
ydM7x0AKsPsthEWA6FKZ+rZx8drkcWdxDrnk4+kFiZ78Na7Fdb85rkKS2eCNnPavuaQ7Sp6UFLr7
142Xq2IVteSiFrnBm7WidDZBVqkS0D6p1YgPruaIK+IpokS7Lp9nhOfEb/DZScsI/cd1GF6SSrFC
kjQhgbonZBRoRDE4Tyrn3kiT9oWqYM20SQy2cSl3kYmnXD3EArFI/WPf0zwnwyLqJM5R5j33Ze9e
5kFcIYu9aCNCjYMBsaGcVXs8NRxCZnUFm5tItdQQPmuU8DS6Ts1YttL509OW9JtE/IVgtp9vm9KR
OR3p2x9XwRRNN8Ea5q1yu1DgcrOGX5YpaNvgGuuNqtOQXXRbMTKF1Ldp+f/j+iDpW8GwfQKEqGYW
aKaXegKcutYV5WxXms6vnD29ksld4XncI0M4DvWz3sMRtpmOqXUaItAGw8KD8zy6P8uJ4Kv4VtgX
MZZgVVQECj1M2nPQ3RPYApEeaFZaL3KXbf7kq+iyHoZFA0z9+w9/JCQ+rDxfKp9L4oS6Oc/7Cqfj
+qhsgaMan+LoiYVHUCYi+O45bWqAEUZZKnw4ZYw3vphFWKRxPeI5WnU+Hm/YSeXmYdGpcXkLvT4N
ai2m4GRpl0lxAKgwqHoBcq1zVX/sT2+8PjLIT4rfzjVdpsM7vRi9ZjD7Se8AaTn8auElozwk36Fa
LZlopVFaJ2B6Iej77BTMVYhCAkehI5vHc7Op+3o1KPjfWvNujLZLD4WbG+p1kN2p7AocILc8kZT7
5xngmnqlcAdJrhO8uUckpUMQC5cdkfY3Z8cn9P35UJ7UaRYlWeBDuMqGhn7KXlu2otZN3b9yHuON
d5pqq76MssWaz+RAPFDpTfqRic4uGNQkuocJdlo0lQaz4u18UZtHbSdQNirQUD96dfyx2ShGRPTp
bo9wJIT6wrWWSAZTLfk2KCxtKvaQuHXYo42n3QDljnJQcFyDftjYKsCLtuvG8GoMbADZU4ONyq76
KFhC/plIENBIbalu2GbTvTS+dihqfQqs1Ri/0Plt68nCcPQotEDj0NAQi5ulpAdWRGtFskrs2d86
W3T5HtEEOHGrjq6k1sxW6oD5LVaw9s8jtPVbY2pYrDYidLrUkRC4FkvkO0tLvQuorhr6EvhijVX3
RkcK131d7Bx2tZzeAzH0S73K1ebacHxP+eGqc0yfypu9r5Y6qdOmWsx65U6INsDKizyrgLBwxndd
GjCyiMs5AwOVZK7+FXjQBASpaieMS2yyveEl9vz3Bcs32HjUbfGsPCqEb2Yl0F8YFOFeZ5K8zVpy
8P3ijHv6jDXN7Dz0dsFdzocriQjdPuF510bffE9B1ZlwYdOl08Dpzry9Ntxi7nmCM0knaPHtRVIQ
i2mtBywVn8ZSoWQkmwMEPS8gp1eYDHzmHIxjW/Gn2+BokFtCwQAWTb5e/B1GZNUv4cbs0q/1b6BW
/8rBdk/Z3B0YRG00BDefFEUiSVdbh2RH3ljje/SrL+d1Igux6UL5MOEEEzmdeIsGcSPR1ubiHRO8
eFJjkG2Ysvz3YGW22YOrkT+n9gCCpip/4bOr3ivwbmPHmgRbqFhb33eQLQFCyHo4TmRe7o7dLnQB
hHyLdT7rNw/L7htyx6VP8VIj7DLh56YGdgGhQ/SeU3A/7c2BZcB+YN18AFi6X2+X4QqjGhsYhb18
ldkfFD2yWuB+cmsIn7MYQGX8TMxTrSX28YTjkwuT9qEjURrzuCblAgW3kJPORWCbrIBNZ43tivvj
71pzTcLoPfhP+3mFvVL4alZEJJO7VPbrBr2Qe8eSEmt6CiKHfdNYLAa7DdiB8GlYIkb7EWv3E+3V
bxdsYjVZlSm6FMnaVM3prIwoxPiaKr2CrQU9vMzIdrz5rnkZjjYodv5E2VF58zBnZXiGHSL+dohQ
CJBkMINstfSwx3PBH+n3vX0wBn4z/P5UlHbNUnab6HmqQVPL5Z4C2XjmOu11ixGCLiVRPrIP/6q2
gzwzPo/Sfyh/8xOfOiEKaPaoLTDRvZSjcWkAd3xpJgliqtzV0DPKvmARP0Hnd+IjcH5LeQxuz7ov
sBf32w/Mm8PrfJX+Qp/SbUXTmzhTjV3hv7jps4Ou0aOs4GSqSiO0lr1bqDU28YcRL9YuwBxaEalu
eYt9plsNhKmZPg+BsSMQz7WcPwC0ZyWbhmlMDA/ppuzDW5kSuboAwa5E5V7XQynWkEI1ehhkhPwN
ly9+bK2x4rlWR/fuXdLpFY0XRxjpzSVIaCEqqCtdfdhxPczLpCXSRHDXnkDVSObJqPZlMMYgVwr1
LhpGJpzp6jEdPOZb/IzDJ67eeNmOfp2XvajIApQZesKda4wie4xzesiBMmagUeBNpcsk6lh/yiq5
678HpBRoFYOwPUv7dJDZtwQjX8vCzcNgc3392Ww6K4emchmybMaskXD1R2IKyED/xi0PJ8maVhaN
XSQTRpEVXtnsvElrqmOKguSBzDhOIqWV3PdOPlEi86ek9hpAng5EmYU3xlQXhB+tZVO1mGUjhP9e
7uqlmyba3Ye7RGqsUYBhCTH6lYMHQrLidLaF+Va3jOyJpvlNWv1+ndtgQbijGX6f0qIA6PYgyYBa
XHST+vWaNXMQrrV8mYANQt7T/Lucht5n1wLTh6fH38NPJtBF6PQmlbJ+0Y9YDsjMvvqoafTT1RvI
b4nqKvm1t1f7ngo3mXP1yT+9uc07C9kEtGF48viVDDzrvUnkyELA3Q4OA/TM2p3Mi8ucWqAeAmLr
du3qMx318biiy2wveQCcqnciwQZE7TldA+SM6RWunMuRh3TuGH6PGBC/pRSsXDk0b46++d1dh+7i
IuUWAGd3YtSZ4Npf5bVKJAC/L30QwcHv7laqYLFvkeZsCW0szuhXxpkOtjS8HxEWUBozWt3cwIaG
oxnrm3HaF8D5964PhaCSyVmiBseAT04myM3yjz1pc2AnqespdES8n9cT5lAAiyrb5Lp3c1r/dytF
PlaTb+qNvcSCodyDaXT0bomShPjcm+SuvSUGQxUnNAFRoMKd3b7wbXlTjQxMp14FWcM4IRkyyd0M
8AjD59Jsq7XGoCgWDO4lodcs+s8PpOS8KiBT+OMfLSd/pGUsL33dEPvUvaX+Hs9F9nW5Tu0s483J
ERT8Dqa0TnCOPdak3nvlstz1ib7DKjg71TQPUYId0nr51bBjGSR1qTzPTXEi7r9nfKHrtDGy53Rs
tB1pY0OVYnxvU5PllyXk7cTIYKReNdPcXUJwy4Nlwng91KJNsB+8sFhmvnCJnBaAkhKbRLhEaqvE
it0DwuxROr7vY6Ax/i2l63t2fef4zx5Hx4jssQiMHVziBkXL4ut3QYKN6cfMDWwFFKl1/mQK+Yyg
RwTvPltuhv2jUfU6NY0s3NYJhJUFo5D0R2Ui1URFwYTh0G+hodOy63PtElHeBRl6AEJD2eB3yD3S
HhysxKvD+tTo/JRfu2eZ8HKqOdbEWWtSFXqmyp4SE+CKICuG+GJiyxILkPNmfcpF0Oz4VEy1sgAn
OFt/azWuij1zn6jtsBBti7HN/eBhDxG4PjfnuYNPjDU/RU65xVMoaNsQ8cFdT5ZqnRdlcRXLcpdL
HTacQXPPQmO96SObYOaN8w5RGj4bA6yeYsLDGXK/nqEVfUXeBQvfpvd10MMPn1SOgDmOW0vuzWQc
cku2zlOrPaKjnUrnaYzZ1sDuEgMf5GW/V/VcjoxVriCuoAZwqtCF54/ZNq/J5MkdMLwcBpNAYJ+Q
dw9rhK5WYwl3hmU9r5jNHf+COgsCxDPNKxSu/2MjGoIHQtVgoKIURxSsJXpEtp8kbBwFF8YLeFfu
URXFW7FcW4lzzT6mHJdxTU0zH9RPXZTU7I3gZEOeh5WvZ4ZxIiLcjjKIFOJo4QCt5GplUtACk+L3
e8YJ7YaN3Ann82Y489RLNb2f/D3zpRyFDiEhx+0XYzMSd2+3CaGR/W88KWzl8o69X2y/oNKl2kq5
+BIH4imW+SE8+Xlcnh82R7KBC0IfVzzO656Q5xCEaSp9Y4Rf0mImTMXl/ZtICpJF+2ChTjz2xJA1
ieIz/Pcf+xdgCSilIlY2pF+IbzJLHZ9Blpt9Ks0bU8htUn22JnDq2MrCN8me+jQudU+DkUDiM7yr
4Xox96ElpsaCGF5x93NPb4LmUB49QYUITTH7GUoRwpqsDhT5PBeHtmgyTnR2io8VoeZ77Cvdr6AS
xkFQyN4PviHQA9gbIKdxyfVXDPvcXEouOOQGYuY/3/C2v6RgV40Bz667awXnNa56FdvLsf1uxN9B
d6t3dfhwYqjtRk95+vLDSL75C176wBv1S65lLGjrgX1TqTgIB04DiOxOiAj661z/913zUz1gNS9C
UJ4XXGuA7IqGI9V/ZVznzJCyDKS5TQSPTGE1wy6xXQ0yDBGP+skHqJ9RnFUcc7eo/Dn+FBUr9YGF
Ua0AwsMBfcAN7v1PKCr3C5fbfC29eDPxUoEhDTYZEwbb2BCyljSecG5DCYDcda57DuPeHAnFFZbo
yscwRY8mAk/Kfo3w1n6QET9YyQonKh2vI9NmEf/Hd4OGjqx+DwWTBpaMbAy3sSjnW46PcGWcijlF
zD+z1vnx97jkZfaUmOmlCkaNfwyX5r6qo7EQhZ3xmnqVfnwbYxtI+90V2Wtww3E5a7bUFwnlM7OJ
2pQ1Mxoi5+flF1EztURtNIm58lUo0ktQNKU5oeoTAuXxQYSX1G6XHqCsHCKWqF2lOni74e9Zrh2O
wK7sJJ09ghW+gGhbDlbLC7ye1nUNeFzpXZpldISDL52udxpPGPCiTneEcSkqPhlQduhzQwmURtdB
4PZsiyXqs0C2A0xooYRtoQFsfFbtfp1PVtLCIoPbBLuXga5eu6FEaowECCkI6ebcwky2azHquQ2y
F0Scc4LgT5Y3FyfG9dK4X/F9t4ppi1i/hDkeZI4LpZGrSVgFrTagPg6IEU1HeNbqipGIIZ84QTsZ
XYZo+BtCcbQiu43zzYI+KXL9h3Np3OOHp3cDFlq9TL75ZkAxYd40EkEJZw7QEi9U8pKRwjD0baed
ZepyJ8T58lmDGhgB6HpjX0QCgyaoUx0Euox3T9tYvdrtrQR9WZOmFwkjMMqLYpF9r/4Sl7qg3iBd
5jF9h8fIWfJxr470Z2o/Ov5vEhd8oNtSyS4aN4aBbQCrbg6vC5pNa/lTnW9eM0awKcMYs8RjJX2M
7bnwMwI2LX2VPPegUxxBo8rxT3akTnTt8T1fdbatRZH6VZAFaccYi4NiF+Lzn9itY79wnzn6Gt8F
92ufDsWzNcdALm/4Qmxqkh1uQ33bQ7EqntrvZxYM/NRW22bWwSWu7/0PZKaFPO+Bn9uU53fWTXfx
egEDIm348+Oca+LTPlM5DLgWmIBbsEtMzr2OLifZJe9g+NN/chGAoX4Yqial2WYVDJLjjE+Fd1H5
fpjj87qLaaMrrr393E23K68Px1Jk3TocJH4gt25k1kxw70ghuzjdKaRuLq2yMPv4b/Ds849wfyH3
tJqDKB1bwRuHtmIaWsRe7numCQX37axi2x/CD6RE0GCD98aUAV0heYW5kJlMIKJQNFGFKbmak0LA
WTc0iwbR5maRAuBz9Ckjrs9Tx+PIwQecw2wUPWYUDqflMP1mo4L0D88snBf9nuaIkmmknZ0CxvB1
Swcg5phL1KPOa7hc6prte43R0SwFjurjBFGvgb+gYvJ8raJRJV0uNpYPIGpAIpUJmUdtCUL+HjzZ
yK4Zw87w+pVY2ZVxYEhTFqme1U68dr3H7Wopl4Nfo/YtBkR0s43YuHiLoidzmKoxttOvj6bimxZU
FkOSRdWxR9IWc6mAVtm6DWj+n9zlohrBSYuxRYR3EqugtkGWWehh5hVU/w1YuHqTSpMOAZdEhspr
RrqUl20v1OpjSSOfkMjXCADWM3tXlZqw/5mx1XGwPbHog3oQwtyLPNY6QUYlfkgeFG+ZKgQi2oJy
ujW9mCLWvd8JcBGMlz2As5wX2Rm0NUuiHA6EQIsBmSU7iBLZnU8zwU9d8hWwx009klEct+FylcHo
q5Cf+/s0bb+Lk8G63503+WDf7vpoe9AAw1APGsAKtovNUP/6yPZgXKzw6FCXlnD+LaejQfSzDglG
IPW68DZu1id56GmBKFO9SguUrthR4BqQhTNPYPHARoMMFMo0oIgRZMElFbF61c11nSpAQY2rL/Eg
k1mit/xS63UdQlF6WjxT0cfW83EAy9sX7/uFIZxPmJEyPiKX6T3xIcx9aALEt5K5u7Mk2UHnajYS
lBvosGt/1VZvPNgoMisNl0xwr/RB4rbm0+IbfojbK80uwKNT/StrdIDFlTRkp2x9NL+NPgvyGT0e
LGxHggy0NKKbKGXufnyz3Wp+7duPJV5egXEgguhTCyqjVzITEVk3MkChivHPUlAZsRDqyQLTExQB
faAOzQo4Y5foXOvdQfqVFJGJVpOUdIKwIf85qZSLrWjTa4xKJPMj76RtPbJ39HYKL1Rwt1ZtEnG/
EcrFq8RkqcyKhIAVHQAy3ztHX/ihIDv310wte2ydQk+LV/FrPAlrcLz4ikzhAoBr4Qao7bPLcGHm
8uU28a8VD4tP5NZeLqMGk46Otnsm7s17A2Bdp0NargDzjO1wGYiR9NvxKrrPZUvu3Ec3mcvDpRek
YFRac1f450MQPgQbPRF7rGn/cJz4TItPuJR2SQf/0O+friqSz/DPoiyMrWnz+dW6N4M9HjlqgT+i
ZJM6swJHHmM4t2lUma2VEFHn7LcJJYQCL8FAitBRe9MeMLyd9Jwzydpt86s5jrHR1tOPR7M+pC/+
orPmHo6Hd1fxVY5NznO1K795KzDVyrsSd74OmhEr2kfhxVaNr8EEMRtclJtrGLrUpOdmP/U2FZc0
XkTFoDB1kJplsY9vSjr19/MAs8kdT1nTx6d7WBIoFDeWVXXEqqiZukn+mE0DhcJLsrTwgyyYib+8
yOtmw2XiFxueZnQBlAvT5kvWVFts20dMpHttherwL0eMWH4y4DkpWzEVr6hthHlmIAgWumyCytA5
BfqIioIz7OrSJvsaQ8X+/G4i2kJQpjPxUcud3jzU3L3Q/LvDoVTPcb9WjmD4ZhG2axtOo+bnOk/Y
hpI7l9QJ1ARjPyDZfMb26m0AWOXkseBeXiWPTj+pj6IHA72Aq67vcS7OgYGz7MeRqAlpdHXts6iJ
fMBE/Can4l8CpLMO4ZmCNMBVi9FEOzClxUGBqUDcCA5ft4YwOXzaUXc3qqpjVJqLa/FvaQr+s/Nz
au9xugOxqPDcu79cYnHfIKISd4ai5irLo1XKCDioTjhJo2VxGYi9kGth3RW/VhxGP/OC0tCmMl/W
6ZGL+8ZyCG1yLHM9iVxkwG7SxTOhVgertgiQcKv3kp8kWb1LWJ8u753ajiDzOCmc39Rq7a4z+im7
jLIdW+uoQrEtXjx6Aij1EnkPlMgZj6iyl2xtvhLMCswx0dlVq3TTTEytVSRZgyJzfJ47Gy5gt8pI
gZpuvufwL9f89BSFtCkYKeZmQMCMHQJwgr13dAOwTZefwUipeIcRwbMVHwnjULLNfmatDWqyCP86
eYfm5BNngznzMJ4FgwJM4Zc/iNe84NkeJy2RWHPcIS52Wn9QPo7ImDDkcePjk4zxfgP772aSN2lz
dReOr2a1TULqz3ocJQ5/Pb4gcJeWa6IwI0l/0KtUq1FiNjgWBJRFcJUsLADoW/cACwHc2sOU9keq
GKAChOVAOBRKLTJdtoWtPAIP3yzgoQgVWSqJMGYRMCVlvjgRzw4fgXuNjob38QYUQmK6+TFc8p3G
CsYsbI2U+1XxhZAvR+wAAMD3RSFNF6wg7bGCE0b7LIqp9GLlogkAxYWGM/B8/meQWWJh7rr8ihCq
2KIczZO9WF9Rzdr1JxyZVgk6PJ8uOm1YV7DigB9Ib3qZSytW638UQNnL5joFUvoBPZACeWIN3eSL
XHaqZ+elZV1mp9DjjC8B88LtLBw5uoP7F6apKdOCLdbeM62F0AqLGM7pXGxToarLszoEUmAVdJYq
dNKpUSepi6h8z1DPJ1zZ/s0Ul48N5p2jRw77787Y1UCsHpMm0YbnZILtGFMvi6LlODyTwLWcVZtn
PJBHp7TgIslUMLdGz0mTrC+Pp0gR/J08LCl2LigUgYSs+vHzMLdb69vVa5CsYBkisG61cqm39/md
w+z8hXXaumjW5ShNyD+9pwl1qtO/N7JKXoL/7ml0khbJaz/fu0Wk4OBFrZPDXT+z1kYoUC7+yz1N
78c4/ZYv8k4dQjpq7PchCjAJfzlCEbtIck7eOBaXq9VTU/FQH5yI3Ww/kRiEIoLtjfhYcWdDEXS+
jsYzPBxwejftwcYzsLAsgbZ1LvDnYmte6ttN3ITJlh5Rm0ULg0OdKgnElPMayQ6mh2/PV7sASITz
YTGuxcFKznGd3jLMX8YQZKZ2JcsXWEWFBmHIqwH8+fgYGhSaQn4SNVtg+XNHthrXsVk3Yz51KKMb
VoCHs3c4A8kCC9889tDNkY8Tkwd3CGdYUMsglg31JGMjcslGjTt8YHQ+JftSA/DU8x9rjWERowpE
CrznD7sIlfBUhKkfoJbZ+g8EAIzrckmsAi8aYNl3GONhaKt8KuNK5KQTRHxBGEzR9oDbNh243X3p
r7U1o69JJIGNHTYoYDpjXAbel3jGFGliUwMhvBbiUt9bNPXiw+xMJhtWQqPb9miYa+Gf4YFMihFL
dTb/n93otgmtmvg+u2at1R61VIhd4ILmHpYphxLlVUzkDU/BEcnBXNVvYqSbE2YkfDTVn5HdDxiJ
+8rLib+nnlj7v82V1ByAd2YwYhCEozM+8EaervCfbYDVSUvxjGdTBERamAS5Pap8MP68gIQ6hRFZ
0kqViK9tA6jiUntayNaVqk7iTQhfoPDift35vh9EQgAB/jF2BPbnp5KGAETm8dnnJJlRto8nf2dy
Zd8atc5TvKZRuo7vPXEUY3r9PK+9CQszCSuIfJbS5LhbgRlJYI/u4LG2U6gpUI6Hewu9rwqyLAcJ
xc/lC5XgOxJIha/WamaY+yCmZ/bhjfRe/uODoPVcEsVKdRPMhy7+z9wk8Wk6aLXn3sjT1xKrtBuJ
pFpzTWq6bSrrWGhoB6KhFLbJTB3lIRYCJdgTIoF5LYKTDCEs8UZUqqnMgQvd
`protect end_protected
