��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���O��xa�=S9g�]5��E^�[8�P`tV�yfϹJ��oy̛iJ<Q��{#��w�G���@�IzN�A�ڄ;$���Q_K�[.?��`�Դ�'>�2w�	&�/�/^���6��8����V6��Ü���خ����;[8�Ϥ�-1$D��T�螸��d&�%�0�~}?9��9�V"�x|ͨ��e�I�����>C�TF��DCLg-sJw6�[��]C��%�-��0��~�PO����m���&s�0t�Ć`	޼�����D�]c)�V�hKM6N��9"|��p� ������ϫ��2���U~�ViIչ��R"�^�����ԬV0
��@��h���Y#.�' �E��{�_�7<f��s�d��.��M`T��ޡ�I���R<�o
�B�S����'�#�Rsa01���/���Z?L6��]s�b��EX��� 5�C�56N�ᇡC��Oڜq]�@�-0�g��ӽI��kr�ߩϯf��`'���w0q5'��	��ɏ��E�9�Q�Ļ.hb{K��k��Q/5�`����+�J��� �!~P8"��`|��tiZ�Ż	������ݥ���+��[*��HĦ�@��a��?vӹ�~�7��x�$-��;R����}�>t��`�X$���m�H�9�Tj�ᨥ�^zo+�lC:�h?�TV3���I��T� ��:s��3�A6�3�7Z���6���R����$���ԇ�[�ӭ���~�^��*�d|j�(��sn7����~����x�P�B=Ǩ N6�+a]<=�h�ʬw��29�CDRg��p�+v	z?
ډbю�Q��4�m~�ǚ 9RS�YImN�x5�.�aܟ<��G͢�=����&�opO��<�C�|��b�in��ɀT%v��J����w��/:ճ`����M�ȪdTd��shYY�Mj!O+DF$±��^�V��!Xg��N�L���Y����:��N� �'�5)�/}Gڌw�_�Wu��/§{�w<K�"E"H��ޞשAih�#�	�W��|8Z��igI��i���n�rN�$�{�z�����������ja���K`t����+�ދ��c#����9bt�i��S)�r���;g�O^*���� �`[D)E�4��R>z���VrR&��{��Y~�Z�
��(u�R ����.:y�x$P[�"�!G���pm�ȣ-_F�5hH� �8�'�7�T$�)Hv\�<:a���Þ��Yt��D��)\�q:�=�T��L=lg���df�<�rܹx}�q�c��K���u���йm�8a�yw+c��3�B�;���c�E�c){栓�aR�O;,r9}����fR�lQ�ά�__֕e���W��L 0\���C�^��܇r��`�@���.�;W�1�o��?e� Jr���N�����y_V�$U(�nwc4�E���V��Ah������qpZ�I~��w��� �<�U�W�3J%��Lk�cY/`X�>	���]�O�
X�珛d:aV�~�_ʄǼU�֬�F���Zq���M���wR�����6�@U,u�T3(EA���.n���VOi��h���I�V}c�4�����CM��B�8�KNˁ^�׭oO�2��/��=���3�jBG���������s���<�<��#Ҧ���^�b���f7H;p�E&y�ݣ�����O�I%����n�2�J#�F��jm
�uԽ�:[t�5���uhb�����ցQ�Y{���(�T����%*���Q�zҩ�3Iv�q98a���g�_���O��V	l�O�	�R�BVg�v������'d���'θ��j����<���'=���7���+��V���1Y�۱����h��+��Q?�ӻ�Z~��������r��L)/���pK��;����L���]-�M*e=�[�K�.���I�{�u+�	H(Y�mH��������e�q�W��n�V��!�A68�q��u.�*����<�ʞ���7��Vu�=�~��8R���_x�'�Ê�Ց��,�>���xQ�c����9��Gdh�%��9���t4zq�G���<��}�[�'o���|����v�6g����$��MZ� -i�[`?�^�Y��#�>�Yv�y��8��L���:�@�� �: �98�)�r�f�B}�!΢ͅr���$�_���;(>C��2B�^�����s�v����7��IF�c��olI��̔�� �ș6�	H��^U����ڼ�B��"��f�7�:��<8%�.�/W���D]R�iu��/� �5����ʄ�������a�Ѿ��ON��$	0�`���P�����ţ�$�S�l�ب~�|�|}~�2��V�tՕEg�$4�"��{�rM�m��.א�=���Xt�����$���*�!�2�J^��i�݆�ǯ&q�#�&C=�A�b���_��P�v����s5���co��5 G=f&:��&v���Ɋ@��]��̝�qR�D`@�n�<<�/z�VT��$i5���n����zL��.���k�Fb((Rl�j��9�4��4鹿*$�;�������i)A����ħBi�q����K�Cp���wb��R��>T��I�������=�9
�A��h���k��Z�_�jz�?Jıv��7WYuʷ��"��fMʶ�K��j�*�f��i;J��4����JSFm3R',I���:�7k���x)Lj�D�	���z��2<"e3�W��)乀�ɟ3u;��&�s��{�R���r��4f�"�XHK�n��H��	yS����q��F!c�
Kbt�'��Vi����A��_p�����uZ!}k�dZ�q�[������3x@�T��4B%��+�z6��!�+[U�����g������˺�u���8%��K�� :�l��ߞR̔b���߱G@���}6�Ū����j��KO:�w�������%� ���l�4�SWzq��
v������)��!Sue���4�D*s�M��/���TFα��q��;��1������@��sX���S���$G�� gᢲ��74G��$=���B���H��g>;$6��njÆ�{�yԫ8-��5ݖ��=��S���d�-�Z.�1�뎨2��M�C^#V����
/��(b��r7�Jp6R4aēS�@��q����qƘGr����{CP�w������eF���$�qd��Z�ܡ
�����9A�Bр��?��kh5�*|�g7�u*1+�W� ��Tө�]�72���\�m�s��j�$�\}sE����%��\y�i0܂��x����s��ަ^Jh�1�~X�e�}L0ZU�P軹��ԇ2Q�ĸBf1�f���N�gn�&���ј|�&L,��I.�G�Ɨ�J���9<~6�q��^(�i��9�s=�M!��=�膊�5o��8K���m�?�2�"��Z�mR�rb���>`��|.���H��i��)����m�T�P�+Ar�X:M�� ���ur���9k��+��������]ŀ/�pHiZN��d��h�8���n�4������Ƽ�*�a]�S޽��p��A�C��(X�䫥�i�퇘f��=imNQ�u��*����y��P�����D��'�آa_9`���3�����mCs�����T��pT$db0@Դ<8Q�����X��s��R����-������y��s�B��KP���f��;0g�~�Z�!䚥< �oK?�@���N�BTZ�]E�~o����(:E�/���f{;���UE�`_���;�F�I�
�"�	8{�"H�x�ౣJ�:���9<<"�C`;<���([�Ut쀹��u�&���}�d�-�8�/%�`�_:ֳB���ˢ�]'��x�,3��*p|y�ymx����%�e�0��ny�r�:Ҕo��n���Wqn`}�1����屈
�AcT���x��2Q�#��b@�
��`����/r�^����;�֝�^�ps�žL�u2|wP1z��0�,�/�ZF!S��@0lJB��ƩN�#�fOe]).�v�4�Sǂ)��"����0R�spq7�D�G?8�Y&9��Uf�4B����k�!�e����&�B� ӫ�
X�)����HFGѻ+#�(K�x��]ӿ$+�k��ݐ�IFFcu�`���f�L?����_&�L�;��ڵ8Y�/�j"ej�z�{ɋ�j����2Y���2lS[$$��RЄ���-/m������羓�t���We~�{�����q��.MaG��wc�U,�S_�l^���D��2VMO� �!󂀾j�0QOS/�N�Q�'��<�4���t���ݢ��	G\�K���Np��z8k��anQ~<�W��yA�G�e����x�8��\���?�oNP�>��}�����d��"|�V���9��;{�fݥ�>t/��$��d�<�l�|9f����4;Ud�OGM�_ssJ��6p����.}]�%������3x�U���3�g��_��^M�5x]�RK�p�=�[�^\� ����T���@�g�"wN�m�Z󨫘��q�ka�f䔃����^a֒ͅ�Io�r��)����7(��W�T��@a�(����
u������|��^�t�w���tg�c���%=���{�^�:�G]*6���mBW�P�|����	�j�)l�CF���n����|��=�Oɸ�;�p�.��vҎd��>�uf��ǣ���2c�w��Ws[K��T���Cg�I��HmNզƹ
���zDeަ�>�X��̆T:�F��:U��kn��A"�]}��¦�ᨄ��E�L3�~B����[�r]R�P�C��;bzv-�N��%�sR�DBeH@�4?j�ɏ�Q� x�| � 3��4�
V؂��\�Ȕ�����9TU&yB�S��~��i٫E�=�A�R
_�݀E��%���k@F�O%��ʳCR�]���wu:/Z1�=��as���V����>�T��{��F9<P|�聭�8�-�t� =I�I	��5u��ڄ�/L����;�<��Ic��.�R��7��yD���/h�֌���O�0��u���ӊ9���Lp��kU��m��(������5��+���o�#$|�ԙ*�1�2��"����
0�2�u���EB�p-v/D�H*�h��G���(Cc>��ڜS+�;�?�s�WJ��'�lRZ���+��A:�#f���X�R�A�p���i�*e�p3���/���RB"����B��8�2��`�+�ˏ[��g阶�x�8��l��ܨ�	tIC]��>�/-&����5F�t�s3?(zl�o��X�U�y��قU� ��A����c�0�����K�}7(�ڪ�F67�������&�sV0�A����\��;^hf��Ȳ+/,_PѿG�C�Gm逢~l�3a��-�������K�N��ƻʖΗ�ӿ�2*"-�q�+�QSc�y;�k��������L�u���R���_H�>�^�i����acΥ�AW<�b�Da��;F4B���^��j��5�j�S�OTnd&�`��:��~+#M8�Q`��߂2%��)�����F;���%��xӀ�U.���O�"Cs�m�X��[9���_�yk�?`��%��~����b�:x��6:��|zz\������ځ�a��!#��2��D�pւ�#E#m��a^͂Do�y�^b'	���8�j�a&�:��M�?X�|�{~]�z��8,.��_�<�s�5�����䑲;.��O X�i~��e؏�����F�%��m�,(Vכ����Z�Ǆ�:79Y����&�Z�Qo�o-b� f�W����k@�٘���[{>�gCF�PIǞyBs=��@���5��}K�H��}PsR$���kJ�_d�+�b�`��-�EB �!t�����[Oa��bZ�����]����J&F�Y�nM�^�R}�|�p�9�v]��;H�x���/'{:�ψ'�h��C���^����r<�(d�c�CB��V�`�|6,G��D���ZYq��cH��M%fx�>莄 �rRsD�2W_�u�L���۩�z'��)����\a�ʱ�ɿ��i~Է"�֥"�vIUxs+��B�J����`K%��G0��@+�YJ	&g�\��`D�ȉ��BI5!hb�=�G��U�/��\	t�7Ƹ1��J��n���hd���M~���֫U���IKz F�K���|�%eW�۹nH��`˗Q��+	��du��he�#H��L(UhC��5���