`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11136)
`protect data_block
lDODp3QSFsx1ZKGm7L6GmfZdxJcwH2aqchRtUm9fpD1SPisz2VGZRHPaWJ0yBtuDavPvZSI/9LQw
iJoFD24R6yrHZA0Oz9tug7j6aEHj0NW0IXjRypOB/DPD7iokB7nnh2GaqrbJS2RyGpxxGlMRr1Vd
hoi9EFdf2r9XDD7Ljw5iPFxr8LK2/85cawE8hfdQhWaFQxnv4wEtyAHA8p/jC8OUzqZnwxchFDbK
+6onIMNyiGEUbyl749jKtFkwPtZMFC3Wxnqu3P8dtVBjqwIDgM7wxhce+hhczycUiK9fVv9Wj9cL
1ImjarHTsvWDXFle6K4tFAn8Wl/fPB6WxopUWeYTkyZI5xjmCMsnJmnpN12VFWqE7DOa7STQJerr
Z9Q8FuUJAJWlE3/1Xl+yFsts+vFFEtZ7IAGLfELQjJrkLUDGvINMN/W9VCAXF1w5m+yYsrLsciNs
P9AGiYmb+1rfxiF9e8mi22mxjBPnCDcU/qQWZZyuSdqbuiUp/r7bHZp/MI6QTRp2mg5MEveH/Mke
WCo9tH5ZU8pa/iOtX13S2bE8C8ejdtEwBv8k4tjAxQBq2O83XZFEnKm77xm5L8LXZxNxcCnBB78v
dTlLBC/sjEgPI5+hg7oehGPeUs3FkBFgcDilAhl3d5wFi7que/Q+ozLl930sxPReI2kEiUnvIjw2
MZ6NRqZhK/kp5237CVvc4FhjDc+7ub3z3zlmTJl9xfy0ZMPdh9/ZFGWSlXAuyxw4PCBDKqTSXgeY
vEaOwyUrZKYu7U977ZhLJS0rFEGgcztVt9BPZII4lpLIWhUG9qH0rvR3vYrI/IO+12Tzw1DyMQ+z
BCmG2lPMC19yIqhppT18opAFoHviv75RLMBpFyk0m5c/23VrLg1DT1FA662No2Y0jm9rG/voOFbO
4iASjeYQXEpA3PNGrHMeLW6Xxq2gy1Ch56mwKYX1IQsQE5D3SEqsHp6Xvy9WJdejdIQ9gi78PZJM
ckY8+HS0cn3q4nr0c33fRIKFCA5J+igOoZke4zLY2yjSw7xHlueXYGyu+JN+3Gfgh6937hEzRcbz
oEASQ2W7vpqt0RaKEQtXJZjVK1Mdv2AAYqoBc/kxkS8XmIIiHCya2JIQUZQmgBcfhL2quhd3KpZ1
GS+07r7+q3nqPI3/LNtzZt8aEDnqCzsqeIjQjhSRer0pVZE8L1zGgcSY4QSxlV107nJQJSJcZUVY
iX39nb3A7WM2apQ6vErr+5+h38HwFoq+fvAdjWQcxwCtHpBhaPrSjsUkjnPri5AkhdpoEfLoie3U
Gap7RKT21AngOx6Dz966bHMu3lwvDFSPeiKYX6CjtmxXOZFH6MIq21EVuV8jn7SRI2nE1peTniK/
gS8CMY3QhtoPOJJGJ0YpV/nRkxwKyp/U+bcJx3CqDypf3ztXaocnbGE5u33MTm8ZDjdGpSVw/JD6
IDWKaXdemmyoxN51F+mKKRyiaD+lqxgH+PAFTIiY50QlWpUbC/UiXpjcV+RsXCpqjeysX/UaOSAJ
Hb+OdW1UlrTYtxBJ30Mfl+beDwieg7iQK6Fmo8F3TUwDsmk82s/J0EQ7lEPtztUKSPQEbFJjd2Fz
aJCLqN2Th+KQCdsJzXvc0m/Hmpyok3stRoApxy/ieS9L1iYcMlzOZQ1HiTlAXo8fiPQIoXozNgh2
bR206kYy4V6dCOlaY5uGJ0hjqiGVaBwmhupl1tgTy5ptcx3YetlVM0hk+DD4nZHiL2oqCyoz0aVr
Nga+zU++57ulwW86WQSgM4795qH5StsTI3BmqFHprNg/lN1hzqr5Kj4a2VOwISrxI0jdu/PSIIJN
wAe9Os/aAZXBRhDf6klzs25Gb++OOMHkdwLOwDAr5jOIpr70yfG75Z3X18Im6KjdxZzMpkdUG0/B
59HLRCD6lW8Hi7uo4bILA8Ku2xJZcwXHjwdzbv1L5o6meD6QTzH6sNx/2pXJQobv/ea5V2Ssd5sn
bQDk1iIkfvfS9ykwWTD0nHUY7suk0YmGmLCR94lP1/JmOF5YYR8gP/SCDwCIkaUlDDlghqKMTHUm
VeLwG3SY+yVd3oHwJZd6z9IAGH19GVbD+/8QOjQeXriQtjOU/rw1Sv1pKSuMG/z6UnHoCEtytSDX
cqQ5qJQnhcdlvE7ilLneunge6NWSVGWAKXTtQjTOrv5oWQmExppQCZJspkRhfjJMNKfhtCRw5+ov
xJIL76HbDLeFQlWmtmKZ3fUMoIsbPQxh3RPGokJ/SjmK1tdlHmubJEY+Zp5ZZ60D/2u6CuAanXLD
P+qxlyd4rp0tQ977gXyMm51KLsHgnsQrIX/zc9dCrUKtJKK8Ydewy4+WRhDNuZSEeESPOw5enpuB
0NEU+ICq4Ba+rchzL+ptonUT5r7WEiqtpwMPUHMt/fx2/Mkt7jjhJz3+jwt3gUf4WSAJFKY7luTH
KlQSKHgFF0YgqZFNC3tpVv5zQhGgczyaSr/ttAKbaGQYCoht9UN5/K1yoY/bMU0jEtsqznSI0WMK
DQj9UasuWsFnAzh0a9CvBznZ/uZK3Ck+jmkhGADIjWcVy55afxiTba3lPT83FVq8oZBkNC2qhlAx
nndstABmpfVEc/c27JGt8XqAcm1OU8nwCPeS4rQCJruUiVO34VrfBPo5YUT6UxG2uhSkvJ+9oKbZ
YnWR5TSUq3LtulSCUVW4G5HdRtxCDAhBvWT2SKLXhMq3xTN1vf93ZRupjsM9C+zfRCe3PP1gnMDK
wNHYx2vOfpSF+Dv7r9l/3rpGcqVLERZvFBwFABbJedGxtoA0a0oP5EAb2QnZe9LIsASTlKWx4etj
Av7ashyDmsqv7hvJQ2hI6lorvPwHIycoYlsO7ShdbHPIS8zhExarKbwuN6Ke2gI/SWUlWa2VxsCN
/tZJYXlTjQMdMp6Uu1NEpDeEJDirc+Fl5NJVYLtuiLFjnleR/JA40sHxa709zNZjerxP2NrcTMOq
Mcp5PYWEDWr6lc7fu/x7yFk0MVA8oowANeWr5RX+af/Ad+ha9YTqmHgt3xAqx0GtALQnVqbI9gXr
taSedJ82D1d8/CDZ3gs3IOJLMxcp7045FYsXCHXnCom8PSkrCEdMYIFY4I5B+7bu1PjFBmFK+A/t
lx+yKWHGFCg2BcLfKss0/maN4VenYWVV1g/kj3rfjfZq10hVg2fEnMY3HYWd/Ukibvv3QaTvn0KW
rPPyLNs/p0Zc/2dHZHXQJkhckBPXxeE409YjgurndM5Xh3zZIKXrisfjUMZn47mYK06KKnYUjIzq
pknKYfWw0idW2F08wbptuCd//ZGMUCcgLvDTysP/qw9hoKvgZsioC3aprVAnUZR0cQzSyhgzyCtX
/Mf52BlC+UNyVl0OR9Z+nLoBjzy44cHEiPWykhUrzk1bgpXNS2F572yBHoj5VnbGqdNVqhC3ksiF
oxpGJAvhT7RV1yRatjbBwFHBot3rZOaaWYKS5VfXhVtCmLiXhdteGi2uPzMJGRIuuYfPVZD7nVqT
MGEF9v2as/tjMGE5ssgNlYFGr1zcPDNbiRDtDJmD00hOOaPBISDZKHRZketo7g6ogfCdSIlZMJc2
hQZf4u9S0TmypT6be5bu8PD+a3K5zrrEEie+3WgFXG3USDMStkmJofY7U02+BsOJ+OkzAnNWGNvu
zCfF+XMMTWqlOXa/ZiAaEcfB9uJEPeBaBmjwJlVkEaBQtViOqpTfJW5NVjmgt+IUVNIMKj2bCzwA
1bdB8XLi1xTjZGyxfnbx0U5BrJVslcOtGmSIihBuTJwci2iBcGEO1h+EOZD9SgeFSLbkr2zTjZwO
aNLg0Pz7pKU6AAjszIGSdHGrrb3/0aX+k0YTskly3/ckfPLORTuFptYLj6PXAOaWhMjA20/MhdX5
tP+HiMUSmoIlj5pfszz6e4cAwYjYSACNuRh3CLJa8vxe2gc4eFLviqJu5Uw/jN5/fCJrCJq2FiDe
pWoKSehEqCFgi1ALyQP2Bi1/7KR5zbElTtLwAdDuybSDJVf18Maw4xp+U3k+WR0U/5JC2FQqh2ee
EErTMQherhBsaQeOwD04EXukKv6PFPVbRXpEut262Pzp2A3ZGR9X4mVRixsCTR8xmMi5S3PvQjCM
IV13vOTnKCumeJahco80R1w0lBbeJvmf6ZO1xBCkWI4bwbdO3J3v2napuRMNAlRqorHttBGDCl3D
DInlQv6SVn9e5EaVW+0N32Y4PMkK/1jqOIKClmRXZY9EURCdizFazaDPQ5mj1UeEg6Mt/CjpFAYm
LUSPZQvkhU3g43PO19dEaUJVGmoEGFJgtfqBMdVzBRt+eJGG7YaQkuRDUnkoKjhpb4F25Og/zkQg
COgRREZAjqYVCP/isKrfCNf7Be7FKognPCTJaT1A2HtQlsuyOZJHQ1RY7gSohEgk93WSkflXXUd8
uEkSdi482wh3n9Tc/ulCyDwl0yXqod6PbQ/TI/LLFa8WVhZeoljmRA+XeAZAMZ0j8Rs+92HgUDGM
y0btBRkdhZiV+SruUaJeQbrpl6nnVfC+MmN4M5XgRLYJNZWqyP0w6nHj++fZI0E3KOwLTVbAWTIk
RbGVFWS5/Wp1pFSCmOR2U36JYzSLd/d87DNDxb564QnZpm2K5mqdqDKnSVlnZnYLC8yHvcK5xUtD
olcu5hwFGPDRJnpNpCog168S8s6CJVBF3ZT2FKczc/QwfqnGHyXry2DG6v8oD2p7iMLmABgX8y6d
XAtQduQGfGwnXY285PB/KK+EU5euj0sRAzxnVefSbPOwwBslT1sdUBxQSROuU6Qqj0zXReQ4/oUn
nOokKNRYqoPiKi9MzX8a8itcNMoPJdlyFriluHHHTLdU6x5Rreb2YIe40QeqWWnIdA036aW63uUJ
ckOQQ8IJxY68tnHU3sESEM8GbI/rYpURAZXYLclHfgqf9pk5WWIgbI81MHiUOpeOOqUdxkW86G4/
iVE5GlLcb1sxDY3jU06hV1EuIaOnfNZiG/gCUNnRWbdte0BEPmNzbzwZMjC/lvJIDCn4/zVZIsk/
TOFS2XwxfGl0ewQ4UQV/021ryGFPo7YCVGOV4BnMUhlJY+XHoWValUyF4fIRVG68IPTpoTtsO4kG
imz0k5oWMlgOw+S0BbnM3MAKQxamfqgVypKByKiN9PCc1c8za/+odKGC3POy+QIc2Vwqzh77dtiL
pAA1mwLMxHwB7KHIO75588JPF/3XRBWiuBa9whxnutIncnny8SuWY70ciIB9EOkzthaB1itpJgoG
YvnjLfXDOpHcoYRHoj595Afg705DYOMIyBZwT/mGvRO7MLFmIwANWD8IAe68TOo5+qbBK9vxVzU0
3dZqyVQ02L5xLLKOT6MRlhfhnTwzA/UwRetKbN+6Y10N46ZISuyXTwngIgLbGOyC9Ws0XYZ+f/PA
11ENJb8/5/9qkcZLjuKDTLypj0MTiPr5MjyPkecotaTVS7CWxvMmCXDvXcv5i7/4NBhilz22gLdL
vJDj2WB3mruhNohj2AmcD1oAIegmaddgWb75W6WC2luw0DYh0uOc1e4BhhyKzzO3C0TGqUVuadtQ
xQn4iAid5F4Iit4V+Ym96bVE3jTjT8y4sFosttZKZq5PBY1LY/bOytIBWEiaBFrJE8w2cU4DeDqF
xLKQGYi2WtR7vU3YBamgZZnzY1K2g65ZOwUgnsvMdCMm6q5bvBE4MT4Z+1wzN0FhDK6VdrPgRo4+
8khW36dMSUK2GX33LXRflcXMnJPoY6KqMkAlyD9PF1beqlPlvZ1w71NenP7b4zntDWakasTWNOyG
wV90GV8DEmvVosE3tpthkejmE3myKYgCWEBqd6Pwy3ZqHb+hDtgdsFIHffvS+X7/cBLaGs42mBml
6K/n1pPWhkitqD6ENyRDVbw5Dg00aqBgqhlvZ9ZBYkl2WHzlDQfnEwbyaRKBm0Gjk9Ovr87w2jTM
iyIQJRJ+y1eiNU7ikaFTOjmghA/o9rho/0tWOr1KtR9E+R1BcW7HFYOeYluqm1KZH9V0p4MdClXB
KG3akFagL5NUbx4ZOY3QdAAC4uVvSuy7d4PTqQG+qDGBf0xWjLMBpXF99+XRfxOQHUJdYu1Kz5yH
5G1qgEtx/UKWFQ9XIYUOiVt5P6MHAkXwbUkRyODhqLf/5OQBEMOoC+oq+hyNtPi24Y0I75SE3dBE
pU/iLlBSgtULI7/09VngKSVGUbQLO3HAzUSVcQ2Qy44AEtEXZCsTv3lcBttJbU9JGpdDJc3iFOq0
alKlpagZMPU4BnEVtiVGNLyjbmj3A7ILXRFRKt/FnNHWx+YBiYmauUMFDrKFOOub3ZGBH8vMYHUn
qI8F06s/G6ni18+QOmJv9F9jSkk1bcrVi8GG3BX4XeQXZZvYPnFpatTBNCOOhKNfHhBiHss6zx7J
TKsNL0L41bjFC5u9Dz0Vd8/JOfAKBCLBkLueA9jjMrnXt6rRDM8cVUUNQGeSXuWRMb5YSjK+VXw3
I1qrma//MpJKVTLxT6VzMJf3RC5j+VakkbEYTPLmqJqiiTRxOwaek0orHW7TsjotSQsIdjNq17Ny
gGg2ikkDEqwqjj448vrLnOSvi7iw7+4W2Jgr0WIwVqhnOhL4//huwwm561DzHWnl8Lhibw5VlR2x
bZlwM0Zy8oyTlkYe4m9BpQb7EzJejFJfgePWVA4g3Nyh9nEKK396+MqmiaxyFLX/jRNjQ9tGvFKr
KGtVLXkcxj/QLaZg2shFgeswSNElTlFf0iwMutZIwJmdT7ROetLRVuPCXnq3+mOeOIIEAwBlPpbu
rP3LxKZ+TYtASbqJQUFftnqdKFWjIWLTGGcxlec9qY1fs5BhbBGSAe+1vgC3yIuVm4PHRYEQY20J
9LLpIlzBDhm3IhUChsyQK+c9qKS8pcClzYlnZcK7zDuIEOO68BceyaG1zNw0DjvePHI3B67jQP35
/e9vaBU6tbMdjNLUvZ6GaaszkY3W6+hC81VVe3brPFmW/rIzHj1N54SS2f3ta6pL0+25aQS4y/TH
KKos3pCCj5wLTruW5J6Z+ntekcvN5vPcmwjWJRiUfge/8Sii1WnRC5d4upjh9bEv0Lcb1W90PaI4
qjzE8Tt3r5mfW4Bg7KySV0ujNn5DJNdDBA2EfQyOFuQm4xZaCS8Ew6S42FeS0Q79DnDU7RTMrzkk
elljQORhf3QpjyvkZSL563HHat079iQLdmt1Pig3h/U/DHjibkoix6hstSC7Bp4yoe3U51zgYed1
VjPN6hlbQ2segs8dkkzKsjM5pB/ehUi8m24CFcbcuAww+hzxdUaYTPd5Cn3egEWLSOvy5ih7FhKx
vfoTDjH8sBaZNbY6PPlqyR3WS307CNyuGhpJvT2ruQrt72EZbdCVPId7IX4x7irR78EqvUf/sMVg
01Io1eSZCUjDgRpKwFOkwO2NrjLYT2nmg2DAFmGRIr9ZINV6rHvrKBUh7MdHWdyjlUy2ApfbNrB3
fjfProhKKrY7hlHdRvc38vJbeM2GRVbJTFTNMaBRPVUd89Qgn1LtQPZ4sLbgiEwPoYYbK8tVVQZo
MIKgYhaXT/2MUkFmfe5hPiXU9QKHTbaRtrA7SftckBeSIx/FABZ8sHlKFc7CC/E1rsErOC5ct9Ld
oqc9MBJ6/TD8t1GxInNRFoWLp901ur0hugdN1J6VaTQ4seLyeLZ07zA0S6ZdrERNbXLQFSodSgPu
c0vfTe3NMxM3sCusenDEqzOHFQpyki1y5lN9RAGyO5Go3VqhL7bxPLn7T5N5RaMe5Gq/8qyp5Rpo
bxAvDoFlBfEnab/tHe+xmHDP70eZg7bhwN9eP1Y8gZet1ZSkp8d4j13u+/HnuTv5CBWyM/L7lQbE
bA4fOeLPzNYfalyUQ8Q+ejdYl+BzVtncxys2A/35R3RkL5ndL4tJ71u0Nro20AFyIAU3d58r5zAE
JLOWyqFzmsaWYQHWmwHwXzG943TvhSeo/pja6dz28BsoVSKIq6RpgeFn7eP1IdDE6rkX/ZR1nK6l
QZrtVJIvRcilI96r+PpVyvBVYRIj5UYBdRyhSyx7CyZPUGA+EfAqAYtxWj59KYJp98pIlFEgzOyn
cbYEuSSwUJfrPtVYUkgmj3AproNAxxNLHFtua/SqA1N08KmKvIXEkLKY2A4VrI/3sXfNkup0Jf6L
+NAgUVXNRzCh7PvxvjE56FCYIgUsOHfk3UWe6UH3GFbkFJcRY7R/u70MMc9pz6pc1SUdkUm7/pIR
adQs0eedwXK1xn0jx9BOcqAz2Ml82mHjGTK6LpL0KN7JXzWU8SXAhXfNg7GYCIO17/oYbyPKE+zT
V6ikAjIqjMfpS12VC0G36qyIMvY9Ysa8AQPUPRe49U8Lo3YpqVKYZo+3ubFIApUsMZbnmNj95jwM
YGpHHwB2rSV/h/x8S1mDE5PeNFBiAbeBawFWZ28oUrAfS0KibYCrz0crHkpUeVGaVSQ+ekmC9JVc
9lSUKI7DxjgEz5wt3xMPfsSE0/PzNaeoB2y+oNiZWSZ09r91HNdddWVXQdTN3cFG9ulOQ2y9+8qu
tRDl7cYRx28uLLXdDATGMjXOu4RxG3v49awyS6MaLwcIfpPKYl/8IfEWJwf48kyCeyEifOufmXA3
vGx8kCHcZReK01NfiBKFWax+HyukUXsLnIzK2eLaeL764jPuUoIJ3CJO1ylO6rMlMSN2ClKTtyTD
fRk4JH4/V9uYnoPMHLXhUgMlkVWtsGmEvsPp6ef10W6bN+DHPhYt+H1I6bAI711MZxTQLwTguzDO
r6Hsl+XxLcM8XsWO5dU1xA6jFYtO9iumvkTmPFXrTmKrWvdHCWK7l8Ws3vGR4abobdR630fnU5WO
D2qsgfPqEWqcY6SJjCK7Ex5gzG3qb2CqW/uddKQU/PBd9gB1X6YInsarsSYqG30Kt3+dleIfCJsG
Ix0d/a84ZMHIj+2gxSixx8S5CWTmJ6uKs18uyhxtYJc9kUYwHPZpvxXOJ7MNqMaUx0JTu5ejFUl9
uqJCXALaC9WMDfplSQaJUtwZ8Sq80e6FpL+qT8tR/eJgANOmmxMaqtEMG+x1Y/X594lJsD61oDxI
97+7yaKTihEKcGhMY/XbhSv1ZQfYZHMIbK0utYL+xSB/GKmIYMwMmVRD1gNrl7KWJEKlRF+s/w4/
TYjGRBRJYZYZh9ViL7FTeiuNb5UJmWE5spyiOxhVsDtP2Np7v0BaJSyB9gJ2Did3tdUMurR4WlQ7
QJX8NZSqone5rcuZ/+05Ands3MdSEtdN4Lzg9mNAkvny7nidccH3WcHMSvRpHU3JGgWy0u0lOc0G
aIKslGmgcWaM1lMDbCcfzimGayPkO08OBXw2XFt8qhKo0HyR2vpD28H4HrJcQ34Mvfd0bqzV2vfa
s94MHyD9knCwrtqdW9VHffi4znnDqTTUS9v84RZAknbl1rVKHulWxs8YwwaqQtbqQ/vxYlJwkjRS
oVtwV99Bh/tMr5Uzpq77M6RUkWT8Udebz18wy2miJ6CRODraA3d1CfwGJO0Qw9wG7lDysqN/fFIz
fPUDJMW6Cazl9RFLaH0SawqH2+9BZcpaPrpHBrdeChPA6XENY9iStBAUNTFH6cC/fUSvJienyCoK
Ku5rbHGsRtMiLR9eL9CKQRGQpyqOIrvzkqLIFKllwpbe6OpkfiwvtYtm39X6XGoetTkkjO8nFJcU
K2rEw18yRPkfTeRlIpGUAi/zON7I9o9vQxz1n0dyKre017mrVqdxMQWlLhIVuAp5LamEG5+wp/C/
4l6WlByDG9E5tiXIq2qEF+mgsCyRdOA/ndmdnEjMAXohpIdYBG++26jv3sB2XFgPuyf3gXBRJFTs
jZjblJm0tXyzuKJZZPGkII29Axr6xoM+oVBXgI3LBrtq877BoSga8zd5Fo1HZvokPdCewH+L5oVE
mx5HW4eOEgfWqiZXN01WUBAxRuL+IVlEtkZw95TcutAPmgxS8U3lnQS+B/TMoZZs/9IbY3m4fsmQ
5X1VgGeamgDPwr7orxY4BfDrUcLMjIXwvZFQyIDkKXw4lTOP8qkrZEwpoTrHMvbcSi+F0DJ0K+Gi
9ptAI5EMu3kZcYa5T5/YufJqvlxCAbeFV+wvEgETtay26K7+cC0k816pLwPzTLQPnPCNidN5kAvL
hlm/AId+/nNu2vLjHzeL0gabLjMrUBEHP3DtuaBP6ckxw4RxycQ32NpL1m/UMeYiBvt7nfCf0PJQ
h8XJZJavRNZ1Qgl2iRUonGxhlhHG/XYFQHlux6ntlPp86qcjGR8p6oQKf1b+6gEg4gLlyO8pKgJS
N1vriseckPpP9a79WHxQ1H+boe4F2KbRp3yLoz+MTyH2uvTwVx+AACUg5TaCC0yEXaFdqu4jpq8G
pKkfZpwz4QfTWR+8pKAm413RYU1BCXajvYRehFpy4DaZJo3FbEAL6rrHki6+HeXh+VCEedoFVjiB
AiYvhFTrvjRuq81ROImL4y+TwAbEeFB2EP/Th6bFE+av31tX8Osyb/8wcHjZp0lfFR4J/C1Y5/vI
I0T7ViSIsr0YLxavEnAkH6EEIJrjD6XqZ7uea3RopuGITk8BmmlH31oZousosqlNzf10bbshedYn
bMHymRyC/BFQmTbzEM7mSc0hA+FU/+uN56UsCR8EgB+2hOozfFzGG2/00gskp0Rmri40f4SWRO7X
BJYPCER8UgTNfd5bxBNLlo5k3S5YCPXQHGVVfug1sOmsnK2laEcSmw3Yw/BCOpwSiBA0n8hY7gHo
wl8jImTOxAWiX9QeyRuhHxMgTKx8TpMdoLy0Mz5FU4OtwJzk7dRdRML0VZUGipkQptcpBNEPesww
teAYBVZONCHOL1ZVTLb9j1rGKfwDEK48Sy3f2b7yw1NS8CwEK7muzDJQ6Z+34ZPAKnkGQ+xLShCp
MswmVE+/OFvyGdTtmKOYxDcNaHOLsuio0SQkLJYxqh71DuIA83+342XU8YQnkXsiC9jZ1QjjdkZD
S0o0z5PAzWyWGu5As1T2HOnOz0/O1jzSmLGxwqsNJyC+cr19nfA4PwisahIICLVoIKtyAzhXU3+Y
JkwgMdcdt8WjJOXubhAWKp7m1OFTE0IC8RN91DR4Sx+n/E9F51i8j5OZ3SSdc6Hxj9iSFtQWzgLO
VuXr+nJptGrSTysIrDa/QKi4EMJ1o8Z+ki2T9z5Uol8DgxKMWx4YdGOttkVXsRnXx9LANE5WYkPU
l8ZEjsY7ygwDYlrlkLtaViKJH8McazLVFgpOVGzy+TZ/dR7kDMe6ZjzS6xZSdKnZEubiANafqRiF
lF7hgDn4sXe0p19guSNAsVzjtM9kV04IHtarCGtW84aVxwnGZEphcdE5iVngMxQlMKf7eVOgejil
RG9gYERZ5yMsr5nh7QJLAfsfiWNXN7yexFoafwqVdWihEfC2efjrUbdmNMY5UQp6cks5YzNHw0b2
9YykoPx7jZVJ883Mz1Jh2gzEoMDdPStHKh06BwZfdXntHpX8kSExb/eghr47snajYPVBfxFcuRR3
xXhG3dqxkormvDHV7Jd7vplQA9NZtl9TtOr3qDcB+UuDwiVggv9NBJCAhSMhlbPuOEHuBBeLyilt
u/F6+6TqrWAVgY0UocgYNeHjqMI0sCrn/TAO8zMxG599VGoXpUzsrnlCZlYsReHvZX7G//KLX1m1
LBR/6NEJ0Ffn4i8y9PuXsi/xj2rhR40SPcUXTQktrpNGwFOdWkg1yRiLxGZFaeE6z+/subaEzsDu
7eLNhlqGrrY0QmsML0NYZXg9gybAm0l6aTUZsX7PEVCzH7z4fScidgQAQIGJt9uwuNtHTNIMLu/l
INzk6NnYRbxYHrjGQnT9x8H/4yyIsMzM6H9g/amNm8g4ZjWyr30h4+2B7embsyVeb43rD0P/Wukm
C5/kl843MX+pi8YkN7YG0o26R1jK19VnmwKXEalqqWh7wRBmXxVWOGyp8D20lIQ1TV2itYkrmLoH
GcWG/fBkSwLut2jKrtDBj7uDK09UsQl/MdTKKUdiJkhamvmjt2qsZE3iYTcuO8eReGAWTUFwHyUC
rMBWtrv65ivL0zy0UArSxBxNDYC+A2abo2L80PgxIazC+qoylGM9YjDbeISv0SGxzQi0fsaqc7gd
rACotC9VQYecB5RshdLd4ePBRPVQZiLEiGfmBfarFrM4yqVo8jvYqvqIoxu8ZuabrG6GJI14iJ8l
+AjwNC7WsqEdP7n47FjK3tXBIEtZi+9U18qAJuduWone90B7kgvMHMUIu1j6JLg4bFbryWRKmLj8
cab3wLZrWpyaFl2iRc7Lw2/wy+DnN8boDkZWkOymyjvNWJcFFCQQI6B/QZS40wfJwdAWdWLdcxq1
XiB/lQlbD7TyMGCDE4o032EADzOO1gYJGgqm6OmOP1DWW0fl24gYR9XcMmX6Up943DVG9vS/SVlM
q8QyIu+gUWiQD1giUL9310tTGzPuzUzKyFnZQup76DS3YAI0hpPXb6E/kmwUCJVbdVgMK80tJlAv
RXOq/SmOi0NShFrq/uSx7S3KqkQ1/Bb1ArOZl5yr9rhJ+AGPdtwqiAXDZ5oNRvJrQvmbiA5T0lvW
vOBQrREdrbX/zx6QQTMy9vwZE18+zHvqnktkefh8lc2a++CrpQJ86IKEhq06T6kFcsij179lpuYa
Jrq3QEhwZfaNSmlVzU8RYpH3nf2DWWoOu94Abg1I+mLDER5hu3IWKcnoGQpdxCrslG6OdtSgkXPr
RLAq9EWClrGaMNnvrl21uAmpKSm/n74fg/25nSbDgcPHG2nTaMme0ruAlOubcgWag+YR8IQNGi3+
es7o9cn5c6o4Ji1x//Vo9R4ubVvAFSRrw2WPAkyWQoG0jmlokS6d/6pHQ8MwS6wsrsOuCroeoTm2
h+MqsNgIbOaCRmYILoIRuKqB/RC7Bf/HaYxr8r6kx08qXZABLgMmbVRmiC888n9vQkzVD9SEwZOt
xWquPFHzC52hdHFet9WQTNayBsUrBqyph5qnXWJjFNKsDbrvqUMW2pCqJc6ow4yzBVKxPBEUt//p
i2CaI5DRu0bExYw7GEWNyI1689LZfggxwMpD2gIKHNoTBfH8TINryLVn/ts/oKEqA+2Y9yCoZVSL
jYwsTcBBBtUYWqtyfXM6fe7AHakVrzNAP6nQ/rf5GfINVkcF4chlKRR+mT7Czzms59tvqkWfdivM
4gy4/1ZP5RhlFm1gZmdT2K4AkwMYwVnR6fuugcZVyvxC6f0WAPUFV+bCAn4JCM0A/n3JVJSpFpZq
Yts9HiF7bdtPituU1VcmIsOEVFUj+uUIZ54kU2shGcBEhQjVHL0GJ4D/+HqOPL/ROQu8t/ykytos
c7AvOQMy/iUrAuF2KAIVVIuvASxVn3Ci8POttBy+N5Ae66mtHi6IKzzSMDGnIzJ5ROA6Ro3Cge41
KIRQm/A7oRfcber7hFbqOngai20H1LMeJDueuatlBshuP7hPwhIz2afqMEXfNDtjudORS6A7tIf5
GkU7ToJqGA+uylJEflsqeLIPZKhmI1C9mXIKcK13zzH2X/hc/9AaNuJLeouAbAcB+5nj6zwnGASq
OpcQ3iq9tIItULU7pwNYBYQ4RoCrcrbbC/hK7ofmVyB3zKezpJ9DqbY06enquHoJSMFqTiMSJ4Zv
cBLt0DMYb+ePXu54840JTfdyfMCiHcvIzYLuteFB2wqj4nITule0ZcWmqfKwCRhgs4RS3ZtO/L6F
keJPXPrjCv3BddzO9aupU+Xxb+py5NIREvUvikcEdk5sFfA/nNxycqrXXofQR5zep/FHvMCfejhU
Xaal5ChBwO5wFdsyqQZVQF/hot0nk5we7RS/ZRX+mhOiunrTIJkB1n/PK/jRWtYh6zUSuUoHPKTW
zUHa8JjTvpaRoVJzvXUvsQwlpJpd5UTXwXgRv9cnDG7KMajcThZegZjnzpqJEGNeLxLE9pjE0Zil
8AYgQGt43E+vuJvgQ9otPQ6BchwrlvjcLPcbYM6dQPVAo4JEyMfg9wAZoCHqdAudgBijJ6XuNKLv
1WwgYpQEkKLVWnodJ7eEc4gAG6mF9UyZKh8HiAYjBmffGRWVV9e61G6zYytVYu0i+yrgeWmZny1V
w9vq3p3Tyv93vR3QiO7frLrfeeLs6u2FaRbN3g+LASGTAElxjG3gGLxpsociywGghRLvgw55lIml
NFow5ulo3ei5Jce0WDdbK+5jcrkmEyaEHqjyYq0hG7kR4gE3mEzFFKu7Bz1hvFA7eXeFYGfRznl1
RYI9JrGSO+OVaxT1NIcslBpPtHMjFVdmHU7rkKXCpf7a/b+P3wRhjoMQoGymtmfVG1ytX0Uz2D8G
Avtc80152enjeY0YJd+4OEu9epa3rePHJzcPEq5V33DiLo2PAhQ1AW6xKtZh0JDaUIZPO6Ybv01F
hZC5x2NA9vsvzT3/zVFCjMCYD33RkDgjJ+FKhn7u3KjZJrPrgC7vS+9N9goZfW/LXs7t2mvBWG6D
2PadtrGH4Lukgj0rv4lf55ZOYp55xje5hJLh9N6jij2hst5HCeF3sbv0KEiw2pJkO8CL2b88kMNc
hsgoMxX6zP3/aV4AjOArl7jZuwUmrhAyiZC7HIMQftuwEH9e0fPQpq0ydMU1wvvoagkVDwVChPLH
bTRIX+zFJXg/vGnkQvAeiJWyuaF/iIMr7+siVVXajbpXraKITyQznonDSD10NZhCWRObxRF0yl7b
IhcdFQbLsTCpWOMmje5rkAaFQ0l28IJVkmT4VAB2iVOyTsozbUu3lTe01MQedNdLaDaMy143OS7f
8BVZS93ZAITTVjfp9j51LPB4c80xCnQZg9pcobWbrrlhmoLUgkFKMb2SjKitXOp6KbBTpbnBUAKd
lEc0Mr4sy0mzzw8lgx2wqI/KbiWP
`protect end_protected
