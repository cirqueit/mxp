XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���0��'F.��͈���x�K�(z�� 4=�(�����] ��"�����,C�t�I!TW�K$웟�!�c{�T�j�WS���w��BCQ%b
�K׵�.���w��;��M\0�!
����^�Z�)�c��D����ƕ�΁j��,d����z��-�-��B��ӽ�d���UվD��>��nZ�^C��U�-t]I�<�������{9"O����H�ϭ�u!&���NgoO��w�!J�0�������������Ҏ4a�W՜�
���_���KZ/�y��ٱey^��=s`G��)U�1!k�)�z-	Ah��e�
����[��ʢ��!:^�@���l>y=�3���Z-PX��K{�,����y녦�'B�2l�2����LcWMl��d����2H����O��G8b��5������?�J�"U%ڈu9�����K ��s�nL�脎��~!�e�`�˖�@Ѕ͹���GK5@>�ā�^^^��sY[x;3�X]�΅��M�Q����,��YD�pY���D�I����b�$~�;H'��l7lt<��~�{lG�b����u�?�G�:�fZ
z[�@0�s��@^_a�3Sp C����F��m�4f&���ӹ�;����F�L�Bd�&�+�Ǿ�f�o�>��6j�o���*�I�٬t$������/���tBD�V��DU4�.0��)���7�D^�(wM�a'�k��j��Ȝ�3�f�ķA��N���x��vA�2?��7ٰ�+Kx��XlxVHYEB     389     180�ߣ��+���m�F}"�QqJ���H���+tfB2E�>�:���{.�� ��l�pﵧ�w��P��1�Bo`�{Ï�'Q��8l!�;���"/(_��&��?2�M�pƷp�Gɒ_�yc�.������3�
2�?�ׄ�GH���1辅ˬ��+?��%H��e�meR$�)7��=-t"1�+�b�&�H�Vq�=� p��O7]���.Q�kJ�Ӧ,�`;۝�\�E��9�"c�}yj�T�\�;�i�������;<چ�����9�KC���eF:�OA-�M��\�\�Q3�%�_�_p�G��p�̲�ܩ��6vO�H0_�@�G��4�Ƀ�=�-|W1zd�^���t���8�9���|�g�� ឨ��"