`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69072)
`protect data_block
S8csX2XLpmWo/I5CFMW6jyQ0BggMGM8R+nUZJPWYe8fnn1Unu7xaEL3lqoWMku/cSGHgCuP1QpAE
6qBNWoon5LJKlaiFHtlA8UY13I9yXnYoXxVzfJpaVfudYCeWk+OdneHp4HszMDTAO6IHb7jxPjq4
xWWZY205F2Tc9VrJ7OX02oVAT43jVDuE/LcctRZKMl5yTJQUgkyqzHSX7maPlHi4NzeRp+TawoCx
TD2Yfh6mnArWZae0n9cMweSNsGgqL1ANk2cEaqP28hQtq5leAiR7dgiKgS583UyDCYYEo8IYf7FR
Zr5Z8IB8qblxwNw69Z2DP2cqxevslR45qn1sr4nH6vy65waIJMBrm31gSf4UZQJFkiT/Wrhapgq3
3QYQ9HSRms9RKaarzcoQSTwg9SvhOTrNSYH9gO/fQNiqy9AH77Bbr5IRRoTyGBYhV60TYqk3xZ+j
C7uCc0y8eMUDeDhowYEIuN9VL38+/HvnzEG6iCjL/Nku8bNMrEOPo7iJjXk3xg6YAbZywvkAIVZj
+K6f/ki2MRQWTdu9OuKXa/qHhU4aiBbiOvfLNONkqO6a00t1Q+u5EiLCfUvy6pzK9d8z0+UgnPYV
zt/hVE/pMNQzxU0y6hm+7h/H3Z4rybTuzxq1YJGSgQ83Vj6TdzCVzeKZXciVpOCvelLRe+lUkDEW
363vD1LuIsB8JeENRz3w17BMUtQ9Yde4O9jYx+uESP0gnAYeDKu+Hc/2QQNyOqIEzvbiombVUoi2
jeW7L2IMZ/yvHgcvU/pJfJeqeWvGNDtxZMP1ECE8rblodtUMrlQiD9RTuoBS/4rt8NNoSR8gbVka
D1kgh8pDfl8TIZEgw+7P/ezbQPU/OEONBWkgvGugjCslj8s/idtXNE4ZpZXt6S7WXzVeWaHV4fqa
RAmZ7P2DYXvSR8V0i5Q7GRi9Zz7z+VRTgMe1e1OTHfvHmzBvFKUuzY4A1x8jdx5inLba/6Zx4Zfd
UtMhDlvprcYrK7HstFGERc6nO2HmwAY+dbyHGa1BY4hIQ2uebDeZcdCFws7BLScibrYqw6okxPcO
dO0GMUuPEuetG8EexK7kriIWDchBinqZz800pU+2xRPb8UEalSpxQnjv5U2Yzb4teLJJ6k7L51we
6SBRQZwEMsO9FpfJP9dqOvf6odsjSfY1L1bv8uyh3i3NKwRvF+qhwZZumTPURAJgyGvKraaM0KnN
btJ3C9mtvtpEZ4GNfGZ7m7xCVZkGQatibKYfffnySm0+MHDfNWnMdi33DiTBo7i9YXrrwBjY0x8I
Y/p9xEyZlB748ibB1FsINrGGi0OlLmVIM7dlEmeJteSCUG7IrPaRe6n5WR8OxPgdf+e5pbB+zzQW
qnYDNRqP9inphO/9qY6C11dC3P3cuLdq59LYTCV/d1vhwjTp57Z6JgA/A6jZQ17OLGLmq4KWQpqP
AJeGrLrd2r5ZbeUvYNTYwwNBSpA1nrx9+YtpMxS7PlR5OqlWI+70J0Rioh3pMN5umBPI/8NwpUBT
P7I3OBCwrQ2GQNwDqhp5evfAu93qj7cM3ejmTkQ3Di+lMhf5XvqilWyD6Fcp8Hy7q4OlbuZGtvbs
xJ2PdXB9+stgPOHFvWFgFHhiGA4N0n+gnJrMhtTTJOGAR1tkk6R+grJWr9Uhhaw5fQFxJBjc6D+h
S2V4rCDduj12anwbV/8tDIqMmJtl5ms/aoW+c3Y71VN5pGF8HrSoJnwZHAnJSBMXGd0j7qHe6FK7
jKXmf+sWhc9mYTAdXhTNqNOx9VTJd9ilAW13KGSEYi88o03zJMIOLajUD+e26ILOQAEsvVJcue/A
M0jCXOxKNTrkLMcClQ8twBJOo45Mz0nuNHzP6NH4UwaVdqcwGZNanfPlE4HrTnQEmqmngSkwt6/q
YI4cVnfuAZViTU9xvdjvs/E6PNN7S4UQkiGDlHlKTeVnZU8/gTh8avWvnVQH+YlXh7Nr/ZWqCiQt
sO2KPoLBPSCCHfRz3p6B/RDATKcHnWhOZuvdyEguG1rVzVh0WkXIBKbzcTPKQVf/eVYSKrjGA0wQ
wQfA3PqZYzgLHV2Wn/0vR3vA1d0RMa+eKevoHdC/0noWzHfezZ+yLIrbJ7jPc7yS4x6dQotMhIgh
PfX+H5QkN9BnQB88VmiVpNZugErvt5nq2SIbf/++9C4jf4Ojs1ZkcAvmwku3KMs73gJEhSFxWKzG
OKYFVf2U1622uHPb98at1+JMYf7Lfr7hBwmqu7oUVmI/KX6FXkfWIKCsal8yKH2u97kDPtREoh6N
d49qBQ/PEcnGwrefjDeZir++w71hEFSis+sHfdqoyl+IibeJeYhx5NvzLXkXsUi198FJxblTXpIu
tRfFqcsH3QuX+SucUPC0zTjHIE5NjRcYxKffLVi+eXuXjg+mj/QuSrLRZa1Uih5kZqjNj4vMeHYn
yzdds40OTDlrxDi0hs3j0YIGBAKHl9utuiTNzyzyvOkQSqV3VgediTEkM7+GtOBWtvDa/RCV1UKI
sMUf5tp3103dd6iwGEuOswFBS0DRum8B5D/dN0l10fuKKtOFLc+tDXR4K7NWCteon74iWwqpwPTU
rLEaSmT9rvUD+Mtjr5vXQwx0EyVGsFFHrRpU3QdOwpTObBxhtl/BZx+irm5S8mnQR+7D7/pUKlL7
ARDZA8feQpzIhQiJOn7JJgarBDNUeY7BIbHguU8QatT5QGo5gtvfSNm87v07ry7XAYDfat1pqgkr
xurDMGQ8Bw4iG6gr9uDGK5GvKY7wfRk0aMRknN+MNy7Kkms1RBMVIChFk1o+/Hw+n+Kf3qH+KnZJ
OlYzLxKRIWlsk1dCrbm1fH2uueZKyhXAjWv13CrBWcqlpGlrr3KYSUsDXVueYN42LYo7z0hmWUBr
AyR1MmDkoP/AQu+Uh5ECR3yIo/3S9Twh1sYgl44HNjnqDkbK6ZdeXkotM4vJ4JPB8Zo10C3AlSpv
EvztYjgBt0yBTf5XCqN0vxCxlfjYhaZGGSGeT0GfhYGCiADRqCRjjDYbVndueH8rYwfQJV3yE5u7
AKOBacYFNKsSyCqzvPftZmRXdPsXswkUg5+IqQh6kyZVtOHcg17gglDA8+DMTQ3MDC8Mx+9kF4/H
3de8Rzur4wlIvEW7KX1SG8l1nBThCvsK8hZJXXXGUlY9iqbuah+ACaPLJ+C0pJh1d/52uXa7ZmJD
k7HY2hhv39QjELAwDDPS3rJNaY+kV5HytQVRkgflvEPCD6lw6HiVehiKC4dS3ewwyYeP6QWuUZCY
70hojirLTxrNs8851uqjmVfPtQxEOED2IegrFxdX9yvnL1y3C+PN4Dyzv4z0eXkBUf9W/XFJ8kSS
2j4Is1FahyNe6IqGZQo4iaIZn6CLDkcfAsRJLCH7KPcyP0dfrvOCVRbR/xBqdHl7aa90WKdWTpR1
RxuecGbf4Pua1uyxZvWMptPqgl5SJa4BwbzE/y6d5hAUCMFb1pYnqi+jppsFaL0capWQRZHWsper
kl+BGednk9B2Esjy8kb3WYfbFMGpJbjHxR8q1EuMFkAknle+fnqBeRB3LYMi8t2HcWIRiA0qY1Ak
SS/4FnKIarS1lrO6W9v33lDFpdB/VW5BhK9qNnaJTbklG4hW/3cV2FiOnv7jw6SMAswXArwJhswm
6bfbJFWBvdXHWJLUTgt7skbtTotjGANKoPS+gEXG684GyuYL46mf/1sbkLVh2hjrLLYjoiZOTM2e
1AK7T+tSHd/df2EBGU+10ZkFCuqxfVgb4104e9m/xKZUgk/BsVkSJbXkL7MOzAJ6XX8uQiav4LY5
OkkZTGrLH3jsrureYI+kNlcSwrS1GfmGe8R9NJfysE/EBC09Ac/ee3kz+ksIYO/vX6KW3Ir8hF5d
TpT+SCC45SbkU1NnSf/m72JwGBnf63pKm/Yl/J8trVnVfWEznGyaHh5/kjVrbPGHW2bldZXr9fHB
4yYTxWF1J0SOuidqs3x46pNYp5bBr3YtzP970Yhli+kraDWBqyIdPxPqREEuoGc3wFbUv48Lsl+7
ZjoA6zACe0lREI/ocOGyqiStuQjcI4zYCCza+6u48er4k2K79QMo0falw8dgJyVHqx/v8s0noZLr
wg9+3dC3bolhMgV1gjGEZUHgeci8lkXs/xIZibrKOazvuYmHGfzMfMrBjSYN8OfN8slnkLbi8wGr
CIyvD6R5ssOViZB5eOd3MKSf33VgMxuvntQrmq47mMQalt2BAIWNGf5052iIjJtum0dhcZICW9ok
OIhc+rMx77m9FxqP34dkfwBombmW2noFEyBMjPXAh8HGyRI6fYQ18/KmKbEQOrtIFwzhGFP5w9FV
t/8ep7j9QG3BWNaSZiEe0wkwWpim8b75d4qrUEq/tOS0oiBuNR1cO18AByoMsxDpX3r4i8k3xesT
9B2/aBEdxkhQzc0ykKEbyKsLXc/8HqCLd+ERcYN7QCtS+p0GpJmeqGVcfpMZhvLezfnMc6ZJ/Xeo
ji72fKnqWpdkRiF/jPrnRF0QTtMalCOwjlylYarewgI0DpBygeO0ICa7LRzPrxBTJDYhsB4rx8ug
Fr6/tVqEu4gq1Prw6LuOv49JyqXpkJq0S7lv4XnbuaMdUsWdsoE01e3NXK+JTRWs5hgiWJL8hEum
NZwjSPLAs4xF6S6cXp+Z3zqkMtguJ8wYVmZy94865ciUscy1ZMdz1L906srfaA0L4QJ18xpTE6Hl
sS3qJ/GMxZjfsqtLW/WKgVgWL6sRW6IB080h0qW7ge++kCf8BLywzaXrtY8Q9TDMsl4OAT/yYlpV
/QboW5CL9IyZIILygI1be2PGBT8hl26F6ogN3TNApbFdGU5pQqCl0WiP59UijVpRmyCzDt0CjlNC
TrbDcrPVPVedcOb8q1FY0LPMxPcU3LUCpyVCT/lZB8fXgmwK9MxTq5AKbRxhxZya8kp2SPQZs35t
8zypDrudWNMKZDr0BgtBGikwWlpCXXIQaMmjf6d51s9cVOnRrPGO5IDzFv0GU4WsGWWS0DU80xqd
YdePLpnXihaG7MXjhJBcAUu672dlwXDAkfC57FOhpgQhPo4c/XHqatC7yP78SyTENQuJxe4FlkiN
cOIjoSjECL6C8CVsT3qkxXS6yWYT14SYNDUdEjm4U2ut04SdLmVk+NCUYHiDJ/Wra4LaOofyqCwa
Qc6QS6hdv9mkCO/sUE6Qa2Ra7hYRM7wvd04wkoG7iOuMQgcLZKC5VBIjPCzaznFwme+pdx+5/JNk
praXd32+fd0eA4p+xR1d2xFzwsCrCsun+esmFAy68Kyk2W6O3+nkZ+rDiV2hkyq1VnAEklpnjMIS
FwWyJL9rTYJrEXJU0v5QDhiM7RIWRKa19Mt+EuwVxZbFdtmoicmOINbbO2oINhx/B8tOeUts0D1h
Trpg0EtTfvi41BhV1hOtprZ1zpZ2xV3ZFrkWQ03EsB63R7h9cfDrm0J7sgvS8XpRvFROPulhZWuj
u0VFlGo5856aHs3SpMagWgrqOhBQeH+yKeyJl5l1+7D4pA7MgrLBmgkBhqHEjcDFv6gtkv5KMZ1F
cVQdBEg6MS+UrljHwavQQfAgEvQ1A/r1Ubf96vDMXb1gGSVAb1d6INnh5DtIcpYdoucqhQC6IDeo
ajL0IcHakTK4AxCmBzXpNmXsMv1XgS83bTg+KJvVYKczL+Iqm9Ar9HFUqvXYs3c5LJbL+jqcFxUb
yzflrK8qDw864N1PCU2ofg5Okr6RvfUFzN/O2sj2dxXxmCR8AG1iB2mLffO90w0lyJtxUSS1T/3M
wVHrOIFgiT3OUvqVArnHd2j2z1/dhF6CJdFAejp+dooEl6smI+X7SRxOhXzpTuJaEpszqjk2liyX
U4iHpDzrLtt9w2c87F4va+YttlPzCupC+YqaBGnAjT2cgjVt7v2uOJ9IWjw/0KGjEx+pWDJvJAH7
SZZ8SXwjofQ/31pe36WzOB/LABecyU17vW1U6Km6n6sWB8ayxJsfZ3infMqmia/jw2YHUR1TMmcZ
7TyXqWlsZC1/zzWS9ZSnwYJTIRKpIobT1j8SaFZ98zkfOhKSiMaR0uJscGQx2e4NGHeeaODJP5qM
wgVOyUGjTJYV52o2I7QtQuLC0BjuwgKFbbejeX4K7RCll2WRjEqMdlOLFXVRx4BxQHNwsWxLw4jJ
qm2fb7fY5NCWRL0gNQPD9zwirVezhJMJ0jYvsN8oZmLl8sCXomb3w2WT3JjpFDSteSYdKjekEuzK
MRINx7Rqih1Ei4uV1wU6jETW8FPaA4/AIsQWfV76vfcq6x1Neznd22YGW4pIzBcUgGs7G6xkRqu6
gzRFaEsUVTDCb5QugQQyrSdWWUPMDOODwaEOASgVo46dOKRcW0/1I/R2nCZ1TIwlCLGDO7YHogyn
Am8TCTdi555AzkmcVCf/6XhXYWehTkKpfUbuRvqgT8fteD7TIpdY91WZJleirnxKZpPtNq7uBsXR
HaqHGobwdh1awUuRICYnKuQndWnc3RsaMztKdnl+kme0dfPqhqb1aJXJTkQJhhHxN24I+We+gEV5
1/VP1lNGh9kR67BJKy/Sf7TghgEqiL4jxVHPDH5vqXYrmRXuPzqcD4YX+q5IZV2YNHhh8uPRFDcn
qIs5uJSNfKnG3cyT6BSJeu8ht72q70ELQLV8cqbz1R6Zuj3TNJWjSOiQVrLgke6vzZpEW7vEF16/
78LBl7/nI5OOKUSL68DG9qsMEv7muEA/zkgLwMglNrOn3DWITOugtblWs8pjs0z956V3KWjN+VDO
O+S9/6/NpFbGkOQWlNckLGHsX1eFnvVHO9jwRm+Aesr2l/FuM5m0O7zRt21C9YdsodSDWO0pkrhk
AHU5gL16AkA09ARQ/eXpjAcjn9EcYynKyytHd+qyZXsKJ5bfoIxC6TDQga8Exbt6PkuPg8dnCaEL
mvDmxsIxu0MbfE6isKvI0u6By5lZkJ605+CEa2YPX9vxRZ+yCDU4ty5vSh5zBs5q+MEcLHSDN4t8
HSoBjWxL+2F57xv3NBgoiKRx3RH2CQm9wDGYOsQPHRscL+hJNRjEtYo6hdyc1IbEY5RtG5xawnA+
840GgyI1SuH5Exsmot/BgTFCy5sVuST7TW0ceJ7ykMcA8CVsyjJmLo2pmzjou8248CVAGybD5qCr
r39scuwfNaA9YV54Dm/s08UsWCL19c1qWC1rMItmsm2yvtLIvjaZNw1bSC7KiHqtQwyuaN7sZTXO
WrvvufTy8i5HIhLv7Q6PxhiL1cNkV44aOV0tlGjv7ukmHgjdSgTj7FI/JwyId2Zr+gx1drD8CAJv
GX64z/GhddXHs3OhrtZLOBV2fTSTbadAXzI3upT80mKMOxyBeAj3+TgHUqtwVx/WzM3kGRBAAcl0
RcF3msw9nZfkzfgmW0PVv349+9Ui8wTlabXqkhGnLsZFoPF1dCcm3VbEj5vRhR9HoQLQHFG/o3yp
h/M+qM/FboEPU+4eScClsWDDn/U/auu617V8Ukxutw3pUHWoBEhv1fi56eJxVzPfKjIu/q9iCySL
bpQC6tdqW51ndEZNPDAblXDZCJ3piZ/Z7h8ls4v7bgUEktl89a3RzJSCt4bVptCEcz+baofRaYVf
rDbQ0Sf3vDckWRBKjhUk6zqO5vjh+D5r3GGdDgmiWntNXqALm1B42tGxuBou2Pr2zTgHMlPDnMx9
zrjPuY2GQTCHX0DwS4IlGlIz8MLudZ4/dp+fSkbUaT6NpzYtXF0Vpo6h7GqpJx1wzd2SrBprEgP7
A+jt0NvPt40SecFhRElTnmNBnYc1IFWH11098YVRitHrasQy4ovrKWKRN27jnxMd1bHA3zykBtTK
JXrMvchNmuass711DFRLRp27jfF9UZjl436jClzDq4LeEn3dIZ0XD6CvAdwGspyjgaxy7nh9jsGG
p5EGsF73dIFcJTugQ8E2t7zhfIUxkUnhO58dI22E7BAGtzHCkvk+U68h81axgrrJYmy767JtOcxh
YtwLiz7fO1hFYeV3bAig/F5RNKXEOKOk3XkTNmkRe+EY53FetpMloat31rfTBXGxXNcMF6YCmb94
WTW2wZ8xqXtdEIgwH9NHkXny5EcW5mqWtlViUZm7M3TURQPnrfy7dNu5qyORokZ8NkHkb7shUY/1
m1OIIplW5ZEjlfUVYUNK4gFVorvVWxWqSq4kkYznxTHXvkxwuz8+e8DunYU5auahbS1U6BP7jjy4
DccYuSJAxbbnNi3wjkohMWaWemHh+buhttJXbo6PF7mmz8B1NFNxij0sT580PssY+nP9tYwKSIx7
l+zRqAoCFOH3Uyj7vrduV2N0EdWy4RyG9XQsfE/cIdkg1WK/dGME9XUpCVoKNzZ7r1DFq3MJ5A6q
tBzfYuj47vi8pvFtwIyKwRoFTAzllcICDr/jeXAs3g7lZzxapvFLMOYtctb+OTYOo/edymQ3eY3M
92+r0rLmUXN1Q22C2Aobq+dCvAB3WnspNuuP6h7pEsdXXXmSwILrOp2EfZcIKiikCJKiz7TUKcv3
5CrdTGsFZKvbZ9fiCxlF3M2jiHhknmPk2oGeT75rEvugqua+yxCKBH3pALWorvVO08LQV9POI2so
3kLMKMdaSEeDt9e8sPa6HdT6T+wWe5KtbrDZeMaepSt2NknzRAXRCqQCbkAh8oA3fpEgPCwRXW61
2Hm/c6G9vWOmRHLZCf0gFxeJ+MjlHSrei6CmGWliXgpX9iOoUBXClEFtwlyMr9v1PktpEdD881vQ
Szs/z73zftFLqO0ksQPi+ijzUGS3mPANeCnscz9OFO8Lp19h1I3Bt5i72BdWsjbWWsxtJiQcUyge
fEnC95vbIDlvYdhArDJMchr+D6LtP1ah+PWEbrNrJiio7FDdPWDHDD5THMIS5X6fDcboczFf2ETy
4C8leE45uP51MeKvgMxwXg+yklOXwq/ByQybWIxqTRpLjJsrQ6ZF3uo2QwkVmLGJFBNFpgjKUKnR
qFlzKfNF8V3gqVWoNuehzkcW1g2NNe7e69I277a/v/pCJ59qQU9CBnHx9zbxSxghZ2zDXcFzc9kM
5bXQBDxcNydALBg41SY8JqRNN3SIUfJdxUnypQsyitosFujAZYMEtTSjVX35dluFKbkhMcIfn+q/
/9E8zsUZXmy+26NfXVyIFHyfPWzzxpVKT4YUI9Zdi1fPJoWBOV4LzZylYdjIMm1iStQa0rs5OVqM
n8nXEJN47Np1vRKMsFZ4I0IRcRMR/LqfMr/rAYQ7nUIvhtMo9qLomAVSMYSFbgBn5BnmK+sIr2tD
6SwGnnOs9/i4BobE1noT1LkjKEjweb7eQqF403foTvf2GTCTQGu6Skkf7byJs5psoMbOc7rJ3KY+
vYQeJr4l87Ii+Fw7HUzdRZhq2oXa/NL/a4cxhNpgw62oL6IH6slXYBuM+Td8wiqKhBgdUpw7GDNW
e3QdBvLLKwCqp8wRnyRSX53y+ZV7T0NnCX2qAE20pyWd18dBhlZ/usBB3GNO+rmrrIAU7zbTU3dp
/a7rDgRAhVaD2QGXOZ+Vc7zJ9nb5rnADGwyWobuoHs6f0Z0kNKSMnzLShpsXeeoOpVloBG6krpC4
YXSgLKFjzexZwne0pSRKZVJR9z8p+NVxmxo1b7BcU5EiWQgK4S8Ha1LJ9nn1WZrNV4FGcPlumXBH
vEika+fSnntCC9U6NFXtUK5nGhQd7pF/ti8tSwgGCCk98+IC0rsba8AWjsI5gG6KXZVfA0SUqzQN
ABrv9GfOTl5wSxI5Br9VhaMitLYTpPUqP47SgooJ2oYQzCGM0h9R3/PA7yc2jBBlYR6i38qAZIWb
IWHkQtnVUyPDM25x5aGol/7ka96dGmYKvxKDb46wt/BYsQVuW41w3zRCMWBQl+o0c4BXC3JpnYEU
jJvBAHxU0de3HHoNwEpGoSaTsAqUj9CoiWDxIzKfRk+5xU7hSKY/AbkIN9oN0AB5yKHrUhwus1gP
zBTHuP/vlwS2GcNzDDD3OQnJCvrgCSVUBTzg+sKc1R7P1JD/b3LZJeiYvnpCHKc/e1E37d3z/vBm
qLPCC5ZikJ4oyaJUIdkscGy8spmGs29Hx9v5vAJsA8hTuxjGtJY5emb0EkFqwSxVWdRL+HtNmSEW
o00PQD7/DO2IGnXW3/Ufd9LUwTYrOs6gO9RNWKs0Z3fPGv2fFTjrmlpTUPA05/sviqwktmG9kuKQ
M0xSwLKt0D/reeTRWZWOW4PS84a1+Ic1Wvr8wZKieLdiCuUGzx9ZJtX1DLy2w0h/hEpx7mKaxMrw
OvIf5VbkuZCeXtRSg9V9kNcp8v/CjwgeEqHTUpTrkwd55e7MEQSoimIDrzyPJsVzL1n+G7zsned3
1rUz/R7EnGHygNDEMYI4eCEzQJ3+gN/LsBKm4cjUt7Y6qvwCIwfFn72t288CoogHZlUG5N79UPyg
LCYzH+mAa1etzgAlOBnha5dpj3hVPVNgOFAxFKm4F9UF0JrNrLWPVzuygKeIX1RA7iogUdOaYQh9
/FF6R+E/ql6uNZprlYpg8Rw9iZDklyGyBfy/DoecA9jZhWlGICxIbJMwPLiV++xEPTS0HusN9SgU
WnABt+ag82HvEPcL1pofLg1iv74lM7Gl18ztdA49wGB6WN9bMyNZ+f/3Nplcvmf7k+YpNzH5w/GI
EAuQCBsDkWKOqRWhgIw0vc9R7ER3z2Hhyb83NtXDK47iRTfJgNceX+l+eJ5UZTeW+7Ygs+0BMoRO
bjtNNi1PROCwhUBilRJfqQpJiPsyp1HreyUhAZA1FNoTd8jYV5zQdMJ8aelWiJSbHUJUNj+KFIkh
/G4GEuujqWuUqiNdTEjIgV9YHitsSe2AcqmkxENmV9Mpzfn9CofmGUQ5mGVb3Aj1TMHqePjJGaSa
IpGEDwtNvGHgbnnrmCSiufL4FjuA28Zrdyq7TcqaOQs5U6KqSitJyUGBah0tCaiaOS5jOuw4771m
pglV+xdUEd0mPQMUOzWXxoIuqn6KUzjHHwDlSBct42baFFnVJVimbrOjEs1UV3WLTtEqA3bcoYh0
Ju7q+dp8m27ha3++5z45pm3SDAyLV3eAQKfbXp4UBgAqp/No6Xmo0NOrxsSrVqJo1ba3CsYfekPg
WUkQ++fkDwa5FahB9NqnGCJlGufoaYJuVC+9/LnHo0ZCSYlmE0+kORa5FgEGrYM1si/OfuvOYmJs
QKA+nNVqmuew/wEOpWXq5tLnj8hQ4iZ3eDcGBCkIozQfwP7LMu0x5PgkvpbLKP5P067ZJe1XdMhO
gmRy6TkM/Wbrqah1aH0RhPjHXklgpGq7YnaDdWnyM7JBqesKJX8VIv7k9C6ZaS0rl+QcLwimYQ4+
jVNOVHI5t0+fbXp1sPlWGI+Wg70vVgcWx6o38voyMp+9kqW+Xw5MOlXtXvNp+t0q5rpYcYyk9cLV
6V8S+/z4ApxIKtI2XyiFRUcOkS52ah9WbNI05ujsc0ZC1u4wQ28AE2JCMbJPEZ4cKI5wQju3pE40
WNDL9QoWrvW/GajhcDhP0D8bG+f7wkdbNOVqZjq1h7C2Lb0N+lRDS8l1doKPiwfu5TEaCF08TNvy
LNWOSV5i7cUi6vaSF/1WBGlrXfowj/OwPfn+SgN6Q1eX7ZEX1WYkKFhPpk5F5J/AlNPwDaDDCcNv
hPW2/xoTE8Ye1iW75+abRJTV/F9yqmziabB4Lq/QIE/leEftxgs1aG24Co27s3AW+WSzv3vdTQXZ
LALR3MeJrwG/IuyCUT66JmGY3SjciOTySC6Qj52M5tYEboea1K7F3c7mpsxKScJWo9lb4lhda8Eg
UY7NCtPJB/VpKhK6t/ZzYYDAb4jGE4K+pP7zloe52TvPPFoAFQZ01K82wPtaTituToBiADN1GzQw
k9aogrc/qQVqFliugfLvIxyB/CxfeTVt+hF5PrJNIa1eLlrLaqmloPJxW9UEr6QtL6XL0zX2i/hE
BEPHU94k0hpeA3FaT10BmYyXTKqtBN5qBYs1rKMGyge95d5v2ANnNT+l7dlbqb8uV9dPjfAhGWd2
HaI7ktmdL9t2l2YQzH6FFs8Fv165zAZF1QA+lKR4nV3BElOjfXhO/xD1Buion9b09ZWHalDRRJQQ
LvSeSTFhBj4h+99qKbXImG/ZifkIM4aVsf1osnuJ3dsxLufnVh11KSiLwNc+dcAdOaFQpzB7X/Dr
CRnPZoNG3Wgh/YkUEVzmW1VwxQcp/DiAAU/C7Jr4Rsltzy5O4/gZKzH0bU1FaIKw2eJ/NONJuAgn
KoNSZevd9qE03Nybfqm41cvQN3VnUVTpoaxrZz/7Q8qSY7uSHgbOCjYB/Rgw5D97wUvmD0Hce2oo
ljpcM1tkbbMLz+mpc1ks30vrTgFh0xSeN1jgO8NB2Lh7wOCZUoJ2JsJYOdC7hfFFGL0xFMFivVMD
LjFI1FputStN2qJF5lnZD5Ab9v+jnrOAqXMi8luG7aqImLsb7BL/AxnWvGTqsnCCTh/hNTvqEJ5T
vcazg/pyuyvWYmNfiJBJkr8NTYUF2mKln2TaQlzjfE68YQWge73fUuy3SmUCUbxDUIKxUbs0eAzL
8n7RJdj5vVHq3L8RGPW6HCBNbr9WCCaPK2Xr6PsMh/28XB1AZgqd2UVypTUSAMX2IxCEbEbrBc12
dWfG8eGCo8FVT1scjLb7jjXVV+t4/M9W7GI9KKceXosGlYS7hnfF/7CbUs8eBnd0TAK40YuyKKlT
j2UmmM1JSFjHq3Gk+JeIcrXQNappX/VL4ih9ow22S0KBrAPNEScOIqqA6mxSGoBT1lmkasXcGFOi
n5L5qjXyc56YHFHflTK54IjwnooHvmTFCl3zXbwnOQSqLHEq9AGCcLeo0GPuVpX4bdms+CB1JSsr
9rIgdc7rpztQDJX29krOmrSZgKT2SQKn7cjBgggbWwzlcLqWCXQ/AeTAOtl1wQw0GDPBENz6YtgI
FIS1wOFcOmDtFxDFJyH0mpty/DthtXd9Y7tsReUo8dsAwMUyNW/bOBor4b40beFbjEhgjOsk1VfS
FwrtprWBk04xrvv6B+TpEjXweXIHmhX1514cbn6rI0aV7b9klRDCgseIuZBAfbH6GPINxHgJUGZa
IskhalY3Ce6KZyTCSmPnbp+FQxGtM8fg3+V7MANU67BlY5Tasbr80tOynT8Q+DI7khU1lFw20ufr
SPmEUzRAGa9+b+3yE+LCgLgOk6h8+l043WpaJC3eotGfW8v8lsC+EMy4f3dz7/4tei526nK++lIS
Hfw8FkMPbTQ5n29n0T+a4j7n/3NVuuj5SDAA5n0PEo8lNXpYesMYWO5slXuAWQ/7WNZE+96nR4oE
A6IMWBq47O++TSDmTatJkdPgUSdjLMSY892vMiDYx1WOi2kDjg85QzQaonxXjCzvpeg/sVRv+dYR
yTZr/PG067SkTIfYR4irw1ecIEoY2JQ1NnN706A/pbTbVbiMsPGAwAOgzuy42u6ZfT1LT/1/VUEx
EQW+9sqadDELW99qILU1gTi0t9X93OJoaIFc7Z0xuC/DMse3apNHS5JRZAmepNe45VImi7RITYtI
9akvAued39d9NKL+9snhuefcUCJaNtvZ4LiDVIBUc3qbqpLBUorF2tchZDYOXZANh7+d+WKSvPPF
Tj7arLYt9lqc6s5T8TdN7Ec7OIB1nRcINvPTXgxxfbmV80L2OqzASoSTjiYBZiYUSeDUbTeMW/RQ
7MAzu6IB2li1hJk5d149xCPSVl38Z2qhw4sVo54z+O+VeTxK8JN/Fw7Gf/ks7OItIwGx7dQeJT5F
wIISOp87Mf2ngMaGeLQ5msPzEanOSZOPJ5/IasLJjfuXVD6oex0ZrLx36Hw7kKKQOYCw/kraqwsL
IaMUqbBRcjakKyXnlSnVRTdiWYj/A+K642ypeLIU4igyXZoQpn+eN4TFUJB18PFnn8PBB/VrGk+8
hz/Er5bL6yHJoOTSvuXY1jArxzsTCcQ2ll/dN79QjLQawumRakwJjjKXbL5IzXfY7Ii6u8tfC08b
cUdyEmbcLvF6lVOadATAbL309sKahr0mHbXIxYQGd1icNYZInHyTVLlkvLLT468khW/5nbAEeViz
8iHNc30/dtxG0IVFoo+ONAJ4Y67fZ7ElIW6J4kEHqEHRKDDKGixbPyrHhzQeLEGqMoSiNvYX/l0p
LCVdNpdAVKhhfNTwMOUDuWFmYnVFgRQ1BPLiLfGHH15qeh1BCsH0lxgxLCQuLafHRWbnPXBFctEy
Ea1a9pgQE1wqnQG4kFR+ipBlPs7IVMKQmXKpaJXnZt9lmsc76VjXTvszd35wKYNkFHQhb2Fjp1Hs
L/doHV5dvv3p4kDtThTMPKPuu4VQXHfJgBQ11h6AhEU9zy17d+LDbh8VLgjZb7qjwCkTKcFlhuzK
QEmmh6tAPcdTbMo4g0TVPui8ECxNikqwPxeNI1AlbSchwEX4H5I3wj6gIyszaaI8YdTvE/AXC1J6
WGaqqFhqcGoKpRy8dORndS/2JXI0/4lcDOA4BprNtnnUXBsjFDu8T1MH7XiFUxH9pmkziebiN4ey
HEPpLV3jeu+ncG6fjWLdpyt77ec3zg8BH7hA5l0TPSdPZszZe61+d/G8qXWG5oky9QZBZf0eKyk1
9Me9ldbP9v5MJToPBV2eU3fM0TZbXGQwLDYiXKYBUnr706uRM13JbFv+JBSBnOHzesNt+zCajjAX
aQNPGty492siA7CnnE/l0GfnWNTT/5kDiyd8/k5XI5crN6Dk6fGXYnZ/e6Pq8q+zvstPS98BZQcE
bf6/C7gKrEZNsLnnWj2uqOdPP8sgPQDJtf9F5qgByt1JigDtuAwVGd8t0OFp9zAVwym8JetrW6vG
RZsbwIlsSqRMVeRfb4g9+CgmCrQBZncKd7dN3/7SlgMd6BYo9xYfQwrG9gcjwSqVs4w1t74c6nHH
qFOLr3637dICJ8PVJxqH3RvcmgNQP4x8UynR3bP0J4Vamp1n+y3sklE2BX8J0ftdOFIWoj6kIGfV
Vx/zIoGKkxQDMF9p8XwlRDeDQ6SHQbfLNnZUjqAawnWa6rPNaJ66Tv9+YHAPARWtA7QmlyA4e/o6
dei/+fRvhw9kmXM1LO8U/F3Bn4cWprEW296FJcDsN2/blvL//6J27ehfdZAj65Vb6mR7oh6NtLvp
pmttDrfm7uZs0RD6w9knSNhvFQ7SVFqb6lcwM4jhqwzHJ0QgD3bj3vKc5XyyL/H8Ty1mNee+Nhyc
v/YIkuaK4/S4p273DuwQELf5T2CenVg63RTTIiFvNbtBMmVPSCPpTTfY6nf+aCdkdqD7e9pJnRq1
+zftbN7P2mzXWSu0pq1eopc7DD54ueVv6FE9P3edc4tUEHZ0PjngnbvVgWIM1GiIHWWMrjTDfOSL
K+odz9yHTFy2ym7ToU7Vn94PEKkbLC0h/VzXIRUlLSUVEZcfMEwUMzuAFb7PuABHdjeg6eMaT5TI
XW9IRA7n+FvF2hPuOpb0/4duzVIQND8zIyCYWwNNM6v37PYlUFo661grfvkjlILfeppHRK5bT06A
8YGtRvyiokjFbGIWWpcBz19TpUbAJTKRJuHD+54G1tAsXnslnZQFhtyctSizKY+K5D1zHPdR+rfv
QIIoGWvYgul7R8mt+N2qHF5tDJLMLd47hdVoO3dEP+XwBy8nx5BR/SxFNDbHQFRFyvfsAFFgdbl1
DyfzSaRpQ5YNlCU7r1LCoSxlrlg94sfLgADlQlYr5tZjnhMn1avMe3cdIHsMv1Nw+3mML4BP27ak
yGat8+fcYTMRWSv8Tvti4u0dqrPpATGKVXe9i3r3J557yMahZ+tIx+8eC771vSxJc1132ebCr6dL
zS8DT61fRmI4JQtJZT1mBt6Nt8aqUIDR0NQcIjxQIlY2ubkfSoLOBVAgA/KIxVGLQQnx7AJ6HKuF
BBVb3rij8PXZ446wuWdinxssUoZUj3JJZYjIrWm4bK6UP5HkbDxzzWisOGL5/+LLs2re/o+XJ62g
ERZ2jDBa3s13uNQV74E/0a10TuzMv9rEr0MZqXn8dlavJl6ai5Qys21uxKEEf0ZNNaBISYtNGV0O
5iMtWBKBHAJzHN5E0e1BtYEWqLDjDjbDM3CQKIZMsH9bgigCwLvOa08MSUEEKjJEM3srNJrN1SQD
OhAta1j5bJeV47Sw10HYi/vqR2PJGFHrLA8KbvU25UD4XsL9GZkFTU61R0o5LIgG8VahmalSzWeR
t0crD7lf4xxzjicHiO1hM/h8REEXdqrhxxLsN84fH27PjxjsuAAue2cAv98cgwHjK7Qt8Pa4zs+j
uOw7YVFGRqF+3Af3j4g/gGdgK11h+dk77XFDk9TAu6YkOhgxQ0YwrHxMKKOLcQL/dNR/k/ISGB2v
jGeskwCGTd5KgOcQmiQHaIISTnzHEvV3HzKLDrL4+RO8QtNm4uE+3bBk2DnWEJ+XgmZs+uq/uts2
ncI58pdC/hrrKrbEQ7Xp0tOrCGUcjianzo0AZWNkKvyeZK0ORmCtxNbcseqghmPb9ULYU73DUC90
h/H+evBfXDy7yMDUPxl4DhSW/LMx0D867FOTjU4l7fe3N4KyXSWc+0O/Xmn7GJXJCfCRWnfDkQWj
V+z+J0ZRTdm1tbjdeJ2OdbpzV88f2gJx4eCwn1ZD1FqVVcXYhxVfd9OTNKJ+2ApTC+kcErm5xq23
OK4f9k4kj5uzE2FTDXAEIumBtKTMAy7jWAn5RhxiFglUoJ17UnaGa1Ffrta4UgaZ5Z5FGQSWPEHW
0NlJe6b5EQka/jx2PMu1iJ6oJsYm72PveSSsRXmcFKVhURf+qvyZNlIMkPYwUOr6MXjUSiUYIPRn
ohdMSFzXuNWccbx5mozMfTFaA95RdcfrpgHQdmwBEn7MmeCcOVodliiZbWp6rH5XJTFXD/A+U9Bo
79K+MGGRNrdM/+wXLP5pKhngQ5XWDnnur2xzqDhNfPpIbsHtf5GAaGFLAHqX2EXRiTq5lutUSH9o
5mhQG/bQlhIWGBiaQIt4NJfq4ATf3coYI46dZ7ulG54+1O95eKJzeWd0FRjTWYjO7TUndIGS3Y3s
CO0sAtlrSyFSfU5KSYEwNmerxkIhUuIR7/eErHuhRpZ8Z3qsv/dCtRAIMqA2c0rkrk+xIWhTrTnW
xWrBQizq4+2r/b0ijb/X+fDJR3ec8l2bXq9n5K/Batf58melzLJ25WfrK+ptijpK+aXBlUhhTPh9
NrwFb0iw8HUdN8UbD3L7RF5/I3OdkF+lPGbIFiWUaYBpSWTG4rlUcFge8j/4ZIMmDtT0QxeEHois
cPCm7+fzyg11te018Upjz0w4As5359wF9ePVYtKvmWtqi79DNNtKWuL4Mpfnnor5o5772zCpNmSy
wwgCbQ0yV+yprjGKpO7sxBAB8dw3yKc036MDhC3JjXi8ZsMiRJ6sPMgWhqIr95OltIuRhdRx+j0D
WoJW7L1PZ0Nd0xZFzLrIKEqsSquYgqOJxqHO+lL2uD6wu28MDU8QUgh86AQaHy01jkaTM5rn8pvb
VULr04ynaYWMzMeylIEpKOnB3fZUtkcP5GVVfsPGoZ2I/ehksswa7SJGW3KRAo8fxhlMIVoonlNZ
ayySNNIxIVdGl0JOGMfGBIKd1IZFAFXkmKIMKHTZQr6nZHwCy8A61A/HAFhC7Eq/0X1MbSnoNMAN
nVy25DMuxWrMsG6DoUkBZX3tlYrxo/BQgfgctysMT+VGPB8fPfR491NPSrvblA8pZSn9a0vfEzk1
NDRFBFLa33lERIgPu4k9wKrJQ35n0gz7XQTkpHKxgRBEsiP5CbWN3Gvcu3oTOmsQUyccXP8ei9uy
k1OH9xwYv1i3l8NvPUqry/s/Guz+Mqw0jbI2CbN9adPBLw81fbl5eyT/zZvvOq5TMx/i0B1VZQkp
8XVDuDByHxapNH48zHepEyH2+PyGIey77GFYZMJhD4BrkCFD71YZ25tSxp7YaukkM6UlI8nI8kbj
8kHyAIgvKYTbyXB1fGU7JkIABhhQTGKkwi8ZzEIWfpAEgo6xAqQQw0S6/JxYr59N+VFDfP2joNry
VAich3hqVezWPG8baXihOaF63acVOcQbatOZBO7gXX2H8CdhodsGd1hKYu4PSy5AqgIHB69U493A
7P9PVPCp7hmBtyuebERONBcbiq+Vr2uGwfTXkizrmCXLXUyPm7lHclGxZ0hamY4BM+TziTCXgfTo
sH+UpIo3XtD9fX3hNGvSjg4wnFxbk9BAL5H011mJQ8so+08ABOcrkJH0p/EdFn+fxWYV69hjlWNx
QkbWoGdT5Dthmukw7iQ+kwKWJ7gERIqHJsM3ye6l9DneGZHft6g1hyqD2TZg0OJ5C5UIgM9PCr34
8DefIw7wmlVlG+FPXa4pZK/q/RlEXFMMPK871+YAnhhnDu1aV82ePoy+qDPbOZadCkTmqrn04q1a
K55YtgvDbmhBPN/VdYFgaRAFyOsqR7MykHHsqGfrw63D6ZAlpmM69/J2MbCCewuTAFBTSTGfMmBF
4ZSmugow+oeU7TwQe2+tAwkU58Nig2h7Jo0CSe9cGNpl01SffAJXpq2wgUzYY9MvNvHSZs6+MKQQ
KS1+lrlFJiVes/ptdY/sDFZDV/hCeHGJhh2FjPFiVbcDRhiRYWit+KNio/HscW0OxZu/638mJNuN
YfEDbFTYRhX6QN3xdjDNO7p54g1n+CLFhfu0OUNgJleTYJ38ZJLZnQZ4Vfg0Jf1OJQFKYsB1aPQ/
UhsUyad9UaEUJ4SJCOriwMe9ze1D3ppPA2/a9RoZlLlMj6uhBUzLeklkLnof9/cvYvly2jK339xP
xViF5rPccdyEuT7nujTF356CbaI3SbJdQuPAcsIPWM0BkaABRmEx/jR849ml6bpR86hoDthqAxwk
P8njP6Dg/Uo/B0VMVBy31JZwSP0ExHdJgtBHVKBtAOwQVhyI3PeJq+ZE/W1PywaXUJB6BGQfeZzj
smoJp9p/+v3HlnNq3lxNxdrUuVj1qXZGDZw3GS6ZPuLU8o/WqzZ9Z0e3u6s8uEn31NyG8N0lya7o
hkxX+vE43SasgNgUm7EiO/5qJbxNrT7uP9LQf7B+QDRWsWbmQovgchbtCBtr3XpCQP8nWvsgMKPX
S/naBE/ctOpp5Rq5ColMOr+X+nJIeFQhZpVWK88VtHysSXCaT0pELl3qoEjY3v/uIFwQjf1Tls1F
lEJwPKzgI8m9m5Zj4NMvCXEAlgcYbmod8mtYhq8tba4qDuKleJXhG8QG6Kw/pV7wkODuBJyGVPDk
4M2kstodXXXq3wz+LNdAYXnnGL8/qTImYhjqTTQq/rFVsryAi2jbTfAjExiO6InzjDu5s4M2fdzo
QyHNPtrSiwXAXURUIPmBeziajC8wrCR7dgOveipbiAKzaH7pzDZ4475sjyXO8KPgd12fcx8sXvws
t0ev6WA7H7JpXgleB/jV9T9EWkk1Ssql51u5U5W3nXADd9SdBKpe64MXKLiRxE5nRfLZibShXB5O
3kKrcg0WEPKREIqSSBuhzuj3HaJ4+Qb5fra29ihAPefrBmDUY8G6AAZ7UwC8Ry+LDOUKiP5Q3cot
a6lRUp76LgPe0bq4RuDkTUrDexnluTFDIFV94MTaMXt5twXlyKBkdNIxti+36z7mzYGW0GuWsOYd
VL3qOwUZLjSCYxaLxLhO3BBwyrrOZY2KenLpu1MyIkBCrcbwFan3J8yG9bl51Kaqd1+2TmjvsS+6
sYsggNO0NdtD7W8xjKj1t38awYsoQIFqej/y41d+gVt00h9fDMfhjn+6IyamPhmPhBlvLzrHuuuG
ePtQuWw1ctfncyaKNQXbuv+dcm2p9oUvoaMnESR9uagdK1+gyyHLoGz+p1QR+Q7dTpPWaaFLJtp6
PKyWu5m7Xz8GQB10Gx4juu/Ooy3ek/lnP60KafYTsbPWvm5RxcwmEPD/gmBqC6umbGQt93Z04j8L
2aTeRxn9Ahr9OxwJARlHzdupirgltHyJ3HFOHHqlrBxYI2638neYKgolNgFZPwMSQS2SlqpCxmdc
6stlgY+hUfRCLYpptWDaT5g2Dsa8xiHQ/zoFs9GVZSnzYIbdU0Xo/6J4LsbafMfPU+3crbHu0DYl
nW5hOL0m+k+oPJSIdj+Fvg75VRZapJDfSKhhsbOHupe0btg66lx87J1aU1zL4/RRjxAFnFUTDt3N
sQ/d2HWfHbMBJwoIRJ3uzap+XvnCvquV7U10qjVLQMofWmyxAVUzHrXAr9lJvJ0DOuK6XsQpfLPp
YitJQJflK4inqmDJl33vYFCWVlSpLuqoYp14SH15IRsFtJCO9dp8FFjG+5yYULWc8jgLNdQp0ioP
RHdNbjlz2zOwnlemIFUpUDGeKV0I96vMwq0Iez3471SnBqTGVJcrge3qmvhWiir8KmCyUj9n+IK6
MM+vF4g8aUwTHwaOsE3ptFGKpS93knMqCxhieszYl0OPkxwbc40k0McQXEkbW17QKphWjpgNAxct
NprgOsLclQ3tt5Wjh8GbAf9CkNEU1yPiTggLBmMj/ZXIJrKicCVY2YeOWefN3wkZhMpPi+lrjI1p
gFksfBdhyZxZgwzI+cG1nGfPUN2cd9hJxQK0xnKMwaz+nKIBGmbbIfBOD+uBXXmP/ihmdluFIBSl
oWWHHkNtjwmqGVWkKoUVPDo4AQu5Idc/5haNiKEuXR6ExsrJwA9ssjZLXfWyY5OenaWMqNvS52cn
6gwcZCNdI11I+KnkG0zDr3MUgdOEtWJgYWMt2b6ut4+Hkvg9eIzBYCrGVRIQcmRXeEezNpFdZKM6
a45NnNHq7yFxZItQ1ljOs85fJrjtGhvZh8TIkVCa6grADH2fEPQ5fCU1BqsFi5Cm3jpdrOn/MRY+
u4VgIh6FDGH9k0yJhzNbDmBg9kfkm95eVQWcvKBJSX86QHkO+qQBB5DHYHxCKDAYsOoAqaXYcRkG
tdS5wvc5lEzDmPeMYoPakjiY4ay4PDrOPi8n2gn9GSqw91gW3NT6H2RKF3mQDN81uib5SGU41RPD
+E9oYHo2HNX747rQuSxpd+AiRzuY0N2MRJbXNWxFMt0PUmKNPcPb1hE5deBZZJItg2uHY3qQ7NIw
/a0rDSgnaAUdEUHTmuhJLfdymn2TpSjlBN+q8b9rFwe2R6kL7xYUYCdQ5cJbd3wHATXZth7vjTUA
4QkV2gK541IsbKTLmB8v60kWkISIVQOsEH2BcebaCWnAitOTRVLeM/pr2FDLq0qEfXgYnuqdcDiw
reIhhLKWnJgyzZ2ufNZHwO/iY5C+vWSVGudAI1CV+wkJekWL/7f2Xevevkrm17Gd6o/wb/+tjhDZ
myRiiR2Ri2zXT/HuKFERx7wfU/bJP4CrRxuzDunduUrkNuv8QTFDMBh5udYRiSklf24/sGl0NbhV
ebFdn8fSR16uWcvbO9hDT7Dt9SdQ+55hwhwsJ4SU2f5ScQpVEl7RRfaW+OKbxyRRZPOzjI/Z2nV6
Rha5Z6TlaHpCC5WQKWUpIyr9qHF6faKBZJS7njNdgOexK4VsDVLY6XcfF9f5eWqylU3JVAUzub6Y
i+zZ4wr/qpIabclxTHJ9sxpQ2y70CK3+BiigCijk6WkYHQyFCrKxWadEbV+nKi5CMmKwJHAHgYJv
wSn9+1/8uLlDxLK2YHC6Zns+ZJvRKJyjCt00UJPmYzf/ab/TRqYMdTmhHMkZA+rXB5NbBWFpS1x7
56wVQb5wNLdx4ER46rmszTSXjyzqhMYz2nj+J8JhnL9+XIAZcLtL79tJU0JfmO8I0ZJJvHpHw6X3
W5CxaiW5nSxuMUppQwzqtl5TsYYtzKSJEpnn0moVnFnXtZrFRHHaN64WQkAOuxsowUDWLPgIgcgf
73GFgbwrYHD6T5PQeRmEFKyRqKiFes0i30N8lUhR5or/bKe1ZuC3LsfprrSdTetHzCuKlEX6G3iK
KfL0nIxcGuLRSoBaFN2t1EcpeIGfG4hw26o3ee8OG/9hDeMHn9rMmWa+NJWDayQQz7tjLu6O9k/c
lS/fxah78n1h/kPGzr15Vj4fstmXSxbN6+irtsDIQGlXOFwqwJdRP37GMkqos0d2wnQrGa+F6yk1
8x0SKpIqe+G4LIEEsmyRDmHiK/X9pPv5hL0wkYtq7MRwRw3Z7CBpurU227vNt8A2RpQz+xC2HWrp
evdxM22p8tAnEZZ0EAzDDmLV6Dc0hPezP+lCmW3V28ucp++uji6N5s1KnoJzpNGnCxAXAjN/ZUtq
aKALfSv52HonUuieoVuIy32tCv1vgXgrwHQvYTrW5U8tDmceKgA5yyL+Oe3uH9qv0xzhFYLxzr3u
QG84EZViVAcsyxD7cv38SrgrJCo3uksBWMuU6RejgAOn6FK9kHjCxsgUUUbMAaddPZYCmND75pAo
3zIzZ0TV2b7Kq/B7GZRmAkos7ImGPqoI8F9NXNmy7MR6If9rgbsC5EsIUjA32YouvEnvp7WVz9PQ
elc6FFkkgtusj1wrzfrwinGmd90BcpSlNgYOhbCKcNKoJF+KWORL81LCd+9bMJNSrRUIzVL+6kt1
PCpLrRFLa9Yt8F59u8/NG+1OA6uFxffxmQLAV7ona25qmFxv/8iMpLlLwwby0nQrNhjUjg3HKUGs
V9CU72WcNew2ktQ1thK/s4M7IoggIlLVdeS0SkyDUjVs0T2DZzQDlDMV9suiS8GgSR7i9bWvTVkV
wuN2ukrUx9JTKmooJcpHz3GFJim3aujovW/iwG5SUcU7v9tlLqZkf7zqkcKwy20Kmc9/fgK2NieT
0WcWqpEZoZq6Jb22gVObbGNwmQrkrhulZEejcDPlXE6ES0+pxpvMcoSsgWkRvBvsN42Zimxi5c2z
6fceXImiQYI5e0m51drK2/rEv3QHg6M5DoLmmeG3NMDFVACUAlMUZMwThMbi22QeSuGrdgVcaQtK
u2O/OF/lr4bU6vJH+H7LL1CRdUtjWfZjO9BmhKN542Q4ztSlKD8Am5nhcA60dbBe+GR029zb8lOl
6kUbSBkGk2/xqL/FCi6VnVkuiZEpjir9AkyENKstjIZjFyVllxiidUl9OR1N33p67KF/0het+Vsm
2bUHDixhwJ7+k0iLo4p5ZXfGYXbUYLmE82lx7rYkGUoFGDzWxK3NoKk6JoWxU2gfFG0SPPJIfNA5
RPA999+FZsijBvcnRbx1PHN0mkKJeJmaGzlOLaKhQ+JR7x4CPvPLuzER9LmALTSDBLFrXWdcx61Y
f3gJK4tz6YT/W+Now5XoFq/AVqDUPSMMs83tK9YFhI4tKPvrSJaL0pHgAe9w/cr4Yd+HpKMiw6fe
kun5N4e2d7MkTxdlWMjCSlSFXwug+5mRXBVGGn3EvJNwNmQH2FDHXdDrsXdwApjuMicirnRZxXo5
OgBrbGxV3E/liUhFnFqzYwB3U1OEwKJfb/VkrAp9QV0LXww3vKjOo6yc3ehyVOtQQgpjdkqSShOg
wwO7bXfIneIBjGzds3zS20k9b6+jIL1K93TycvODVyu/6yZUInsYpnZ818dMKZaMRxU7UJUW242p
la9N2xS+n28SP7f6sR525Yvi+3B6NBY9GF80AEJVAyZDCiqJK/KTJjz2CtKvFFap7vGNZz+6+6F+
tEyAygU6L1C3bjVEpBR3Z2QHYWFZISpYAID5FjB/LZnsBD39dOTN1huTmqWhyTvxZ4ZKS5hCaXLN
5RVki+jelhjF72jKZ/DsUv6lpXdpHG80TeO0yHndQA1t02D1U46Xn9vmCTsErH0qWFBO9H/3J2II
IcGeC+Q1yQ4tZSIrLy5yemMwNExNxINtL8ZWAl0ktThBmunw8fDUFO1iDuYvdi33bDAQAxq2HPzr
+hllgGrrtjPKy0HqFThDyr5XJ2jhQS/1f2nlDyO6PVQVaSk8yfqy+ub9wWRUMN2wsiNaNZ/3Z7vO
6tGjNJXwb7lRos9Q44beWstptnMeJsAEy5JnV9F92XLzvbBDzwKbZy2bVaCudCva5ciejJ2frqOq
mO6k86LczM2SqdFnv18NUeDog1iVnBjV/8XVW9HkGr7xFkbT01ReY6GSMPnW1psqSImBO1zhEVle
ZfUnTMolAdRf5rldQxmuTcC5rQXQImn3/IY0qAQLnGaPhj+VQ7y0+Z1HTjffstWCB//tdklDGxyL
W8LlNNhjtrkJKMIvFNknPJIWYEoNUrlB9AqscVw7jmBDPycbWA+1PU0LbFOWIRZ1zDq2y2xLLqI8
EeqHMiZjWM3nh+VhwmyaDwTL6AbYV8ZaDTF5ZTiwZspZ5/rfhw2O6/Uh4mQwEj39Bgnajlb0EEmv
BBjJJFZL8HWT41MEqmrHcPjn7SikzRcIHghDaY5l8T3DjN5VW3H4Mo8cNdHcY5Wu+5XtWO8OZMmH
qSHQbtHUunJ/CTEtZUzfZC9b07+x3Ad2bvzwcbzCsKxLNlpIychEJcWCCl4lyrTnT+43wUQ4w2+E
A50v/7dig+uwNw6x5JLDtNUKPWnGJRSYPAAg9RdxhLBII1RhUhPaQL+/9pKUj1y9Y+NTK+Fz89Pk
ilJQ5LqfoFKpyAJzFA1OdpzlFIXSnXJc5tgBoSYXOjAeAaDCMl+aY2GdU/H26k0mS15xiBItQXJv
tiLkL+KO6hAfItp+O/xash3SFVUGfT4GPyiQSdwEE/Av/LSgg85uDqQfYuSac5RNWRJKpYQCDjwg
6IzFBFkFnenRqzV3Jc0Q+q8f97WlKAE0WRS6A27aHcGbY3MzwkLewdLeDyR1gTbFhiZANPB0hqfj
OGZMVw76sehgkGptX/8XnxWTViKjClJZKOB3KOGljF7VX+AqhmMOFzOlWTEGJPjFhl0WzmxZt5Uf
Vu5i9SvqT7RbzRhx1LGLCRmavh95aTcCujfDbftBQ7cj916/lx+ERP5ubZBgj5nqBp3Ha7uLLCZS
63qH3ap23ngu1QcwBM6zMIaFWaYJ3MwjqVuotO3bGnYXIhiIn7+to82KYD/oRzCY+ssxm4dFzoSH
bRYTfO97VJkFCKmp4z5zrxA21Rv7V57j3LqWfLU3wEH3hY1Mqj5oRoHhF+mZ6+1PHr59y1YOJYEb
Cp8hWFD5bjcNI3KS5XleqdtTh88/xBQtJuO8n/0eNzWM3VZhbFwpo+giOV2PoVyCOS/w3vjVRHKK
ZpBroC3o28NWttd1M9A2CPPR3ojHcnAMtsuje98Dl22G5roUejbWQtJtdPRKHj78k39t76L7SSPm
NeU9/j2IEXIz31qeBGHXoddP+C2pGvEfSawrqGsop8RiCGRifIGH6JVk4NZJtQDBDsiZNDQgQiij
tqd2k9LNxcqW51H3oLQRVxjvJxPYyfrUefCvm/OT4xL6gc93IH62tl1efHV2dQsezzt2gIUCKoDB
v2LkaJPJLrHOUyqQSjIi1QGzJpuRnpAgW1p3PmDZkAEuLS/XSAkhkh4+fGFDGHb1jVS3barbhdZ6
HhK5J1djMSRDqwb2zH5qlIDF4D7/nu0ue/uRLNs+/h5fMPw55FQzsAQ18HNbHyPauvWE5RtzBHB6
80dFAfgql4iZxApufpc+559T6QoqtQUJeUhyXab+boaa1yviEnH6aQ5QO42EJMsV/R3tGQ3oA1Ht
3wr7sYvKkyuhXvooa8JOMGst5iwWKZDvPbQzK9L0CBatMF6GFzMPOm/dcVAxEcJSJi/R+6UCxxgY
vIFkG/T5K6AmLmiQoXSlmTZaHnhPVI/lfxW0A9qaA09bMuf/EnaeZrTkaiSL3e/QwBflKOthodLL
2fTV5GmlqTJqARJHucWd5/lU5Rny54BjAThu1PykvJqv4ONsmi3oElrqco8mFVT7E3Y11W1LmzZ3
fnKzF7PKkzpUva9nickTIfCf+g17ybZDxs5BzaZJKHt8LV3b2vV2X4c7SxqPcfOf3PjJC6huNEA9
G2E0BKANK2FmVn17eUgV82sTCuNE3c2JsWYsJrtGSkUiOw+rdz4EFWU18ww4NjI+kXxDDpil9/OB
ocPbJBYBYQkFue2syJSSw/vX0c87N9y4KiWMVh5KuGFn/qsuZ7F0AEoHjum9xkQ6QJPH/Dcavk1S
YGHVEpqm00wV0k8Ku1uuXNSOTWzerZS8qAq9CNwlXJKWDK1XQcLTudhgC4uvJJASmfNPgW3BtuVk
BZiXTcFoaSRwDV6eLc7efBjd1n6Nkr5QHYx0VhPIIAJ7lNJVsG39gBaN1hwT58x9OoC1O7lFMPUt
ZGuqsb0I1RBNdZIBl14/6Isdxl6RRs6oyDajWPSaeuEm+aJUAlpHOAuSrU4hXERmrjcVXAfrtxW1
m7npjYz9ruROI0EEGqXJ9OH0B5tc3Ljgxssluf5abFen6h0mQeVWPBN6VlaRUXbtlFybY8RsMvjx
9whUuPR41C8qe7auvyzd2ptqL0JXNNDYIaOC3YiqSBCabjbmecSiqfS0DyK0cLcRio++OQXD5sbh
5vjI5ZGyVkrzclwc747GqeqnrkVgLm912A4WQnPAy/0hI/v/kuGwM63OQ1RZSCkO682U1oTxTQ96
beXTlaAIo+x+/ooiCdC+S7i5TQo8DeywBu7J+FOK109IBB1Nm0BPSwdAvW7yLZHOCQi8nRtV3UcK
K2qLZs7rvNO7zF/tx0Limfk//dc1qI3rXVy2SXro/hI/USB5/qMLO2ZLZ9n5TVQMU7/Hcf/j56o8
vphN4zwsHq6mrwqkKXfKM2N7b50UlDTqWb9+XlBUjQCnlqDiXO3JzAxqKbODjNJ6jsy7rCYOXpKt
/RQeYUi98G8M52nxTkXFQSLRVlNS7UpSfzdQO8HsANsadAsts86YLoVVkO1TxeLV+IGbmY+6b5I9
RNzEFTDcoQ1sNghmft/HM+M3VC9b0avPTt7e3ycAGZqwRQJNjx6/JzkLpScZ18WGzmMu8izNBYC8
/NApXDn01b300v5v3ZwMe1wZooKhMajWcPyqhDn5Z1hlRSAH0vxCsHJHx5ZWUj9Tw/Bi4cC7omWd
aa7WUg1m67s2iuvjZksmEv4gSsCZ140ZzZGuaT6iGa4juDZgP6MaQmSXNrX6m5iUJYmAu/bhqvlC
ebY/KwE6dzsaJ5wWOUrLwBpmk9+QayuVjH23edV/1EQ2HqeZqEuGC3BCZYCxRvtVT2Uo8+L8xDXO
0Mrwuev+t0zgrneYynX3H7SazmwR/LS4q+DP/pb4yp4nOWU71mgPDqn9tg9ACwCpp0AQKE4laGZW
6q3o7F2UY+XQMHGRpS35sGR2HEf8nzHp1hyvf0aJAHR0eewJpuW0TjyT6+8t7Qr18hsmYI6xfBVn
RJD1h+cW533Lvr61tzEjdxgXwTa8k7dvWJb0B00500oZW4dtduBxTYdmAS1M5pRl/CI9xxbHaBRl
SCJpCHf3f1hmpH1o9tCk2ACFL4SwBkQp3xEf1VTWr8VWs3Ihy4ywBpoW/l0xyld78qbud952CJaQ
Lbd3XLcqYrJ/f7lyc6/ugkAVWwdTc3LWY9dc2l2+alnsik2qJmrRGzlbW330g6E6Q+it9SY50aA0
yCPy3Rk+oIhmNvdUa5rTTToeXIM5a6Z4Wl6S0GtYg8XOCO21jcMUPcbAoHVRGEFzG7Frtr2OytzH
kv5QGhCnJ+29sa9vsmQUtt9vj1xFWHyXiSiSQy6T+YBdxzf1bLjTChXo9/aXCYuaaQYO0ZidvRBJ
rXKbIBguQHT2fgTCWTnhFb2QZPNAnnM8MBS2i9+X7s+Jxqn4CaXlOUGF1k82TjecYGC4z2+G1+qC
CD3mqv3qdXs8aiymRu81IhykMF1BvKgA069qzan4C71ILML5Dg6jo0hhqYIZtfoH2EjOehLd1CR/
835L4Bm/okbMeUUsF17evwBP9iHxb7DG8MU9SrA/3qeDigBMwjHQbNSQk0ThLtVArFPPhxN5SoIj
s6FOSwdfv0+gyA865KXUA6Ml4ETJu40wlIomNtkV78lSlnoGd2tV2GVzXFM9LDkZ1k4IZm4FZNSc
vRBFgvUrY+RhZytNQiRBCqXow61XgA0OarE5hXf+S8D0HRJtmQJKbZWyPo6aclWXl6/B4vwtdBSa
yxs/ZejfGkr6eNUDbOSKTVvBLqlFJOqXnk3AN6Oo7BahxCtcGwOuVHOXdnGy3cEjOp5ZNMZoOr7R
t55KAg9I0b3wk8S+muUAWSzMuwNzw0/S9e3Xpo18Py+9RG8TvLkNHb6EXi2ZchK6S5dR40vrH6Xl
RAY+yhvnu5n1Mgsu/fLM9tQcXw1vmbUZr8EI6adwcSmN3o8F3ozD+kDRttu6gdMob1E6JvwkANQu
5fsOlRNETmdhY3INZ13j5Agil50a7D0UQ29UjDRNZBLKlTRqlxuRqb9jXMdnAw68WFPHystchuoG
wMq2C7ZK8qiYV3hggDRNH4dtG1pDjzILzQN2fPSR3H58EUlQT2Iffb4BEoGMvU40lks2HHv8CLS8
P1klT/zphAothEuSPcPa91OvpVn7Ai+Rtdy7974RoxReTSWGj7p17WCMULO3Fr+9vwCMePv59yZc
Qavl5BI9dDDFDzDYiEIytXNG6vCI+j/iXxETbDT6kzZ3JVvar2WsfHBCBCjAF8Jq0DSYOPMCYrO9
o4wIIvybQPbDbsD5GktJG7m4ytgAv5WCWrTc3iQBaJJ113GERCSsOvtOh49LoatETBRrDl6S4b99
IQCg1U9WluB7KVH/nweFbdR310Lng6SDc0tNpVWLOKNKnRDYdTUAMfiakNOtQn7hnOz92gTPGbpH
UkuKRTZC6tuZmUhsxujfDub/tqq3YESCzGzvEMp2cmMyTkgh4MXUdLuN+pcGQjik01+VYCvjzG2s
yUisGOh+4TvuEBCbgCnvPTvAVKY2JldCBuEiif6Y4T9Ck7ocMVQsqHmyCwl6SEXJEwbsQOV8AsRA
HI2Pq9N8ZMMU6OzDVibQqcwMSoREZskOA1/68VfQoZDT0oUr6RI8rjdC+du4R3RhQ9xaCK3ik56p
hx1366Ve51PMJ8bE0BSTbTtW6/jJxCZp0ywJFMSSO/lakWApS5QhOjxzNvgcrciBNCJgijrjyPpt
TarTqdgWQJM0z5A7YNkLFNBnPdxS+oMDhENaBv0XvumCaRLidWQRnvQXUAf7tUEKKjxxuVKPBZC2
fNskifYDcDIzHS6l+wlwZ+yo7CHhLqadft6WzXNbFoOOXNvdnlKWPySPIOpzFWnTxoX4tSlYe1lW
NXY1Iy86LDoUSzu0f8WVKjrA+nr30Jl29vYMMU8OSw9J2XH3m1eIg6OG37YxfXVZEOANWS2RJ2/g
ZrZOWZjYoBb50ofa88ADgB/PNWjqxi85LP9Y51FiyzIGI2cXZOG7rVT/GP270x6gYbcA8biFnOmC
EiaurzEmooG4aueL6qrdMo3byK1FRGe8Hmnx56cvTo85+b5xGI9qfQowuZdGpL4aXQ5OhgGS6Cwi
Xcwcq9L7BsKhnEnHCRZN5v8dGdfAa+fm8Wu2sq6XctVBN/xVU+6JVJ8y4qMw1y5/uwpdlw53UBhH
YedOOuixB3ddckM1XF/S1r9A8UiB94Szs5SHWs2T7ZouhqBUt1iyGN22nTwrI8yuOtPzMuq6z3nX
mlsTGM4LPb+RIaCsKSgtGg/O/IzZqP0Y3OM+zHrDP09Wru+qNntKmJq5jAekt4c0iqelRQYh0Rgq
X7VOueYmEvqcDUMPyx9njwnWEkcnX287mLdqmN+VAJUPhT6GMWX2Yfst1UKFy0axRl5jUROrP61m
4o6llZP1ZBw7ZvP4VSMZHJ+TpDVoJ4aNIi0RFfdpSMVj6g704ZMb51N92q1RfB3WW+HBpV7hoI9a
HQyiJif71hr+lByLDkYVQBy7mwUk8zgORzgUCvl1hl9Is95QWBFwUIn/IZ91SG4K8yp3HyqlTZBj
bqbwPCdsEfJmETUMRrJz/vf22Bw1/On8IvaDRD7J0/0CDut2C85sapxfj8DZgjCv8zeME2XzYG7f
eQAs/umG3p6Z3RpY+dEb172lXu3/1xVrEXWyU8KTtoq4dRUZiHTgeKX2iM6XnVrU7OcHrCnvE4d6
26QRl4+FnD15tU4f8Op8IusNPlYA17+Pwn+MB+QCPhD4SHi0z+iPHVOHHGHF19YqZPyAPxS8Itup
QmShXpVUh2+MTYiL5lAdztn6t/JgNtusSnaKtJATQ7mcvRGfahxWAMU3pBGVPayzsG64dDFtDLHX
dp3CBIhqktQGjk2LY3Ik5AMTqsiPnNuicJd2xnEOz3SQRtuRM4+xHARndwXbQmb2XNJ4S5ju9X4L
5jTo2gWgBp7V9ofJH/THba6GXRDe7KeqhOH0uHKOXghvpOvlbU+KEMnp+SmmTXiEeyZf6pLetyJY
uZQihZE4/hvHEoTRKQ/5jRMFgynTe4eGAfhx5oFIehUSso/UiZkaPh9W134gyND+l/jS4+c5cJ1I
72iMAvbAHs20/5dm0tLBJrUhXx0BBJDl0dwi4y/h1KeqjvTgDGKG0EFVNoi5RyrmgLUEWI5FLQtR
gx2m/xbWwoqGaMoT1TP/hCTctWJyHsZ57JZofYl6dklgtqkG0flQDdkydAV40YqvTTA7Xr03/I+Y
dW8EsFbXa+p8ukwPT+BlL7wjUx3eEuM9gISdISxoOXiahX/Wc4PLkoT+fKwK6tmiakUjj3KMcYIV
Sc7bgWlXVwtieKKVDmRjYNGVi+LVfg1TzB7cel9ncSDxg8TQjk4BjEzpKX93iUWZL1MNk4FR3w7v
rA2MyHJg122ilHuoXh2hyUmx8r/JTX/Gu9mUro0HzLE4duPvJh5zE23/suKheolMPOlzKA26lnOj
pjSJQ4KDUHpD0MgFrEp8iF/K0+zye1hKQmQZzgrsrh+u00SJvPbmrWzn/6K+StXdt29U/trc8yUP
qFBKfpDKewxmt0ei4jlTNKPC4XYLl0Okak9mjKkFp++HvQIhEOH2vzUH6eqt1gklZP9JpsRrmlAN
yOrnVXTP9UQI+9mYn5gtfaIFvRwAtnSvdsYJJ+5Pcvg+NUN6mK9GNWl0/KGvz52c5kjAjSWI+L0U
cWjgxIZsBAQCBw6pH/suQWYpCyzwFkgw+E8s9fAc/4loFgq6lONd0s0/1lH8McROgd+WxtbTJYY8
AxR8Y/TKkUd24nuBS3bZh1oqgVX9tsN/C2ucZG2ik3Q5FYGkTVVRADGhhBMJOaS8GJQS3PPOAn3p
JNdj1E65MC9DxB0nQtcduauaQSlA4CG1py+XG2ye1Mv/PwZ7duPHTOnpQcYDmSbyCPTfJe5QJ+dL
MYvBcZTNt0xDD9uBZoDbaQV1vf3k2bPns1DkY0HGf+0Qq9+Xmcwx/rV7qGNztLVUJS7kwmmyHcGw
t1RY4Zb1tU1UUy2VoJ1jiSayNNlCAVPXgmkwhwbjwI7SFJPoQNX3BdsmbWUkhwfFlfNKLdCR28B+
ANt1uE1UJAUKhWUvJJfXQZNpprU49Q7S7NN11N4dFBiehzVQ3qsCpts3iT8F32ynaJauRhElxfaP
/jIJ6YY3bLC08d6nrBj7jyzQKvEeZxjGlm+ymjHWxNJwdGubkfdYlhbzitDZ0RAl6DTnzlrgxVvh
ovQ5E+HN1Oge+zdAHDcZCkbGhtFnD1MG90ElV3yj0kPGU+3P/LTtIQDupGdESy8y1Yv/Ais+ANr2
SoPZAUAxM/pdNiJ1EMSu08FfpT2QIDHDYhdRh1u3IZT80Yj5omkY9XFInJAn45PmY0uvrcIal7m0
e491IL5qdg1BU+vFxsaZfEroQT34knuDu+py39loc3QiVO60VydeOkfKLkG/ohYVMXxe8EZPQIzf
hfskRH14JKBQGXChUvvhDTtN9VzvYvOjWN3GdjTzaI6m/uY5qcZIgqF3eW35o+Kpjxi3ipepNJnC
Qi23+GrS3o1e5pFNSfzKvJKqKhXreM0SOTTsVmOdlcK+liRJmINDVXfFRzvslQSVScuStXDH+RHA
0pjZFBBETi6zvHCLG8TmPDWhcpeCvyULA1RV1k89ZdLYq7JUmqBM78E+y1HUaTNUR6xramuOktaQ
L+US2hCXkP4fh82YsGV3xcH2raRaeefaJy7LMWwCUQU1vmCLbUEMp1+JMmHbPd4EqtHDbWjmPRBl
xWsPtRlu022CYOlSJ6V9fM4HLwiq13xA1RLO9btrsTyIyA6GUPzq8EJnzqcd18hzTozsoQaugWSJ
rcXYPQ/wKASQXNkkG80W+5uedxcRuw9mE2h5Pdppi32nbeyAPSH6BU9BYwpXv/nLlvuxdJbzGVx6
Z/2cYKkXO9WzPVMu9Ch2XmerpZe4wl9QpgraK4dP612pbZxLFf6PoRNkrsGWdvxk7MnxntIaS3ps
kn2lJLU8sV9dlfeMuZ+pU7ff3prqnY0JYmucbNIoRrW4E3NhgcGT1lcOa1gHJ84beu0hF2bMPHVT
NoO/qlLd72FqzRs927np3mtl3KpWpHclz3MwAU25blTQhtkRZtk54KpxaDVLNwsoU0OFuxLm9gRn
Ad3Io3AIYltDxryDDlFcd9UNBj8ogVt+bwaAefdWmRo/kP1iBY1hBJ6mB3Jb2GNuruOLJxbJT0e3
Jsx32v4EAfD4nKrqb3UihskH6j0wvnfOJw1mcBFb9JltUNpKgZQnO/1HA0Q8s2clRDa21TtzE7tN
0dskdBxQEaxiIn3WqwX5ssnsJycbALQR92K0tIUxMQpmDgcK7MISMwBSMVeiQWe36OG9IB/FUU+s
xGB7EgT20Qmp634kD8TejM1sYnVS3TvQCjE/r+m/7ps9DoQIMwrUZ28fVIP5orYZjSMw70geSQEz
7fQ+thzqhpGwKcofT7uUzg+NWvvOdS+OTBEaLr4vHjP/+p/6MciT4ghE+MFNZuV3MJjWfOgpNh5d
K6ib6umm/69cO+44nFiU3lZdvwvRNzFzg5nmyL6cKly9zr/x15nfzJTiz8mnWTsbgTp+Y1PwmHev
hrHYQ1gK9NGdcQfs+Thc1n3uxwMdeXdJyhaEfw8t6h7unoEfH/T5IZUaSptxftIxDl+J3oV2iFOE
Lz7qKI0CTwSJ7HyjYQ9mf+sKjH5yusS4UXS9w6VrRxxlWVprzrIG7weDqJ3pwpoa6TY1+jKuQ/R/
Y992wmS3pz7j/TztZ91zMbytChR4clY4FvdURe9lhPnoEWwq5EnXlpMx+dl09ToEsP8tNtGJiHkJ
DG7v9Yk4zF2TLXZrwVmlMko3Bfg1/fk1DMfaX+6XRtngU4RvG1EXWTt2N5ROSIsN7RF8aZp9Oit5
o+Ifzqbj02uY4UYuSddNbuN0+FgaUZqqWkcYCJChAENbN5ml/AtghtH/MmSDNcG8StVdG3OhRiLC
hjZ84iT7IXfixqnWLzPvNGyI3FEuwBvgU3nLm52+M4Ff+21TnlD6FsyXewG00kZgQ1sOrgr4npMQ
YP/a8Y8x+LyS0uVEkOExrjLFWuhMHunc579wF3S/mR4CrcJmdV7of7OsmJIfhr8oAkJeuSGr1dQV
02mesNLtz+wrtSA6AoRrtu53pa9A+ynoWJY0RxjjmG/0n7/aoNj6cWEPGdT2xR2qInUrtAMcauVW
go7bhyPoYUZJs63TFjQOKeJB6gfR8KpXNjVNSSpl5wp7nCEYjhXo16abINS0SIktg3W6IDqLoP+s
svdJ2WHbdSFkYPvNp1v3agiupCi8XOTNHxZRBrCDUlx3xUWE16EuECYNPVlMDEPBVzkvgwEop/Mg
7gCxYfg2uXVE/bQBqEvgtqiRwsvLulClLH8TnuAIpE8TneouO0seH2UgDKCGb4J86JBinzO/hETD
5k8sw3LeGZDc019q++ooulHDD5ow3zxO+Zboilqa/b+OEp9aVZ/p0mzpludRVcwCjM4vEp6Zr00F
E49iTFKF+OQE2zaHxekjU9zCmDZQhXrPkBiM/4p5a4CLoPiTcApK2Gkppl3BMzn17rO+9akjGt6w
gWzaeC+xIqwN5kO3jfFBPOSlOL7FYlO7I0hqtl+5eSxlWDMhSktqWyCtUTU/L+YIlEVZs1Or+MCb
d32soRnsoehO6GssquEi8dZ1IcqmY+W29YjiS6EGeTBgq1KZBTsPnqH9OFTqPeCamWH/UPG6gm8g
rjObpG+7wnbCi+2giVi45Z5X7/RLK4DqQWzlwXb749b9mNkbM+yZIva1MxAKJl7i2nna8k35IJiL
TW9UA56z3XyIGMZuQE1wSuLhyL102GpJGpFceLG6dMTov6UYCll7c6xC05lfQUf7sO0lNdls3H/W
kj83r1HmPs8YlvJoeUH9eAoA1KsSi57X2GoFGAKH9vAAQXLiSUnHfhYewHF/QmkjeLj2YseWMjsD
RbuPDCNnvcUfpBjzwtNrlDHFOfDjraz1aNSTo3o8eF/cUZaY6hj9Q3a6OsVuUML/5Ehzp0ysgIXL
v22VF9ntwLIU+AtHLzdlyIhgo1bwqLIWO1b+WK5rvPs4W7yGAIKzJxa+dMCCwwVZ8TwXiJ49VfnH
sa6H1ktqgJHtJnLdzMcdWeFGlQHypDhHafIENI1D7UudQgznd8Y0qD5CadM+MyQ4VNcbmQxNbj0g
LICAgrfv80a5DXCEXfmsAeGRZ+sZAKJ66+orf4K1havV9GaKRFT+Uc4Bm5D0lkFpuJtniOxEKBNX
gB1VoQ+FKTxcioWQeS7EyPowtZXBPRE5usCwhI7VkJ8g3uNkAi7mI75wxPS6rExjjxCWurlSdb1q
KzYxdsThE7gaXnMuLLYiGcTfFmva/tlh4ZV683KByG1NkQk+VO52sSKSB2aKZPA5rrKhtwV1uZOe
BnFvWmbCATH+3MfxYfX5HbnZcgWQC4obIjZM/WbC1/St9krvJ+zHpyF9kngF0TOvIbmLG0/3oI/j
nshNxhBT/IG0PHalbYm46T+IYHdntaOSOIK015mVq93FJO6Zipi5BUgn/rjkrGMEp6loRoCdZd2t
+HYe0XsC1LdmV2OVu8FCfYmaSxTEPw/44UuUlyiaERovmW6/J4Jhz8fKgxt+tnrhWsgkCXUvVEIf
BGHbOJGczeFHjb40kQwNdsdA5H4aP4xA/VHlloFjwzo773ZsPI7BiOwU3Zed3t1MD7nQZrClVXYy
GwCgU6gSeT77E1X0pbCYif551eZh8G6zqs8BuiUV3uTdAJP3i4HzgSjyHwHO6+Jmq4IGFOOnxOLo
W0uairDp0uPOBOhEkvGLvUk7e+1RHOelH+N1ulP9mQ8CzFzT8ClYzFZYHKDx5tOa03zoSAavzeHD
rNRsIrJ/0dhwDQlgFHrJzasGiupPuqBq+fj07pPZVuRcUHwXL4p1f03aeod438PZ2J6s4yU2FvGU
urdOVm5kq0HEA5S/5ElqICl9P9Uq8gAeQDqUb286BmliX6hf2ftCmUNGkEQM/RlEw3jOl1diZXU0
/M1D4iuSiyq9SUwYoFH2UPcCLX+KrksWyOdQLODcgoXR5IgWOHCJOdHcgBqdhp+TeGaNy4SfNuNn
hk+fT4xcHa3+5yebLRXXmzVuZVrLFsK2oJyTIsfTCPG+KNsiFgrjqGpkQJxSIPsBaJoTyu4Nyxz9
HFkAzFxCudXLFSAVaRWqLr/csh7BByeywDG6Uav1MPFMMbp7fopnB5zdicuzOtStmcf832I6bu+C
ESJTbkif10HV+sw8nIqxA6GQjPy6+kQtYEZjf4D7ecWg37jbOT5zjOxFOBdPtMHLs1LNN16+5Da8
BWekEA1pqX4uuUtKxNITq68pwsOT+slHGaUTrToVNFzxbK69JsWOUJnS5dboyYVpiPG59TWLogjx
/7P+Hd7tORmOYQ62wWh0j7FZeIkg0+kOteGkNRD+GbpQutLJJnC9rdoy8B/YkbgyfS9NGLpIQO94
Tgo/stT2rJE3WfNbYSGnuxDG8tp5szhk32rXxWKTbmFD0hgVl2SKpuXoEkzUsLKMFIzo3yV74qEY
Eta0GGNv2GhpExC3uRxAKJpZm+WKH1sQo2L1+d1Tcv83HbUrHOJdqz5e5QaLrpPticZelJzWcfKM
o3ZpY4JlsaDg/ZB0El+P1Z1L+qAyrAP+4dRK/qe5JIEc91HzMr18VPnYD2pUvs/4Mn5EYXlJC2yQ
91LP8gaI27ef2fzw/bGfAzIOwjm20Jtz8gxkUXO46BFAVO8dwT7t3b08/AW9zlAGz1GdPUTOQffI
Nz0zfYHXUdb1IAtYuMAAG6MW23m21eq4Yp8Gj5nWjVqt9m5p8zO6uNCRBao+oD5IfhTPAEjtb2R1
CI+lZx8m5ObpWisLcQ016sBvkN/iSzzLB2Xo9Ihyr/4AUZ67YoUc+RZu+vhl4xb3fc9ME4M8a8id
ow94mBqZUGwY2SNxxtvX3abnzM4W9DCMZ85FWZQARxnyGzGqN20NAbBcFSo6nx1/L0KAx2VP9xjF
QiLjAiASmcHIf2Bi6kjPPj9Kfu6+UoAZ+rqkjn7Ee9QKZChEeCnddhfRO+OwUv4lN7puNpnBHj33
rgV0SuBqMOvSdW2mIwJDkVwPEVHNILYtzQeXRkkZ8TcURysTOZhhs7U/bseV/Ms2ln32TogMTVDZ
XyCOe9M+k7KzA/vZbxwP2GgYTXrMC9i+wrt+v+/oBX/6Y5oV3dwl1RW+vEPgIkvqTHQDaWhHjzxK
rCzjK8BOK4dSnvNZwoHHAmcYvQGSNgofbmNAIADYddG9waZowYHt0rQSB+wheE1yxNZ5EGZZqS8Z
+qKp18HulxXgwNbeBAnh8drNv0oHTXOAWvkaJl0hosLYOU/zOqmwiIO2+pUUoXly8YetIYzc0qRd
YoH8Ha6Xh+VM9W8h7zB/3sV4Jh5vUImmKa7jmOV7oiSqYSe1HLOnIH6lRugdaKSVVVUCHBEyHBzx
chLwmiEsplnRpHJnY+FYRmwCRSZeI34WUwbhveEJS/Ksp/M8QVxGX6KwkIwzhtnx5N3j3EEMCkBN
UDYUZ+ORnKsO/np582rgPS4yE7j+yvm2h31dcpM5yHKPJHqkHCScIWmc/5xoBPlUCQ4dlL16P70u
vt0Gi5L0Pxz8SEqpYmmPLp9/Sg3Otn54ymObtVOQ/sQyLMG1M+er+FrG2RjQ8FJMYomHFaT1H7Pe
ToPHoXopAx+jbpDayimPAU43dWO9Wf0mPcuMBKvFib894ABLdpDxajJ/7CENWmqth+A2xkz09nu6
dwhjzpKF0Vq34Capf0LtSObU7vjfPI4p0G5JM6CzDewhziGeerFBEkWkULx5M0nq+FCcqhNGbKP7
EHui5DI5X7p7RuZPCjDtCNHSj8MjaLhxAx2PNol6ytZPoTMBvqAqS6fkq+HCA0eDM7z51fQCcRis
LkrIFemT8g8eqc9q6vqWHTamiqYW8U2PgYKdIts/9qQ3mGvoB8Rt4ZrBvKO8gcmJli0s6NRzrPZy
G5u7CZqxw1o85gMpHSXCv6kpy8S60XE4+E12xLELkn2CQEzSpuH8DtkJyy6XHne7oJ8u6dhg3Gsn
TSgyJfRVw2FWWYzaZ8J9MspNrwbFR1O/a0tt5XVfGoN1yijQypIOhR41gYUCcJ+q1US/WrctBPD4
f1zm6pQ9OdXSFidOmgjDnTfuVYQk+KqAn1ntj+mVvvGR8ZeLiJ+7sHfbB+5/ApRSnN4SxL8OHHTp
5rXuF+Fz0ywzMYa7LgZidiq/SytJz+7uzVyOwHJDK9oWvJk8D28ZtHaRqLj/HDzUb2TiyetXSoj/
RXxRizI/OHZlz83TsQ5M3pflPABzbPMum8+p85Wnd87O6RNPfGNxvhx5vhuO9fdBIY3vYuy3kLYs
MkxDeLfOJT5nQQ3/fm3UQvo2scF7XJXAF/6lMMt4ArjP5Y/wF8boQ7CLeDPDGkNy/V+6jK8x68lq
opPOo9Cxi9wAvFOxAXnbnIp+jKK+bxyVfF53buITpm1V78Ux/dVYL6NnQQPpr9xJsX4E2ZBapvqh
jwkHgGn9iJ88bhSZkJwYDQ6NW7BehNcTf5cgLOycWPwNIpHTl6k6nsE0sCG7/m8XWRQBUxeeaIng
bk8bclJqVKbg15IfqZqH2ZUZ+wQ9KBDzJKamnFDCvwK6+QyzidUUcJS4qwNrd+lIYsBAz/FXl77m
PoJKZkU/4ksESzg1r3FSoGIJNtpa0PkJxm7TIqwPsBedXCBbjkgcGW8VDnAYNKEpGAUtPgbjpEfA
ggPLfuolA/Pq8rOpNsb++IpEDHz8gLO5dplT4UuxVwYxxLwoyw0UceJ7Xe7WQHoQXnqRgjpfWC74
ZdDkua71FAnYtEvR9j0xA6RoLPeraRZBs3VbHyJI43RYYj2ylZAcfZrCxHFNN79ruYHdAeS80M6s
uo9nKcEXcDRpuBmM0SJ0OIgYVNJ5MMu6u50I61nThxlyGYMKcgGVWQ2xcoaMOydPf9yUAnGKxB1A
WMoyozT9pNwmrR83xoJBFDL9zQqBvrIfd0CvkLd+XZwJVb0Z9BR1QVFdNtKAKRMocL8/EtnIx9GN
XKAnk9F1GFMpd9Uha+928sOVuKTLRi5ldU9+lkqK/TthXmau3DTfZkBzIv+I50MVTq5sWJo5T8HD
vTvk/2VF5jGuXgq+jV6dKnN83hEhOBr5eut9Pp6UzhN00ts8n9PV4p/i02iBJ5h3sFX3gDYNwqnZ
V0OqqP37qe75cBIGQPrGpjW+MT90END1gDYu0mnvG/MjZaozwrRR1h3AjOwUFj+UqJ05LdpBtZhf
Y9fCupRD0DgMBJta65UoR//V6VTSC1gZdgv7/ybCNzYbmTcWEkNVyijCAfA51b+kgB1quxmVKJP1
KByPlV0SZsnvzm1zLCkOuEFteDGFX0QZjm+6JE73WVOnHGvUIMcnMcC9xv9HYd5nqvyRiVbawsxP
l00T1Iu4VeolTA7ebiWox3O6UL189/iIDTfM0H5dgXXKndrFJmYa6cMcVtYPHJe+WW9VCgzwj79c
LjjHme6TIp4/5HAUJc48oJUgx8s9CAfRa8xcskGOZgI3Q1Hq2s47wSLJpqzEtp8YjTYl5xAhVSvB
Tonz8j0zIrMXTShwsGvB3lpG0pw7JcP1Db8tSMaghval/BOZA0kRJV2Dyk4WNkOhEGjcXdsb7TO9
+nKpaT4A046/5sdgnGBEgVpS8AUUNuzAGD1r3WszwrkEiXZ+SC64aDsSYKkjxi+FsuqpCqquUXks
1VVJB11qFUlA1rv0luJlPDcaKHFDxk40ZietKxio6WX5tf+9wayigb0Cxa2geqT/GAp/I/rpZApU
ArzY65qsvhissvjEu36G+U5+SJFFdoGsnA9KTOVHj1eSPbD6WaFpGgD4h1RxTlWqdd2DjUDmdZiq
sqf5lbF76bB4qeZZkN3+Bp28m50zAUuhBzFlglceyEZlIH2YKvhVRkOOb4UtGezXlJLM1JB+fqi6
YmpN3TfLQXT1Z2vx2EvITHVsUUKZKXi8nbU2SRV0sG04AlwQdXTd74N9Rm18NeoNrCeNQEEXA6DK
vIUs7JPQMA+4KOBWosPoTbVQVI8qcXMs6ggC3rdgyPBrr5n7L3++wBPVi0qkumrqHB1HpL5uHLIS
7yJxy69/rAjBHiD6mHIcgulDw+3u5CEdp9xivoGrrMDeuQ3G43dtilIQ+oyyrKe+Xra538pukDtp
663GcHwN5pWbg9SDu9nQeXt5vNCoELOmLBygaoLRDo8UgOBS7cfKut0dnH+DVJqHZGPBkXjwjclw
cihKWfYCVro8nmd9xJNR/M+H4HARP2FtrxV7Rt114Ct5Lbu0N+hJAcfQOzVBEc427m4vpL6SeRmb
fTTZB1RjFDCbsVwjTdvTHyuirUjq8ftQTxkU4SsdILw2RYKkYuTkBnm50In71c6AZ3ORc3Z/dK+7
kTeIx1WV6bO/VdOUyUsEecLh8MiKYBYSD0Jvo4kebE00CPqkiTevcAPuUCfG4sjmlXTE0v3+oxrX
jD/0u5rJtAaft0GwtXrbFr68kdQ6Zva3+jnyRckkLWdMUKOcVZSn0+jMlLjsKD+YPckNiF3oor0K
vJ8BH+6fA6iXe8rKcJukseA61kvlS17A0KrE8MGNePZU0OKMkBMlugrR0y7LJfi22XTf6CPAsKyB
SPjgSPoT7uuUygfmteVjfOt5zwYpUCkWz0atx7TnO+pMQrGNmSvApy//RgJOf5ZbzTvQYIolvo9O
BnpGQBy2tHrfBtjuxe/3dWZfMXmtV7CfWmTiQUU17ejCP96BtucWoGD0Tr6nY1EBqr10p/1Q6koN
I/wSaS63VOTkAoZ2eyC+ZmorDyqubjnYF/L3k/ZFZ4ubPcSqwkaPEtxTI0uLGknHqT9lL6i+oBTt
rpDUBRPe+febBPQwnxISyPU9inIaVvHFC9R7KS7VQw47TgG8CuedAnzKReOg17Tbxz8UpvbuqZ2/
5bXjrkwogehpNzLeZ9lhMXFf2v52CYWkwRbK5DC+0uoV3+mw3VncTvBbID12TFH/FqDUJLYwvWU9
7bsDHxEbuXd/x0pBgU375dBgoKnChekdQQwiMsCzqYeC2TEFtzimT81eRdQpnQHyTKhP3QVlL9t7
2CNCmCeE8ZcGt0KEcIZs0TdQRQdyVeyK5hs4isotLnq0Du8leOTOAQtnrtbd9Gzlxli5uO4lPDOc
DxIZsmWoBG9nB01uXAKKB1c+JpnV8ka0aBGmZU4Uvuwb3lbwUMa4wYJfkusWDpPZgHLexA85I6Vn
dxTuRFIjhCHqb1afwMYyhJyTy6doAnnPFGfqj7NAElkacOHXStGPYsYYtTJ4tiP08dpfAnAcb8hR
941X+i8Dko9Lan7AUT8qEFADVYdFdUOnZXMlYLkgkI46HqXoj0VyZmvS0UY9Cxiwae9jMGh3Wyfd
ucCPrzfMReT3xCdXY/CTn3ON12UF3UAo5sAYq/NTxTP714eyetOuw9tzYHnnTQFru6IS5c0r7wqS
3+JsUK3+nOBlEgPFmA7dV/6m4NZ5Xt5qfZXQZlV7R5JUVxCBWYH8f4FeeeF3uzWyKFSHVO7Wg9Bv
30reZzdzVoFB67GKes+GV5NtX3fsR7Y41sgrfLnUnwB17k35zGv4iAOIpOI0SIaGwTzxHE+asyfa
h3D6vIeOvEgZY11lhJ8YLxOHHNr2DzmPVim5kkGPo8mCFRVU6bUrxak0b5qL4NYjf6BdX39F5k9E
WbD49rr1O+j/qv5HOQnKgKC2R+UQCwVjJEF2zeCCZijigZIl/KRIf7g0pzUKPMdkov094va4U7yf
1Ru/bWF+nJnbcKpjjgY4gjqVmeiivAmqfcJWpJ53tD9veXyZDxRvjtREbLLxJ6io8uj/PU2JH+ul
XS8KKk1UyiTZO5jGxI2EYg+hOltqJ7L75JnJQaSAGv/p+ftadBfxzMjQ5J0lAhps1Ygbme0JMp43
AZP/W5NPsCOb7qZtextAG+JAp18yw4WMtzwo/n0x5rcRq5VirJW/gk7Dh/hDFsqPw97197DyeGck
cWjyPGaClZvb9DPyq9R/KWfF37ocErm0Yub4DDvGIzNwQiu7A8Wd/TK+r+s8NVZGBi2D0vC+RljF
nK8L12fe1uk18gqojcocZZZFzDT5MbFjNpyBezB44b6lJsOv1KTYrfpmVQUmrLZhdKqFXwMUUfVi
3fAPJi1aD0ZZjY3um8jpliLbb2xhRCz/oLbpjovcvBmzU2Y/r0KEUWgP3YkYaTLN4pdgUnof5H0d
XG4l/fBORlvGObwp6VaqzfKBQ58Ku+6xo5XUHoaZiwDK46dM9tlOJQuCMQLiJ40TYEvXzLwaHv5R
OEGnsReCN3SC8IyslQmy5rqoW752aRZYu1WRaCZ+xZViOZPE1bO0G0xKCClOs7AgUyJmvBFmZi7I
HNGCQiPLXes4gFdxFe3UE09T+9NP1mHfK2uT71qBJZdTg9zXNijyBNaD9KGejRtvRYXRRQfXbVgz
kEOqr9W04MIKGf3mcd7em/bGsYVCoe75s/v6iTrAyiUL8yalw2JBYfd8lb83l5W0mPsDC80OQaQA
xe56lOeqDrfgdXB21x+PqFvcdJnac/dQRciu2zhX6rJPuXl3HTe0LuvGXyD9OCAQEbINe56/CcJF
aa00xfHApe/o4HodSNFE2NdTFxL9l3EPrCsBhpgqhbx84RuwpdSBmenSlIMWP4oxMYg1yREoDLfB
WsUwMILd/7zdUFRwjqO+e75Hi/IpF1tfd+IsmWnfDZgndAI1nxiC2nvdRzW33ZnUrXKtD6DyyEwt
4JbQZSmgrUy5JETgBYLhpXlYcGLi1pR9fZD5Q9cdUxnH1wt2gmmqS7EOe3Nj0KuVNhbZQFLwlQVP
XXqQnPfBYWY92rxiQcHb42+ejHf+haYuzlftfJzLlVEXoLcNULOEDSc91LxSsyE4U9nfrcLY4ufJ
tF58yyRL6jncW7qaOMR5yHijvSOd2eh/D+b3rzcEoxs4aHl0dJs7+wnHbq+Mi6SdRrBSt3HXZwDT
qpNMZQ40oncAwqcpihdLW4HNC1HAtniLa447FIwJOVr4wYCLnYqCrF6TapNCxYCC2mLIGy1R9aO2
qWv4fR630qtYxZbKmfO7km3ahiZHoTl7UUCqEeCBOO2t5L2ZuEcl3CKWOZyheNa1pB37AiDY7U6X
EsG+HTg58mTZwlmA2mPSglBoS9nRhBkSxwK9cKm8M7mmoTWbOfgjDyUu/tSDTG6Fhe+eh8QyTrME
c7crn+i004dCDqUqPLaoFEIJHbMnYT4hxyFzL3E1z8XW3B2n/wut0shrNvrHZmtaGL8uGEUadhKB
GQz/5oMZgaFtIX/djgdQgYmw4JeElwo0kfextKcNVvl/pn1m/72NYkUhIQWFKD3nmoMOcNJ2pOq2
7tTxYdmUkLOu3i4hlnrYK7U8r+0zCCPzssbW/6tHhy9tmGN8RD2APP1LdQRaVUz/uPCn0+huftud
FUvJrFWuqX+OySQaDb2dYdY2ueSpoXJHPVvuXMcwKOjyY2V9DmogL72wV2wTQmUQJKSJB1ZQ4mSN
DhOI+BPOI9SarFslmErB67eMsmoqLbR0bZrOtoKO9ufLlKb5wpgRVichrmqz6I8/90vm1wTkkiJc
NUJ7KQn1VIAhzOtdbtvHChjAT+bpJktfDQHN7N5qrSjPVoU+6UXxxyhHvaAPXwIbLpiAGLOiQ1lx
zK0C1VDKm62agyH1K4v2QdcoL5chb4kduSkMMJ5fjv+8w7HYzva3d4tljNyYmcEhDyJDGMS+KTYn
WzwrFiugwlgSC1WCxazTOOhe04xM8x3m5PXade386HYp6bYj2flzQSHbMALufTKLKqTxLZilyCc9
fzRMA2v0vogE4iozId2versLshzeeMxABt3xpMkvvy62r4/sOdHNBUGE+RG+IdKHNamVZEBCZ7a6
xAcfr9p5Aqiz0Lgdu0lZfDQszf/AFJVxCrtymXBU2gNoDQmvk+Ko9x7ojm2hsb/a6hRnTNFFpUY2
u90crcW/Eih4GRN3UxCzPKW12hDY8nLZeV9L9rZsZHTZubvHR9GeHY80cFM8dJOOQ90PqvhZVzsP
xMmtrExQOt485iEyVa1dPSGb7ZqBWhEiJ4X34Cy5gdQgq7wFAGr9FIQQKHpoelsUIB169ZXBeE37
W6yHysrCgFH2nnTvJ8TDP1PK0XVe5c9ZFliy3oeoR/pQ70ZpWDZyb/coGH2suCho0rYVZzhIgtJv
1fOtnQpJorDfnM5KNOCODhSja41RzcDXGlIWvEVytRVji2yoHVQabGhVkA6Oob8fjtxzZp4TZHxk
GTUXSjds/pEwccaDopVcmtV8Z0lrOge7xlXJ806ZuU3AzVNUCoi/4GC4X1v0hbCF3vmesNz+hKjY
Ppd0aLQj+QXDiBjtgkk0UnIukrAoKLVRReyDwN10Dy2cblRTV8k156a/o9+wJNbhxP6G8vCWHXEl
U06vfmLffnXVi/mKD1pZUOsaiP2P91xf/lf0bph5JvWvWQaCcVaSmD6DjrUn0PQ7tOqmT31svZzZ
rEzKAx4a8TB1ghqFO0i8PUmlIBEUZGfP1dZW9nT4npb4S88SNdXrc7tafgeDqHsc1nPqfwFevw2c
nB1OBeQ8Lb6QnMthLV+G+mz2mY5luy9YHbY2OcCMYUn069XiSUtJd6ugY6hH7A/JUSHXoqdMXNuJ
aFoWreMB3t+zeGngZtNWFD/ILjAw89uUtTN6ryec+AoTQxwrQk8OhFBsDQqoU40RwVAvO4ed+0BW
Vz3EUpG1LEycR+vdSoWpdERzZuwbQiXFxErLApV6CFdLDx243/fHAPNEJgUB3C3jB+i1TrNQekaw
Z4axApibhxAQ48pjElJ0TfJpYDZPzdPiMsJHN+Xa6WOv4xmIFCX0zs9OzjVSf7VuIvQzZ/1fJO5p
5iShVrQkXWwfuLHjA7udY8zzGsz+oM+K3fJSx8RF17RA6C8pk8z6T6J9/j33Bop18MYQZ8K6tj8A
zOs9i4yGEvKyrK/89nI2Gntrnw/LxH5sBMyv8u98bGgQfgjuTTp/qhb0rJLd0FSpCcbutBQuavHq
Kgcb59e5uHDQDqYiohbb5aPI2jPaBBxxxbKjR+48w4s91fAuLaenHNw9SFjM/NfKNRfhe75IgHho
VAPYsyEM5ffGgpoxmwGbtnapKNj62Y+ZoC39w42DiIu05LXbGCxIIMnXVu1LjQqCcBEPwWqwvQbP
2NU3XwVhYuF6B1gNTThqoSkiAsjOn6KZyEEPpjNBmN5MbJAoAFYrP4wlpU4ejB0OVHiQiCsLO8tb
8BpF/BPauMInjOp5P62m+jUlp8vjBjXUEUFJygNWydM6cNbfxCIUYJ0SHa9nV+GFEeWBeP48sao8
qccufYj3NhBhrO+nio9R2myzQz4Q4zdJsKe6c1woZ4AJChf0DRCRV++zh5teM1F0738ZvNxu1r6y
+A9FBfJ14B1Gsd4mz9/o0xUuQAHYdQu3gr1OCMIwzedVZWLlvUZ/Wh30ewEDMnrHoUUHSRjDrT/o
I2Yu6CgxTkkXzfo5DFHS34IP5sAhjcJQrNvL58ahVENImR+aBDyK/wv8jq2Y8NzYsSJkbzDeyABD
74aCjyFTNohGUEOdu8oo9dY2Hly6WB+6V79Jl89MyO2C1MCqUWHrphTYPCM3zeN8syThbe61PglA
qYQltUQ6TiwL58jydQyrOPhQdXlk+PXbmEmCNIdXbK5IbfMmHIYIfTf2oKWNqHivOdvFTdfKy+U2
cb+xpe7+ngKA9fCR+Eg8tlnPhPOcNZ2e5dQzSJdpSJs0D9X9S6N5sc9aXPoyGDhmoRqMelhT2VlQ
R4hp73wqOoL5yvtfg/JhVKuGq+UWyYI9VH5Y61pu8Pbc5QFRGr6CthS42KhdeNvh0R/bujtsQuKw
E4xfJ4UFJMpdt5CBj/HPBP/XlwfZyhWFDdXU1H3Bgx5XVm9gd8ERPZmq67QQlPwXt8JnxnKgBYDb
f3WH76W3IO0yMwVI9zqdczrGFTS66Qw+H0qpdEc9o/FGn5czA7uAeqyKj3M2BbVcFtiaF1aoPugI
NR67egvlxqLyMoJ17bI7qU4O1LvSNwdxEBKTEuMajZjX/eXcQokn3F5SGvtvj3JqRP8COa1tECho
7GEIUkgQcwCvykJLs0GalyOWLT09GSnaoWF6tw+aoEE/lMk+4p8UkFY/EZwZ4yCaWne/781/DBoC
rNVjv2QtU8K5Uq2BCn3ofyv0uGGfeJa9T1Mnm4pcTFGRR7ERLcOQSS1UeGDcNlQLx8lbObtofSKe
/ETe26hFXKLmHlNllMITkwsY6Xpb+fxrdLRRuLCnd5R1jOM/Bnqto0wUSf0HKufyPPLhPXszZLrU
7xe9WGuAQv32W+nUkNZ52OLUoY5BlSBA9a/vf2VnZvZyrGYSrQQFe8mb/QNEm3QUyinalXDr6xij
54PHc/dbIiBnfNsauUWi+eQHOCcaChmRlk/Ef29qpRGebIM7kWDZiNn8Vd58OO1GLahQg1v5+C7O
zGE0AJ18Uz2DbgTzNMyFY9yD+SgnT4YUSyQbMvfpxyoC1ijJ/e0NwifFVJZg507lAOTXST4LAQFt
Yy8eGH+E9ENtaamsB71E06Wm0Fjqcc6MCdxcGRVQKSFFQniHV9QrvmVy84DqR3BDOp+yjtis2vhH
SjZYKv9diYc6Nm9icJEEOTlfUFV81WEosW2VPQQRM52rfOo8c8lWLIVd/emG57t9mUyYZFOPAOxm
tWGsHtgcFqwZXY8IYAsQWNesAbNaaGO7WBjTiL5ZpjUY39RTmDyfL5tptXbTN12Iu4HnfQQt2AoF
1JzZ1WaZrFuGt3/f2rUXFXpZXd2UnfTVsSIoyxxef++ow3NRdSMXSMWUEuLXVxkDcsjxMFjhBhak
3PH+Orjz9N/QTQEx2cl0SXumleX9AqAMA26h+txNQbiZRD/XuBKH8PN57Ye0Rg/9tOannsq2oEzI
hH85gRVvnuyGiXZ5Uv53X3F1UUhkRiNLHwdD3toKTYjlfDzkX2SuyIUJQZUdc/YlvfXiXUgRHKe2
CzLVuQx2Tig27XD3bYQuZbeag2zNR1Bd5qpDvkoQnn4YKhfIIdeMHv10/Sx0c86Jn2AbYfXFuP0X
jsng81oXZbLS7jUY7DKlgajfhhjqJTEXWD/KdRgVDHCW1Z4A6GT0OgyCU4LbIhO5csdLqXm8Fwc+
whfAgeGs8jNtOjB9+J31csBYnwBGB17Yk//sPRoiv2jRHGRV2u3qkPME8YcPWmAJh+V4NwKgjJ9a
sMo+WzMHpoEZiVmoBx1tv4W4tvcSVyUIl4cUj/VEjSpa/SqjiBeDrFpUYt/KhFZlPBQcS/HbRidr
IrV1yJdLK4GbFsAlTqyg1AM0uupJTgd3CYqPCrLlfmUdEnk495gUadofPHf+Q17X6eObVs63ahRG
ZiakqaBmJPsJxeMbSlr4i7sfbN9lr7egRP9zl7LQAFcuSR8W8xHeLO/SqDbeAihCy0mWX3toYmbC
iqRpzC0gVCOSzB5Z63TkFY6Wv+vT5qMrZ0JbOoB7WLoGUd2k3g7m7MDJaRj264pxaZH2ZFvGmMVw
k8/EHT69PuxlQwAmiqgbv0B4g19pZvxcrY3vyx9ccnlVDj8ewT9Pf5wmF01Yo0GugzAMopUXaLq4
toGX1ElISjrecFUVNHApWDLBFOJ4NKI1OpplFkQlRhTN1wKr6Xi6gi1cZ5EhKNNhzZzr+mxqW09M
lQRbwBYWJ9vJWLlikikCB9VL4Flsl3Fl/3X8gsOAfCpJ8luKLQsLXYR8uuLRwO6Nz3e4lvmVC/QA
n09pRFdGjcLF1kXNUi0RVyMqloo9adOXP2cMaVbsHhS9mxG3m0670cGwOEKQKbF4hjIoWUgIkpeb
NDKWg02Ba9LbDlQs866Mx4ntvP2NjFg5SfHltH1khSNsdbORXXq6t+/eiYhF1vLuEJNhCUKyFw2T
Yq6wfXb87Q1hLvUCAq4hTTA0pP/GtPAWJK4wvBliIewglLVa0AR9Zqf2radSQxsisA3eT6KIMAzm
IlIh7vV6mtdyXyzg5k3OstFQDaPEzPoRtm9amHO8mDUzDWW25K2ZdndKk/veRpcTWyGvsdu7dPBD
7Zc4AFcav3K8kvtj1SXm2SWCnO4kuw+8YWaiV7FzZtSJKLEW2BmyqLDytEp/DA7xKl0vpB3YT+KC
VTpMStKc7SHMcXlMQ0xMNEx4IQyPnjEjZfEHQwy7ZyfCMVu0qqFy32fFWZObgpLwHZQ/xxS1FRHr
4cus6Bb+nbQqVbwRXqK6qQuCdiMzrS1aSuPCh0zxfxZRKOclB5cB2y4+t1r2XYefRwdqz15GtHPv
z0VxxEGM9NB4eikV3zKqe1QohhEfZjeeJ8EfGdPhsoXsUNS/oui370howJZVL8Ntp5YPXC8iwT1u
5I7l4Lvt85DddphVQL2ybdbMjB4nz5jOW6oeezuxM5C3mBAu965hfS4yjytITqPB2cqAuu2OnjeY
GEixKCMALH4dO1kU/d4o1oODhJH4JYHFpdW9kTODRAh7cvE1CfOAtOgZ/iQbJQrwuDlCmPD4Wtob
ONXm7kAByiw7pMtIDsCos92eCiFiQoB1MjC4JxvdB0vd6vfBG/8eY/2iqxGe0AFXotwEcgeiJ3QA
iIvPcs/TL/QTrEE1IzyzTUHk5R2s97fcpIfY80wFjbRdY3qmyw9N1dcaEsYiAxsPm8k9RWiAX6ic
URelLxWtsq6X1O3gbEAjoeRip6BNmrdHLI3VYpbuWu3mAHN1lyJfpHHK2qteY4oao8rFGhV7cUcB
pRiT/FRY2R4czxQ2DRfPHVZfgBgWNlwO+at2jrWBDmUkik65bV0TOTNnLbnhMikT2e8qnu4wqEam
IaAw2F0pRd2owPqpQUoVYCxaHKI4dBvv7CC6ikU04JPyX1H+erhLmcVZ10JEw3vb81fBxR016L8l
M3yvS3LQ+RpHoH9dmpDTin9/hvtunecNWHLZnVbC2xvFTF5ueVQmkn9DS/+l0jTrazyQfQcvmk+Q
XozFLyphQ8zl8rBTyAOE3adJitz+Io5CMAeJ1vamwSGN5ARKuT98W82lmBcPmBcHdh8PhHNTvW/u
xCrYfOHmAqOnqaG70Jj3t0QX3Xq0nXcoFJEKBJgAcsJol19CSXJ2cLixqNxYjcCMc14z+XkvBMxi
LBh8SKG3xSpEE4zSSy1i02XFqbfLquHubnLLKYSQfCLgfmhuW0Pqoq6DN9jWb/Q4jXKQvA+0q828
nkHZUQwsqbAi5xOkCJRPir1LNCe25UIw5wyhiWeYlCGwb3YIw9Tb70trTmqxwiL7Y8u1dBOtfdrP
GaK559Xvyl/x3CaHlt6FEfra+ylWY08v98DcIDYL5lKi8FcaRqRgfj29iiBDtZqhcEiP+v66Y9zv
LYxP5rafYA4n8rH+WJSlhmrfBOSpcC9wQOB4cVxXMEUjIW8eq8I3Ug32vZ6H4nRYeJ8j/W5lBSUx
BS1Wj4uLurAgYm4KhE//u+zrNW8VtHqpxxfg84oTU3sPzLWMqXKgNwS7UiDaucaON4innYBORDZS
vLPdHjrpAt+kCUEkOvVQ/THpV0pR2bLnkO/lZnMRWCYzZa3ZaZqRV1WcxwyCDocnBy6ARFC12bqA
7LSGOTblW+8XYr9X/Zz6T9O0dzZ0hVjiShCivSiHd3CrXtfPl04/QVCse5etUVSx9BMabej0WEpd
rNvtq5hROlyXQDJ0KMrAeKoMuzgK1UqVTV4loGjnNi2TR6BSeSzegxCjxtRs1bcSOK0D6iNpnU8M
MbH6GoDsc9v2lyBEAYV1S7S95NLxpTnuxUd105yHXEFe5ia03YxwlCzD4I88uFIbdjBumD8Kt8gA
GlHeGsNwPrDDP6awHnFPSc/lSaKhlWg3va+tO0n+1/bwry9VFhkrSvW9QnETX4WzXZBW0mPjEd2x
7tHoRc9trmNvEEFqKGf+u8FmDU43Izh4el6nNG98jOxrbv0sItKA/TJhBur30Co4qBdIas1i64fU
40GKuapwB358bSdSkhOvJID51yr+j8qk8hv/h+rBuXYcrmYEjSZzAYn8k2glUAUlXGkDBZscjC8F
y/+glzcKxJuow7tXHauRxK+ZgMPnxWp7TzgvGB0DyfhnU5Y+Wb1dbSB0YP3Sq82Ab4Ut74dGGt3f
jH5OBlaAoEf9bM7dQeKTBrC6/m7C3VBAG9TSqjS2DZi64nKaUJvo9uB+3L3zU49nRhw3TgmGW33I
Knih8+K/FIWFV1gLVyPPSqN9wsDLMuAIaYvYqAHBWnSSqkA9emzsRW4cug+CbV+nWz4rNK5V13wJ
yucqEwN4/ImjHUaRhzCKhPeF/fvg8K/zjpscuPTzbMc8DEcUOeTcga3xp31O3jfdMIwun3kSGEOf
7y+w9E6gP2FVYbWfd6V8N0ZU8A1xPRUZFNKJlzHiExDpa+1BVM0nY5FTzvrHgpaC+cvXmm7H+gFK
xSca+1kj9YSMHYO4YXyOPSn7EagzFGmx/Sze4q4FQXmJE+Hj2gtgEtE4B7FovaslBFD7az9c8bOY
k55Q+C6NrfSzonYyGTBDqufeKENMZxSFyVQ5lHOTuzIWom0shK21lnfZmMZ5rsPV3RAu9KT11g+V
JfNoS1VtiLJ7dvbZZ1FE4S0TRHYcVGaNXEk4XUYhatioE5sr8YSnHZ9lQhNryJ3zB184yZvX7hyU
c4x/g3580ok+x/1J0qKXInSFZOushtxkNfUeEmykgERtRwbQ/IAEfNa74GQrZkqlu9rEpjPZxL58
YiQBtiDL8Lr6MBTeHCMwADdYeldVIHLpAXvVksPp+95h/yyefSzd6zMyb0O/HPKvYrFKqCdN/rBN
cl4AWA3Sn54LL2WnRqcZumTGr8Tpys8dxJm7Ayl8IkMVnOrkV+ZTTG5zST3BoSLGwYfhpGYSkMU8
XQbJP+yTTECQdxIqx1lNnNZF8wm2wzdHlUtVg8lR3Nu/QhI/2guDlGHBkNKqbFOmaxuV6kvmij84
coqqL20vS+J1d/wjmzJh9vsTKxJUb6uGja7GuDvgj7781OGbXncCrAUb4NFR2wHj7Lyj/QEMZGHk
gQ75MNszicEnSIrkqleXf8gnk280j+ZUWelV2ueHzGu4Ph64uuWbMVbG4NUp/TCM5inuMbvp+Mu6
GSqH6uLN8PoAKgtPgQSzaHXCXzvl1+wQdwKkcWfoAV4CNfz+Fi1p27hZEPB2uFWK2t6yzoCQwzz4
vbhypplWImFIFw5pQ8CiievvM58GvyDaqISI/JjS0OSgXpobqHhXI44WbJBieomW7N1KqHhoCKBU
II5ieR+v0tj82ExVVRBvAc2OW2yh8ePrRn9lHr0A6KTL4Dtmxh0u6gHViIpOMUGMd1l/Ium5q34B
the/6LAhdD2c7pV6GTdMOdcnxBi99w7ZgSipWd5soZ1lIjtKLFdLuUvjFB7eRaWIRFSO60+hVcbF
CSX6aPbI+BQyvFOs/4HOQFX1cM9aR35iVWN0gIBLwG7dfJTjE8Q82pZQd5OjqRta/X6Lt1YXqkXK
bz7AfpRvFrro9BjBfgw3ToJN8jnzlemDE6GZ0AhPQ3FaR5S5m7uPV65xgqz6L1JtOG5cFAyxtBF9
QH/1pwJMIiiH0eLmcym6wdZCcp0XrekhfFprT0aUnpPa/f+yu3KOTbIrvBbP8Ei/NMEfapkxfI6/
/uF+3fKlM9PDdUqtpYB+D0XQMcDN2nWsnqZvO9olCDOSSD7A5L5DdEyFALgPFHgQ1P/Q+Rmebi0n
CREEtjBx3MnGmzSn6+bPpkXJPDJtLwta6Ef+e6Utuk3A2rHTvcCjn7Sq6u0rmjywHI0r5aHC/boR
Wfle2DHE85zKMqSw7KhMxbwJZjHSSqeJgH621FYtVxva+bFSUhAN1fQRlOz0dDjV4f0jvAcPWm9H
MNdYyWFg0evkVD5skRGY3sKMMiaRW/wTucked25190IR4g/8waKzoStJB8xwqRWTzpSXkcnOxdEQ
umUdORdzkkqKlQWH5eLTcwaqTMSqQpQmnhEj+AVVUkigGWSWU/zndzX9SuTDzJsYCxixYGxBhxhs
hKKmL9BFcDj4UjbwFsk7jappyO2edj5gy64F/Nmr2gkAc+iV955AppRHvqtitu9rby1uqtgfpGlZ
ZSXZroTnD4j243Ulm2POJTrJ7eHAeZjO0GgGQYXbhKZS/MXULwpKzrIenOgjXY67Za5Che54D20i
ZMZ+66kxOMSYLICNvCK/x3xx01LJ16R1sKcKony/iC0Xl+XzA+m8Z+TOvtqIkAmUTF+uymgJrGWO
uMxvlGHH1k1Q1mjBytctx+9FLtgScGXXNL2VfprrR2RNwL0UXgZdeBh6ha0DIHT1cv3rGNk7+peJ
C1oy85gdBbJus8EnGqLxW2/XVepRgJxl4rqXxsjN45H4/bukdoSVA8XLPTtuLzdkSfsmWrWFktGQ
on1JrAmABJPHRcl2f7IUD98YwakhXnHgVanxht3YIdzC7r9LS5B8B1uxuKbCo9HDrIQSOCiE/urO
r27EeAuww9MfmnsFT9w4LLrYccZUfzO2UCFswVgnuUbPPnzpZV5deZlpXf5jIXEIxaoe79YiXOXq
LRY5n1MkmIYmZ7gaoSfKr9ODkwhOE8lrtFJb90OaD8lryGBItc5GogcYmtkmSd3OruY8ifLSXRrI
oPBbGlTGLlUCVgeqtO3WPZuOL8w2P/RX/BbmfTiiV1y04TUAcPHyWGlebxcJDzqTGkY7WBr2GlGS
KTEpINqlSbG3BDSQRJ5Wuj75mUBgARer0i/mBZqSkaE/FPBBcDNsVfknQoHcn9YA61I74L+mR3PZ
0uC988fVeuequ7wc9H7XFAlpQlJUkkzu6Tkrwnf7X0Xl1wDlLOItW0sxZ0A/NKpfSIfy/KM5G/OP
bKA9XUx3pXNvhqBli7Wdo0fUoV0tk41qPNJDkOgrzVa5SwqdHdi2dzl407QMTSDJ32akr0Ba9yq+
CvDES/OgUYpNCIK3AfuylbzMkfm+3/knvfhcK0i60PbSY6Td21shQZ8aYWjOQfgxXZMhTgs7AZuX
LqB+YrYp47TSEpz8SaWLLmDYo6Wb3M289aHPriLDQKQAHvEg+CPk1/Jqr5sCL8XofFbitI/wnM8n
TQKrcjS+2ZBfYQUOlEY+fyDlzkAMMtB2s7GBRhINTOghbPb8TuIc/6REDFgM66bEtz8vkN/mvdYm
ar1OUZQzXeZB/6/L3RW1MtcVQHjwGAZtMATsuN7MtuGbM2YoX7vLpm3oAfkqAhs/xgto+3IjO11d
aCRkP77wm824Dkk+sCQ7PEL0jckokoV56DgTHoZhjaCI0LpS7EXIY5gWUF7cvn/idwxR03wD+Z+4
AqL7HZwMQG4i3wxCVrIeX33toQrl7UpsZnUHI1F/vUPG2YKyvNdBNPkbyrTuQ1LPtYsyxdTs1a2A
jHq3xVjLrYg/EOtxRdumLSxmupWKcjI5RVLx+uBMvlw1o421mHE9zVKtTe75X35thq7lvgY/YsHe
zF/WzkNGuSRTrAPAt3YikCm/ciG1p3vi14oYBCX8zB8OTbRHeDYdLznf7VowOG3/cRO5Hw2AQgDL
O6CHZOtimrnd0RrC7Qup84GJZTnQxmpNvNKjyq2qtP8i03C8kKMEM/jrnG98MTnBAG3/7vvL6mM5
oAw50q1PQJFjxAnP02Z+N9uSydJ8YrzjAfceiiVKwi3XvgR6IVvRBtlL95+EJMP4x2O3SPwCAMGV
Y4uTMqyTpISxnkP8BOM3z5C9X70hzRj/qnW5qP1wJxtFh6rx/AK4TVQtlSZIo9hZ5BJH0fl4nvPc
omFg+QwIcc8FdlHneqCvG5dR5p1u9TWDpiJH6Nxiw/5qVFznz/pM8qVqmMYrQlbRJc5iSTW/EeGI
Cm/CNt615ms0tb71FMOd8qFhU+ymSQAy5kybNsrlthAndH/dqlyBrJM86ayRXXATMX46fAZe2qkO
oqrJGxPgDY5Tlr8Si0wzvphvQXOlwPIoAk3lI5K0qK6hfP7egVRMw59fE8nnebUoT8y1YbfnGb9a
3PD4TAOB7ogZcC9tk7E0r3gVHDbQm6hynLgKNBkT+7eFlz9W1Es1SXY9aBLD0613PsidA40ojnZ3
bhccUFa1WRQUtaLK4q5DPxxxLYO2T3P/R9F5N1KfdDUDqIpZg947iIO/CjBTHXSlVrTswKbIb+Gs
VG0Vh7WQrVysa7vntwpOENIaW7DzCDneDWTYIF33k20dEPJaY/9oO6uVSwzgnhfAFmkuqrIsEMqx
9AHcZVzGVEYvDyoAwMwEcer+PlNZQLN46HIOKe/6To+rn97gCXvEnlzfdfcETuxYbn8goHloaku7
zCjR5qTYgr6WAuHSdZ0Yau96dQE4XE3adPWcLmb1MRblE6852GIj8Z2b3TwipONHcyTFm+eajgsc
H0avrovBJAbORnr5zBNLNPiK42IuBUstksgA3QNuD1CQZkg4tifYw8J84qvTFpbx152JRx+rkiTA
k9ZJE3UQUAtDmvZr9ksx+I7gx3iAY4IqSz58hqawDC7PzgQj4n4ebKg1GPj5pYnvjnfeKAnA1sa6
oOyoCQcKJubHih3gDtXj5xEDJVHh80oHg7GLSBKF+YZhDm27SyqpIM9kU9Vkmd6XG2Yc0emvQ6a5
f1nQIrKV7Gz1BvVjr6SGx8R/4XZPaSvHPlBoEo1Xuu2eP9+iCXv7D6PcCY0rBI5KlxUYUDLIxzuF
I0QoBDCScJKjuhU2J8SSXNsV5bLgU9BCGTX+rFsTTfTQGzYKF23UjlVAZAlc1Y+saY5WBGkl326Y
eGkaQ2q1W99n8sozl+57urKsCvcbkmxmS8we4dtTEB/t4pynbTIqOIa6F/TDQfTp/rW9suRlPU/2
bvOyML+9sCAVYLZSPYE16Jb2/y36qLKHjCFxItUOnpIAS6PM2bI8GQg4j2Trvx4eOTwHrQycYto8
ZA6Oxw1lRW8onejJxxyOtmdNc5thEgWtO4DO6M37Gfjh5VhMNY7EnLUXpvTSPGZw9vyhKIm0ZeD7
qE4F5yGwSyMwarYU4NC7OzGib2QGoUhdthzP/ZkpuLthEZQ00udChAhug+1HZUsQW6rM0ML6rA2I
lsGeDhgZk0WjvYPq63QEkjvdjt5fi7RTDo8ns1qGmFpgby6XrtuWlcWxEyAW4Ncfoh3btQaUxI1q
T9D3RfxCSZYQg6KUO4CeqRK6jT7zTGMbs2DvvstZi1mtFSdp8WRmiwtJZ45CsHXDvR1vXL5IKCTc
EKZp1I5Lka1hNffoWjyRg5yydTV96A78nBHgfTZLQ8kwmV4m7w0bl2S73myWbJ72MwUDtHvKZcJ7
p7bx4z/Ec/f5zvQ8EBimpEG0LsYPMrakOrQluahxg+7AhufeUMI4x5up+Jga6MZyU6C1EHIImBt7
TyoxJ1P6XPRKUDdoprTGrn5AN+wEFryXIzeFQrcoVyAdd24qm7l4rOomIONXFdfW6brmJnx4biMF
FcIiYJite7adL+Z8GnSXaNUWoy+cvrVLun6ynNXu6bbOTxa/z86r9UKViklz7ab8oifPydgif5Xy
SsDfjq0WrvxDxa7xvDThDuXXL1ge7Vzlf3SHUpSSrS7CTDsjRuhsr4qOFt4+YCTrTcmW9E2OQM7h
ccmrOz3kBWEonS6+NHd1IBsr+Iu9FFEs3lBp+IIVWNTinm/iJW3lVEB3MpbUTRqg46gP0CMCZxeh
LRdl2hsari061VirHi1FDLFuXuWxn05ZaQAbUfX30RF6pWr88l/JdBo/1NvvORzELHX89nb+VnKB
G/6PFX/kxcVgf7g7GiT8mU/ipjeU3MhX+wVRVASpvkwttJuJSK0VJZqj1LCsj2Ek6OSplywBvMnn
lt1M6Me2RUIg0S8NhGeg9QRmZ7c7rXCW2IH6K+KquQOYM729sj8iU0fRQUqu+fkR29pPm8LwCSQq
oyykR48J/G8LHypuvZlIlWyjqv42zvT3r5AceFAF+3PAti0hWPOrpUvpD/+Ib4MXkBDJrRSdzaWG
WFg5uGknslikaEX0WWJSb67mrr0wAspRupZyGeNjcCgbUjWdTgmS3A66Jv3mcScZuEKGDpn4yrf7
ib+/G9UkkTW+L3aek1MtRfeZSa1EjW3eeJo9QFZ3tZI6XzuxHCeTlF7d1/Fw8EeFPKNhRKrLH35w
h8Lm+2azi56u0E3fjKqxlfN5TSkZ/OJ32XMSruahWToKbZhc3FPUvG2IPreqmJMoKhLjbee1TPyd
sZ9AuXP+Ygr5+APe4ufwy8CjBm8dnFURp77cq30+rSKPNDgTcnBoXH0lcm7v1mrQdUo6YqwFOObP
cAqSQOYrMYpTYUk7qHq99vSQXRf8Dt+nkaM5QP7iW+ahxmqsh1CGzvzqBn9umxMnR+IsaRCYACzL
tLlogbZwPBK5SsHAfk8pOiBu1+Aqn3ii6sfGZdp7kSLfmcUgDMYOvBmHapSQPkk385pzqxBcWZLz
ZaX2cg8Kyp0OdHLdCQqYH8ru3pnwthQfEeNgqz1hqARuO2F+7eRWKT2UfNIA2rnlNOcw0zAeUwk8
ngIKv9Y7sl1+FEzgMXZpFXBljUsv5bNny9CIMcNVULtfERJ2H5/Szf/eoHFDSbxnjBRkI1JMxjaw
AsdHuJr/zHRB/8Zaok7K4VUNfhR8KlHPvuhl07HhymVuBMaMphBrCR+OyO6usKyF4MoczSPtxpj2
s+7iZyOH18HpfkdrmTeLoubKUDcUpyTtJUbrAMgsWCBdFQJXw60ialVDxaTjDtMNDGtHBl0oRlmq
D1WgsKbCRvHTkntDPEf0FqodHCNetwyJWVLn98Wo1YH2lioAZ8o0qNGduoiFKffdRNHsu9vhZymF
OKuw47OwtmT6eLXT4v9BPahDrTxp+vYwXaNTM47aBVAZUeq3stZxXcI2jiJ9pyx6BpRym2+9epGN
X76wBkh1t/a5qrENzRdcVVbf2yHI0yz/uG1kEAC1q4sJmOMne6C9LmAcR3yTzzQgQO8ByS/FLChX
POXwYJkoms1h/NZjuBXDL+vsgG+x77zQzT69FQTekkhte7q6xcC2xrqOlfa2oK+X+n+rZHLedRzQ
5R34aZLyNe+tsMC447yGcRv5MTJFIqWCRYcQxG4TK4h0r9bTzenSLokdAu3blfyBTmTvdE1z84fX
wm0uWUkhXxUr0qQ2+dcg/If1LSjrXsVZ49bqLsiKOpkHtOwJE5pi8UQ8EfjWC6ilGwDJQD9dzRzg
ShinD2MQEJZakQpvUbCiRaojxIfrH/hvDXuG9ceczHurOfJHK2yry/DlX+3nrSyKO/E2IIPKlKr9
jgCK1WQ04Faaf78uy+5l6V/TyBOCBgduh11OQWFUDlLD0dRMXwfA4p474EXfDP1GcI3ZYUsxlGXB
s/U1jy7bgqSvH6S5CzNwnkoZ4061YRpX7auVHtRnI/abxwAx5HkNYK7oHG26AZ3955N9KXsP+Bek
oFTIuLVGXt8UcjhB0jT47thgAsiI/BJxeUBTxy7aVsXbqfH+OXgDu7dSIWekOVKMbV7lZIMoTAfw
F5eJ9LTab+6GmRmIhBoGBnxcvf7DbCOjiAEmRoVzQ5A7mqi99AAcbHLHV7sLufRKyeLaKFQupWoT
3XRqLLSg+CKn2GCFjo1MUGbGQN2S+6RIF8PYK1j9JkRRHx02hDT58X+Q1r8/I5576U/6oPwzy+Nx
4min8nCChMgHzW8qNxlRmqXV7Srzt6iV+/tzMqluFx55B/cJPT/EEGwopmzDStPRndvcDdB4NFg9
6Xz/cTn89KJ9ljN0cQNxMFNJrJorUx/sknhpcxL6lK9HSW5Q3r3axMrNppBNBpivdhuvutzk/ZZL
nKXGK6k/9COa8LPZT/heUg59ekYVs0b7+kD6JuhfyRe7ajOVaR/X8YSzbQzmEV6d3nZUekDBCk4u
r+H6/XDT+n2t23uArET7O+4nHVBpbJr97NY7/nFJfVNZnVCbLjWc1tQ79R9KhEt6so7NUd+8FFL7
nY15OGc0kMvyOVq/D+QUhI0h/Bea2a5ADj/14JaT5V+NVjnoHWqO7GGeyMrPmN4u36pW8nT29rMs
WpTSvamUWQraMX9bKnaTKRzSrUrd4sJxV3uxLyPpooXBAI6FsUHayWVP+e31zjWQW9k01jHVQmhu
0tiQQN5vGjdYph70WXHtlTFpVIuscCX7YfVWUcBnJHs8jDICLmJNlrLM9Fwfcwy1i6RJPUI2/ueA
WiNgaNrYJkOS1qFYlOvuReaBAHWC4bBXhQdFIEEbEBNJGmtU4ugjx5M9tbmUycYXKUFcxDYAvxFN
CITSaNliIk/nMaeXA/ai9J9scAmck34h4xke+GLd4G7hK2+2x07qRzAIapgk9URBJiVUdFk6CQ6X
r7pU+jvm4qw1RWbFPGJlJ7Cv8KTo6YCeruU/zVIxBJczi+UDV/ZwCLWHjzC3mWX+0NXBfvUm2LTO
vNM/nl8ZUTdhXh/Hd0ebqBcY42YNZ7l5TdJZsKbuPSsWVx/mT4GCy6DevE0/3SGRfnnqRWFneXBc
B/e1iZeG6ex7q/OKZc+zRetMeNnk0xtGmiqu2GYBTD7zowbZFIeYFX7n06fG5+sjFyfTTpSCGtwb
skygvu8IL/XDGcQXXiLYh5NK7yZLSS+dvJlh/Ix0SGtjWikTiz4DEppYKz+g30GhO7Sp/++GmmpC
W7xKYPdT4UuuJnOWUTVk81Z3UUZhHs/lHF0xnewPd9ssd1g6oC+eD4qb6Usr3R9AcWH4Z+MRzUbw
7oKvqmQMDYzTKXa4SW91IYJ0vMeMZMXnyo0yVx2azKa8gLd6Tn9SU5Y0qBrcA/5jZ0c4McjHkDsW
mtmGFcmSHnumoI/4lazfatKnoL6yC5By9KVJJEauvEbHU8If+0PEIUO7RKehF+i2YGNdN6yAQv3Z
mBrSM2RTI3ETod0bM67REchbq2PCiS4gMLUzxk1/0yRKX6GcYONoJt5ctgC31zD5DCwiaz6g97Wu
My4eaQMK8ondh27nXaybbDwBeuUF3LU3BCY8xRydqzkq09fksWJglCLYW5BBnBSOAYyF4SDc+KnH
auoErE3DWqUYNF74GEOV0NtPj4q3oxcyF+HvVPMs87ZLXsI1ejzhLLtfcnqE0xsYsdNwYgekDP8P
223hR+dNepj1TLGrAn1Vfx69HS11Wmp67QFBlKpcLq+CGq9W549xKi9qtzvGN9EscXyH4rF2Q7gK
9Ss7Kmovmx7Q7d1drV+nEdEaR9lJflSpzMR7Dk1Dc2N/jOpKRJwOABW3yLN7Ct1M8//pvQJNqDF2
kYIq+Fuf0aves92eChnn8zThSbu0jn7blcmuAC9oshkPv8Qw6qPyi9pkrJEsJjk39ry88OMEGDJ5
oeZ8GqndDAQhgpQT7zGjacIr9c3R/ooPbPqyg7aSZspM0ihr0yPz51+/N2Wp+AvM4cQf76J0doxt
eGuFvGJDxglW/jGBbzuYDCkwY2PninGwN9AVBn3OLkfWgiuKE2FG1upULZPQuo8Em9qzWywOhEwp
jdtcQQqQifl3FKcIU9LgyZozo0neBKtYmVfNKc2qrNsKTt/3jPXBmJfn8NI1ddW6etyzWfLN6SHO
WhwH9CgQlHN/u0Llw7gGv7B1q1yFwqxhdDWPjcouyGSo5GMOasqsyJvKXjbLbrAYaDNimZ8d1Z3S
ydKaCbhan3P7awA2OwyzOs0MuuzFtmJT6lnxhJd70Kh/0u5ZjA2FHkz2ZTczjlzeVtlhaSNG8tHu
KrTkGQHysdz/NlL7Hn3SdfFF5rX/E3lmg/uWkO+zcfBWGYZ0toleco0OXhnFKsm3k+3Kf/GZpsbj
1T9+ujxT1/8Vkx+uzP4IzW8ttMuml4U0RWBnSQBGc0GKlSiaMFt4NjXEnx6kkwLLDzutblXxayzc
K1PBdUVtuJ7JOLEOR64LL6rvJXewcIbilY+h8Xlt/z7jlCTTdA4O5YZS+TlLF3EEHE8r+bK+qZdz
eObpP0o1+No3hBgh1NChqu8oW8AHIPzyU4rZTtreLV2UnRFemSlEWK2/W7zixF0sJbCMVwdOiu+n
0ENzB5zmjAki5DoWsAggRgrdcVnvpAVq0lu03V7BWqIg50KNgPHJjH0dlJ7E5G/kpm80r6IJcZU7
Vnd0QThL4Sy09OI/AnBL0M07yvHiOWuNo4DOmL9JxKrbRW4si6Xp7zVhmC8qaYxVKKGhTFZ+vtKQ
Oqdk7+uhkWlBQrzJhaqkD5olbu8CkrCtB2whGFhJC1wLh4vPcoNuF1SdSGTSL5Teu+cOHV4RC6Di
/OZ594GiNBTMyRPZBqpoLyY7ttq7l/0xibLHoh80JG+IwNy/7hxSJ90OqalZ0efjTNm7LRptMtAt
ze5apc846y8D0+A9+DZbj5TSD9yreT3LMHi5LKcXH9UA0Yh4Q5gHhN1nIh8GJ8pvWm7rZl3jZOuV
T2wp+cUiCk3M4uS+bj/Jv+Z4cODgX4iknCkoKoO/EXwxUnYBRP+gWwhZ4TodKGa3FiuMJsIza8AQ
ciSQYYXw8ohW6oV63gXjdpM3wxXoMYv3rlcemk8/fHGGyYc/XBuI5SBXyD0uvsNmVrDwbfmgCdZN
RPAVPPYZfhLiRhrGzeeymxMjdtQzctaofZ+lelFN9dcVcgJn4wwSwqPoUKqb+1MAZNEKwHRDIwdt
HsFY83hNb1LpjEwm5NvKggxxzZE/7Mbjh88SMZywHEV/qDSJM9NuE3UydiqbY0kjALoUslJc0Qp2
oNAso8gDFECUMxT/X2DYlZctN9/xAexD5Sp/7VcqqOtvrujlsaQe2EgaoiFw4utif1GmD+nEsSGG
1Bybof+J+PQRwLx8PqHQzeFhgFzPTHdWpnf+p1Sk4TrrSMO8K6dJLZrkiNTUxSP10CVXtkYIbHGP
x21Bpfcl06APoxiOrcqVOZToHKI6MvucqJyGuusPTWjJtqPGOypKGaKFgknkWsTXKCnj2VKNVpbw
ZtMtkQOF/dfLY/eC/FKbD32+ILQAVPQzQ+k8KtQuO5dz87kHJz40gbGUFhK2pfBABhtBKp3eFBPo
Fk7ZqeJTNkw7bESM0MwIKnL4YUIohOH8d/gYAxY4wxupWYQihZwC6ZyO8nUBp3bQuJD5sKX+nRpD
ZbGY9N/0z4NmrWBbbQUjcSFd+3lw57UBQkyAmT/ptAv7zOjrI+KeiwrZhpQuwDXJ5FuqcKOyPSPC
UgB6pqIV2ldDb8f4KqNSIOikdZi4wYIhQAP5Spry6Cv98iuETck5Ue0UrOhgiaTmy8k0En7TmnsZ
KpJn52hjSDG6Pi6KXfK2sTfu+1b3xyz/jb959Kd/UfM/SNrzX7RRHz2n5zvoefnCvuSyPNG3BXhh
9sKlKNHFXZ+lUmqfySrf6v6olmo9pNPH8GyfaeD4Fc6gJBp/wX3iiK9p5Ff/SNaoXxOmuFkvEtNt
tg4AlUSxIqkWRUzB840cbOOWT+b/iNcWHtSwZR1g8M0S9N3huWw7Sdaf+4rpN6HXZV3CoCczZjmI
G5qkpSNDWv+d+FrhgO2Ew/X/6QMa+HAhxbliAjsybaysRhSM5cIJbLJxU/Q7pJrnRsxfoKwaE+Dv
lMl/6aqLaLBabXwTrrVDomdmBKkzDT9pbrbOvzNcrafRjWC6S/mbRm/YNa7uKdQGMDOjU57brFKg
s7b3chnez4IA3S+h8H7TKK+LYTyitXao/WEkQt9h9W5ci4zoIlsNZY5Qco8Uz07N55CCeMrDMZkd
wbvlfJtVu4cMf5tNIGcg/4cKlKpoNtpE/3Qncx7AiJo3xbPiOczcURmsFaKvmOJHApJRAk4sbIwK
xa+mmqQHKxEVCTlcZtP2iI9E+cNBHqsnD2W/qYDK40lUai7qVq3UlBLMaLwkmob449Zap5Kj++nf
2T5gI6zknmCRuxmuT/OlBendCEYeb4yBnYlDYyfh7Luo8P6ePeGr1hR6brVAsJBXZeGNfQ2HlJfl
oJ+Q4zmRN1b7DNoVNcq6P4g/S00BrAymlLxfcDxOPYz6ubfN/h1Y8gQS4sGzdUD6PjNi/8mGsqNA
nTVtcnMOLMwotTiXlJEESNu8kFVzt3YeM58Nhn3R+P8DrE8J81AQe6pCnKNOvvx9tK+jv/b8wHuj
bOASuG1PC5CrsvcTQ5G9t95Lo9qaihIkn7mwXLDIFc36K1b/2Sv5/WBcjnw8pLstHTBsjXvZdHMA
ZQ5R512/UYFMSuBx7RisMTmiRd3g00s59gs1I/GWVdWMsXdj5cdX3HQm/7hK+S6Xp47oK2Bp5Od6
toV0ChJhe4fI+tRvRZA+QxZAWyn6aD0fw3B4ZYYe0Su0/9vQwOr2AfmSk+ptx93bJkIjXIdoglX9
FY7kLR6TYQuNu8lZ1L/4Ai873nP4g+RvNGEJ0M1jXY1eE9unJ0D3SY6jmiIlTXXGy0ohOWM/OmO4
/IYbzI5K4T23nsMOW56JSVI7CEmJq7kNM5CwRhHEGHo2jRgLqVzXcjjYyUpAqEUwnZvCU1Vx2U/s
x+lUm3g7kQfn10bzm02zfFZmuoIASrJ2GyI9qWEhMm1PE+eMV/ftl4GmSVE2U7Au+Onh4OYFiC5D
Md6ItN5DRASA9y7QttDkvY3yFpcAnET5YkZcKVy4++cIfde0Q+79gks6/wBJvWORfRFxaTxuCcXI
CnbAEbo9JT+So8esWYIOIZoXf+48lwNwtWHEneTgMhGmhEcT/AAy/S8kcq6G+SIRGGp7oQel6fvT
WT5VjKESNO8oNtMgAFT1/nhvAbGi9EF8ci7UaKhO0XqMDWhWwuvQGSUwJtgdPqweZtGcpfIFDN7D
KZ8W/UkLS+ICOriF0+8Fsunb5HkZrnGFji25ScU1waTLnbSEHnXdXkOP14Bmxxdlys4mimsX1tmp
vORJSz7JWnwyVaRlN8PIxbc2v6OhtPXQ7DguzyFPlQgYw6IH/77E9gAXPi1hhhHT9QzN+lonXt2f
YLGb/StpX9YByJwLPX2DRbowzW7zDeQk8xMESvzdyknZ6pyoE5z/5rmVRNhFhN5ZBzswMUFUaVDx
OFUsLD92VdT3WAhhcUZHZpzMZG/mslwyCzeJgF8+zRFlD2h85XafXDQtgiWxE5z6MOt9Crrgq+O5
of3o/wbuBxnWzv6m6pM6UbbLDf5splNNatebL1m95Lpak/N39t8Qk4gHhkZLwGOI8D4bxxCaljYL
XmyPyYFb9RKHehCWu8/reUQcwCV4xvkWd0xN6dQue2B6lgGPR5LoiqbAj2dNeKRmd0d6Rs/y9wzC
1sV/SojMDweUNi8bZN4eQzPdXyS7tXOmVWd55biBuoMHqNU9ooPkIMO0DoY/CFFI628B3ORZxTfe
1VcX52wGllJTIRczlRHJcUhtxckBK+n5aD70Mvs/iaGjo799Kgu9JSNzDWuWFXYvokG8i7jd7ShF
UhaqIH6J67kYVeh+9s+3Etd3s2pfk1yKHmcCqmvLK11p02Y4R9GB98rMYwHhh2HPwipkl1wUqbkJ
hJVcQo/cdeUsaEMKvstJSyjyUzZo6REQrDmSOnuXliQcTFJUWb5K7XLwQ/qHolMB9eytcPDfCjZ6
KeH4Er5NhwOCnOuLQzLCTEWAUSgOCxvu/Bu2NFqmYE5gYPIgH78C5yxLSo29vVRLuJ5mrV+p4/Cm
3CnWZIkwDTl2qSDq3NBR6O+Vzc7n31mMDLDFJb9RxDRNCKlxTMwRmsiDmQQe1QgzmIW90W+o+DyY
d1U/0NAJnoQ+GoPDd8nhG3S48ExhVV2754ri+UuPSO2VLlV7ntOjRqkC8qj2x/Dh91caGKGOhiYY
oiT2VG6VeKBUoxkA9b/Df54yl21FlNu0iyfUU+T2gCeIRQ4beS3UV7K29wIwvvjh0wZqRkNSlogX
CeTIPJ8TQSZZ3/H8F41I9yZ1xIA5uqXyrm5xxc0zaiHNRO3m78b4PmnA2NvFnTs6mHgoU+Wws2h9
3/JFAd4RPzVf8ZtYPDjQAXZeI2KAR3B/OCI06c95Yn0gYJ0Ysdd7lSAMRdl3bqqc9WvTMd/7gq+k
5uodHpTtuoUZ3mOP9wGsQLs0TrN+GKImTpYU6sfJL/8dyroSfhipPSuibgtO/eMC67PSZsKUkKri
Lb4gz0t+Cc08Wc7oqZVITWnRGQSykPEv9/OIiAf1OH4M+EgrOmwSfNk09IlQECugiWm1dKE7jXzi
xWxJG5Pu9JEcWQ/77Knd0kIAw6ZsL6X1ziyGM+VNH7kJ3FOdFT8bcmj7x+qJ2yvVMkbmR349IVPA
ZhmBJrIj8nJdA7FagQHMQesTDg4wmbSe0Ugwa2upqOC7Drgf3DvD73wAVi70Gw3+ZOUVgmlblmxX
ktaopbPaIEjDFGig2mMNyztNM4vmNQglM7JUQetoq6yYBBtGs9zmNMTSXDxvghVjB2LTOJ6M6rwX
Ilrvxx5TiBMmaMTiaK1nFUupwAVq9U4mbJpcdy8gY88LlZZdbFR1SZDqOEU/2ipOJJzkK2bmTejz
KTc+Qb4QSf0uWWNIE9WhKJGyC7jIP+wBu3V651Ln2S/UtkEytkWoUiF9rguN4xFxLeEBhTh5OwIm
lV2khRDvjZwLi66olivOl0aeJQrI+Iz9uKcZpdfSDpLod1ohFv64hJDnP8fA9Lmct+41WeKbJMEA
Ti5P+qSiBsMGv4M+p2/ckp+MA3B+AZWgT8iRCAL8hSJsMA37K6IgptTP71wunbEKgZsrFybB8zWE
eo04FRKl3VLnAO0dHJAtlKBcrCisnyARR7jpcd2cr0cLsIClBqDxAXwHm8zyoeTMZuwIJG7/ViXg
o7t8WX5QCj/xb67ec3lDICMzJ3C3YqSew/s7J1V2She3DPLAspFuw3IImnVHRmjjO/cDELQK5VsU
rsIRpooTNx8yAn/XNfw6HwHkcyRPOIeywvXZslq/3iDcmZ+Ad433lsIywe6FOabf9mXd1Xm0MW9D
d71ufNnSGTHQC869CIzoFjA+wPR3BaaeYJFkZzX8F9WjOlrln/2gKdKIbPvbzUEw1SqG/FheWQmm
QiyCtcwZzJ1gBrs1sL2T5F5lyuy+IqitQov2I/I8qttYZeZL9w2spIctwR4GZ6i8YyFfig/p2Iul
6pKAy/8CiHcWYPcl8UwkKLg6cMKj/fqX3cyrsQTs+2+08eh0CX3v5lNVejplB78ayBxcMY+N9Kpd
ffnrN+YKtAkRslBL6V35h3ID8k536zgGsQXDZrmOgMge/0SV/f/eR9kxcuqrpsMMnMVWjV2OCiMG
7lB6SyqG7jdsgVaJsSC4bXbI2NuiNYxWEfAAUrtzTX53eEQhk+ESrv/0HdLqU4hGBEIUf89TOGgf
ywpE/30I6awQ4xAoBzf6TxHZgSLp9xgJ4HC+lKL1JPUIeGoLGWR1OP9nKPwMbM7rYMKIQ/0dg0bP
1xY9dQ1iMluq8BA/ZJrXyg7nWensKbXh3ihHtoNsOBHnjPkwMt5fuhIvyxZinZoITSsH34nkdqht
ruXVPJ5IVDlodtLxzLoBiRBv+BCEUjpRVMkpeoufxg7fi/6q5qzOuBE+tN71ayQ0XCrLmWJnWopl
lp/Wi2cbWPMNfY0EoXy28DXNQx+OEmMLkTGiPQkTsTG1KID5ny45ppLDQQgrJaR4QvGJG85X7Jz1
judUfsgXOvvjxnDasemWglFcMFcAlzMlhsFndIFhP+1wr2dRr3wKRN9qmjYCyFaDo/FwAvXiamCe
cxHR5i3FZJDRS/HnKevDjU51C9jPl0n+6xBuxr9XrkLIH/rtDEmjvwh9/Hry6g/IIrkVyucqrhGD
2JEbw1dhC9UBUZvNQ4T5CgyTiWaYqhXNyKdoLoXlxQJZrrSUQ0s0yoJLc4e4eNTk/Pd2NuRi0vPZ
39ivPcHW8EqwYI4aSAdJIdkjpnwcA6k5NujpBdDhKNpxw5j5k9E/149HnpSboz+YO69ztfZUPrJW
p2TxeSFEjy7v0HG5NH9NC8s8RRoP1Yood5kq110zSP3iBekvYvHjm6xZ4706rkQADxctmvNPtIy2
ur+Gue6kzoRGqIu5GTUusoLOAGvLhvdUSeJYZwNoWlwuvPhAKJdIMkwOxt7RpgfWLJ0/jeuQjpru
rSR/q3P6qLQHKaizjImCjhqoahrTXZWU6dPbxWm0PrCYt4A1qF81zkYKmuLemXWRqMPtOp6QbtWb
eQrOpiVIK1SV5UuYuQv+eCqG4XsBOCok/mHXAD1YgI/+y/cBN/DMyfcNW4D1Sj17Tz6XJRVGpEV0
ZDDTFS135mGdx3Th2Sgi/Q/+MCY32EwMBfzz42CCfX+O5SoCJAqsVpnGABqCr1R4dLHtlQ/9Qi7g
2jYRJjZNTt+T3kvTXWS7gne39SFCNAtO89fUpVusSg23GkBmr0jwh1Laqp0Le3292g+fcZo0u0gC
JmY8aQBxVO9JRigGSMvrLastyYojzBU9DACCZ77T2Ld+Z6J2r9nZDeNdMFzbhmYk+Kdcje1isJ2E
0cl9EEPeBOAb5iFGZq7flb7XxPK3jDqrtubGH7t4xmChJIqEelp9RZ9wcEf8Um4qOQPAlblzxVUA
/4B3gtNe1CnYQ2+VMh3ljV9G8EcEdCcoPKDA6zXFtGkVqKlizaD0aiYB0AW1ur5fmkfSZ5kaOjGa
drtMN3JdqK1QaxdYJ99X5LD030KxvIxr8TFTWHMruqf1ycY3yjA/2YyDefzpRioTG4eNKoK7yKKm
DNtAnsQy/HIG5nasGImiPANBAd7IeuirE3wqBp27CCau+CL6ONzopeMzMXi+gI2nRpCV0gK8dsNl
ZknDc5D8FDe2PZg61xYPM7dtf8j6DaQzXpAlqA4SzJhBcB7hT07WqFNA6ATWhdufaijBf3wvtGz3
MCD+tEqnHW6QbnCoAxcbozcUV2jhbT0Ny3aO2Y29XXPROxhhtJrL2r5aE3dALqN/bAmLGQfPmuh2
Bbx0JaMi5+PJ5ivfAzt+76KE/wibfJ6XE7JRR21bKxA+J+tCyzrZF7EzqN5Yaaym+deARJrUQMFr
Ndc6uuzmEr4ZCWwYcolJaUR47M4wW1H7pmrm8BsDe8TN5WH7ULyrRCCl5RnH3QllZWifeJEhK/Tc
CourAMQH0HJm2Yi3GDRigeceK2PlBE+C7K+yLLozD9a7gmVUwfd2Ks9U7SsxMCsaH6NKbBtNfFXK
p8GrSubkHSHUjEVX63mPB1UIFdPJvVcoRW0uY9W899EUyR0fqL/iBXzwQTkeGHJxsEyAIKGAxEj9
7gI868CXQkKY7PRdlPTVXnABb/vreBLqxCmmLjA3A+8vs7ylPm9FrRapFB9LJVzPnKF2A6+Y4Uet
9LGtFkSRR826RySQb+EsUxT9PlbgWvYVDhcyJ79ZHV2h/541mBR6Icm4wiZEv+KCVRMONOJAO31q
r25oEKZB0oe8ss7O5fWQpUqBnG1PX7JQArl4U0HiDOPnyWKKQ2dZcmF/gvWKdBdN4uHj8n0cmmTb
wh/4OGA5QRmPoreMqm7au4yCZga+AcIc6XcGpUt8OXU3CUNQID2QGMFI9J+pEMg3B8XgbPMOz9vB
Z4dw4VQJEi2O5D6ng1UIPzgXqOZDlKYItCzCDcFl0e/Fz+nAIedc9x3WX5GBEwfTJdkTX+fwL/d/
5QzeWPU6qeVGYDC/fOwqJoc3hz6Vt6CeeJLgpy1DosTlc+/DLSWEokakRP1EoqFvEnfQRvv+ql33
Jac83mWWiiuvqaXRXD7Dlc2/UCDgCYkMseJsmcAJJ2IGvlT2LyrUjFAl70LLIMfYlU1FRvencA6I
BwBb7M3NQ0xb6s+uWjEyy6nWtcWN90Y+i9UmUFDvUwY8ju++n25qroJfoII8plAQs73YndRPuuZ9
ZmYQmVU7CSucpzpwfLzhpMcD0GVx+h/TAPKYGZvdwuifA4qSEGupap0Y3G6CqIIFAWL3zGBlDHI+
64cLi20OYlnAuIif12kGJZQvCMuWDGhFQgtD/ghKe64ez+x0Y5BAsWmDDFx6ViCBxjrbbzK2o9KG
Rm57D5lcmmafaQe+DloAwMsB/Oke/WslBu39WXTYE4ysR4WQXGXy2VFYU/E1xenjrzTi1XomrOVw
MH3+RaelImPBTGd2PruOFvmGFjB8ovZytWJFZpX4lQL8bvfBORM0T1dCt80yoPYds3SrZatrpG4S
2xqbpNHJwYplJLtkGYts1fmVnMNQE0JETVYUgUOuS1fi7KCkyoeSfa2o18kCmpIOtMhZgz4LYe4V
0Ar57Jh7e6dIuszvC86V18fxn7Ims7hj97AY3Zhr0IqJRjst9n24APrbHMEipVivmNpm6zA0lAvQ
Sys9G5ZB1qvsFYFPiVNLpfrWbGzHpQdk3tEkb4yJGK+lyx5WSo9XaoIhNDZexxuzxq7rzZ3McrSq
EVNAg3px84ToXAWENz9Hps8uCMFFtzhLDXAND9c0teJHpM11XD/kbidZgLHxixwnYmI0828TcH7R
F77+mVZ/c1LpPby9GGe0lLfjksrp1bmOCDV3ZzmDyMsDys3N4KyLU+f2v5EJVvobW8D/DnD1pTdS
R8IbUJ+Qjv2ic1bbjORoIipEkMaef6rqbndi7qrsuCsMivYU77rWOnBwKKQXc4R6tWmEqs+5/F0o
j0WYJ5WoGOriOtMVmZULE0BSB11cHYZ5yLs0i0G81VYpYBM0FDFxJsH6bQS2EQD5RFrUuC29QwkT
D7O3NL0IdORw7Dz0ks+TCDVGX/GOUo2RB4eOQ8d7WyE7fOy7zMARQfggHUtStdki7220om6JXTxY
XW4hlNUtLALryR1m88n/M//rgx/9sPyHTvfIxWNjCkxoJzyLc7yWzjTPWICEWb6ssPwCgeUi9Yox
JZmjbWSv68RrvBeFSmSn+oo8pNSddY8geCRdXyBGKgFObXd9mDOvrwMcopj5CUGwsBlrgzVG6htr
MqvW3vtq/bmLch8NN+l9Da2M6UaPSpT0PzhYdthkWuJ3Lgn/PTy/kF41h2WGPaQi9JLahDb+3jqv
o3br15dv5KUabxeUIPS+PgUowrWuDhVTTDrLdTHhJEoXSVBLFcrTcYNTeLPIfKs/IInvT/JVm2cU
M8FW6A73CXyIGJ46oWFXgSPF4yxBt3XoSZluBMda38aJNpXG6pBE09tLfvMXdMu6KXDRZaFW9ix4
HZzbwurZ3LtizTvq2mEU7N+oXJpFcMiXVE5O6j4yZnanL4zZ4q582q88PTDTVGOijwth97mhPpun
6DPSzPRvkSDzVcHzxEUJ0a3aNQokWrZNjyzTVddIqnHxI2l8cAi4krMvMBVa7LA+2yCoz0jKtPEq
nGBGfj2M1tf8a/wjKh18p1bpT0kKnKucjY9S3/Dp+XO8HqDVk0AsbyACORpcqLjWN78RfaELST+1
TtsQ9MX9Yl1MtaoHnEEWuyc8IgEptSru4gT83w8mqDcjih1ts4MttknbhfcEeOtE2pdocRlL9nEA
SnFFqLLAEOgde+UQG1ukMrCRCug+5tEb9fV89WMcqKi4kpAd+Kh8/0fmdqF7N7sbdsa+n/15luWq
EwHWttW6Gb3SE2NTqPBDffxwJwgLUxW9YxEionaAC8zI5e4IvnKUWjy5KtHJWr5ymcBiAR+j1Yrj
OAp1N6TasDKEtDoKG8BqdTGsMY0gMNcYLacryenJgkWzG2SlTxuCKNZ3sqtwFpQ8uPFHCL1n57XE
9tP3puflSIIAgSS0CYffzToXKcdVv5NnD/KZv6fWTr5Gd1EICm1eXtnL2AhmU4ywCtZ2DjCSac13
Jo+Jo+755GMmanjf7z+R+W0vBBIEG5tfTqd1q5iZS1TAEkSLaTm8BcALWMb27f1omn2RyMuwdPh1
LvVDsEAUd0JQ5LLGic6wJcgIROA4fLlRBVkcTHjk+lt5N/I9uz7dTBYGzNAPgxsvpJn6LTcxLxmh
sfjL2VMI7YcM6aApNWXcJ64XgOT3KHrdwt6d/iT5bORiso0Tg5Fqc1X3A+EFDdDCh2WucI73Q6zR
gOFzZ+IF7d1uYHYnkNOeox/gsnsBaprp1g0d2VUZPwQrldkoPevQooZbgbb+2U511MWtDlRBzOFj
MdjNM5lzdIKccf/pen2+anC8oSnzqUTVbhEXMCxVOKJSOyKbt2dvtWmxYxyKBg2BxRFiBZ+li2f+
d9po7hl50TYWseaFEmncE3WwVfgOR35dKOP7h/pbZ+KIeOtLFQ5q+I6aZVCMNXaequD306A/PZYy
mIaJ5IbClWmNlkOPHMN0BoI0thB8IZt3M3CkBmF7Nr6ZqybJ6Iia3lLE0BYZd8MVap92tgReOElC
q/0NSSRP3jKvjZarwFyRx1iN+ESPg6mx4w20vX9bHOtyzIN3MKztTV5Dw+PgLYIdlXMHMgG2De2a
8Hl4pXX2iuj+cXqSOOWZYL8MLhg0CjQZ3X/7IwpCXvuQwHZiID8k5pLXuqgLz96zAp+03vwqg++d
Ki/d9YKE8FmihKF454SGfQTikty7gGSbn77uIXy+lDB39kKfyjctxm8qWmwz7uCeIqbt+bWYHpB7
gTuTy+tTtyB80bhV1BD4NZkxhwLM16KdQXeNF9ekdPF33XPvFyZZ6We4LWmg4roo3y/pe+hGKkZ0
UkcvTCcDV8HFEOrkCoAGO4SKI3bN293jouGY41UwammyCbb3BuzbFL7BunlSousJvOf8Ne7V5ue5
wKioRJxRFLR9hs5jCm7gW+r3dDBWHLj5BdTxly53KIrCfJMVAODyw9BiieYvXV8HHzWCqFl16Ctj
mzo9TaEH3XuTGimx/e7SyVyemX5WgESXkpGCFGOQ/VPg044m53YHrmo9O82sBOXnle4WBsMpbdfL
ZNsBgJNx0ewH07fBamR++74tsS/EN+lRWTZAyJAwZDYEqS0prYPTfr/eibQjUHzLvipqFymB2+3x
iNrur6ixJJwc1Qsg6PHIlyDR+Q5CCAeZHCw2lLmhwvyMZsLWBr3XWa8WRFGzgw63fEJBh0mdWBIe
2+mbGL0hqxHqcJXtBsk3+WRkXITgmGaER8TViWkqvgYsNC8jAlopcmJGFmT5l+H9Wm/oJY6tnTTa
flO1ZPw0eD7o+QVJ69Wz+miq040Kg0QGI9FFFUieMznbW5xq1FgGRpJ5BLZiQ1/oqyPvqK/sYDsL
+P6Nt79oj59z8Q/eYKGrDXYyPsq21xOhUtMbir5Wto3H9tSC2SylNcRP81NMQ+N5TowYVjSO10kN
ROBGHc1ZkiKat/8tKmNpqj1JxQH/QHFs742RVGGDytr9a1xlYYnxlEc4FVbm9guYvaKAGSf3zVjI
Aao+2bzIaJf5bVSUaoiA0UcJg0eD+pjDPodrH554APBaUyo3tXhI6R9y4gIbFBG3PQKCOTvqRq1G
w7Z95+MLD0LMJLbDOOdF6GQJ98Rc6l38F6y9lp+1b1T0v0s1JVgyEoUtzYbnckzS/TcU62K+Ppa0
zXdaxkaY/6ODtHRZ2G7CgpUSQG+7wV+p5Gu6R2XKe9p2+pFh+iej4m1Mfx2cc0LxQIavDWx8HvJz
Ni4lAW4K7AAebWaqL0al/+VpFEdxxhx1xSjrbj3WqKGQzlFByQC4iuEqiD6nbPLRLx/FhAGdYELc
5CvyfBe9x0eCNVtjJYK4Q/p0ffv+VwdJe8zopgldbozMTpDBK1EGBt/yjq1cu4reiiUVAwMn4Ntp
xn43G4B7wwy4fIMhLhZuRhokMtIWtiTgg6rPXYXlxxjcBKiBRE763sJrMbtpnbsCpSHlp6wz4fZA
OZgiZKMGSS3m+txVpeqK7cYjMnNQlJ4AcGlNciwRR/JwnMTOkuuR90n6SBYJNbmVeI05AAhAb+b0
3FHemj77uLzKMGmR9v0IKXsBUZiUsBYuBrfT85hfXB+Jon6UOATaUR8ZpsvB//l3LSliJssMLQk+
JARh7TraXsnX7G+hg7kHIvro52SJaJgoAH0es03im/n+/EASZkf4iDVg9I8yBX++jL7WqYTF5MAI
6/v1+oNs6Ry0wkNvg5suezEDSylWjVaH857qku72tETAAMijnn1CjhUXRPI1ZsPu2oCbCdOokl0Q
rfnVzuwcPCxbao06ogFU++Raez0Da8c0+GJ20E+gMc9b23F66YK1hRrwVRMMn9L9PAszy6y1ef+x
DZx4Y8evTZA/IPw+esmAUuEu89RVEVHAiR8qYU9uXHVO3PBhDwJL692q/Z72cfUPzrFOcZjJqoRy
rnZaisBEz5961IXRPfEMNN7NufjLELNYeiY8BMD+Bqn5myXvSB8spxKirA1DVcO+tq++YeJN2uLM
UwrEJtZOhFq7VjFivt/JFuJBERvmYMiGvT32rOA6z3zEOb4H+Xss24mO5L4f3spOOw10n6JHtQv4
U4kx923ZOekFi+0eHMkh4z8Tvdce0OOf2Kk5s0SY0rEciL4B7HfastyvWN+2T3klChPV5/69q5lf
HGWHATHgJEW5PsTVaCCr3xko09XfCx2J5Pg7OSHYBvJG/l97C/+l341GSFPNIW02OXDbSWT6dOeF
aYeBCJHzeBHatI7Xef3e8ProbEYyf6cwdUWSvQ0bAlMHlNftf9UMy07nBzh34aNouaTLyPoIZIV+
PnyewyJDcgnoSKyuzxJtdwfdDWzXieKa25Aqw6s4JY3VQm2MfO2Snq/Tq2AH2P0sUsgOUVlQqhIF
hbjD8G7uTndmor7QCY4Nmau1Frb/heOwC0D3DcN5/Zvf8PFtyD+OGotEtsd7Nx26hGoynv+nrqRP
vM47bktZ8tE8KNBRUgT+V1ZDgyyFRyh/B/FAUBMG+ZA+i6wV4jkwkQub8Ze30p/Qzmv4rhNTMCZX
kal0OlzXMNkWOkJeq69L2x0AhTF5f3JJDb55oY33AdsUlXVf1rAIPkyRNDAc/ttFESGR582usrnS
bOfNeQExiAPcLOK+/5oSzYn3pHbWhfxqaOJplJ7tOC6C5VWl6l/5OY+ZY8SIXlUBJliHo6zM9yS9
VsUkKCp7QhEGKi8GJiLlh5XuxDB4XwZk3eB9U1zTslPAsNeTti1BjoVG/KWERNdNRY5JiPEE75Me
MnofdT8DEhx+n68taeEoJWgWc88/vaEu1oY4a2hTLZYqVeTpSX3RDe2zCorUD486SlpsgJnpWLKa
1WymNG9PilPS5Lyb8moVosvku9dcSnG3CtIvekUQ37cxOj86yf+hOdmNYQu1CG2ouZuPmKWI4oAZ
OZmN4jSx2JMnFm1vGxhqQID2VXdwDjvE6pVlQ/hikeCzHg1b6RXxVvwsgpmZLCziU7JxwkxatwJZ
He/a1pC/kPuTJaRCSP1o54gJZi9DNVqSb+gBG3o+ga21QwyIMEyLBRrL9LSMn8OTgZeo28XeG9aH
EyRVJs3utnjmEBAQjbMADlZ/Q0Ew2pfTK4w8/cXyxuBtZ78dGQxGVO+cPm0o1Ca4AsIGo3zwtLsZ
MYA+Cfm4Bt/MlE4Jc/dm57ciWEfzOIXZLoIxHC+iNFF5g2gzTZEo6bxuc+bOtSHY7vakuQ/XPJ0P
0XMpy3t1rf3NOPvDj8SdQITeoAcbBQB6QbUKNWuxpAIHH7iCLcvsxrZAF74QnE/roXO+LA9bW3QW
g5H6aHM5BCTU2SBA931bb5G+LynuI3aWCunvLzqy5OeVRau3VqNU51/761NFBZi/OEInfJNJxPDD
+sB+lp41A6G84ks/nZr9p1ukGQU1Cp1rLLx/Od3xaH+/NSglIBiWVoJpwL4MccZcJ0awWIEt0oMk
8FTbf2XmsWQYOaeBEqTtVCAGAM/N9c9ATjRe4jmw1ty/f+QpMib6q0h1QriG4hORMOjx4UmhBfCE
pRP0m/amAazuORAaIJYLop6aFTVwAgtbl8IpmV9CSOqKHXaDqRL95FiNxB+QiBDQPHMFhZ8mYSib
RbA/mHfdPrts4iK4/RDnybNmrEsrLkveWrw6CYCf9SkSQf02u6wTA5nTADFZmSLZNo8UjvyPXQdq
1wyGvgfqCnpcTrHI8kNky1cBDliszVvQ33RG0BRBWrt/Ys9BL5/Zocv3tfV+Ow5s/qHRCLozPLyC
L4Y61+yHHQ1UCQ0NeqWzVEdVtmSOUq7O6oWe4KdW5SOF9u7AwNHYbNfKc5yocfFwntL+H+Gqwbhu
W19c6q9PiCgwd57Wv2haeCxhI4pqL81Vqm1aUDa62Vd/BISavm977Wttmptw0ySapGCFmHglIfmk
xImH5GXIVfZ+4e5PsTQmEpdRt7i0CxpBN8ot+O8b+58sFDQrUwoJHwMnkkVbo8OUcCEmB6WOA8Jn
ZmeLqoILNgjDwcDwdvnM/nKvpailNni4Z+2JRB90hr/s3NvgJyZOoqM/mE9QyYLz4rhogsvP6dtJ
cPVh9lLlAZ1FscOLp4s5ppfpSv30JzQVS5DobmII6MCS/ZrGN37NJCGJ7ey9k4BEZrgMbF9UnoIW
yM7v5m7mxj9ui81yQms1G8F31/852uXi4slMzcVQ5EjuHJadyvcTwCOt+ucqxqsJDbYWxysp5dC8
zlk40MlKtBPt0loQ9ffbm89GoufX5VaUudkPav/Cg7hhG42Z5Bp15VV/3wURGyYpvTK0mRBwBECO
VonYiHOK4ImC/zjc/cZg9hKrF7Evq4ezumaC8AEQq/4pmXy7lZ/DGKOectFda2JosT9Pok0FVng+
h2qBM9/bOYl1/2LUjWQn/2yeBjMee3FMx2nWOJB9PUkrL6bEzfb/c4eX/CSDd5g0kQZN46jn8ctm
0Q3BeLSk8aKN2UsQ4dgv3kXCBafhHmwcGTe3dAaYouluAMU96cW/+5JB3odR5gvSVCPrWihdUGH5
FHEuuJpG7u1NQNc1AlR85jsmPTyS7V1bkkvxhOIjWGKFVZYQfvEFbNQ2BUDEgf9wd+5byYQRcJEU
KUe+m/ELVB/Vy2xi3cKHnBbmkTT0f0f/ACVgypGvTjsQuAieBlFxTsx9oetYk58DvSYK7kJwkPA0
2UQnLtg8easdtX3lHhOQnYDsS8OyZqIr/8MfULMRHfi1Z/yxjz6cVGuankpMYyDr0qlavXeRgJT5
wtxM4/gvbdcdo3O1BLzEBVKjNQD1AaVbpNRvSQ8JkWEomOuiZihIPG4rrgHClD026ypq2Z3xKzfy
QUw3idSsAupmLODk7ebB7QyIFWjxlGFW6PyIjtNtL0j2HgzyE5m9XZbf2QSOpiQUX0QfAfgLYWES
y8fAIXMa5ZMSsgf241a8/uSWUxV+d/QqCnvs/PL24AcmnLxCWWSEVZrze3z9MpzPYxcd32/aFfdX
jyyNybIUn/QT45bAl8tnCAiSCPSQueImYCxPECTTPl/jbGWLYZMCFMlFRFjrNROE/AnFFPYZ7SX9
kKhBRMIuBd8IeCo6JOIPRcA5HSE6NgSskPBA8Scx0pwz6j9P40dpUu2uhArcWqMbwz/Y7jJSozhV
1ODy+R+FkBEE+ciO/3/0CXcPP+oU3TXw1B+N1eyJH6WWkY1veK9YLmIW7U/V77w8B5uvZK8ewl0u
otr+7nVZW35EmtsxL24feFyIJzL5058jNaUlYW8OrTvF6iDBQDvhd37916j4913LnVDDvZ4FQcGq
U/9Bdeb+1/zLCGT4DZzjnIKX857a2zIdvV75T78yLEk7EF+JDQ6WkkKfJvvVLcf3KVWOelfqJswz
L648mleQWVhqyKEr9b1pimOomuwJt6W1Q1BByB6LVWKjqGdbCPFMi3Unu7cOYk7Hyt9wgcRYdjz2
MkW7tqTwD9Oy2ZR9OkyBNxgkmASeLH0z1Q5RyhRGOdq2VYMqrpOro5kSNqDh2mLy2O5LVDDruE6c
D2Lx/kUocwz0XK8BRhYJyT1C0xMw/qK8F3s6QB9Znjjvi9hEdEXZVWvvWw9JeaGhUb7jf7W1M5iQ
nIt9FKrMs3MjPou7WzBCAeHTQ5ZTeOQ/E6UJDXcOOGmEW+eGxsdNrjQYL12yiM7Ll354bY9KPWjX
p9tjktuYlldlSRdh2KCKaKftd9J9avsbF7fdOnL/78dfypeb41Dm0o+l8La6ZMf1AdXdOXAPdfxi
4OkFJAohPblwWZ0K0Y6tOHRQm/R86X08wE6QLZ9HKg6OEFEhav0/slzZMzFwiY+1mG7uSgQlvB1F
2f2L/9a1HHaicPGUfS/5rJQG6RAk3BAuJYQxzoJOStCM1KPaGycomMKXVHwhW7CRuJ1Wey5Sre9a
NySsxNpCGEHILKE4kYkFH08V3cfUWCtv+aIxnZL7SCWEqreOgaE/+o60V7E11a+qJfW2l8RlTKCg
ckbnmY/Mp1GyFkcc9kY2R/m1cWf21IGp7qmFlRKPgSv8aizW80czwimsdI+hRfkUjPMErUMW2zLD
B19/JnHR0cRB4fBwPMrfZ84wPOFS4cf2iOkqQoGi1WdVvx/3q2qzF66ET2mI2pZry0i0St7et0BZ
6QHOusFg0QO1SXiYRv6HsmbOmFYSRBK8sFZm82mpSxkiAvAkl3cs3Pww184ZBGRq71nB36E6BJje
YeQNq261EyMy3JjGwbQHO39FOTqnF0+IwcTJb3+H/hTackPpyaMOrVc77gVYGn/Mu3RD0hX6ySJ6
y7H2d8kNzYgVkVBj7VsxF1FldkjnMTz/a6s1tO43EM/R5MGuUiu6H5AR7RKTw6R69qqQAzqg9f1O
uXqrxnuqbF0c8lPYQ5jVzdcTlpR5xFf54o5JxfYdd9b6+hXPDZ8/pbx7RAtYSBAzW/cXXxcHzHsB
o0aSaVo+D5Kt0Y4fTudSFX4SAy9/OMz+1FSHoNzdQEFmC/kT82S4NiCAJqKOf5SRiY4W4SjSxy1n
QBN6cCqW400N8Ty/LAYSj/Tm9bvu7pkKrh3cJ3O2tNG+WJlAxEzUVVZbpAbz2b8qx2QO+uDkGvbp
cg/hBjLO924mKR619lnHY40J0ZRmiw4cxcKpKgcmUIL2v8w+lUxrWLYaouiFUuDi6juDCfVy8PPi
lhIPwLJz4xep4JP/M/dkWKQNJfDPJLf/kcd5ZNUaveWVcytVqyZnec4NEVes28c8ur6d+mViocT2
fDRmIu8Q+5SLFeL8RrOa8AixyKzkgEtJmWkjGFnNWOL9ghIPnyZPHdzB8Lq1ig78b+14IW0dl4g7
lReyaXCwdPbYXHhE+le8beLq+8fFBip6VcDVum2Bgu/NhueccOvMvEUNEGYqdXvDcVARyj9b4RpV
GpfZ1cg6Bre5mZlH/gJGj+T4oFWJAMuLRP7it9+U1Q86EpUYIWWG5Ui8SZIEGw70gwFjNZutmmJQ
17eRpyBjuLgpZileLggaYn6rmXHIaqz2bE8uboF2ueNsSOT/x7VwgLAjAcfqgvBV1wdeTJgi1lXZ
74FKSlqvTM2++zIQVY/Vx5DblhZ0LxszaJAwKw9UtvbJlBjSOeHorf+QxKOwgm24R4FjFCh0tpD1
L7vt9dVr5WHCIrtuxtQL3pgZhJvwVY0FL0L5XeTmqd/QUj/J93puUuJTlxK/4mF839ORWv73Qo/U
uNSsnsnSmgXECcFc8uTm7YoxH2X6V0/2J29CSivZzfoq1oOPlIvcaiwi2LZYkwrX2RCw29ILnyDT
2zE++WFKhyq6pnGFbx+SS9LCV/A7jcFVUjrxKQKeqdJR02BzNOqDSAP/MozeStu394ZfDZfCLzXd
vVPhKp6mFthrpl48L+5IFoUHu8h4o/bNyhw2JoRdKpvNmu6E6ZQjFAVDZBO75Qrvq3Y1uwfac1LE
Qpx4KQx3oLvO3V/USmR/0iJbLsl8jAfrwy4dMo+1IFr8trG7PKywaNil3LxIKVhjftb2DaVT07SN
fpRfxbp/fr5bMvzqVnTBmFUnOGSrHV585O9GiK22tEzNVkv6YRrGyIDhFFY3gdc7sa4e0tzQ/MGz
HQz+x5OSkQ4oxdUlYcF3yoKXiI/BrAndIai8JL8et5FrFfphhG0RukgR36FF3GgTYiBaY8BBu1I9
IlLr+8hJwJs27MI8o5vXShkD4/rzSkWOsNKI3v2dyCcHBmFT2MS+5USTyXA6/Itv97u2xia5vLnw
HcbrEZ9pQEg70QB0WWMx48w8GtCavgtdwa/gjbBEuWBmNCtl1RO8Tx/TqOn38kMW5TGQvCLaR6ax
JQXqJGJju3gQCnIQHdKphazhkiU5Hqmc+ycoZk5Yl1xdIPGQXFcUj5L+kwGygRN/6cIBQQ4djM8d
wY+loA1b+VbbJFFOU39+C/boSEnoZabg4Uvpg2ejn6BPs+ZpAbtSShe6636+7Bdb7g8pfs8unJFE
38lTulVQk36mtjUxBeFFnK8/VwnH02G10TkBVPmwLnsHixaw+bkDwVeT/wirmXDFNxATGUmd+/oG
D3ye44U7rH8P+o06116FMhSBMvRZHO5hW8wbn60utHr/IGE8VGN0MGL8ns4Xyr0w7/XUitaYfu20
NoHZMlBO+3nf4grD6tdNBIJIhqiQZBtD0nWNKEfSkYm8neZ97jH0Nt2HjocZTk29QtiYoFCPYedc
80Me5lp/I24Co84AnPd14hWGj/71+bMm/AOdiF7ZBd0bAUoN1jwzuGfhXFAvjaU9qBXUUYtYQWCZ
am98QaIeNmqTEEF9w3N6yMgwo3ZFF8mJ0WKr5eb3qpbXZPj6sbmWEhLHqmsFuBhXX+Bq2sPV3p5J
AKFh3KYhKlGxPYnsM34O7ZepvtYxT7MOJ5WMxm/tYX1W4BH9a++CtLiUW3gbR4Cm7kyYdXTW/SkC
sJdMrvPsR8Yxq8XY7Sk9Jd/r7O2gTe7vCzFuzNqlZ3sRlvUXBSbrz7ysMMX8gsWPgMz51FdX9CyD
u2g6qwwARapWlCrGT0gnfX3TbN63mjQkbEIqLxrajCrWW25+008Z8+DjBemoIn7LK2y4ETOQ8NJe
n8F82pN6bmxzTXBU2XvkO5V30k6NFJo31eC7tZH1J4CnpDisETp/pKGxh14mzeY14fGBvCrw+W7Z
vtdP8E2CgfjyyhAei3t6/nK9TDhudUr5vVJguBB6VNF+Y7u3XJqIw6icxOT/FU0Kob6GO+SoHhWL
qXsehZQHbljhk8DXiqw4pC3S1krl4lMhqjWBQeoToUuGlhVPdKQ0egt44xLPUequK6BvVy4Gem8N
xDTmQebUuPuMBJ3ceROze5iBs0qMx3OziDY1PIjhjeP/JXdtXvQyw44wYTPN/Pj6HX27kg6V6Scp
y3fUw1TGv9SxCwqjoAPOYqBkaLbqlZ52AU0WX6RQeEwN1VEpT/MQD1a+51getb/PFM8irgvLCXw0
c2I9pCEs9b6K/YVZBg6t58YItLmAZjY1ILO9nSwbaMI53wNs2GekSJSXxgf6SuU2nhivgt0eEY05
cH+GHomo2l2fzVnSjRoUURJMfQ0SxuCC4/hQquAzK5BDbY4okaIHALQFWA/VK6kBemPuIDiIQdzL
5p2Jqod4Jin/YnIJpe7syrO5DAZ5yb7qNz9kOOmWq8xzEbD/gGgOTLT/h53hL2xg7bCGhQ2TNn6w
gP48QDRPInOjDJDaA4CtLkQeID9b0dmzvwfDqCoWqP6HYLFlfeaWvNFLd+1CbQRr+IfP+fyXtNnv
MQ1UAhbcKu5VX2zfVYrRQiCDfilci69YgRcMsA65pToIH6OyPHqrIy1GFkXiUs54MzkMegmfrqf0
LiVqbgX78efboL7Yni/YxdUuUCQ+851hJ/eZfWp/EHkZugiNVl+3LGII9t1igdNgDnqS3hrJk4wX
ZtFJDQgz46yz+fmTA3Sw1iLVX98rqwuskebMrGTRuXgsfwqZOksyTnNEGtCTAQEm8cJmSLOS8oA5
aYhvvuqwQy46t/qUgfKDi//xRf9vjEZGGB0xPENPJau1YMDBKhMdvbQgPK8NhifXLjnWwA+3ezuM
SoisBf7mtAWUatKldy7kO4b59ugv9GUFLMYFllOYntJahN41n8k5DK41wnDpxDsqbfJsdjopgLHl
sfnd7gkpN9Nkn6OcX/pK+t4K/8zxbfvcVHWPFhqtfRNkEp/hY9V7BgEmR0UYNE3QlYMapXBnP4aZ
ha0IzTltFDq8RMwyPruFKTlsGHpE22r0R2+eBGZ3H18pl/pfm5w9/5Dw8sLjVACuRsmTcRtsGrRA
/+4GFOm5y4wciODCoDVf8BFV8/WXIYUMUru1/v+Ueyg3KVKjmMaEgk6PteOkXQhGgJXpFHEuZOat
wEV2KpptXHFiyHY+9ZpRYhI/3Xm3hG5VSdvrjEzp+uOwP9ORtEYYpkro7GdVvbn2zff+zreOX3a3
ZGqmeleVDm2Llkk5eH42Szq1qqwAzJ0+yPgZKDiCXABM/a5nFiMUKWHZ4lYAODdNWbi/V2ebw60j
+fVhpVEKwmbLeY98DT+yPVT8UYPOhgEYPxOJG393Tb5hRo1QCcv3sD7mfKYVmRGmAIYD7vpv45Xv
l5Gfs/P0DiA7cwre8PbV1hM6/GISgIBPl5VNQlGQaWM1hvvlpasBQwxRDpU04rLwBjSIlzovsr5R
K3tg6Wb6M9+AUNXKZcD8SxM4L2F0ykJmJn7cNbF/mbzKY2+ub7OhYm0swBxaTZsVmde9YuHqdPcL
dNnnDCJ54pDMlDMONe/EECYbMbRGHlh6b4JNgHVotTB8cBz53lMPWHbfAro1sLKGfHut78caIqQP
2KHHga1WCgefrFvVDauKqUtJuMOUNYZmxdELGD87KOimT6103CE/SeGGZzwjM7Sp50PA3Dt7pjU9
ni9tcCk8G2PN72fPh6/VZd8UiXrLbcbMYjIicbZDjZN4cx09REdO6wbhT4iQxv8qWu1sq+Sjs33q
GO0X0oDjaTxZBhztIfwhvWOQOkF1MID9Zf+5YlgkbaLm4cq5Sk7S0BiGa51C6FepT4GX8qiDB/07
/6xdkjR87+rpnUNxSLJ0sMEvwV6UOf3gdYRK20vk8yvctGFVtElQOycPJ3NNBvzWqvg1pjKU/pN4
nD84cbBYUY86nYkqCUpbPFXgx2SMNVwLViyVMihQWkfAweKPH2axrHAGvGxGAcHKiaGMGY0MbyyL
jLzCkwvD+trTQROo3CF7kIKQLZWVcEZ5Ht6s6q1VG7qkxyo5dLAgCih7HNeOzaNMEOoHC2l7J3rg
8er1SzRRX/9RH297wVurtMwrhM9e3DSlT7tITOMu9AzTtpZCbzaDSrZJF2+HX5DWi/NkwB7hOupj
/J+61UozqfPC9/Vj2uA2KPf/sjLsdqSjnMI2rjfXEEYtyP/AulhYPYQR+2uNZaCuy6H+flyesXvg
TMI3ism6Act4+sFpYBH3wb+h+TCie99iNevBqyOQs8hlrMiWWqOZEw/qfa4smkMdA2dESwBMkpRb
HdheB2YRhk/CoK1D8O51QiJxrPTVBA39MBy65SfO7chndon1MGPtzcm7Xi7QAViMND1yausxvy3x
ltvGLc2dhO4nI2fNKCBq4sgpVBQCQ5K7hxdJAF/NgXVTf6pINEliWjOHQwY/mWjbhqlcoW4q38gq
aNaVzIK/Hqgbgy8GqlMgcFH9wvyabLQHD+qc7U9ccGX2/ayXUopuBLb35l1SF0NDxpV6d8DB0us5
7p1g3PB3rcmYfBslB9ICN3AfXqbHH4wJRjkDL7hjpk1OBVFa9SKSjuJJIaSRdkCoPZYmPlbACnrn
HILCF18zzIKWzPAF3CYpldxalA/fLpDCg54nv19MyO2cnALEadjfXd4eCs+OR0DVi3P0dYzPEzbB
x0TD541wo56QpJbPk08F2RCBX5268xCmPgHFJbRcLdJTA/tJ93PEOnKwjbHpNKgOtV6SrfYCMhkf
kRj/a6h5fodYfewfD977NM9a/tjnKxHYP8xaYvtdJrN/IEyxm0YeI0fh255DMfTHjN7sE3Fwo0lS
TpBR8A5Qe1+THRZxcoR/F4mPrp2VVddKyaISctyeY8e/3pXoO4ERBBIkHL2zvz4Uk74NrXm6rxn2
M4Ok+XBRVsfjz/t/G7ND3Hs6sqWTrOQVtOTf9iYhP3kb9YHqWE7acXiis2MeA3b1ZgZfbLjR+xAU
w0S88LmL7+JTCRHN5fswipxUts3c+dlQA6ZaRhit3awHaYWFPHjr/xbMD56NQccsTgV9IDQ4UBjn
I9WO/hrSafG7iV/wRQbbKxEEj/EgbVb7XKMF9bS+vNbCQkO/sreulZKcNthO5qtR+0jY12/8ph9W
H5xyMKzwG2ShovCl6vtOuLND3wMdS9D5W/uxFm0eUnsTNs95cun/X8DVxez5cMa/GIcxd/4sgayj
NRyv9CE5InsZO6jsgXl0zZYi93tjYyvdd/NXCbOzflv2UOISMhUa+a6KRbyAvsvP7PsdE8iZzBqd
r7Q890WXqSEim2a+OG/E0rBjnkLSPLJlqw+SzBM92jPLOoCmI1ce7Qh7I/5gv4NlmFRp8q72RR6D
C1tdKoqUuxGClMGvljetf7UHyQnRHWCiJh3ltZHLWi/cjLvgTVRI8YnMkOknK+Vgaym+4UG8AR4H
PtSgy16IgyymtdAZ282Ynvw/u3zXtEvw1MVSk4xJVAC7G9u7roARvg7Tp/h3Csz9cxfPpX2r1Joq
cRuTrKbZPbz5xtfNqjm5s/BHEWaRnRgPIIHRUDLBzWJ96guV3VHwQnkwneApi9tYPAHfhpxjbJ0i
9YnDncNOtG0hpQTX6k+lD6mDiyhT4KiaYSZ12rrrR0tY49+X6kpZw2NSfXQ/tRvWis6h6eh9hHtU
f9URqwjWQM8Gyc5NvbE954ZYiZY0nBuidNFhHrl1N+wBjPV2A5oEvg/818xKAIRFM0BibP1XYkaJ
SdeJineYvJB/SBtzuBKXKF4yxT6kwHv0nUrCTxPHiPbCKFSfabXWljsDTj7tptcL/7Uineimt192
wtWFyLhw5wOFWy0+xUhBQ9yMfXMUqJ8QUtlsIwzC1LOW76vljDGw3xaEGvZqNBpqDKQUyKNS7r0U
X9NBuUd9HxhFQkydT41XagKdFJO+AsA/j6wAQ6wGlJnoTecgfuw+bpOl8xIzSrwJT4w6Oy0P61fT
H7XOT9a3uqC0z9mxhVMJFQEpaPXgkgwd+Jsm6eIy1twf1YJtq5tuhlloeTGZ1c3OjhYi5vacKn4Q
dL0yBF0IvOZNQ3yCQMGrMZcvzbycFROxGHfhvohcw2tDG7ybucQk80X2SlqU7c5CxWR06aoomxvP
L89PTlE0/nKCUfz+Q9YDL+I/50O9YL2BVNh36YXyiNdN5+1VyN7Hzs5ixRv7P365uCwbWrCeBBYq
8VQXtcFzDhRAofVg+JDSrfaze3faHwNqzpCpz10VEfeP0fqNMTmsFBD03qdZPK41AhmTsiq8rYan
uhKEe1BIOyloeaNFXLvuNi5HxEnuav0sSMDcOddpvE6rKQ+LXZ/A+NJOpUM95UXrWMXQIz0Z4wna
LgLSJvP76bjlrS3cEnPE1kzoslmonwjJ+t3jfDeyaHoxeo9qhkFvjXr5XJFvGH5/d9vIBjtd3F7l
pn62Hrd38G9rm06JOpPqWacl6YVTTtHf2tg5eDUuwWNoh526OejW0qB3YHiEJbH+fb7cVPX7YqHx
hvo0LJ4xw+nC7xSD5nC4nWR2wc7zyUWbVq/baO0WjIS43BY4nv90vWQSMcouMtA/lLeW1afUs9aE
fjvl6neFrgRPQ7aMa6bH8C8ljjEJubLl8SRSL1Rto8roLHgx9V4AXPbSUKyGvVbZefaEfdvryRCV
0TD5anK+Jgpm+H7hw4xvFkAq6d4JZViD+DsEJuNeeRRTVuAgdi3L8jgfWXVY43zUXxacMVLZEvAu
XMcaeTdXsH5b3OzxursFz8YxlVaa/Hbr8NA/N4/q6EVmcSNX6LfHYgSqgd5nLyQpTfsiiwv31Nmv
7kJZmcQ0iT6vuFuNGrRp/NAYbfsaLw9S0FYm6uoBUONBLQurbx8lvpHzRDLZzgDuzSPtCkbqbXaZ
s5rv+VWLiy8PrjIR5ASNrFWUw1sSEcl9f/iOtzgF93BMWr+WK8Fd3YvWIfUjEPNzw7Sjl8gXYWXE
4Td+0UBDb5cVw4E2tvp6OqHk7QOYTob3dpxr8JMXwAX5voaaXxavfjUmYbobUxRPTl2ccQfIaavq
Xn8j1who9ezbrjLKjkGUcdd7QOlrBJ1PuuJwG8GmAsqeI9ueKttwei4tSyCPmJTfT/mzRAo7arIz
I6uzleYayLSr5lYT3gApjbU7e+4LoB+lLQU0Ym5BdZzIJeqQp3dy1ErTbGv3xLWsIpXO0n2mFT6y
bt0R9IUIxQiGOFNUW7oMGHdSZvkc34uYqX9OWHvPb6ducFDo11X7HZK0nvoIGFyCriPhOXaw3K3F
Oxh0s152UpN+NuuP/ecY/DZl0k8J1doe7Xj6/g+1ZFE/aGks7NoL/Kw1l4MPq6C9pM0/15Afbyw1
rv77KHmlhrxZbfNmzGrP/T4npfFsxnkaoR2PuRHfD6jHEshnNtmsQaFWxwrM9NrBUPw4WgIg+hCK
k6xbCVwgxJQpXom7SHtYSymQfXOjSfPmQ7fW/GPUFo95S+yZRVgWzY04U/LatDgiY6IO9o4j3sQ4
OnwUQDuFtuzVTNLWOFHo+XZuK000Qi927KQPOrkQFdzBBQyysLKm1QXRna46F5Rg5FxovWwWN4VZ
i8qE9JQsqCWS/MVz149ySJOimov4jvHFQEmKV+3x2Rln6YbZ86aY0TkabIuwoqR0OoyX9gAmskCc
JU6k0nHCtYGnb13CRT+8EPuIR3R3AgIpn3i3R3/qgztvjIFnh6RMHPF2uvsfhFFj9Fq2guRKR8EO
l3i8QzsMlgtnucpPRcXWEXYjL9DnBDThmT0RcHWMceaimZerLprV6evp9eM7Wx5upbTypf72amRW
5rA/Mqw3qSZDrbH6+qfI8avkjUoXk+Xg1fSKcn2XfunIa5cdiNJRWcHeZUQSTTwTZAgir/yoQCjv
xVPRr/wh5SaL3MFvySNsZrKrAL2n+i3rD7EFdNMb/R672DQjWxaMy4OPwNXGAMW04u2U1m4gLf+0
3KaY2PFUIbaWvgILNZW8HbQfY9v99UnvjZyGSl1yEqZq+iasly0ZA89UO1HpKpbaqdCof1E+5DhE
xvVTnq2TeRkDA2s7+jWhAkmhAjwSNCReDhEsxVX3KEtcTLkmj5meRxsu0ZSr4fpUBFXjHNktvvnZ
AvF5heVbETlyO1dg151WLSMBvd8x9okmrb2XSE8VViJuffCo00M2lY6DaPH7WwWvjbxDiNizpjT2
bzhTIAM0PwhkI/oLjOHhZvYfFgyVrU/6BIOYjVId+CMOmck4B2pHxSejO3PpslqrfLgYOSfgm5CV
11kYsLnLHDVxBexDspnQBC4avdQo8m/Ai3LpuVuIqsPrxyZcWRpXC2vmhEDoLmc4+GFrZx2fMOIj
gHU23cd/YadVN9spcH+8zFvARWaBkgMDdiCpzTakET/h6S8E3Q5aSyHv5OBTl5YHHvMqz9/K22jm
2f/CqQRalX6AQ9+k/v+XFfjUmxWiJNvSd2SD3OsOGZ/Oe4hm1ZMC3zQtMnis/x8p5jPJdQBToNYM
UTANFpNKhU5LfgcGNA9MrpLGD4Ot9OMIgqBPe08fFhoPEGzLZ1K8FvVf/UKx8WI//UV6xwVOyupt
0rBZJFwgUEGVdwwsG6ytrpKzd5e8CSu153Sq6cE0Hs8DwZFuqiXJTzfFGh5+tZ1KBdd+z8Z8e7SD
2nKJpG51uTpWKThx1H9rZCc/cmPuaR0iMUZhnOBbShvu/ef8SC1A3obtXO4XdL2u3VpRi+xikncf
1Ef9E9QKjogDB3zy7h4N7YjRHlor/HKflWC6TaZS7+PYQyH1iBiAfoPXjO+xPA4ChJ7CnPWfMo7K
jWKFa1++ms7MvWbvB8W2DZ7EfXmOHLNdp4syn3a689XTe1d4EQpkTJUDHh/8cat6folOl4sEtI0L
fuQ6w/gcsGmF4iU8zJQYWTcSs6Ek6XrkqBLS/49lmCC67cMHc8LVFOCOlICcY/D34KppU9z56l9+
vkbdHRqBMWufYjj5HmAN64Nbv5f0zcxLiRHfGcNoKcRaxfrikKK2lYN3p3jBDEzR/syuaKKGYKP5
Hl0yAd/JomYvswE+CmdulVQXyZ1OBF2LEtdFPOmf4z5/t3d0fOLpXc17sVLEAQlSkeM2wEX1XqsJ
hqTZOfBXToj/l+6dQZk3EoRNOi5BFyHza6QBPmlZDDYZ8paHzKfA+c6NbxY9LSqsiiLpzEtNSYRy
WQyytWV5XCXr0VWG6jdOLuD0UusGE5LogM+f8zepWV7dGnPgOaWpXEouo94QLXvtZV0dklXcJWyz
wthf8tzmwh20gU7e+ytmLYnJpvfLcoxKrPF7lDRNh7D9bJ+PFIgKMFHns2uysx73STD+UxnpSvfc
XYKUK/a5rgHuF3mYCL99WEJs957TwEj9Q0gn1YuoEEQhhSNOhpP28n28mMdKf9AGcvoETD7ZN9Wt
moJS4X6QbbWxPkH0fnnfMgA0XohfsgXcXh8tthEbpZRE2yGmWeLHCXJSM/WhrAPe2XUNIEbamKAp
Dh3KEatGOd4jgT5wyVq9aCoyALjeOXl0XInYU4BP8Op2Opmp63SRO0VSl3plUqFt/hIW69116eLa
/TSB18YAOI1Ni9N6rgGqPjJsJbpZwJb9HzFVqLkfE3WLzl6oHDGwkrGH7N9NG13Nn0OkqFE+pDwy
rFaWwPxxL734engBoTH3A+pfixOiyYZyzMe5M3FfUYx/J58i8uSqc8qfR3l9o72dyzyhoFVz34nM
Rhzxy8ntjROOOtRpywjNM+WKs15U21+MhItN2+fyIquI23HL79NbgMf0O8Ly7kZL6WuKTAaLgSJv
aAlysW9vZIcMn7lL59nulntd7X2DnZ0O/bEzo1v5XRgA8EBErhJJkv3gjPEXGdvrvnnWBZHwTEE3
gPCMCS91VJwxoDgL4QE0HfzlhEYhXbo0iU+jKMr4VUFrX5RgIN2XW6Vbwrl+3aAgLHPWkyNcmXze
fQaLOFa3wFTvfSUKTw7aO16hcgxXe/YYCGe4GtCPWxGwhaBaecwnYqRlRM7KdMnCdII2lu/sTdPu
OHJGqkSTwYLZh1+eEDHGQHyOH0/9TqgccJ4FIgr1itD6b2q1mJLKvlbv/G3E/HAkC+HUhAKGvPpm
H1B3BTFnFDalYdOUeVlvCfu2NJCDpTNvefHwrul4Ioa35EmCUx3eY16x/90XjFDOdcvwAsnzvcEb
/x+u7sxM5M+xH4vfnjHPOseETSr8I2/F9uMnr2W1CL3n5YBmGJ6h+BUbqRM4rWKRpbAO9yBZI2Is
0r6MMAgPjplzhV0T3utDpLYCEg6QNd0F/jIC/RSRwh7gO1Ow5XXRi2ABttcH5jQIlahio1qZVKyB
B0UJmfWx5V+Qqfo+LxtUJLz9lTwxr/Q5VzxSFJHBU0dTcbnchwqUDfF3X1GBRAqdtw1euIwoyYXu
LiDp/sXuwV1zcR0zuKIrMQR5nWhztzO1/MxJxpVU136sZKEG3lUw2ustNbQUzOc7DomjqsPYSPLs
G1JIwPej6sg2T+uWwonTPOEcZcyRmM0NxkZFVmPQxkN5/97sbhA5TN4cvaZDcQ+cJhLfHp0X5lRW
bGhTd8IbPecrvMsj1pLp5g+cQLYF59Sn9UL4jaaesOa+jnRzpu/duqv0/XcYorgzBLGb9Jrl0Ekh
z4331fBOKmWnixZ1YfLewyf+0R5mwTNlBfgODPqxXd6MKitWA9E4ubXgApgCOcFh3EZVRHyiGxZr
sQTcSqcS/429Mv1sVyzyjd0ByshMVZiaLgx9JK6OE2TOzfKxZpehS3/XsFsKs+p42Ul3y+bQrwGK
oAZLIPFuCiyF15qDFNd7c2CTiMrtZfH+ct+zMpn53yxpZMoJT0hj8/TsJ7bVq1RhRbnMtD443MQ5
C8LxG8WoETLYQjH787Af15ToI2aYHmiyv2FE/oSVUPoJ/5M3sh1+SE8l8laVAHrMXUZXn2UjWH5D
n2O9sUKuXVkCazx0rEcOvvrKuhdkmv7T6UcvxbrU7f8QddXtCdvDIlWDS+XXV/oDcIy2AvZWI+PL
9pyjcDRx/ms2kpAQUm7P4ZmLqiU3oVJ/tYZjgmaOEAApAVAIjB3G+pgpMvMx7C1CfDgFKloN0sad
3Q9OJ63zubgpSTQa3Rck2rMpeM9AMmk1ugas7RveGtu8T1rdg+R9Ec7frxuSkyMhmMAC1CHBiaro
5hDiiUZOVGv0hS/zuVuzSfjBzhk7N/Uw3bTF/fhMsIO5asmSzNzxAi1RqWwixd0BeKzUi7DfRlT9
czssyXudpUoJi3Qxphp3cH80nKMfCJaK7cHL0iDFm/cjHUw/mnyHR7jPmWhrZKAW4zPPvyIH30bZ
rg39OP7siIJtINcm/lptvUqJuYPIRdbZlS00nKQ2KHi94yN/9qMsx7SKDpUCD+S4dK/y/OuL53hb
6heZ+OEUBqPhNDD67fWEctJ90WtzSabLaFahzhub0olV1xnOPLq6SgCp9esfUrM2Am5WSOcze88o
Hv6oBKs+TK5eJEw0ZigonaPjOk+SCVBqHen+cJNS5bFFpDdxj1Qc6bdu4Ul4cgtrGjFIXjf5VJ/r
LirYOfdpumrIB62JJ4Ut4ClCtg7jH5rSpwvDJnNQEytE70LqUU0+HV9ir4A8SzGEpmjJwwoLuAaY
jMegjapI2aCsEFA7NjOtYEA2UVWrWydVQTdhuw5Qx5vLCUkP0wt5fnM/NAsU41hbvEVeVkneaPgT
z7ukxKJ7C7WO9hiuX4sE+ZM3d3u+pv3Ez+f44WelGJ0p4A2RaP9PUcg+wU88dSJ1wLw4xpyX73WW
VpjbkM/wXx/djFHS/SRux+o7czZsoNcnxIripEonwH5a+ZGjNtS5Q0UDr3ZwSmxCcJa7V7OEzk3C
30RWQbH6CP7bt4vPXyKkiKr1YwJbPJVyN99foo4FOXjEnzSHQGANAydDMV8b00qKyfX3tiZmAw96
rb547Xiu1c/PaHlj4mBHbrwhEAhJMaVZEqZQwcf8q0LYgKnCu4v84qVbO+DP8RQg2kXb8h8eOZq6
QfpSX7dcMsZB+iio3GUZOdKlXlYKyXytgTMv9fOyCcppKfzieeCLqTl6/oTnhBBYRufAdhluQhW5
e2BN0K84YOTkBy2m4Ijq4gnmAXfq4cy8cEWEmPsuMvF32fPTRz52Soopt+BnVj1HACOLjcFzth5H
qZwTrkIKduuy7unzMse4CMZuq5EhjR4DynejKeYeQrX4eFU/4gZ+6J2bUMsZN04jjNilp9bWImcs
OwQZ2WVNubogKliraLC8M+lIjxFZBJhrjGMZFrJxPbrd691/z/m5MkNHBvVKVdakZXTmAW9FGt0o
QwBF70xCmVM/uWvOBEHpr43l0GhkGY36cLEA5i/HGkxHOpiV9+OpWAET7b8ftRPcyGe9EyaJADvY
7VxAT3ieyuYBJ1UOR+L5TXKe8vje6z3lOp/9kIfnAkrB806+kJVvI8cNWiirFEWvcKA1xcHGKdCt
Uqp/hwYzu0uhiZtYvnbotxQOdwNdwxj4ituEBMqvfK6az8oEl4lCLCiQm+QiU5JQLne/DTu4ja+9
YGJao26MMLtjoeDN960Em0Yf5t8yVEdDUNTsS2gTlR8sZzoOltiuoXBK46gtfhElcDtnQSzgc5Wz
aPGzBM+IMr4jFWwCoKcMbakV/H1bfT+1OHF4ztu5JSejZUor7Lyi4aQzDKHVAA9OVw5nlfrQfW7R
TminFxW3mlltEs/KXPj4jyD/Nj88WJ704qUcYAlV3cv+5Wi10jtiw9EgpnHZn93zupVFjmH0IJZD
9lDvd6GjuVowrYwYppJy+wJRtkWzhpbX6qyK0yvroVV5RK0pQOBXDHVffFPFmhPdyyNZK6beBeOI
m/xbCrUFBONPLwfpKwXJv/BRyCDNNl/MrtS9+em4Hz0Np4moGiOP/pXmjWYZQRjvEXFuYVVKIgGP
3MaZRV755OduwISsRZxGGx/xdU7+E82ltJB84fjxUlXz3peZyTmiTb85or5lW7BMMlnV8BK4/tZT
Cfm6k/FF/bJlz6r2qYNqZ7PvGIU0z7bKOgJLAwniND9zCF/k5OpHhaAs4hwJYEltUHJk7bNTbtZm
CYzMDiyBcIo/ikqlOGBR2k4FbY+pmHv8RTmPZN0ApvQkABk5z+frpD4nXaJI0rBwHPw6S3qSCfb2
usgXbWLX+lZ6PqeO3mgGKJIj8aC8OE+BIdTOWVrJlQk4uN+z9WA/QyIe0taVg2ex0/3hq69NsVjG
V7HWkHf+xf/Hu8jW/riW6U3In8fAslKLTTW5xX9Y8DRlMN/wwl1tBLuw+YRjLbdY9AniqyDf4a4K
UlJw5A8kLqjNSkGHJUBik5o7dsz8QJKTzDfZY5Fh+C1TNHfQ7R2UxZdGhLg1/gjUPI8Wd2QWqeE6
WWOZUxLrRtxDTqYpZeWmNRw76GUHUKkuXOMiqdiYAJiCfbshYjnModkg4dKsYt9HuMnVvH2uhT6l
Pi2B5MhOuXi3ndPjfSd7CqrFozp1eW8PA4WTN4Efcwn4Yf8WpFnBg3rYg1hDHHFdry1ODo0/grIu
z73uFtLaSl/BuBTczTKqKvvyp6bDSOmA+wDLJoICiDinY0wdTmodgG6B5IKuPiItqXN6dd9j2nX5
og13nnaLBTAQapCYcojAraZXt7nT6suNlA4L1wLTibNxCjNefUhklkekd+fOTOBj/Zc+iyE+Wvpe
IIvBi1VfBG8puNlzut1pmyB2c90k44J8dd1a0NqvUQqQVzlUnZOFQKHMgJRHjSZwOD5oE2UzVCJT
S9EPVvO4LglYlqa8F64nXMtl9N3KvQCCHddBQGmZQhN8HmkUqgA4XvJW7zUw5UC+pLD/NOj78FdG
d7UuuiopvhxfYcE9DoBdoquUc3riVxKmuIYdV1Oq2rK8dLgkvVuxLohi/ShQTKRd3icpaxtLKuhp
px2AfJHqGWay79TcoHPEIwmflXNnHuQBXsA+ZQgYWLBqAQ2yk35WkGICuMoS9yiSt4XZuX/G8Qi0
GBE1RQoIn7cYqqWggvh7bTCKWadY7YKbfjtRoq7lfdH1CahC1Ty6IaWAq9MYIYHGaVJq0+a8TcPH
HJujo/EAsrP/WXFQG1poZhF83zKIGfv+UT7aEDWUAelA0VNzS57YGbthN9ttderx/B27AKkH5eA8
jOO+GPbKiMJu8Sgl3pkNN9ulq4q3cuvupqwYrhK8NkIzuWhY8P0xwO8hNZC2c4GVKC+AjVmkS39Z
6N3Sg5+8HbXv3hjmARQvKC8XjSv0j+tC20Hq80kZthyhu1ONL8edFlWaV2Q3eIX9pvIVg/pE4cnJ
nkTvSa2DCIg0+fVB3HA6wz0tAVuCrLotjQ7J+E6vl4UBetJXdR5lrJBQLaMZf/GhAywSsyOyEudI
m3bksQEBstj8ZiyRPjJjJCopY30mZDflg885BPn9DRlcwaKLJ4sskGe31g98ChE8Fv+KpJkaIs8R
2AlOk/7RpuQRSg9/e2fE8nzV5Av19mYzIvzSGkI1ow8qQqkS69J255jhOcHZ1Zr2xXhsEIHLOa9n
C7m2oUwo/Chf5P8S7MdzSFAZ3zKoQiMZ6+QAnbXUVNYfLn0SuRkkjHwk2CYLsz1rgBZd3I6rxnKC
ILx5s/hWXbbXzYtGt0JsLIxnsdkHD7WuAj0Se2cCJwKCQnKm9IYMSCNmVQ7ctMFTcxi6x2HeW+0V
ljvuKd8Y4iCIDF0thJGB6wzX7tLh57uYHjpE4rqm+tga9U8pYqERi7b0rELGI8vamZutRFK4h2ja
FyoxlY2A4zM0+Ps6w+EQV6xjBoR8dji4AnXqT6YYCnZKFW4TRq5f4W4YNgMYErxDB7v5gqrFXsLJ
KJHe0Rlvmdmq+OgSAyCtk5PfF1FRozdLamdH7QuVYml2o68rwpvUKVO5/u71HMxZs+NsF7ZNe+01
7sIb71jsGDTTUyot29FYbsWFXx7Vq1W2OMg9r4adV1a8znuHBzSs5dvFCGkp4u1ZiV07b6CgiYnB
BqnQEmuIAUjevCiNrz3unfBX9kZk7Rg8SQyAWVlYOR7L9hCYllPv9Gwhvo3sESFAusFiOQtQOgdu
ewwNt7JkZwinjsjURhLF/Ym16pBr1ThAFkp6nBYiokVdRjmBjkmKSnVK8L3YapEqSSCJFlKnDFtJ
/4SadNCIGJ6PjAgSiYHVMnjWzaFA0BZfDyGYxic5zBmKYByN9aVy5sQhTD8gcsclGQ3Hdehzl7dt
Ggi6vizNNoutJ/zdq8visEM7jdHUKQEvKwBswB2QSFeJzw/ReymCvED5Ha7jMdwHXpvA/KQIF5nI
+HCXhDZU/1Z4jCJF9DPFqQxSlzKnCaAOCBMJ8FmeqxOLCldqN5WYnKRmhhDrVmzJ4jjO6zUaVKLQ
gNn9S9IU/fid3mXWo+X64L2mcVE2PRTuFGTnsUCnoa7/6EUm5TE/9eCGGFx0d7bOdrsrovRIUGke
X+AbBUVZRGqfLd7d18ITYNUmtSEFVMP/L32ypwCcCHftR0oqCzRG7nIlW6UhrFM8W1WJohG0mA0/
LrC71GC7m3QVy5SVKinysDfa+CkMD3N0DPAcNgeKq1u3vG/m4NO1zHjQN0DP+CHsPwioNnVEX8nN
83tuh3B7gnoctGY0GYArlSawNB22Rjv7yjRyIIJNvu9qoZt9vBfmJKkZFy5Anl0kvM/M8h1g6q5V
rIbq+C7wH8nCFSYXdcek+f6uUj6WvJkU6Q1fG+vafAywty+CTjuWoTdD4kdeC0ycTDH+CQksOxu7
rHbwsxvDMX1eYcRmrJc0na30Z4cyJ3QjoK1P7b3r4b7TQbQIEG7ExNlJfpBI2GsGPuhKDseBBtRk
fQObj2yCcWBB+2XIPWtmsYKJXpPIZSCgyvl7xlcuXgkTrh58Tjv+f4mX52dmrA8OIbsdHOuIuHfx
XpLRccoXeIWKnC6ORECnt26cWlPdwZ117mKb41HyfMHmDM7pfr0tGvyfD82Ukm2lpps8NVuql8Dh
FAt0wBqjItXSE3m26FHfwIRiiH/qHEnBdttH0heN+Z4puV1m1p6lY9mbjlSe
`protect end_protected
