XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���d-|*_�l+Z�q�c��6�P�T:��!��[�U}$��R&E��~��rP,�oܬ��MT�`���3��@�Qu0��"����l*OZu�3{��j���F7�O��l�:��hWf�4��\_-�\b�0����@�]��P\ԪN�.����1���n����-�Ao�X�� ���-�=G�?*�h�`���{D�3������5(��קk"%��h+};vy���L��\E���$TS���f�<��} ��O3�������_��;4[�C���mCq����h㷊�:M�j��!�'���A��;�2�OU����?�|��)����^��ϙ��Z�� �V-Ei`�dȾ��#Kޞ�۝�'5&Ȧu]Ŷ��_7O�ހh���~m����W�X����*�7sF�r�.�0()F�vR��/��ы�!1��W�Vx:c��B2��K��.�#Fl�ރ��Z�6m�ާ�9��.��B��l�M,�x�h�`�� 5W���1mk�FA?�{���*��[��I�l��Й�����j,q+�X����UY�j������ڮ�&���S8���J��ȇ�v��6�"�Q.q3�@����\�O�����p���yɔUn�R�j�Z�W9/%�q�JF�Ґ6���̆����c�=�AO|H��O�F�_���ym���Tp^��0���&2��[�����p�~�CN�w`[H='�Rf%l�%��	����Y'Vjm(�\�kr��,8�l���<Q/XlxVHYEB     400     1d0�̞@QC4���<�E�I��	Ͱ�[JB��ь8�`wX:�,������HJ�v��1��y�/>����;r\��h�v3AG	*���wH3�F��"�}A I<����T��RD�E���.�����c`��l[��-Es��_���gϊˁ[�j L����@ >�z���)֡ J�
�P�F�6AŁ;�֎�&e-�}.��_��{H��7'��dw;a4d����x�Ί�Wn+ɀ��	� �1�ȳ�`�������mڷr��:�1� ������0La��w��oK[�m�t�p;�/��q���¯�1��vOl����!k����uc���6\�z;���m-,�w��2�?1'����w/��8�Vu�����5�T��#�����T�{��Z~|��N�c��#i�2��y-(N)�˅�=�8�^�����),�����IIOC7qI٘�Ķ�XlxVHYEB     400     140�>Q����� �6�i����_�~ !x�-���l2�G(0���$�Y�y��n�`��S�T���b��������#�B��p	E�4k-b,y����t埤�����������Wj�?�u7��i�c ���F�wxH2T��b�S����͔�l�8
��t��.j:���6_�����XxU$B�A�Z�])<W��">�;먭�\vȥ2j���m���U^h�#�B�_�? Ž#M�"�����]S0����zY{�H%0��@�|8j�kj�-q��q�z�*�%	�nt��}י5|�	Ϭ����(H��pk�5�-�t�w����XlxVHYEB     400     170�<�%�#����@ە��[jT��	��H����.<��?��(<�����cFL��cؖ�{)�~2���iIĿ�rP��q���`}���
H�4��ZC���R�8�dA�@��`�I7�o���E��(�ɀ�R]��Z|�8���) ҈�����T=�������=�"L��9	�1�E*/bY��� >�%���H]4�o�*j�������n�A+wb�;�ϊ��K���g�}�����F����� ��T c��`}�z��(�6m��=���J7%�c6p�ǸI�Щ/	�ះ
���N�h�c�amd)<�)��j�+ba�(��Z�x��� ����b {�%�槦��n���r$jL>�)XlxVHYEB     400     140a��n�=���ٗ�r�%T���pW�%�`ld�x���b���X)���]����O�Ӑb��p��t^���s�$`v<�"[��z�I�!m#F@`e�������+��N��a	�kqq�&\��ǘ(qd_�h��J������;'5��!G���=c���ܶ]�����#
�Ku����3o��pD?#q����~�?X�c�=54<���M��M�ep�n�w� n�ss�z�݆��MUd��[)�L���>����0Վ��lMs�&?j<��S	߻x�5�]V�u�;vW�K�8���n2!���%
��#f�XlxVHYEB     400     110��9Btc��+�<^�s�d�� 1�d<쐃���;�ʷJ{�-�u�� .5�[���}����IX=?�����[&4����F��U�}+��UV��OP��uv�����P����X���D����v6�F�H����B�pĚoX���;fs��'.�P��
Sc0��z�S�e���~�DJS�d������{�����%Ǜ�]�3�����N��[v��*bǬdU)f��:iq6r�p������k/{%&�޴Un�JB��J�;�)v̻Y��XlxVHYEB     400     1201YMj,Sk5Q�ȭw� �hf�bhz���{���z�������ՄB�̱:��VlF̞���%�Nf����R�6�Ur�fp�*��-���(�#Sn���NBx�	��*��"�X^s�llm��J2ڿ��\m�������S���v$�?L�D�<׌��>��E=>[E����e��QФ�����-jVbʤ�>e�c������A���/~��lW7�r+��Q�d)��[�S~�C@~ݙ1��+Oz�kZ8�ƶ����d��3f|�s��l�o?T
�-��V�XlxVHYEB     400     140*R�q.O-2�T(#}���"�>�	]3�N��⸟K�-����	4�2bGEF�*����\��s
��r9�Ғ:����J��Xo=x5���ˈ�F�u6% �8L�v�Ώ�3�ʀ	��;1��0y�H�ռ
"'ٜ���9*D�6Nw\RFQzܴD5��-ă#��W�}Jon�P쟐��(��r�]X�A5�R�K�e�ⅷ����E�!��C6Df��������)�9�����mS�e3��-ِ�4Բ ˕?���Q���.@�;. A��YR6��P�g���[!h8&�T���������q)�XlxVHYEB     400     150.8D�#�ހ�Ǯ���i�h5�N�fu����+-�}�.4o�K�{�n�����1!pQ����b=`��*�)1f}h�W��JzQ���%˅�)�|ޣ�:�Mѫ�q�,�"(Z�p�O���>& �ܞ��l��8�L�h4�(S��M��-��*��Y��7��JU o�j�n�9')F����3(^�~��fkؐ�IY@��9���	4��r#:S%��Q'[㝊��3G�p��$��F��Ym#%[Ⱦ;�e<�Y��D��e'��z�~x��,ǎő�?ಪ���� ��QX�;Q���;~�.@o?��2����� W#!�B�sXlxVHYEB     400     140kHE����c�v�ˠBe&�u�� j=�e��$ޮ%)��!:|5���G�r�����&��-�(���h=;�À��+�4�l��e(�'�gn��]�����U�/��P��&�?�tw#��?mu*��nZ~�_�������Z`�Cf2�9�S�·��ٳ}��P��5wVFF�=-�몣q�m!�
8��}��@�����G�܄��%��Vm4`�����)X�V��$�Br_t�k��$��H�Y$�RUm��,�HjAy��[�_&�9����gh���''��b�ޔF��3(����e���c��Қ��7XlxVHYEB     400     100�)�|�ܐ2��2枷�{��+436x^.H��:Z}��ьf��_}��~nR��3��Vqϛ�i��.m��	����,d�̫�,!��0�"�_L3�g���"�eD���Ɉt+�>At(�V�-���~R�J���wp	Ǌn�xk�������i� j���`[���Aݫ{�D����0�I�9�g��7�������dl�r��>Rt�^β4(��f�PŰ'ϳ� t&�h�.H��/�A�i}JN�fiO�XlxVHYEB     400      e0NL;������r_�F����x�ذ������nB��#!��m�aW�S\�&ֻ���>����.P���_n�%��l���U=i��w�ԩ&��c=��/߼:�Y�ث���p?o��\�fq	���LOVx�_�KL{3����hǏ��Y�Ѽ���5��a�����UY�<:�E:��ŕ0�5�z!	eq��Ϊ\�N�*�n]�1)r�^t��y!WXlxVHYEB     400      e0G���Cv����N@P3u���^YRFYFO)�,�r���]ss��8�#-ﶰ�6e%�`Ԃ`16�o����Ec(�}����;��E!>�`�{Z��JC��&(<�� ����|�]Sy���~d��θ=�s5s�*����d{��g��Ժ��Ϡ��׵�o,4�d݉��2��P.�[������A;��U
u3��\z^����#�|���dc�W��ֈ��4XlxVHYEB     400      e0���H�#[}*���<Տ%�Ml��n�vP�YV]��)d�W��Ϊ�3�	-N���H���Hޮ;��1�ؒ����4�~�ԉe�2&,#%� ��7����۬�(�?Yyּ��z��rxǱ����n�ƕ��s��i�g�ވ�Yw�7�$��G9��=�n5/嬖N�M>�+>�e����2�XL�]x0��3؃=s��p<��io`2YoO�|c�qa�P(]XlxVHYEB     400      e0=�txU{�-�� LUE�U۰�L�Y�CpuL���L�dXY�������&�C\hD	.`��b�ҥ�݊9��}Y+����I�M	,�9
������r�#�٠�f_�6)�{x�D�E��0v
��6��׈�'�`�e�wЏVШ�E�5��@+"��=�Sæ���뽂"#+�K���O�4u���I��@��a`������� ��9�σ��kf��@�e�$
sa<�k�XlxVHYEB     400      e0	�6��Ѽ�Ph��cu��wl��
"��i�$�/��yL����?�	#2�%u���Y�/'������A
M�P+���M����S�kK�QgC�wL�k���G� ��L���.5���� T��b Zx��_����p�ۄt�/�%wi���V��$�r�Th��>G�nW����P�G,81� �0o�
y���Z�pI2��`J�7I�l--�����fjY�g(�XlxVHYEB     400      e0R����*!?&l$uܹ�Վ̏��Ffe�mQ�����С�!}�ւR"3��|�Y ȡ�C�IM�c�̙mǪ�>�� Vx�蹗J�V^_&�
׻(� �v��E�����l��������ur��Y�P����h;bGjPӭ��vI�S�S���ң�B�@�R�c�8�����o���m��W0��xmS�qn�-���u�m����A"��Z�&��XlxVHYEB     400     1c0U}�Ӵ�,Os���w����L��o!�ɣcue2s�-�7 r�������?�i�u/��W�j�eh�O���Yu�T�Jɪ�C��a����ȋ�玷}I
Y)Y�,=F|DI�����Dt���:�Kl�3�)e��m�vw�'M���e1�!x������E�otok�Q�U@._���ev�����bE���I"/F���Q�����JrĘ�p 2��G�ea��CP?�͌;�����^B۔5�{g�����$R�Qrs����rW^{E��8O���m���s<_ex�D�f�祔� �z��]q^]�"�Č��-�yO�'��:a]I[�nũ�3/=��Km4���+�FC�"A��#�,+/���wA�t�d����s�>
c0�BĤ��{Z:௅h�\�u�6Y�h�)��WV޲�)�����T���B!T'�;g��(�KXlxVHYEB     400     130cӇ�>9iD1��ş]I+@�+g%��I_��̥����s�ԥ	�leh�l���>˛��?L�Mm5��#e��.��y5˒x�!���B�_VQ�;s�L��i�p� �IF�3��{8`�]]��VT�R��ޚ<~&A��_)�Y�@�\�j��̡�X#w͆pj� ��fH�ӄ�/Ђ�����P�eD�e���\�%���-�a(&�(\��n1��~+��&n_¶��C���P�]�a����6�y��x�{[�	�U��$�(
E$C��K�qT��C2[pⴷ���ʃQ��|S� �ڔxXlxVHYEB     400     100႟Q���6o��9j�F��E�\��K��A����+�Jz8X�/C�M3|��'�+�}�9�@6�k�t������_~��xi��l!I}e~�'�gA�j�xl���(�w���Y`-{{����Yy�d&�v�i�h[ZVmi�^B����<tW�&t�T��n�0������/n��Lp�D������%�~�a/'��[F{�[M��6ı����g�4R�=m7(L�U�H�����M�!";4UMC���������XlxVHYEB     400      f0u�0���q034T`D�#[��*!�K���_��y"�$��J*RMw��pyaͨݜ�/��6g�c�$Ҿ�GN��6��V[P?$	CPP�2�vf�|���s,�d(|��P����rXP�/%&�$�W��.�֬�P2�S��n`�q��i��;�XI�Y�@���'����+-�?��f]P~���`�E�ڲ��
���{�^�I�p�4��c�*���-�qĆ��6k��e���XlxVHYEB     400     140R�P����	�W�;��ٛ	����O���u����1�""|y�o�;�-��2]�=!5}�b���
��d|� [��-҅�w��@�#����ͪ' �4��r��'���U7<*a`9ق�c�x�NM�"ԡ	�u���>�i/������`�AM�&!��04��{S����p֢د�3��B9{�F�����>�)�d6Z�R`"���}&x3���`m��]�X\4��=����f���x�
��*[w�w����|c�y�<�ܘ!H����ׯ����iXA}_�G6�p�7BV���`:IXǛ#v�.���B۠�s�XlxVHYEB     400     150Y���h+i�,�F��4�O]�;�m9��5����T\c}�A F�7�����O�M<*���bƻ�5bXem���JS&@�r/�<`���ȗ3Q��CG��8xL�K����:`�K�Cͨq�剉?���g=aB��cr#��D�N#�J}�ۭy5���u�`9�A�˄���űW���AB�mj����ȟ�ی��L�!9K��r�Q�8$���]��	=�t���YHï���̼��W�ц����^,�E�Yuݐ����q�J�s,s�]3QI�����d�<�����KF�?�M�.�*����#-Ȉ<�m|:D�7K�XlxVHYEB     400     170\OӽVB`�kq�H�ՏC1�:BjW�C��i�>X�������Z�h��
i����?^B��쩏����U8�����D.์&,&o,�n������ʭ!�,Π@��վB�M��.a� Bh"ͬ��r>�3!��<���>NŎ�&��:���H@^�Eoɢm%ޥ����_sM��6_��:;Bc�a��� ��V'�z�n�͆j�Ka�7ĕ�_=p�J=���� �b��@�2.c)Im��m�0���	�%���_�W$�t4n�R�NE�\~�pV\\ol'Ԑ��B����s�	x�}�ձ��N��p�g�H�C�54q�E��К�g��/k�,D��|�N���7��҅���8�˵�ee�XlxVHYEB     400     160�8z����z���Տ��t��Sk|�g���;�Zx]ȯ�G�hx9?����'�D�u2��ى�6��y�>�M2K0'����>�cR1X+t�-������_�i�TySn���l�ӴqK�y��jC]��븼(*V޳�g����w�ܰ�H�#��Ǧ#;w�C�EJ�@_��sv�I��rH�޷�
`��0%,:�G�F�?wp��;k�̔�q
Q�����϶��M�d���f`P��q9�qm�<Mx|���,��}C[Y��Sl���'� 3�2$e�
�)P,�f����J�o�,-w�X�ew�z+����7�%�eT� Y~��,��h�Y)lO��XlxVHYEB     400     180���Y��N%�Z��7I�S}DMԏ`VF��ɟ,9,|R2�ޛ&	-�\t����h��|H@�qH�;j鸣���Ti�s�#c��Ju3o��ƺ����5צ�Bnʷy�%�)��F\�{�r�ŦxNYV?�+c�EZ���9(�m��P8��%m���f�頛«k��L����륡������Y��ad��� �'���֮��!ĨH�,I�/���C��xg�Ǣ���ϡA"��A.�����Y]�$��z�6�<������E�_X�
���6{[*��0i�VL��|�UI}�. CtI�$U�����8	��Y4���:ܴ��'�	V��$�}tQ��Ŀ�- P�s�L/��/�Ęt�Z�����S�XlxVHYEB     400     100ȉ���Jt)��7$�ż��\�(���;����};�#~�{1�>kתR6b����`�;��	]����<,�N��ֶ欄A"5���%���ܵb�tK:�yf��k���Y��Y��/�76ܞh��C���cAQx֑!� �L��9��!b��<uO�R���7\�<V�9�BN���Pw�dFq��#��=#��D�;���浘�5oU��D�g0�JX�������5
���$�����LXlxVHYEB     400     160��}�'����t����?�@}����^��a�Z��h�_����A�}S�L�/��?���i�E����;:0��xKY�]P���kHqAM�:v*d����HCx+��u��4���G�5�)���%@�
��K7��e!���A����A�}�le:bW:k���"���>ʾml5�5B���o<�%6=#^�2�
WHLv˧>}6Nc�T��B���6Z9�7�
]#�Ӑ$�3RRƀű�v6~��G�)?6+ʺ���yh Y�!��h"�U����X�'���;�"'a���cq��!nǆi;B��LXaS�̽�x���*����4�swPQA�֛β�H�� XlxVHYEB     400     160��>b�-�g��57�r���?�|^�fQ�E!�e����m%����H#������|=�M��	`�l%d�P�i���$��_�f̄.�W+�� ���.�_�6��Koi���P�'�rA ����
��sT��Wߠ��A'���*�jۧw�DZ��[�@��Q�Ye>w>_�S���C���G,�H �L���w�9�g�7.�="��� �6|��Y��22����_y����ȩr�^&XX����Uapkp9k���m�Yy;u5E��5�s̑I�]Q2=�=�i�V#�u��~*˿���պ�k,6%wȠ�0�_ksLJ���9�u��p�k�S=Z��\�:H��_R[XlxVHYEB     400     140���ٰp��n���?���x����e7'Fm��8��wi,?`H�SF���-%}��q��9�}$|�E���g���N|��ǿ��t���f_[���d�!�*�<~ds���N��ގ"�ݐ��i�q�����ՆȍƢE��:M2��o�l56��x׸�3�kLL}��x�f�����+��kF׹��5 ԙe��v�51�x�c^�]*vF����Q� 1�xE�גD�wB�U��!���A���	FWl	���N�*Hg�8
TQ�)x���G=b�&������m﷏*�Z�������Fh����a���XlxVHYEB     400     180�c�\H@#�f��$�$|[y$�$�C��JeZ�3��9n�X9��t1b�@���r1dĖc�Lt�^��C7��N?��8�$�iҍ��ȗ��P@M6O��Х�K�⮊�w�-Gq[��%���5#���Ծ��x�_���Hh�AHdxhN-�`���ď��6J	�Q�Oۀ]��l���p@ҙz�1%�e���y�&��R�zu��9�N[H)��F��Q��Wi<��*���?�y>�H^�|o�".җ%��_Ox��Q�����a���t���爱�g�1��
���3�kn1�%��JB%><[ܨ��~�O�G�*�����f�\��2g�ڽ�"쓖�����Ok�ݚ��Ԉե�'��U;[�!!E�0w�XlxVHYEB     400     140�xt�yl�����ܠ�S���p�1F����Ik@pJ�0��7��m���g<hl��};>k68$��	+e��z����',c(m�F�e��t���z'J�H�p��G'�ѩ�	k~�/&�<� �vҮ$����3��3�C]�q%�6F�C�S5�ktM,[nn������#o��W]�K��(M��T;N%��o�^�� {Du|A8w4P�D��o�N,�R�t�HO+yh50�gmpk��}���B��ѝp���j��vrq�k0����1]�D�|F�DT�A?_ZTf���~�HU�od�*)��'�XlxVHYEB     400     140�D�K�9~��&�����f�"���A��c@6�0l�tծ@]ch��c�<qӊj,V���bU���Z�j��{d�7׮����Q���-��;��|fo�;&j4���VKr�#��\'��3�w�� B�_>B�L~�&��&�������]J�MҾ�ac�!�c[a��HƫSO���#��$����]��~_U��%^t��`E>��g�����]�/��`uDMK�[Ϭ]Y��L����z��Iͨ��[�'�WNA�g���h�H�g��H�L�
� 7
���Uz��,o��FۣXlxVHYEB     400     130I(+r�$tf���� K=hu��ޱ����/��/��rh5M�^��2�Q���\�uQHr�k���9�RJ� ���4��6����'�k���
�nUM"��� �7f2	O���ֽ �.1�P(��ZIE�43x�G�q���11鳉x�xz�\���}��v�Rj~�Zo
� &�3�ӌYc�"��V``g��֝��&1����v��_S�# )�}�/ ]�x[Ŧ"�Q�/t7��Qqq}�E�GTn:���}J54,^G��S��b/ᬪ��B~��Ul�'�&���Zux����'G�y����9*�\�HXlxVHYEB     400     170�^:�U�:������K�c�r5$0�!A�R碶���!W�^5�VP8�d��
8���)Gq����3�o"�.��X�;���� �*�����<Jb���W�B7����/|oFS#�<��}�Sܩ��:'�?-�(Hƀ���
W�gr� �:��^�a�����`�q��g}�
:��f2M��r�HǍ_F�,6�T�t�4Ώ����3��7�b�{<�Od�"c�Y�}�!FnD�����*�h�g8
ݏ0Xw�]�Ul����I�JS[$E_%�����J1ۈD\iT
�~�.gvJ���_���_9�}�(�E<�͊���Sf����g��^EH�s���'��M�JE?�OY�HO XlxVHYEB     400     170Y�)�n��̢��`���ɯg�]!Ո�"������ ?�c��O?IV��y���1B���v�f\f6����U�N���b�d��+rH[^��`���	�T��P�F^���kG�χGؗ���g<ej�����Q�+GZ+��ah�2�Etʱ�Őנ;��!U��i6s�)ֲ�8�gw�oL)t�l�k�R��#�A��z!j*����G�:�H��ߥd��[�'�u$4�e����n�[�:e��Ʃ᡿��Ô�b*�h�8?��^��(F�s����8�����`�V�tt����'(k�-�vv��V�D�ш���$��ʅK8k"���#�1��9��#' u�C��0R��-E(��Uğ=��+�h�XlxVHYEB     400     190Y��� ����@�޶�6f��1�����v?3���%l�s�&��Uٗ�z�gaS/����p�
`�Fr���YM�R�f��!�Z>|�U	�B�+��Z��:$�}�86iJ�d7yP�⒪�A��nbN���5Ʒ)�]�w4��/qzD�`8���q���N��������p~�,Z{mT.y�	J����y W�	�rܲf	$�{��U�	۰��wK��-�̙����A�־�R� ��::qyr ޓd���J�X��U��)�1j	�Ɗ֘�Ǫ��	�4=�< �ء�U4V#1O�V�"V����4�*Mӆ���غ�6�1z����ތS{?�́��i���bHй��L~�r�~n��Ko*���@
wu��h�^�2XlxVHYEB     400     150���NW�o����и���"��t]�m�Ca�֧��i�����|��"����r�չx���<TH5$���O�{F�6 U:ۧZÃ׼�����\K�����H8]]6�hU&zƪ��%��j4���*~h"�ap������x�M� 6E�H%�AZ�]��D�?AA���uA5ݠ@ /4>, Wd�4���Rtq��՞���s[�L<��J�\��ts�Cc���^~<hN1�n���ZS��C�7�a�'��q�H�b�r2/����&�d�m���;G�� c�����1��^����UvH�&����U�d4Ai�׈�(Z���������v�XlxVHYEB     400     150#�,��P��|�-�a���g}N�<��%�SlWV��<�4ȟ/�:'���z���4�Y�&�Vώ-�1��f-��@�+_0sd��
�{Y�B0TɊ��/�E�?�6�LTpݦЕw��M!T��ek����|y��T�4�����_i�O��D�~'zٲz���xZ	no�����KƇ�pڷ��� =@�uj�t8S!�nE$榪���]vΙ+6�j{�;�/�gŀ�wX����Y���@��iՀ�!2�̬�=�DtJ�S)Eg]�7����!ӛ�>t��C�髉��C���a��)x��IQ��:�ʸ��Yy������Tx��V����Z`XlxVHYEB     400     160\���bOƂ0�F��Y���AͰ����/S8l ^j>[t���Y��G{���n�:H.�l�T_L�c/��(�ծ�	�Eo�L�0�J�Un��h��E�:?&�}z�)v�w��Ϟվ�䄇A3Fz\n�K 
u\�����ǝ٩���0.�Hڜ{.e�)�(�3�*�X\}�LzX� �����d ^<�T�8i��/&r�C�a���{����c�>*݃c߷}Rag��ފ��+}BX�jRWA��\�P��jk/.݋��1;� �U�]d�~f Z�L�.�������ژ�%77G���,P��Z��|��6�l�O��^U%����G��5�ks��"�60X�XlxVHYEB     400     140p�na=l9N�B>�bk*�¼ �g��d�t�vG��'k
�qoz<
�NoG~�Q|J�U{n.����=�p�# �T[E�dQa�����{���	qZ��S;�Hm/�K}�EO��^�$��w뿈���n�@��*`�4��;rY�&��q���P���&��%��.秼�&`iV(��m����p�o�>�8���dqY�{_��CdX�/�w/"�k#���<�۹�r����l��t�`fX�k�m��<\�e?��-�F�@+}��x����a��D���BC�c�(
�
¿)�3��X�M$4�D��u��=<XlxVHYEB     400     170������+��%q(%��%�k��U��C�H_Hl��!�(e[Lܮ4�m�>��!I݄ɋ��xsۯPI���<=�$}�]�R�k`y��TC�MX�@����6N�F�c�y\�.3��|*ĨQ�*-@�PvYo���J��,��܋�c��b Z���F���ϊ��� �<�w��/*#˶��֭'[���/�V'���?}&�U�;�����)��T�#D�sU�"�9�<m��&��E5��Sͮ�IX��L�q��7.6U��Ҥ��J�Y����ۍ��NP_�4�b��d�l}�0d9&�.r�G�.I�"(M�7�Ć�r\���(+��
�9��d��@\%#׽��L�]��dIv����A����T��zXlxVHYEB     400     150gȚ���<?ٸ.Q�F��"+P.J���Gk!{���=KQ���M\<hf�R����,>Ɩ��8h�ji��n>�7h�T�m<iz���bIx�>���N�ͦ�9���0�-I��[�%��̐�C>ē�����9�C�C����}f�J0,)�y6jt�pڦj���K�����i���čX(�{�DN��Ȫ���ϑi�o��4	�KB:��^|��S޴�E�������!C�Ms�?2.�t�>��r�L���;��Z"��L�O��Q��^E�cj�J�(��#vRJ���{�����<[j%ڜ*�����:�i��,
��֢�	u|e��XlxVHYEB     400     110kA��L�x�P���H�6	a�PA���x��"�,t��'�H-Fr��z��
W6)��c<�hE����w'���җ�<� t��L<s�!�3E�c����<��d�Đx��]kIxI��������x�?���\5.[D���&y�IzP�����xWae�ҳ��1�j5\���}��,��h��@"�^��a��͵`n�3�̻f����(s<f�sk�@��
	��KulE�H�s�V=o��$�S�`���#�����r��rE���LXlxVHYEB     400     150�>�2[�۽U�Xc�LT�
�!`i4K3#r��*�
1z����շ� 伺�Z}ѵ��a3t+eW�֖VG�V%B���=�Oot;�yb,��50HS�V�[m�A�hkuh�&�g��vR��{@��7{�-��Y]ӏ6A���4"��4@�C#�V�>t��swew-?�`)�_B�Ek�NrS���6J�g����cƓS����G/ڦ��j�`����T:3z7ڴ#���;��,Dc��^�_>��q_���V,��+�Z!��:F
H<��7�B�&$3�Ƌ�-�'z�r�|�j*����s�	��$¬�C����O<�Ef�XlxVHYEB     400     1a0^�oС�Vй\y3�{�TGJl�c�-@^�bۺQ�k˾O�|w�q6��<*<בz1�ɞ�n��M4�%�� л]���0�G�A!�����}�����wm�^W�e�.�>�|�#��YY�΂�'��#�7�J7�"��_0|��h�`�T���y�5>Oǲ�'��	�FI�*��M1�G.K<y�S�K�%?��'�ؘB52|;��C
e�z��앫�U&�N�B͕�F'�g�yhЭ�hGv ?�*{J_�����,�<�w)����������]����B:3�o`�ͣ�:�e�v��X�Ȁ3N��}�X�eS$xIW�
�J+�a��M*����RI(��p<��2��B��U���<�X6����#�<2`8�������>�XH�0XlxVHYEB     400     130�>�lF���WlbE��F�W��4��4 �JϹ�.i(�3��Q| ~��� ��V�	Є��ya�c�:�P�io������_�Aj��ɪ��|z�i��n ��^�����$ �y\�qt������z~zw��7�k�2���<77�9�����	�
�f,f�ɒ��rt�O*�,���D������&�M4��SOvw��Ʋ!5v�LFYd!P����dϰZ����%x�$Q<6As�rc���:C)�g�]�qy���AT3���ݭ�?K�[`��:�!��&́��?"�Y5	y�XlxVHYEB     400     120�;���&���Ǟ?jy�����|N�g�l�t���?U&�<��i�d��J����&`µm彌��e�� �-�����V��	��"/�_,$�
s��hy��0�'j0�wA���I�m'�Ğw�OĂN�!F�5I�d̬bУfi?�Ȫ�z%>�ء٩�}8��&	��9�j'�Cm���S�j�d.����x�HC+�3{!O�Z�Qb��������9kL���NS����
�)N�nÍ޻����[�ic�3�W�V�/,��2S�%qnB��+����B�XlxVHYEB     400     170�lh��i�>��?I� ]=b72�b��i�]�w��քo����e_�W��Dً",���^��WzD�[� �׷
l�!�sұZ4�'�U�(7�@�]F�$�w����5aͮIPA�� �����)��L�6z��ϥ�P܆L���d	�_b�ٱ���pnj��O�ʄ�}� �@y\�;�����'�cJ���>1�����ȴ�JF>���
�1�<z�&*���f�(�����.��:�)FeN�]?B�(R�@�\�,���9������7�Y�N�(��l,�'�Y���5�m���p���W�c��OI�1�*����N�<���l���2�=�?o����/�i�7sP�XlxVHYEB     400     160l�vL��]UC���Qt�)2���нy�Wt��ݼWMBLv� .����0��>N�d����נ���[q:���ŕ���r�V��T��uS4����۸�0Ӈcs:]��d�JY��@sW�V[���|5��y�~�����L57$��g�Ȇ׊�� �
�jh�x��#��r+�H�׳�F�q�� vZ+Q��ZS1]r��8j!~�s�);a���Iqי��3U> ��T�+d�$�x�|2���t,%��S����:qg��G�����s�>��l�H�e�H���#n��L�A���1�7����bb0%�uv����l�keRN��J%�f�_�%p'M��fXlxVHYEB     206      e0��Ͻ?�!��18�k�&�jm�|���k!0q�1`W�f����N��6�%�5
&��a�����5���3�b��e&nGj����X�Je���c��f�,��w�h����*�-Ʃ��5?0C�h,f]�"��
���,ְ[&���#t��]�7Ĉ[O1=�O!�Z�r*�x�u�u�����`����gɽ8�qx6๑2:�
��k�v�1�}��