XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&w�%+����G��`~���qR�9E�i:L��5�����,� ��ap�����].���>A�!(��9�Fʞ4���/72Z紙�]
P.5�Q4S����½4��88͉V�ױ�̩TM����v8J��|Uc+����=�e�c�iĤpo�	X��Y���P���{��K��8�����,n�����Z����U���a�C����}��-���WF�}��*I�㋏��iC�^���\�V��];a(�-�E��]Tj�8"�AHw�VJi�,�1嘸���&Vϙp17� ���7W[�aL�AA�W[,6�j�!呐hA���^Uy�P�+�65�0��ˇ�c��-h�m��[�{u�1.�g��N��:�y=/s����q�cN�-�a������P�g��[.N��5�\�b��Uu���U����]�gA�|�8&�Yư�;��8�V�� ��)�G��+0���0R�� �l^�3ސ61�p�SS�I�C���`Z�+/}�a�NiQ�!���q�A�^��y�̀48��c��.�CD'"d�Tr��^W��=�.b7.o�����%G<7&��ґ c�}n�nJ�{�U�?C��-���=�I��E������ͧ|0�2{����q��Ƀ���e�[�|�is���`�e�?��6q��I9��< ߌuJȡ���������O|����.�[?�NB�����:|� )ٵg�ܝ�H^�8R�j��~^c_eWѦtW��L���`c����Gd�,�d[�XlxVHYEB     400     1d0Ҏ�VZ� (*Ԣ��T#B�#>�R��:,���y�J7���߅n����Q��?�G����TW���V���w�����h5�]S��sXG��)�pqF�D�VE� ��;g��H� �P�*U]\ϛ�r�����f8��@����ơ=��S�U�%��,��@�5��OT���:i�!�׬-@Q�'�r΋��v����G�(\�)�ow�q]���!|Z������
���݈&A��v�����@����{�k��UGH��˙T�ʗ�U����y���3��3��Y�g�i*@���9$3?�$ �7_�ߋT��q-�DhC٘��t�|�)4��*f�ەce���QV+X��ߧک����@����S�O�Q
?�x���ř�|� �s �8��C�PC�4��ox��.�u�ө�ΦR��A�ơ"0ͻݵ���3��G���YR�@�XlxVHYEB     400     110�Z�u�-���L�F(k��(8f9
�+�Jk0[�O�қ�6(OǌCy�x�n���[o~
�������T��0�π\�v��t�W����&�O}����L#w���I�N{\�H a�yh��/�*r�ԩ�#�d�F���
��-Zp�DcM�"]&f�;�#M\'C�ֵa�X�n�P��`M����(Yl�/��+H$�7���5{$�@V��V˚a�ި�A �,�n$N����v(��K�1!��x����a��~v����z�XlxVHYEB     400      f0r�Io�7����P�(�_��!O<�[�s,�N��qihh!V �
�&خK{�8?�F�_��ɢVUC��s�pƏ[�D'0��|��՝Z�`�c�Ob�,恊�R�Nm�ƽ�M�8�y��ms]�(���=��Y�=
����.���&,�z'-��,X�^�Øl:8X�r�f�mOw~�,b�ە��MxBS�B,`'����]�����D��u��i��7�P��$Hs�?���@XlxVHYEB     400      b0�	���b/��%��Ku�X*�:����Rp�G�� -����e�c�J��������	�O�>So���s�� �D��5������7�㝞L1W���=uWϻn��~��rrpYܐF3����q�{���޲R��(�nȵ���H�[�|�ߜ�
��}�k�C��-����rMo�4�XlxVHYEB     400      d0m�&\`�^J�x/a���D�Z(U����q�	�59)8��1Ì}D�^I�I��ŝ�	�

�֏0������a܎�o$>q����J��u��v@�R��ɰ��?�U�N��V
b��cϝ��]��gK�RpVK[WDX��^s$9������r�d���|\p���0d.��m�p��)���+O-�e�v��������A�t�XlxVHYEB     400      d0�	u�PO��"ҍ�d����vQ;��Ȝ9�k�������J�F̫/E9O��>qǻc�I�]���^����@o>�E"O�?^�}���ճg9���I8C�c��R�3�4�;��C�l��
,�������K�SһXIU׀���X&r) ��=�LG=5sЄ�"�N28��S����|�B3�k����3��-u@�M�,ćXlxVHYEB     400     120E�(+�g�͔\@��x���e��X>߁�$BF�����-US�Y�lt$�O[� �4�bY�!�	��E�t6���%��p�.y�R�Q��=����WC-�˒��1JU��ٛ���R*+�@T`>�����W%�\�^O���UsN6H�gK��~c���YM9�,�Ӽ -�s��E�JDIg�?����p�`g�M�(���WZ�F�|�Ϡ;�X�Z�S>�+�r_��pŒx��H��l�>6����,h�˥���1cXe9C}��Z�7f[1LT���4XlxVHYEB     400      b00]��8���ՙ��HO�7 *���1Q��>a�?Tjx�, ��X��z�x�(�%f+��羷k���v�{�J�i+V�r��:}2�	& [R��W~�	�������)@�Ϟ�v�3���j�3������)2� ,�P�,�r��JloèRX+L ��1<��(�tg��XlxVHYEB     400      a0��ߑ2�	;v��n�{�R'	�[W���d]�q�F�Vΐv"����k(�D����Z�P�Θ�/R�hs�IWȡ@�m�ʶ��J\�3%�K�
�E�0���@ܝ�iVsj
W�M� �/e���&,���`.d7�zh�"|�sOϊ�q0�C�����XlxVHYEB     400      d0�����5�j\Eￌ���B���Pj#�/">�n��.�&NG��J�tUHA3��g����4P���g.�F���C��t[��4G�����k���.y�O��k
iR�jz|
I�Q����#ڼ�V��y���\/,�*rUA4��As�_*ФC�Fz"���@?�� ������[E7^�~��<�	T��KS�o��� ��==��XlxVHYEB     400     180�[-C����.�w_s=�S��t��Fw�����p�=���!��$޳Wp��J�˥�X"��Ȟm�Š��@�3�~�K�	;ށ�uy�I�a���;[c����^�����[��;����7E�B&(e!~�c�yr�� -օ�|]!�0���*[�
�|z�/����?��L�Δ�pA�}u1��O[��B[&�O�hߪ�wz����ʛ��e,�x	�1�GE夕uA�ؗ�n#��e�0�D�6~Ų��wY}>���owceD��������`a
������L(P_ߢ7�ȕ_}���
���s�P��T�~j���w�R+K��$ѿ�05��CWi%�Y:���LM#��J��x,�<|����j��~� .�����v._K�{�䌯~�[&^XlxVHYEB     400     1301�d2�f�{�tΖ5~����E}�ΉB1�w�������G�SR�$�Pѧ���7μ�Ӹ����g�/ޙ0,��x�=A3wP�e��;)ЊE4X'��G 6;��9��QX�~)QMC�5�;����&ʑ�uK�]i���'���,F������S�3��h��S�Y��(�U��?E�Z���0"vi�������O�{3��k�����}���E亂��U���/��'!	�����u�Gl����L#:�c�	�.ٲ6�K�2ld��uE�����7�bc���؄!�'��ꈵ�Q_XlxVHYEB     400     110>����� �z��Ϝ��nW�#��/��::�8�B�\L�xG�8�a��Fb�ѻ*z�BQ���@U��6 '��`��	���u�P*t��EL�l�2D�FJz52���������H��5P�k$��\�*�nk߶M������z�ix����PPת��Ǧ���Lu��a]H��81WK�n�/��_3�����fm���T��Ok�t^�b%e��(��4­�� F�dAw��M{Ƥ&
� �'�ăL�8�s�XlxVHYEB     400     190<o��5�q/G�� Ǖ��N�ϡ���v�L��ffa��^[[��~wM;�S��=B��:�V(7���C�`Jf]U�!����Dz�>hӭ�� 3��r��2 ���r �.�Ia�XMچ	��*�؜�ڗ� `J_I�.��uA�Ox㎡;`���=ZAtC�XƓ�c�|*ڍ�w�ǻg�|�f/���sMu���;���f�0n��X@'�;���b��^]�F����#�wπ�w=l�<���Kn>� ���� ���x���������C�m�!����Q����%�h4�<����f�R����(#&�?K�Y3@j�o���e���?����^���Y.��	ĵY���q�̗���Bik{�G:��c��{��%윶�_2�_mXlxVHYEB     400     110%~���#�[������J=�^����b��!-�+��͘]��z�m��4-���r.�H��'O�Phs��7��H��+�Rk��Qb�ؗ�B��P[��Y�O����j���2�ک���~���Q�g��
�\{�pW ���r�`��ρ��������le�0;��n9oGK�/#9=�b!X���̐Kp��������R����2�^\�C��:������Q�I��hD��v,�i�vݴ�>�N�x�5�]�������h�H�1AA��XlxVHYEB     400     110���n�r�����pL�\��ݪ��X_�Ik�@�KoR>U�̶������Q36�8c0$ͨ�s���� 6��
-\[���5'�
K��A6���[GAA$��;
>����D���U��}���N�8�l*t��Y�y�N��me����Qp�~�@��=k+vk
Ȁ�'�)J;�5 ��3�1M�4-�ٜ),�A�6���U-0��s� �%�����3�"ß9�a��}���~1��ԱT��v��k&�}�]��:�?��H���f��'7XlxVHYEB     400     1101�&ג$[�ǔ� ����e��.
�d��)�0ؕ��������
D�|��2�W�: *�(~%hK�2�����s\��r�/��Sn�-F=5��6#;�P4�%rر�<Ք���Ӧǋ��gY�#+�!��Ng!��JU�H�;a"���S*�!&�f� �c��`���o>vN1�Hr�*}̖�9�1܀E�W��y���%P�Nyj�TX]#q�s&��J��������۬4���� ���U�e8Ͼ��!�c�Tz��8�����XlxVHYEB     400     100�7�>�^����R��s%��%�B~�'Di �M1��~���M���q�{�W������l�V��1H � c��)��p�BU5��>�}	�<��\F��E]}�4t�1��e�U)(�� ��}�h�И�3gDÖwZ5�&�N퐩|;p#fLQLpΔ�(7$�%t �T�s���j�����#��  ^rĹ`y��r��G�&���^��0=ćnf�x�oR�N��~0�.N_���8��}o��?늧���6�:��XlxVHYEB     400      d0p�8K�N��a�ĠX�0�\���G��]�{�������>��P���~�K4�r<Q~ۙ��a/�O��	����d��g�t�^l���Df��%��C[�i�]v�vA�mx�#40���H�f6	��'��/�������\�b�,�w,wt_qgm��;G��8=�B\����iq�:C�XW�EmY��/�z/T����D]�@�XlxVHYEB     400      d0Z�=jZ�O�|�|*+�e�Jvkʿ�mNF*3]��0�Û
�C+�G����X����3�`=��
�r��޶���UL�+\�?���|�6Ŭi�r�Ke;v���~��|�Z�.�M�ӄ>sD�3*��?��A�K���gd��	�|;���]�"h�X�Sw����m'|U���A�f��|��(�L���U�K�=ƛ��i+�XlxVHYEB     400      f0 b
o5��%/�`/cU���E�����^�&�Kff�(�N��\P��-�Ny�k��D��F��x�9tA�;N�	�R1,'U]��~;OV�k!l�X�y�k1��-t[Ղ6`�����R之R���q�O�!3�NL�Ƶ8�9Ѓ*�\p1�-I��}��d;��`�wh����?9E�?K�s�cl����z��%��	zq�է;�S��`~K��\��`�֐�vݥ����@�]lXlxVHYEB     400     160\��z֖��p4\ܦ���:���D�z�S_\>�u��<L)���r�fq4,��z��A�j�����N�	��G�ݩ�t�%�G�t�����_�6c>�g�{���O^�_��L\e�v���v�����XՔj��#�[��/9I��XJ�/)�a�
��s�n�:�x�Ne��Qg��Y���)&.;����A�
�y���A�z����
n�(�قt-���82e����9�za�W�q�d0l�8+d8�2dp*��9�F(h�i�H��X1v[��1fE�+�𥞇hW���������Ea� =���/����n9�B3Y�J��1�P�J�r��˛�2
I�x�Һ�rt�sXlxVHYEB     400     150ui)ds�+\;�	0��3~����Y�k�Gt!Թs;�^(��H�S�&����Ô��Ys�E�+7�P�4��۩����?k5��3��n)�ѥ���اA]��2�ŝs�C>�]��-4��\z��d&7�q�`�2�.�	�+���4y*�T<���$a��V��Xa����e$<O�P��fHe��}>�����������5D�YT�z�{�b5����.M*H@�M���-AqV�d�V��0ܰ��7���',��9��2e��O� ��9�iA]��7R�Կ�@i��t�*��������7�t��E`$�H���$��8��Zd	"z8g(,.��E�]XlxVHYEB     400     100�qi�$�3�s�_�۴y���C�?��9�� ��>�TE9L��:�]�aA�}Z�q�[��H�y������@�&�T�i� �U6�ƻw�h_z����\��̽΄X���mӾ��0��� �Ь�v��=����eC�$	y.]��)e��9{<\���:��ҩ]����&����RCi��-�S�߻�&�n6	�:קJ�rI���i ��/d .籙y�3m����:�b�@%J�-���K�ta�hxXlxVHYEB     400     1406������u3Y�2&>z c�j[��w�@"�\��Zo�x5��/a�x�U�D�oV#)�mo��H�|�e'�]d��}��\�u3_Z>kwQ<�Y�E�QGi�(d�[ͅ뽦�>OhH�/���;�h�O�+�6�%q%ZD�4�m��Ƃ���Zy�� 3���e>v��Cd��pt�${�������8�O���R��DLy�4\��k0������~�A}��2U��T�)MPhM�]�	)�j3����U�C�N|B�F*��}��2��}��֪N8�ڰ������@�f>�L��X$N�*Y��2�����{.݆Na5�_�XlxVHYEB     400     140T��b|��/H�
�
������bں�Tί=����"���1$���9�b��Հ�mF��b�-�5�l�V�XKd~�?�מ�_�0"`��"ݻ FTpr	8�2���v�~I�Y�c�w;&7U;��/h�1���ᓣ�����&��L$�O�\�9FG��+�݂s�Wh�w�x�"���ܝ1<���i��5wR1�/��.�$��<ZS�Ek����k�3;�;���N5����>�A�8|�n�%�kE�{^	O�0��8�0��"���ڡE殫���M�=�� ���sG�|�~=��r�
m��#A�$�XlxVHYEB     400     130	�w�Q[{sh�Q�oX�~����L���C)S�%�$|] ��r���fP::w.�(� l�]�mr�}�J�O��1"Zwڕ�5H�%w��t�z��wy����<bq��k�6J�=�ڷ�e��*J^�1a�L$�8����ض6�u�}H����7a��~5��p�OAdkl�}��5'�Q-��H�p�y��L��2�0hȔ?�,�W@;�{�J��TU,��}�͟ʞ��я����v�s��40Yo�a�� /o4`a�K�ZP����&!��U�{�����@�g�EEu�J���D"k�jXlxVHYEB     400     120@ ��!ݹ\7�8�SA��Ou|����U�Y�uֱK
^�R�פ�3�\M���ڎ��6Q�V�8ƕ��h�X�۝��M�Չ�綣O���	K	�Q7{���WvpTqG�I���qV�?��.{�My���Y'F�5��e(@���B����v|���9J�~�Fv-<q�S{� �����J᫮\q|��(X�m{��c+C�d�:P1�鵔�4��ɲ8p
�s��i`L�g��� ���l[�8�����gԎ˅Q�I�2�?��^�������i��f��i�5XlxVHYEB     400      c0ȕU��+�$oFK�)vxF��x4\	��[�@���,o�||�V� �[���
�,�o;>m��ѩ���z1eI���a�j{^m�Yl��k���k�eT��PX����� �3�i�09__#�w����4{�;� �0 8~��pji�X:�U��k�2��5"�4q_��s��*ֻá���0A�XlxVHYEB     400     120[���_�m�}������?�q���D��;�=\s'{+Έh�D+C]`�F�v�J?1�
�(U���T BF�Lv��v^�79������f����R�T(����Hyp*���R��"$��^,G<�Q1W�~�IM�=6՘�I�ӎܥ�}��[�,���v��EHg4��c1�e����E�T��>���/�(𦄱��~�,�A2�0��D�}�z��ch��'+N��APv%YM9��� ,���1 ��\w�N*�"�k�8f�L7^�:�G�-j���`�߯�OXlxVHYEB     400     120<3n{�Rn?/�}d��b(Я���*c���tj��_�=d���ϓ�]v}u�����I��#	R���n Gc�d�$}d����&c���eH������A��^�#_e�_�M���������d�H1e_u,�e����7>ي�x?\�T��B9�ـe0A�p+
��,`
_4Ř\�3����m� G����SD]kη�+�~q���9W�A���Z��l���,�<ؓ�;�S�e	���6�ݾj�T=��nH�
���ݶp,p+aB�<���CXlxVHYEB     400      c0�<���gg�<9�џ��lF����Q#nb��b��^��Vt�9%0�C�`65�d���߳�^����{6��ߥ��?;���X8�ʦb7�:�^X��P%�C�-�L���?�o�T<�c��@5
��1��:nJG:���О`Ξ����M~�`	��nZJl�f	�븻�\�{y��MU��o�z�m|��L�QfXlxVHYEB     400     120*R�bH.������� �+��yvG�����4P��8��k%��|X��W���E�p�H'��z�A/U	��[��b�������,���ּp�����S�����ϡ�N��ڥ��u�M�?PdEȡj�d�)��' o� ��E�K��d�o���Bu������dh���:��V7<u qA���V��WR�f���{����;��N"�	�z�Е?�G��.z)� ��D��~��#.��B���$�3�޵EvX�v͹��|R����g�C6$ƙ_ީ!1v�XlxVHYEB     400      f0u�N��	f�ΰ�qs�@�,{���w*�X]�tK��%Yr�J��Tu��r�<K|��)X$.uR�J��6!tC5 � �	���$�,�t�|ET^�d��AB^�dlf:��sM����m��>{��#-e��� �EÕE=�Qп|;��MBc����&�}�ls�o�L�0q?�]Z�<���i�A��L)-��9[oFzk�(�J%i&ܟ����Q֔l��:8�1�e�&�2z$XlxVHYEB     400     110]�j��L��F���ÚT�h�NQ��V����nv(O�̨?��N!�BJ.�#�N'e!�Q*�g(bS=�3�������N���C�}��}zw�22��__u�~D��{���uD��:���Y��O6����w`��y��N؝�+���6����e=M���:�b⎩2��d���`�qK�'x���a�4y�Q�<m$:�2�r.8%ƹ5\�.�:��@���5pw�,pW�g#i�I��<��X�R4	�.O^����^M�TC�9mfD�i/XlxVHYEB     400     120���¨����b�f%đ�Z��\�p��)�`�`��A�s�6���{����>o��c�S2�� c��f�`|�ÃD
'=EU3 �-�Ώ puR ������:�X�|�ݖm����p6�]�Q���	��Ѵc&�\�ǟ�ڕC%�.��<���_R~�,vv��S��`9��}�3M�����$h�jV_s��ޭ�^�Z~�P�mUm�k+�YX'�����3�6���vE�+�NN�+^�szj�a���\�8*Kه#�r����_=2����F����h��XlxVHYEB     400     120�i5�,���iw�^�51��Ҿ�K(�/�h�X��s��2�-A�p���@���^6˯u��$(�y��Ŀ�Κ���	8:�{�5Xm�������
�C� �
Tn��_O�qK&�̡����/��a�ȍ��?��"�b�5�����)T>v�� �)5�����	 �9t�<�1�4Z!u]��)������<ʥ��k��2��U�o_��X 9��o�d�W�>!��߽6SS2���zĬ�/:9���#+�c��������rH�Q}�%%���;F���XlxVHYEB     400      f0��l��_紮�2��Ǫ�j�{s
*���s�_X��<vTn~S����9sE�ԁ��7@5�l��|�JA/ϧ����q�8Y���hRj��|��a��(�-���h%��!S�g
��;4�����#�
.�*2��T櫅EF
��q��_4ȢR�<#Yg m�#Ewn�x9
~��ye�V�y�ɍ�;��#�F@ye_���J�seBK� �5�����皷n/�Q�p` �|!��r�XlxVHYEB     400     130�ym���Z<ޜt����h��Uc)w��'(�Q�m�ۅ�fdCa�g�W��1NBb�O2����sLd�E I�����䖋�e}��ث�US��]���/~�\�I���ƛ<��J����=��\��@k��AԠ)c� �Zj~�v�O�vt���/ަ�B<��繙_U�B�q��n脀P
�����Z�~:�a��{'�C�-*I�4�@�(��;\�07=�Ma�40��@>h�S�9�5�@�9����FW�
���L��g�.Z�46K����R�����#�=�]��=l��Qƺ��l�iv��XlxVHYEB     400      f0A�ۧ<uYg�[���&B�u��M��݄#��;Z4�D��K��yd��%�P��`���C�?��q��,��_V��������ʤ���.��D�m��+P�f��d����I^����t3r��k�/�x���(	�׏Qn�� �e6��>G��l���[�|�KKۇ�&O�SBh"^{��Ǧ��Q��{ti/�� �@��}�םRY�����xH#b#����=k��	�
-$ә���K�B�XlxVHYEB     400     150��:���J'��&������\�m�Els�B\~y���l.���@m���?�G����0\5�el���z�]&)S�[ .�\�z,�5Q���`�2L�hº���e3?��bc���O�^ȃP�0����o3Wen��� /�l]�f�~9�ڲ���މ�8��fD��.ɭx��7w��ꦒ���⽝ǀib����y���	r���s�%-��Q���{'���JE}*U�qH�w��\܉�>1x�.!���/�����Ǜ?j�ɍX����&����Ґ�a�X�Q�G��A� .��0�vݑ8��T���rPo2C�W�|�N�$��DZ��0�F�XlxVHYEB     400      c0��A6�={~��[{�%h�rtM�w�t�"�q�ht� ;�>�yRu)�M���N꛼�Y������}�����@G	�{J���W����aGi��B�0��yf�]���礙�COg����M��F���`,��ǥ�R��)ϪT�G�ŷ�p$at�qUjȽ��5��Q��l�\��D�L^��������5�jO7XlxVHYEB     400     150�eD�$f�38�Dӹ[��ƛ�ĕ�|�in�C]� 2�;��o��ݭ2r]�E��%V�[�=�� �Kn��S`wEz;P�9v'�5�g�w�Q%�F���
�7��/��\T\��
t��J�exWT=��}�Nw��H�w��Vn#�T��ؕ�O4�����ѧՓ�vn���k�-�����Y?�����Z��e���`�n�cN�h!�t���|c]١8%�����@ ����OS��	t4W��PߺV�q��D>�js˹���D?8��A���;�?7�W��p���X� ����mL�%;�%�ܔ�<V����_�6h��/���  XXlxVHYEB     400     140r�N�vN��%���ti�`�	��Z�>7Ԥ����m_�Ϯ��*5D1��Ef���O�2��֣���I
m���m��nU��%�#?�:F�w�G����(+KP����'�-�s�*�#o�6 ����FP�M4�:����"�|_>�PNnF���� ?!��JU���(R0ѷ�@q3r� �5�Ⱥ�/N��~�YE4da��q�~�]B9�#��O�U��
(��.Pi����vSj$��d�@3��,�>�}ko�ȭƐ�w��}��8eβY�|��1YB�|x;�ǌ�A͌Զ�����M�%�1LE<E
�XlxVHYEB     400     100� u��җ�*��c\_
d�AɭrB*.���A#�C�$��0a ���48�xs��oFi�@�o�=KI���ߎ�ND�u�⿧���ƎS�[Z��ͥ� ���A �ǖ�ܬE�x��
ز8;��K�
�[��B��%��5eG�{��l� t%x@��ao6��b���h�g�.M�X*���`���{o�aTۛH>�W��=cc+�,���!}V��	�9KZ��{?g�x�i��͎o�j}VKG�4�V$XlxVHYEB     400      c0B�wk$���y����C���9��4����γm�W�/�� ���B��U�.3M��Ѳ03�ط ��NQ 7��A�CI1�+�y^ ~Yh�)�Ohϴ ��Wz�����i�Ř��}1��((���E����贽��~|���5]�	�Q��"ljx���cco;�-�ڋ�otp�b0)��c�{����qmXlxVHYEB     400     100�]�mds|լ��9ZG���
~\.=�7=�Vd�& ��4h~8D��m�,���u䍸�ޛ�h�B, �s	a��.<���+P�<�|�%r��n�M�f��7Q�;X�^��ph�R��7s���ua&{EM���n{m��ћ&Fn�<Y#!9i��i��c)�����[;�d��adc��7��������7�U��%��5/����Y��d���}�cu��6`[�X�Ha��0��N�<rӍ�Z�4FXlxVHYEB     400     110�`� Rmu�0��t���
/��">�a7�fQ��j�kGe�����TacV���0�DZ����R�Nj\���-1��Pb�[5{ګm�;f���d7�S��{q�ׄc����>���\��Ng��5�Fմi��v����[��3��v�2�=u�5��oG�������JSܦ�ڙ���`ּ����ےJ�j�X�O�KYBr-=�U���2|[j�$�Qo�s������aU�΍��j$��h�^ְy!G0�g�&�����Ad
XlxVHYEB     400      a0�i�=�<���~��_��dY�T��^��:�_��	܂n�o�ĺ����4Q���-��a!��=I��4�0�f_���-�&�(B��ڷŲUe�3c�b�ٖ�]�N�B�@�35�tN�����+������z�J��
�����	��)a�i�XlxVHYEB     400      e0]���{Ǟ޸(0|޸ӹ+�ҧ�m�	-3~��_��鯹������� [b�}FOt���V��[wE&��U[���"�1��8�畝��>i�h����)<�9�� Fek%�%�g"�'`ƻ%��p�m?�F�P5��ѭ~kB�4'��ܡ�w;ab�
.
x6���X7>�Z�QOֆ�y,ͻ�O��4�1'ұw��k3�6�ᡭeV���Y�t��XlxVHYEB     400     1a0�_�Q`j2^���ݴ/�]�d�� F�U�]�v��-c���s�X6�� _�7 DELM_^������Xbm�����fq����WMj;4A:���"c���# vb�,}_��\%K9lɧ/T�vT�Z'�5_��(�B�J��Y�'G5 yA:>�D��? ��
����2B��Ԩc{|���3Veރ��i�����^%�?���>8G��97b�����癔�KG������0W#j�ms]��v��m�vj!���S�?���6vܾ�o�&�ܩ*��ʠ:R���D���,V.�����0a�����2MT�W�å�[� ��B��/�(��J�B��a~ONE�Jf�Ȇ9)divx�c���l��u����*��x�6{{��)�r�c��C�UXlxVHYEB     400     150r��S��-Lu����֎�^[�X�$� �l��[u�>_��A��PV��I��
�J�D�f�����\,捷�~�D^��t4�.�1���n�'�B�����:�$I�����3dV;H:��I�Ȇ(A6@�;P�K�#kUPe�q/��q��@� ���A�Iiu��F���4�[<@�����I�w��D�a�>�J��׮���LIe�ϻ#'��ƶ7���"<�@Ϊ��m��DT�Kq=��[\�ř�(\�	c�߹����GVŹTb`��7����#����_:3�S�O7<�O-8�k� z�MYޘ��+(t���a/�XlxVHYEB     400     120�"	��'DM���*�7��M���_M���a�M�v�?�����P��)O�R���N��RpM3�hC�&��3���;g������/���w�l���Ń��I<�:��@����]�_�}z@��6�o�؍�Lғ�82�O���7G�_��b_�PΜCշ5���А��#�D���-+�����6�}q�1!C�X�O��Ԃ��|N�d�NK��/`+/+�ַ�˲�F�Z��M�@���E��P��Z���q��(�lG�}�C�~����N���q�e}�xzXlxVHYEB     400     1d0#_�]�k�U�wp���xP��S�Z
o��Ӽ�
ICE�O ��N��ܺz�l�ݗ��*溜K/���D�7ʓ\�+�ǐFgA�D}f�ڪ:�F/@�;��
f����.�7\�.D퐴 Eu��,,n�.T�(���H�C���Zb�)aMգ�Lu_�L�d��.�An�Ħ�Gu�Ƒz�9����	��vC��ҡ��&i�3VBm_�
s0��a�ѝg��#��r�/K��,a�?S\"��F��@�}h��*ؾD�_]�~j^U҆n��xm|�F�9Z�k�dn*���]�Lg�C��I����^�4,��,L��J�}-�h�ű�*HO�����g��؞�F�8�m�qx��6Ǆ�~�f.5�e+�;!K>	��r�G��R���*�t�H��1Hم��"_�x�����܇e����loJd� qU�	���B�Nn��XlxVHYEB     400     120ゞMJ_���io���M�P�-잸�yY���T-�H�Ê�w���d�����%��_&>��4��O�J�7P�\܎����w�DH�:���E�v��jH@�=*�5?�P�[��|�ח��5�݆�7���\ݺ"qiҵ��MɆ���z@��$�F�����:0>A�R��rH*e���%`.>�p�g^�c?Et�$�N�c"L�#!�U��ҟ��γ�<u(�#tCR7���G���f練��i/��57qǀ�}��]z.��	���j��%���w=XlxVHYEB     400     100��S���� $���9M(�����K��3�(+�垹�	�:ȷ	� ڿRQD�1��Zrq։��NBF�|I��
�QUJ�D�����`���
�`nlޤ��a�{�����M��q�g&sI)���-NS��$����$���`gp���)dШ��3��øN:���bwyau`���!���H��9B�#ɿ1o�S,\pl�J�Tƍ�OC+v�^,s�]��Ov�P����G~�v�$�v�\���(/_�Mp�XlxVHYEB     400     110~�e�os���'8��#�G	S �!��.��Y�vݏ@�L7�]Ѝ\�\��@��&+(��#�g�d{�^S�Ӻv�_t��^�0��v��]�+��&�47&55��̥ܙ�Ow�T5C ����b<��P
�@���:SS�Vw�5����3���!+���Lp�M<<h�Yh]�j��LVlY͕x�$ן�AD�{�7�yY<Z�I[N��F��D��kQ�M�L�R����͌'g'���ئ�Uʾ��t�{��.4P|�V^dXlxVHYEB     400      d0�6���^@1��Uq|)���:�J�|倾���o���$���eo�����K�@ �h���xx�e��G���|A�J=죦b�R*�eكl��~)|' �`����J7�r�j�'X IƓ��!��#IA��F�k��{�=�|�q:U�4*���8��+��S��ĥ�
8(bbJzF�̋D�B�q-��s���+G�M�s����SXlxVHYEB     400     100��f��T7�0��q�(�hig�����˖��(���z&7��������O�6�u����BE��z��\
Q��&x�iDq�i�����u�׊��n���)s>@ze�B�q�6Z{=;Mȭ�1��V�'�q輑2zIےl�>3i����]7�V!�GTL�(�@��S��sZ�Z��cK�������qTf��o��Ո
2h��V���ނ�v���B��r�$8!ȅ�ѣW��@w�)���X�XlxVHYEB     400     130O�-Y��{��a��f&��/܅�5c���y�'C}�V�p���{Ņ��P��y��a��j��c�,�k�Mo�)4��*�8��i?��7e�*��4���Rp�����LF�o�F3����]�SM�zxb
k�?v��SE~z9!�q��ߒ(��"��,�jӰ�_�� 0{q#Y�,h�:�[�D?	dP��U�YՉg�ʦ��%nc�h����:��S�W%�,E��د��i�".��=����, I��ڕ���@pKh{��d�N2����'č�Mg;�zmz�7'<v�:���+hXlxVHYEB     400     120��0K^p��U�Q꾃NP�x�� ]E�#/� �֔T��M,VM�דP�7����P���T��M�|�s��$�\��
�\bU����u���}a�[M��o����Nd�T�?I;��s�F�.O�Z�nG��o��=}�}3���cm!��۰�0#\Ib�\󘷞O?�"1��޿Z��:p������=��/�䢣�K�������.�1�iRtO�B��_��Y�{�P������.:y�_j�x����ď�	��D���1��ON,�u��j)IXlxVHYEB     400     1501D��hq�V����י�{b"X~���\�@��EU��%T29�;�G1M0:����o�	o3�.0�8,g�~���i���#�FZ+��8Մ���+v�����A��Wz��PJ[ٍ^�p;8K^��8TJ�fV���f+X�k��]�	��N�gң�|k��/�Ul�~*����<���S�vN�g Uf��R�gHs�W�mg�8X�&_\���O���d"��z�Ƈ[�4ÝR�4 p�k�($��ȣ����R�'�گ�)k_�����ňІ��-�GY�:�����Dُ�з���.��Ј����*̠������6�$\���Q(XlxVHYEB     400     110 �"��G����+Q�Y��Fƿ���iuʲ�`L��Qǜ���J��5��l�9:��?����BY&�Ÿ��!�O��R��~�Yu0_�v��:�B0uA�9e��7L>��7ݿ����j�s�J���F���%M\�L��иz#	��������#M/�rl�� ��д��x|��	�K�L�����dׯ������m����C�p�5N�L���G�߯ ���y\�P%��V�qU�pcV6�{f$���O[��m��<����g�XlxVHYEB     400     110_�8b)/�j����h���y�@�q��������`�|g�k�%&tF\*J�y��9*�2��28�:5����ʻ	�"��R�$��`��I�x��s]��zG*�r���*Κ��'?�v�]}K��n��ʅx��;�mNs��v�4���	�6�*u*�-G���M, c�%jb��2*q�U���@�Z�w��F�/�&d~_�Ki�E�b����1���Lwj=q�=��[ �"Iύ�Rj��,>ܨ<�%�b[��	焿b'�kXlxVHYEB     400     120���9�� ȡ�s#u����I �Y� ��e.^����ٲtj�����qo��/1dK�M�/�9����z�N���i�ݹ���'C�\��s�	�P��@���Y5�7�O��{>x�]j_@A�m�<3��y`nJ��}�p�ē��q�L)��FY��c��Ja��|:@Y퀥u��0a���d5�¿��tq�~��!�	���c�r�BsO��b�]^1���xC#R�����i�[�2HUsV��]��K:�nh�h!�O��v�{�-��l�v�T�E�jTs��XlxVHYEB     400     100hGP�����{����{���a��UgD8Z?m�RyPL�`g�D�x �-�dm�GJ���}-��z�|u|&�(mMLT�^���4���ҡk�k���@�:,�%`�ʽ����ˍK5H7�U�]*XY
����V�L����aE�J�h1��c�C�]%�����}lF�瘝���F��Ѵd^�$L�"m��d�N��K	�gw�����*��>��5c&*_w��'V��?O@wj�bS0]ᴔ��HI��9XlxVHYEB     400      f0�	�\���re��y;t��(��@_�.o�N���_����K�;�cNw�<�����(��"�Z�O6�_��8��Y�/����^�p%��dv���R��K�X���I�i`��xJ6WA��~5�X� �6�a�T���r!�|��?�&h�:p4��9r5T��J��wd�`��ы��o�	j7;	M�϶-L��Kh娶��
���܊�6g�O�P7G��_	�皧��F�����nߞ=a^XlxVHYEB     400     120F��Q?�v�L���|�32yIs�1��4G=)���w��
�c�L uCPDw��@l���a�	�o�r���[m��8u"�X"�7���nhp���ˍ6��S���I�n�Bdv(<גRZ�e��q�����|��*3
����_�ȸ��݊=
��
(v�D�r���9x�_v�,��e6�r���D:�!��7,��l� ������8|��VV�X��ը��U�A�#��������xymW��8��-�X�"'�����f�'w	�.p!L�c���T�XlxVHYEB     400     110M#!�랋T5��k\�*��<Ľ�Ӥ���}�'.�����$ː7���w�N����}��%���S���l6�~M�{=�}� Y<�W��H��vD⯗���gW�5�:�i�}�l���pply��ܖũ�S�&-�뀀s�ɦv��=�+\G,�Lz&�7[[-��~���5�ȓ�KV8'��C�d[�fQ�j�^G5��AO��������R@k9��鯬����Θ�<5)o�g{��ъ�y��vv��{D3��s����@SXlxVHYEB     400     120RB�iMn������Y���j6g�D� Q��n��xG�~��a�������%��RA��_%��B�&?�hSʉ͉���Q����K9��*v��T�y2)1�ݥe��l������
��:�>?�C��#y�E�ڜB��Π�!�'�wN��!�����\2����/�oJ� wO��B�H�Mن���z�2�I�� �����^),�{h�Q:�X�����ߘy�AGX�H<.qPD�7B��8��/O#��x�;��ۺ$QQ$�4��`��^n�ׂ�����9XlxVHYEB     400     140�/�g�%���#%�U���>��U�r���tu�$B+��!�y�6ؖ	�n�җ�*�KBi�"��E��.�
�~2
.U�?��J=}k��m^t.�Q���l��52�x��eU��Q�P�������M��z[��l��E�M��Qi�j�0��C7
'�Ղ;gw~-��:)�31s��8A-�&5��P�n��Ƃ>	���.-2���>�2�\�sd�Ҡ��]	i�P���V��w�x:(@�	�X�����rw�����k��uOÁ����1&&��z&��6*
�q�����"h��=��
�-_X~ 4�|�c��?.����&XlxVHYEB     400     140� ��C;�0�rq����VcC8h 8�@_��3\
>`��梏,rD/w���V?�Ħ=ڴb����uˮ��a��(�b�����r(�\�hħ�H[Ќ�2��J:UE�p��Ro���8�_�{סt�IF%UT�����q�������*!2>*���-�\%c��2���|%(��]���RV*{��i�ǖVls���p�aPϝ:�'҆��*K�'�>��{j����D�
���������kq��-��b.�$Y�����7��=��.�l�oA��0�_�,�#��
�W��$� �>{,cӢ��-PH]����0XlxVHYEB     400      e0�=�*t1�˷�g����f�]2�Ӂ�6[�o���S޲��:"�ݥ����-�~��Q�����,�}�s!��(���^KGp�����wŭ�r&��1��a,��/�ޚD��h�1�2�����8{H�<B�+s�A�B�E=�]�������5s?^@�ğ��'"�5d�;���8:b��%&P
����7���Y7S��"��S�y*4���(XlxVHYEB     400     1401�g�����'����� ��d�"�����G\�~_�<r��=���\��H1�-�b��E�!�k���;�)ZI~q+�q ę����w�ė\o&���菡
̆dm��[�@���|�W��# �y�H��A0�^D�B�^�������et{��O�- B��;�� U�KG|�t��@=�Q�u��Q"�*�AS�SFGkp{ �u����3a���ʼ�t�e����ԁ����\�|�:	�)���PO&��Q��+�3����~�-�0y�,0�
h���,T#�>er��!�_�eu1 ��wc=@�-��N���XlxVHYEB     400      e0�t����Ul�FS�s���3�����Q0���	���8��{ ����I�0���R*j�vw�(`E���C#�� O�`�4_!�}2���q��Z2E��h�J�s ڛ���v-%ҝ��|��L�/{���lO�Il���O��[�:��1�^pq��{L̀��������������Q��'�ԫ{����d��̞=	SG���I��<B�?��v�x�XlxVHYEB     400     190�r��<�U�"L+�ؕ���RnJ'!��NtN=�@#o�S�����]�O��;�[^���*4�2�o��(�э۩�RĆa�s��cN���^�f	�#c�1e�W���55�b�X�u�k�o��R���H��	cFi��Jt�br8���X��%��^�/����s�~CJP�}�1�{6�;�i���*oh^�-8�}�	�u�;�+8�lUz2��Z�De�qt��X�@,���gI��	���do8'�%�V���Ǡ��ǟ�vO�_�Jkװ��o�6�\r�ʂm�e���\�����������Rc�@Gz�N�$�"�@��l���F`��`�Oز�F��1�=�z���B�a6��,�����U\���������A���&G�Q-�H�j��XlxVHYEB     400      f0�/{4״�,�@P�9�=��� vM���N	�v�����`���1)l���O�n%����%Ե��ᯂ*��e�/k7���ؽ�kz'��,M���/�#^�zl�����k驙t�G^�!�-�n�Hv6��-ͽô�F��/��
��
�!	v�:k$��+�c�+/�U;Ƚ�![ؚ/�b��}�ڄ���㳹�N�H��f�j�?ާ�,t�p��4[������XlxVHYEB     400     120���mK�j�O�cZ�e�qځ�|ki�=5��ϯ����j\��}��?��7�j�:����
�">�7)GK8�0Üu�F���d�e ��� (6ټۉOa��E�RKZu8cN�\yj�b�4��'x�	�j�c(S�+^u����\[��X�H���� ��NW2��Z܌��ĴҪj��y'hqŦ�,�ю��n��=�w�^"�%���J��M���g��wL�ctT"�>l�[�D���l[�%��h=X������HpE���S�I�XlxVHYEB     400      d0�Q�ʆ8F�˂��C9�x>g�+Ф-Y��XBa�}RX��\���S�7�=qñ��,r���-��H��ʫ.����{<�b��Lr�8��7���d��E���W@,��P�e�����:�,f��·P[��S��5�ow��ߟ�BzB��r��ab�bs6|8�w�;����!1(�,͗�*�E_�����e�@uO�^��XlxVHYEB     400     150$7��"�@R3���jN[w@P.��ex��$Dx;�#�akg�\��8v�s��ߤ��\vrl_C�c��q���8	tK�;�z�WOt4h������$��/��͏x-O*�4zd6�<�dM8yi �U�D�~@px��Ĩ�ʷ�[oT��M*��%�67�G�����Ьs�-/ � Fd���ɧ��L��I��)_�t�kZ�����������H��}5p�J�i���To���3{�~Nj���t��2�L�ݨ��p��T�,t�y��x���3S��u'��7�Z�no��z�~_Zf
K7������Dϩ��Mx��"nEXlxVHYEB     400     180�F1E��+�rx��ou�=?�����ʁ���8��N�8fK���#��ۚ!��U	��B�]`�?���윷���XV`s(v��"�4u�����9$!�WV�&;�g�NuS��KQ��Y|�w9b`��c��+�[a��<������.G�b���|1#���N,�HA�E@3/�]��l�'�-��D���G��j9��EY'��*dJ�lO5M$h��b�^���nk0|��Kx��a�<�p�"尵&~`��LͿ�w�w�+x���Da[�_�l5�̣�v��g@����֙�r+ �����p�����y!i��1n�NevM���S���[�lsTL/ɫ����5�;T��1!�]�=c['}��XlxVHYEB     400     120}��z+ר�`��T�gȑ,���[���A��$���}>�VG&��&qڄu�T���QL�=:�<�Z����>�`vR\6w	@��������D�!����.�J�e�N+�l�
�!uv��O��XG,�*�,ʌ$�ݴؤ���Ş�әdA顂^X53��� �q�Ȋ޴ ���ɍo���z��3��P�a�� %.�P�3�:S��NW齂�V��v	$��?fF�g�|?�WV	&�z���>�Cy�p�׮k�6�K�]�1A=�s)��:�f8��>�u�XlxVHYEB     400     180~��N�;1/ u��F.p�H���ܻi`�s��ۣ�C���c?��c�� �6z׳�K�t�#�`�bB��+�т���;���B��^��R�Ҝ~u��"n�B�h[a3��-���+Q����Nq)^�q�������TO?}�4���F8��8b�vQ��T�A���{'w U��iq���Q	�T���
������*[S'���X8i!��ޛ�����vl�
y�=�Bn�fr�����񯬀t�Z2Q�D+��[a�A�x�I�N�3��=s����ٷS:�8Td_�܍𸄤Ǘ���+6_��&DE4U	U���Hn��_iv�.��o�bb��L���bN����ޅ�U\f�Cv%�Њ����!���̬���%lXlxVHYEB     400     120��Vy ���ދ��X��*���(~�4'N�0R�O��8�)Bj+]mM�It=m#���G4>�v-T���<E�&/ģb�˿6�����0��>G�irp�qX�� %����z)�UB�yB�y��o�}��rKI�PSg�s�7��]`��Y�R�K�
sb4�#�l��k~e�~{a�㯑h�,���0���}�s��B����^.P⠎�e]����᳅��%@
�CWA�FVu�N��ӧz��Y�������S�ٰ��TV���l�3�K]��&��XlxVHYEB     400      f0l��5d��|��c����Do��� ���V��B��O&�����;��ι��"&DNbQg���`���M���Ƅ�2��
=�;���'m���@��.HST���0��2��!��
��rM�.����!�X߇Jh���&Ԗ4�S��c��`�Nkm�Nޒ�?2�3��K�J6���M�k�>Q���#�q��%ߕ��;;�-�Ē[�7
J{���T���y
�Y0l[Y�-X��)�3kE�XlxVHYEB     400     130y��a����uX�oKbNk٭���K>�U�R�>-�=r��q�F:�Y��&�@\iS��ֲ7=��fS[���D�$��4z�o��Z��i�^��{�Lea3<s8iEUh��:�Ij�a<<$Ē����|L���ݖe�@w]S�gw�cba���]����b%�Q$����H�S���f��aNa�0S��_��cz���5
�DQ=p�b�3*J�p��U�h�����r廼f�s�3��Eqd���qp��o ���y?�H/� Y1������e2�7ZIބ�5�AN����hfC/�s��WXlxVHYEB     400     140F�eS�\�(��ʖ���!�:�q�Dp�Ql��K�0�c�7���}D���P�Ų�� !��s���v�j�;��gg�_8F\�4)�`�$O����	gΫv/sj�xɀ�;��
�!5�VRZ�eq��F&��7�
}���<Ԋo�<�7��@��y���a9�m�t��]�qE�jKJ� ��IT�j-�����M.]���1�',���,��{r�MO1@<ɭ�1*��@�\t�����sHRR���T�����:���QO�W���~A���#h\�I�I7}���e��1U�AG��967WI�tȾ� ق�XlxVHYEB     400     14038�}����CE��cuz�X2M��ƻ�6�'>������ޡL�ek.���9fC�A�;�]���s�M�H�����c������;BiOX�a]_iR./7����b�4�!��	x:{�}.O������U_��se+���g���,]p֨g�R%�C�d(fl#
���-��6+����A'��c|Յ�Y�~�����p������%�$��M��X��I�S�H��U�4Q����(l�ƜV �*x��
�h��k�g�Q��@k@���Q����m�x��I������	��J�7\ �r�U�+W�?����+��"XlxVHYEB     400      f0wmX*+5tx^�z(������Գ���,s���8�{�]�թOTG��[&1��G�
����A�Tӂ�V0p�l��L�}q��}ALѸdCN(��i
]v�O 2�a�I�P^��zsmګΔEgs��1�f��|#��Z @V� �:��!�Q�B>�6Q�H5��d�m���D�f�H�9��uf�uou�t2���<�����9$Sc�NN$T  _2ͼL�Q{���Oǰ�XlxVHYEB     400     140-�a޾��ƖI!W��B��
~<��oIɣ�{���i?*��h��LE�d�[oв���gw�P�>��ԧ��ѵ��4l:��~�ro,�@'}iKa�M�$�����R"��L����&�1ܥU���VE�`b��"hhϓ/�y�����VO��Y��f=��gD��e��P�^��NV�\�T>	JG�C���V���I��;�GÂ e��_�3�2�E�uT�e�;?�gdFUU�Њ3�8AuQ�4���B���c汕$���	ŧc\V�f'�#=e�[>;�m��|�ܩ�(��q���P��9G���i�XlxVHYEB     400     120E��^�t�z��؟ԅ�'�1�'6I�0J�W���ϰV��L����6�jt��KiRm�d᯲�os/�ܟ���ȇa���[�X���;1<�ɗ���?+�{",��@����i	�{��Y��Ar�Ѓ[&��LՒ�g��=X>f���]���	ũϑ6��j�����H.�dNUM�������u�I����>'��L3,�D��.�\"�0gj|c�a��mE#�%���<����T�h������Q�LB�9�>~O_��sL�&�7T��a���L5Gc\XlxVHYEB     400     120W�x7MUR?��:�)�ۭ�������G�x����|G�'�e�2�|ԡ��5!��]6�9J� l�鬧�&����
�]�����4\���g�)��Ǉ�AAe�l�nU;a��{�#�+/��J��)�u�
���@{���~<�*�(�� v�[�7��Z��.�wya9����@�=�d��R���RZc�m/�h%0A�V��UTJ� ��C�L�+�Tu��^�A��QB_��(��<~�RA�Gӷ:�؟�]���sk,®���s��zc3}�tM�&q#p~�T�
Z��HXlxVHYEB     400     110X�1z�S=?�*�5��Ԧ�߁��	�wo^�4�[��PY7R0���G�$��0L�1�i��%����\Wiu�y��i�̼�
쁺ŉ�M���hU1�X m�nZ����/~����w~ĵ�N����{������C,�x~����>u�W�^��o;���)ne��z�A�FH��
L�^�MT$��
e%�� ��-�x}�!"L�߱2q�{7��!����Q;<(��YmoqL�4EPL� �j�C\�@�t�;�؈hW�=�NY<sL�h�>XlxVHYEB     400     160l#Nu~h��1M��F��5����L�����:�iF�J� p9�K
tbw0�W��6Z��%�0������(�L�c���O
�m�^]\�٤����-CM�+�s��h1N��?�Ы���y�O��T��/+�� ����c��$9֐���(!��e����ѻzu��s���D�O�� -7נ|.״��R���rU)* �!��B�/K�T>U��
*�+c(1H��"u���>dA�chMxG���u��K7T�D�g�܌�{ajd�,S����xTe���8�Dt�#���Md�{k�PgS
�;�(�=��[a�ȏ�����c��=��O�*�<M	�d6��XlxVHYEB     400     130>�A�!����-������UN�R�>dW�@������_h�q`/O!Rډ�ɏ|�Uw��V�S� J�	���!��q"�<�vv>A�*�4ǊZ�� 5�
�� ����滓֝�2.�8�S8�K��s(K;_a��h����c͊yw$�S�u�Mn�	^�=߿�F���9�--��9n�2�U��|bEP}|r���"�;!t��r�+r`���
�P���C}se<vp �H�M�JN9�삉s_�����,_� ��|L:I^�.~�I����Q�-��m.� s��V;�J6i�Av�浨XlxVHYEB     400      c0kws8�3%�����m��~���hb��kJ�c�ɮE^H kd�1&�� C��܎HU������H��;�^#(봷�X���R���K�΀б ۶��#Yn�6��o��G6�
�:��w{�L�q���h�b�F�((�b!y\�)���5v/>�t��Sz�Iގ���g�����|�թ�W�@��w��XlxVHYEB     400     140����/��=k=Q� {/�Fj��Н�t��@i?a��5�7��C�5��٘2�뉒��񫶓�}ƉaYt��tZ�Eg)�~q�G"gȦ0���|��@k��&>8Z�
{�c��{��J�-�����0	Qœ��2\C�*�C����_�E�oT��&��c�d9M�?_������JB�L-֊�o�'�Q�/_�����;$���A���s��������Z_��R���#�b=!2�� �����v����
�!	��m `�U˴��"%�>.���t��NI�ȅ���/$��/
�5`�M�nGv����)gXlxVHYEB     338     100@��wH	�[�������Y����b�� ��HA�5����(«�T\���[�W9����k�N���p�R�u�/�}�<O����"�|���{U�';�<"����p���E�'@U�Syd=<�E�cu�Q��U�ҵ����s���٩��*�w������<R�x!ﬃ�h�N|�1�CǗ&pN���/?:n� ��$�|ױ��r��srq5?{� �m�67�1��iE۞Ǡ�Kϩ
&XR)��