`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11136)
`protect data_block
EuVOlWMaCaX23WqTo56ig4pC7p2S2ZbbuH+C+CELqaKfGq/uiiPvmldNF6zt0fr4O/o7070fMDH4
uSoDAVE7oigrXjBk9eq3cHelqL5uwwTKRKi3QbQmteAR+fEKkiKhGU68KhX3WevObkoQx+hRsSpT
fbqGvqCt6MKmFuKVHTP/PoBzMA2K+XkJkHrBJWdnid7gDLnZPSg0bd+l9Mo+k0qsABQRWn/+NeR0
88fJEKAQA7UayfCJnOuzoTYaLeW7vEqTFHebRmQ1nv1WrsgOPyyW4ZoeBAe3ho+eP1sW9ouVrSP2
//1lA0et1TP55aW7sFxCz92uWKg/eRPQ1/7xBCaES6xkeDMxyb6RXLJF8TuoGnM+sPgh01Q00GBY
H05Bix+EIJpIfSCnNCmmRyYrr3/oi4vVl51Acr9Y6QLOYQH+zKsb826BhEqbGPfGIWDp7sw+wjsG
725UPo9nogUywSa41SVGxwzy/4ruiZD/z0ho/o6MiqBYck0NhOsPR3mCxvUIsJ7PFWoYwFIvSxAh
tW4T6mPY9LJPF8pk52zoaNACi10NxgMIEEqq+D2zuAxx4vhfW/q7v3ifb4kKjcW/5nkZo5DUHLIx
1nCOk2HVn972MKxYM+bjZBFMRnKQRB9f8dTzLTt54OCYjgQST7liPoTsaKYgtJeW0H1BVMW05XMZ
Ou8TA7emEGsRpuVeCqrUj9yCv42XgjLDkmhd9GJLO6opgDgGlT8VZ9aNh1b2y/FdrhekW8BfHVnA
Y39qQTnYsYdYJ8Xj/ksHQZ752hLqTzTf9Hw8/9q0+EyFLnoXXHfHJV5cBQN2+WbjinZg8hXOEK32
WLv+HI5YFd/LywdbOfAuoZnrEVRRjZU+xrTe+HHNWnGBqdHrqQYGnp/EqRSgwyLsiR9WDHcBRwY9
0R/kQNGs1g0HF27uUnNMdY3nKKxJn9vvXFUvAzfcpU7fF0q1iV/+M+AqHfx+vCHycWe1QSE5RTxp
lgKmIXDel649JYfypa0w9o2+Uf0eIp4CFM0HPiix8ANV0hhOwZ+GEXrdp4n9JjSJjl6Uoovl1T7U
NbEKfT/RLBssJmakALPFik3Hlyg+N6UicDOGW0yxe3UGLhRTdNJzE/AnzmlzNX7K1eGxq8YLl1EX
AiOApbrAM6vjPWqL0p02RZqchvV/6PVxq6F84K8qgVQFUah45p/HOIWuFua5OXs6iHvii3oLLwKy
a7fpacIWezvGi2vpPCSEjvWmqlEvdkC+3FtiXza9ijN65ubgJEbAhY/No8Li8pBAT2CiU3y8sCqh
C9JIaKR074V9aK10maoBh8U2/Sh7v4ehmuKORrL9XJI2aXsxEci2RujvtZvh7ZEVAUPx4pGFohqY
ZnvrZrXEnm2Buu6TDnWmGuzfFqKZb3wsb8a/hIPvBw3Tle4uTyd6D1EXw98bLDCQ2+Xigi6heia4
Ej8GyLFeU6uBk3z8Js+srzeUFqwbVl1FPWW2SsamTaXFDmaQpA+z8gpFOiPtSMX6QlVfq+q3djUv
7tS+ZJCzRvae9kUOPusDVIcIyTdQUgp/ZaPak4YlUIanlZhKDxX8rCd8WPoLQZjq4K98ZGxbQRfh
qUA0+jtr/zGL0v3vmjWzftRV38AT/JyaafvWV7sgQiu+8FwKBPj6iN2gfju88zXkBdyKuhsGjBCz
01GAp877eMADjOE9KxfxupZ2bQqAZnUkfL+T1HOd1gGwzCo1wrOMW+4S5DD8dSXP4z0TwV5uJHrC
helvrsBBRM/HZOzPjnXMzSpNGxj3nJ8+Y6E+X+5xDwv3sX7T32KInUMNc+pGt251GEOuemoaW7k4
VzDmx5mYCwN8bdkfAenaxSIp134VLo0cwFs/Goh+Eg04Ql7S0YectYxbqmxCophNXDTcyq7rxK0s
kac5FqqIxbB7APHQ25S0LBK4KTOyoWScSoWlxcHvgUh0JNFriMGM28+MkzMKo2fZgfR8uWQrLiiF
6y4QGiEkjusGfWvDvwHACaHtKzmfqeG0227KHqFLtwZkOIQ4ZksVy7QrQB9OK1iMzjv55yjnMmhp
qFRZdqsNlPvBeubX9kkkegE7ckj5tunztFLLPer2IdC2NpcXB4FULmC3suEgWzyI4yifY0waiAQx
OEh5ibAnIjkrii5AGATSpP6S5O2k/hSlBw2+fsFB1+re4HKP13fZrU2uR8WCW3X78dgAHoIRqtHQ
20FxRW89rG6uUWhoCCjnCXi1YSqDiOAs0ydgaVNgqn55tQXxkr5wNcqCONvMQwLicti2VzyYPliQ
ULvAuMGliRIS+j/maTPIO9FvlmguF3RvdI1hpmHPH++Pz46+rJNmMvEhPR9laBdRDGKwS2JeCpo7
pFe+a8TZF3PhIWCCk0si1LezDkLbYsTLWjnUhSLhe1ChdBegUorWkp1oZjfx+FLjCGUHH+MbnREr
+G7N/Idmm/7QgvEZsQcLgSAC67OFFc96hVc2+xWoFPXp4NN93A2QxupD9wluHvvVyFG1LTK8G65L
jG0vZQooeuuWm4xr1uDIn8gwqMU6r1VMIF7WMeVOdfYgoGeeb69nsGZSSL5pslofJeDPSrMplzMJ
cRbJ5tfwus9uD50s6qOMRA/x+qf3Y1bOCU5Jk2g8nzMxBV1UyTc3ccEyfZLRc2aaXM1dyV0lA3L6
dMvMJ6Gu2UgfrZ39L3+ckzFwjSvgu1gTs279YLTHpuUnascUPbV55PXrelrBLADwipPORmEa+19c
lgVmvw38kgtmn419cF/4TrZbbGBhHVYcMXXUcZz25265Wl47RdQ+6+61Guo6FRQn9p6mhITWSyU5
37MZRJKdOCWAKjMFqlM4xpPHIws8n/nQ0nzWBCSz+kxET2xhwT+KF8eXhNF6XiAJa5Lyk/bRGS+n
1YOf5azCBqQ3FEyCkUJ8rmAEbcZrzYUPurJSFvyEMIs8HNLZikMENEZGvMMQ2aawphWskGYueC30
VQ+tVHE4h3txaDJYYIz6P1uY54nga8qorziHEiYegUyDRCsIXl1UlPlp71dZLPJx0UN0QWUf3EQl
IIgd0eRMH8FyzVa/bYOjpf/hqGSVfePryJRXNDQn6PKT4YBeXJ8deWEH52LlWJ8WT/KRotNwF2OG
cOEWlVNgQdX4pqvoUW8W2T9FfaOwcJxSaWdI/+JUJtpVBjbRdGAiAKWHKo5vGz/JM2hoZngeskdi
qKPVbcZqzNxqrHSxk98cpXOG1OwGE2efAEfEhy2CHZdOtCSzW1QIkBfqoeFT/o7uhAy92AFc8kSa
2FIWL+lfeMEzAsqOoKiEdN2/W1slb615Qt7lIW4Pk4vTIHBC28k5Ay57MwLxqoVogaP+0mM0dXM2
CCH05l28jL9XMga7lxQE++5ImP/cPTcsChlQBsjy5kdmHbMTyDix+odyAUHEK8yHv1Vq7L68K1U+
tDtEuwPexaGovvnJ6d9PX8EHM6ZqADhx+ThiQaSsNcDdy21xGZEsjOAxwuL20tZdXgC//hS7ZCBq
1yO/hfIWOo2NS8QZP3lW8CtvqpFCkMFMfJjqPYmCYdatTnFT1vZiAlWXCCNU7IPT4IiHRVlnCTY5
3rW1/6KSIuFEXHC71Eb4z6EzE8FFeTEx9FW4KJpaz1RghxTWdROGHCTmeFfxpDEFATbSSO0upoj2
4ASdv77MoxbsNwW3Y1bxno761ldilXcl1WbTlTTT6etnZz4GE/fWnWQTTrleQGDxIyNrsq0XPuQD
cpzlQnNvTc9XtZEsUg7/78qkPyZb27Aigl5qyGfe2VWkHUjnK12Jqfx0cUMglr4kXJploPFwGHYp
73aDNd/C1/m4S86mVFfnrhUqyttchlbOUfWn0lDhFbWLurWeRibq8RgMlQovuV0wQbFkUEAp0MYA
8E8q2FLo8JhrzwPh0uR3CHszU/PSGGL9HloL8YqmfQBsR6g7zlG6ua0UKKq/vG54f6gr8XEdnyUL
QxnhXy/4QVgjceEa2NI5uU2oPBVoRn7lWGgVkHTWwM/1pf16EG2pehJD6fErH3RftgrJTN+uJort
ardvjRv6v07VE2bp/++3rgFaEjGAWrA+Uj2sVRZmJA5Rlg2ct4q2HqFXzDSIK8L4c4FHk0gojSy3
3FHX3nly2tht2NbMFbaVsuzZ8AM4VpoCxUr2UX0VuhyFT8dS3DMnmWHFfEBNYLxQ8ZBvxC2LByCR
RbZS49VRnVXMmQDaxRc+WvRqbruwIfpsd5pnXBkqA7n55YRGLiixZTG77G/GdjoWSbGfZ9BekmW3
V6/T/c1yaHVZ5p/VeotiozM3RcDH8iEfkYSKuDBcAqHreTajGIz9+ti2lNzeSXki31ZjYzEai8jg
C+rRHIVV8eKQetGXMfOlH64MPSTc1V6pICUU3rlgq/dLU2RdJ3XGRJQRsfupMW5cCG9B6BMwN2Zb
wjQShCP6E3j8TrcM8qNQAJYivGOCPCun6/NkNjk3NWHqEIH3UxIp5UOwks+XktRNu7J44XJ+bMcl
EyxLS+U1vKWX0kKhKvFKNl6QQqtAPLmgoXMljDsKkhoFHoBjRSogW6osY+VfTx2kNv+Z7fTN1yiC
iGOrUlM9CRhixRDAPwq9mqS5lWo9S9gLOOCZo327rqWS76nTWhlEdUKYc2G6WaNKJMaZX3QrqMlW
s5mq3u8p2Ilar5hwNNZScmrAo71o+zNcyl9ApgtXrT+YiaseGdYBH9CmwJoZR3YkAxw8k24s9V4V
lGibUgG6rXh7ZbJQfChVwtttKJfvdRvtrEw+Q9xMtNsdvjGi+9HWf+BfAtdK8kSR8YZEhzl4gMrA
eBvjxj/i7WiJFQ73uZKXMqCodLOesjCBrrZlDnbfeqjLKAJK0N6RRPAFw7Z9QQbJeT0Ax0U6g3FR
WDqh/+tLgzURhljvpoDWafkUZShLqgnXF1vweERAvb7YI/mKrswgJtYrj3+TCNp6SNzLlvjkkxQx
shleYWE/BSc3brXJO3azpQoGnd9R0b5wn/hWqYO75gm37lcDrEyHqSpWQR0GmmuYEnJnbFHKfqJj
CpjlvTdYsI4rDlxfpGDuiv69gJG5AkXEQMoJy4xpuCmkvy4NQrWzKWXdJi1jvDOgowWtCKIgXwb/
XIQGFTsKujgkNku5MOiaCrgrlAs+WG/aACERlCz8d4wVhrCYt7ltalT6dW706vcFCrZOHWccedn6
HAqJS6xUpbr86RsGkDOR8w5L/EigZ6OBPLj4KvSQkmd9fGohszqCPO8qiLv2w4qJv39SvHJ66yGu
usFrFfbGQYHo4qZXOLgufG8S1NC4l69iDE7es7gwWUK0M7HOaFIz+HJT8GTgpUXipbJDQfmu+Emx
+Yzs/ySmCc/PASN9BaX4WD5I8N7a98iO5QaSETm/rfmkSo/L6eD0AYcYhOW6Okd9aMhRQaulGuwU
/vptZLu+ZpTwe6MQdVEdcvZtBAH9EJcoppL6zhhSX5fei5+RBdM7sM6SCHBxvjob6xmIaT6qilfe
Hrj5HJjVo95x/9h8U21WgN/oCohDP2Sj1wsZxDflzmUq8yVkX1OFm7Vs7EEc9p0gQ9jaKyHGqcAY
cQRnxISa8QvlD3h3qy5/M6uUk7j1TZqvzJctYrG7feOWnicRxjqCE5Lazc8zYDyuUhrBznhMRmIT
jVsK3flYtCGPrd/ExQ6yEm20FzCiqUU8rAnPkoZOQGoD45n+XMlWIInV7bAw2dWZ+jeSidUPpH3W
ecKY4hnzk4A8cR4KM9OGwLkJabxVDlKKNqWvH7f2gYNaUVGSaaia4t34JT4tqwEWpzIOVqMk7DK+
/P07Z7BWni7dyyf1cgvsFZvpz1Q2uNAZoBjCGbAb9LiRJPbt2KTA7A3u+cqp/khW+x2xYHBzuQyV
M6ogTEbAqnRyXAP/0AtXbM2j7g8xpTanZesP5TYozwYJoFX+bxFe9iLKKw/4hkrGH7cKOLAB33eh
dIzVJr11jdSpne5McxSX4etIKi60lLSFDgBw817O79U2Htl71ySg7J3p0947RdR9miyb6ye9XmfG
hE6petllmevtoi0CZvTEalJfpnNxV+w2P5nJRxxztpsmSOVeLThpJaf2z+tsNJf3UFbKhiC22b2W
ZlFCInzLaZaX/fsfVzyipCCvWJ3g87WVs/Wz4q+ckfBh/qrtReJN+nmabqzH6qJpmLwed730RSyS
BC+fRsemu5YiEc9ro/6c4Y++s/LOJMXiEMmDP3DVQY8iOVYHNtPo4O3vx0VX7eblygTil5rykDOL
yPYma0DkNrxCNFEHhGm5h1x/DiGNTuYRDrl0uXTMIqMpcfpoFz8wFVdERq84qTA8Abyv2fvSGl44
j0Kg0VbhSTmDDfM04Xk2YjLdi1zqG180hNEeDdRH9V6at9QzJeJFZKrMrZXWrvIPa8Def4srmdxY
egdBfG8PODly7uqsRj+ztg5ZjuSxkuDgOjBYT6pXh8lZPVuo1YQxHs5PNuqOn6LSToaSIxksQQ+p
DjVryokGaogZ9hOw9zF0S1ZjXgkSKGW1RfHfutr4j3cVmBifdcXdKvzd97aqh3Ar52VvA/IqYRgA
NtEw8R/UUgHRZduAohSRhht1nFQlxNBabE0O4s9OySnqbXHZ5RzwkQMHc7OQ0D/i1u3k+LnfPqV0
3S60JIU1VCp0J2AF1owyWghOmgsL+aeZTm8bEGUAikXeSG0RVBhVbThRqUlCeC1L7uGXWsnmY4nZ
zf/fS0UZA4Zjq2z8dpvbJDWmMINe1ffBX7T7y73Y6mtkRjWxJ6kZZ9r8S7aI5ihohjtIqmcFLA6T
To8MdTda5bHLLWxGRNOeOELq4bRelqF14JNZSkOk7Rzu5fyjnjjVcX9GGQoKmnCNRl70XqnchwZf
yKZAaPNc08EkCxfZ9n9HqNuY/QahljncPmjszQcB9dBvDw+s5tDLslinUxvT0MMClxAjwtXNdkTe
r0Kp1l1cfVKaSaEF7UtXV3FtiZhhsGo53SSzdcah1k3/xLyioMVfSFKeE9YH62KyXLK8NjnCu29k
Tp2XkH0HA9ip4a4h2YjEdss7Np332MGRX2Gvz64FdxjvCMmDm1NnhAcOG6kdeY/SCkrHF47za8pc
O/p3Nj1+hiFxsbDeiFnbv/uO1lHZb/V/gmigh9wilfvxgngq+XsvKZXNT//HygDyPd0XvYrXV6eA
W2WcWbrvt4w46r8hiJGnny/NYSnGWstNoeqwMhRbxyH/HHEAZ8arPkMg6NVaB4AZvUKtmx97WLV7
onf/uA0s00ka5gJy7/kG7czOXOhhEycKI4qlwuCc0WcW7DoCf3E4n5Xiapi0R1x6PXLwcASortPK
ugrgufs5/FdxLS042hdNMjkL/mOtKtiK3hovNXWrxWeGHczQinv1mwGQNMTuS7uCuX3TT2HFNooL
i/lW7nraQekcms4SM/wkbBmM/+i7MA1b+IkB1C1m9dvXquqyZvXZKbYyAT8+eMR5NRCDqQgOMPM3
b50ckxo2HUNf8d6+iMNWwY0sMQ7yCgPb5VBDDDyeAwCyOxgikOV7FAi1lDbfWEcW46TxQoK4zUAY
hFgV6xGMk+xIzhiRs6Tt0r6Vj8cFJ2d6Vzqrh7EApUieyAf7qeK4RjDRP8pfHa5iTu8nD/CFy0G2
9RS9HyrMy0aIbOCk2/AoE4CsOGz6kge89LDDOqW0biNs5a3k6yAFy+kAldKsgjx8WehzawHBnZyU
zF8fTcsSNCLE7C+lrEPKZ7shkMOjPtZzb+Me6l4o17TW7KMM9UKTjET2nLvAdEmpY1xTDts24rA9
yiMthRmVOGT8fUPJQobfT+VnrOYv+R4/Ierb7Yb40tCAv46ZZg1mnBt/UZ3Fp5KJeTklskmLFTjA
Nv0v7tHzEJakxNu8zFrGDwGv0iRtRQlS8yl9GtvapaZKfT/qgeQqFrNPC/IZ55oDG9k4LIJg2xUc
d6xSQrcLUufhOqe58O8e1QYrgrCcIqvTsMZQyPW/QI2eaTDS342CRJ4edgovrXF+fFk8PyKHyPGc
tqwzJ2b+82OHssAcSXqohm6ZiPQxEgAwKZLtcRO27nrYjL7owf2O6YVJq+eLFM5duY/2fAmqrdcv
K2bqqTO2gplvfO5lKbJOHM3xVoUIZGMWJA4NF3D8OBdqG9Rd0A7J3cR4r0yGFENRSAlnIOEDn1KI
1LeiY2nFFMIJXkJLyWXjc+Vig1HZpPLPCsh2nIGJ+Mq7ATI0fIytwtLMKncVHRlZl6QgHphmHBtQ
OSvQgJ8NxOvtsg5uv5mcmyVn0R5U1o461sBWtlbKA7GVaIK7OSe1DIdsCYVxntDITUt9/f8ebnhy
rNACci9biQBbxk2HxXvu+wowLt94ySf1Fcjp8/PVpxhwtXL+1mbNSCcmqWkAaCQdpO4znvpU+NoS
mO9s3IcwH+vYMt+LGK8xWHts28Oz2lKYEIplK3QwKURwsFsZRChNAdFuWai1MT4wWKRhTeV0GjNv
M89CbmQurDpWspzCkdpEvx3po73WV8f/+XmLpqU4ZED5lKAAm0NXkld6pmNzQcYd9EUqPajtKS4S
RfNjQ9/mo5GuW8GfwA5cR0rsFmak8ADg+I/MNENUBRCGOu13CHtwkWTfVvLIjjN9twa7ksi5CPCF
KsRMP9hSf7Rb882wAHXIzgRi5Z8FBAzmN3iv+p5R//az715OPSbO6ba8eo6BBDdvTK2CccPVmVDJ
RW56UBjGcqMgreWk6A/U8HQprTKlQjjYL6Yh2QqgVPDsVKQm9ILVlYd0O9c6IPPMmzMNOXl5VCKe
TPziu8Peoe9N9GnBCyc7K3c27sBgojZHx/fifsu9H9CGZ6+lPSSgLuZK1nhOiSY3PtXOUvR01l5J
jhjVWMCEfRWgd2V7MNeLjLggCYZvNrG3iIAlckbMlZ+4ZWMx9UMX32wHDQvXgg6XtzGesAlU1N5X
53XuXG2gJrC4e8HKHJXccf41EWHh4oHs3bI8FVSN1iYiy99E+BfssNo3qGp+H9Z306gXZW7jYafK
ALzRLJm+FZuEtrzegfAgxevHUAhp/bsdMeYb4IdLpfKaxrgqQTo3yNSEfWjXE0oI7PaViZoMk2X1
pt4GMm1hC3jdLGtonWAzcr0sq9kxZ6fM+RFzbR0P54MK9nrGz1FDyHc9PBJLr4HsFu0fNrhVbtRQ
m4u3I/jkECjBy1qLYHXVbY7/AeVq3wjrYEnDaZDbQvVaFEeBFepf/N535M+8j1ksCV3rI9fUItb+
v6MuEIPd2YgirXgdKXiF0bxV5pAB2f1mbVj7K0Rg4I5AObdMEDgEsetXnEiY9PxOxg+oXDANPY0S
+rYauJQv2Fwae0SJknvHWk9vnny/l0u/U22CMNr9zgJE8CGj0ZGO/A/kjW9lQqFRWWrWVsKzeyfl
ekfStmyxyIA/0JQo8/Tp1cjF6/zCHIwd9N4DJXsvpQB3EwHxwcBkh62Y+WFFJcquLLo6idQ0vLth
ion71DDcw7pdEQojp2G7uGMACLt/cqE5WpJ4hElhESW/A71DQDRz/nctyKyv5nAf5kc5c+SJaTvs
tLl2+FA5qOLXMU06q6D4oS4kuNbvAlTc0NpvsY+vzX+AjPdsOKaVS151Wmzw54H7tHjegpAhgSUo
Kj6XJYcA1IRzI+g9/s5iOH5X4dAieIKWYr8YziGN9BbdeaeJyVKkozOUDs/xEZEdzcyGmEle20Pz
d3B9G7tGh+yys28JKljDw9yq6+xCZj7J+0Kan3cXFQ/2y1DHjm0AzaFKyLrTHH2fWr3QfZp2wfPg
EQOAjkq42nykhgqPrUmzn8cXvYq/oaYVX7mqdEl4NTAlHlAiJuu5d4A2aDJDmxKlaoTFwnCNSwYi
cPvzlp7Ggbf/CEvSJF3O6uXPrdHaILsjIeTgKdhXUQOCu8jApnK6dQKuG3hzWPay2EH4Wld5nyaH
DnRFSxv2l19EZdjiV9kLo6tfz52Fk15qun87P0xnd76lZdPbSIi7w2FyzViKz8pvYdq3QGQBtBpw
D8KuNX/Cdl7KcFTbZV2l63TYL488+SnZP9Roi/XrouG/dzsds5/cHeG9HO8OQkhboKxZwCKVpXjY
bap80LqpOOKXv+8bCZLV+44wGEUWirH7yXdslSDBCuz/orvJQ7JVL1oX30cjhQNpDhdmJcKvDjI1
PM952R39BY0BIS87cxDKsDytlBa2K1XkmkGUz1erxBk0YGeXd9cpGeczDFk9NZBfG4b8jiIcQmSL
GIkUeClnXZAVNZK0dbDDFAazssWZkjQppamV2RnViFk+BLCCwziB1cEf85OoAgf5LwjWo4B6dm/f
+sK5kOveCdETk4PTntonSfXK0qqem/BXJ3JL1mjbDas7QQFYyReq11BFqa09OXeJe8mlJuMsjlzk
0afmKHXPquqUlz+/kjSNCNy3H0fr8X1OSAdU0vUlYL81zgG8PxzXs6zKuUaVOMGQJvsaQDBGnbur
WIXyTQW2YSQdCC/m4DKjaLrxZdqmHS0TR5BKO2ZFvDlnzpnVq4YXIUWR+1+1rBN9LMFQ7eKA7g+2
SWOJD0QWCF/lNx2RgEk7mQkv0kBaGPCaHQ3ojW+7JRj5CG77Axdwe3Pgp29ilFr+QR+elVhIgEHR
zPb3o4TO4EqtrZRgDFsprukLAGn8XHB+1KQgv/vmgOIWkTPyPhtxB7vuq+2SeJQe3kNXmDvY+v8I
fuxx2t4cdgPNZYxUya+KRWy6tdX6Er4FthtuRzP+Bk63njJt66AjeT6qprBoLBg78gOXADvXY4sF
X28CgePgzBAKvqRVHWWJVTLcjR9rko2pgSJCgOK/r4AsWzuU8yBJ+nENWASoxRUTBniaKJQ/F6Yk
s5fX2zFJLy8GI7sNJZQwxFrP5qoJ1x56xVuz72Nnqgd7JZhZK87vpNcpWaUm2bP6sJ47wJZAg2Cf
jm10f90KNl5uuX+FHuEAYitOEHV8NDP5VC92FILEvy4E5eNJjWtRgN6ci8NmInJtOQXYb/inRFLm
5Ayn9vRQfd5V+uzJRjW8Fl1P4UWdL/HtY4SBmgBOjoR9RtIR8GDBTk9J0herElSvVcV1M5QcbuSN
7/18j98J/idarzUPisUgvWCtelQ1MKLIUGvPAMTjTSi16w8ikhE+D9cbvM2sdTfdQHmCzl5u+7VE
mqpzhE1f/pfiW/rR+IV7SuJnf3ZHGbR6ES9clFBegbuYe/PCNBy7BFjywxAYr4zG4ArdxTcGMSDN
OZh3ZVgXptaOG9ShjnLJcg9JFUn9spCQdGTCKv0AxC7SYndfZ2YrdKZc58GJOCfsPn/0qqfgx+Rl
oFCnOZWhm8j5sgJ9+oxPMSk+pluK9m6uNlmhg/92vUuFEJTuIwk2V0UrXCTIffI7chCe4gKtrre9
FzI9F4P1EE5Jr5fDCVWFXa89nCFMev1h1nhzc973AHqh1MrPlipkYOSdc+ScxSd5oiRQ40ZAYa7S
ltCO/70ZqLHwoOlinu2sLHq6BWom7StgN2MSM8qq0x9co1wdsC3e680f3dTzZF98hooGpSiCHh5H
IAAOEPNCgJJVHtLC/UNX9yNIrynjLHLrkT4yk1CrOndNWmG3TtcSO/zoIPySpKymQvwQj7eMCff8
fTHDJRjkObOIGMJSfhwPTTTUFl+CLbBygpydlszrrEubrVgH9+jIKKIqUtPbx4TO0fZ5F8Pm/rI2
VUkH+kR9/4EUA16OHVSPuO+QQtcm+Zq4mF38r+LbaAvqR5x70gLWrnuVYKZCENn96xfw1HpGS2OK
WDKuC/X571HiZEBKPOZ4Fv71epuCP9c/thC5cjVTru9urTbdhC4oM5HnrHURkmqwsmWjrVw+Yr9n
6GWB4lWyrcs4vgrR69w3DPIYxe/NTY/p/rSj3HuBR95Rmq4BDUpJMsFgulICEPuUforoZkpt9hW6
uD0KoBbhvK8Yni7rOSxa3WmGR7NBDdowdAc/+t0lBEqQYRO9fEBBz6W844CxSPXe3CVbIKe772lL
A2n4UQFGnCa3wCc39NruZPiMKS1eZSge9qVehK9elSbehYwm/L4OqTm1vtefxxHiTW3SXXPIz38v
H0aWylgpbxeme6QAblUAMSojmgQA150WZuGWiSzbA36Sg/CQj1n4al20hlNB3kPfb3BaDE7j1CRK
CQMIUk+QIvWO/uMpmXVJxDY1nDqPnsl66//76nDWlYLlrGm8e22oRQlqgPAq9s2kOejYf9FSoSP+
DKO/wGOkSqaSXm+jD8fbJTo7xayhFhLH+w8TSuWeS+KrnxkTQwpN3lxlyCJnB4sMseVOzGH7NMeG
GCaKzlTMZkk6NezJBInRQmY94k4NdvApoiPAn7HQ5vHKQRxciNvzSADsbvduw1NSG3g4XTv2nps+
Rdf2i4Kq+MiNZArgt8f24BRzoqFjtv0InWKdseBkrIWkAuCBNcfiVhj/D+M7KEVoUPB/+pVnLHBQ
pi5gmnWOzEclebV7tsfbdC1V1HAEx9TRzNYUpYEh2k3sqpPcCaoysPJdZfEqaQfMYMzK3gpGRB2g
uDqhkwqsFn96pib+fFLwOtjt9rxz7ZseZi5SOtoWzamG37vGY34rIOqJGZ1qeQ7sCOhailgJnLfn
AajkKa5goO0GCO4+axw+wI+CHhIJ34KNAkxNZFOYqNplHPB+gOSnjghwJ+Qanz9UCIzIO4ABv+mE
TvBz+wrJHm2/QIuUKNjODQ0rD3b0N28RTozmZvO+ObyF59L9UWR/IRK3DjIu1NCyaIP/oAK8uQ+a
F+IwhrkGCD0Zd20e1PERLxVt/8QOvAqnLWji7Sw2wY9WZPpijDRxDs6gsEveaX/8BaL31WrgLy/F
+V/prtimcn6rD9MlF598vdpQV6NbXPi0c+VTROWFD3gUZ9Nw537Lsza08UDCYERlQMLkCzbv8/bw
Nvvm2c4H/0ERGzQgZkWZfCFPxTbulUBrZANqatsjWR2GJkBsFUCg6bKz2z9TSgKKD0rBLx86mqsO
rJUbfzphu57fOkfSNmdSiiSPE9kCTDty8KdcRnEVH4IKr9wtMMuhCNNg3BuwdAiC5vDeabrTRf34
tb5JgBJJWPznh9Qm75R++ev7v8Cw3DwXdPP2GE4b33Kdvr9al2ta9bDvGb9Kxi2Qs9qHksN2f1Gb
/Z9h84jTTNTwpHIG4YyrcCsZ+n7pZLf5W70beAMe70pzvr7X4FFSlHEUCPx8jBQKb8g6vqideYvc
b2Za1q9SJh9XaM9Yu97oXNRlN0cQxdZuIr53AQiPw18Pmu4KWhOGtqdCJ0EE20LQJ3SptcR+NXOH
ptj0U6B96Zy+YDxmSeaOzlhtH4qjmj6VCo1OlPqiZc2V7hBv7mLy0B6YEqdtqy1+fQrAXK3TSmm9
LvQoXfy2/1ttxGDi9eDAabLBbNkD+EtFjXHmbCSgeT3N82PTaZ0CPulBgAP+6O9WuEf41CvovvP6
cEIspqRlqJe/fIRMcQJkaxvooQ7g8UB11AQvU6QMDT7/apNIQgehNUumV1Agukv5WRNd27JA8N1B
kSQI9JSF20dnWzHSt0AU1SYVwHQwrl+pVAz1qqvLHg4FMSRTvfH3yO/fc8G3bfJNfP8aTnRwjCpg
ngo55Kyym9IKonZdGF74erbUhRm1rCX0K2RInNOgGGEQuwz4f3bn3Opdq/ZULpasyBLt5L18cUPy
zQLQSO1Xl7Vfyf21Xlwio5h6YJWS6uWxgNTCABmPM6OK+micAAa38rGP8hoQjEkoJMPdMWmv4C/a
XLh+oCQrkvvYUUq493WJeDepRe0ZH9Pqez17g1PGGMQHhxcCDbjZHPDxViCotJ0gVsxtpYNJAfKH
0sTeKaR9XW8CbAnzqvOliVg7mwVxsYscPbzLwrf2dsin8g9YiG/JamamTrCS0FsppW41bx00k91Q
igc8j+k7itIEeZus80UvSGq239DQcRhtpQEwPB+6ZsIhmlIvW1jSlbw10YQ6DZZjvPXdpzsUrWf/
4CTDKZxH6Agg45FlxtZewaX3eKhXRye5JcurXWMe1GfeshfUm+DMU0eF6ZHb5u1xmMCSRlbj6Mal
dVy+e4DnOkmoxnGWhb3Mv/dhon1p3JSOtxgCcGLIctbDWzwvZPoL+vTMk5mYSBeVyN2YuC7aQ2mV
5mRw6BVo+YZeJ84lBL30y0WTHjz7c0Yw92/+iaQ0b8qwRlBPOgSEP18FFEgFJc8SGX/Cb2YcdTUX
LpyK+9j5MKwcd8epOWsR4QMm+c34IMQFw9KEQ0JZQ5T0zN6ORG/hY4sCCishi9OcHBAOs8zo7WGp
YtNV1bfhi2LNERMXc4RFH8XO8HCGYqrpqJ5sWBfKvr0PLAqV8Zw/JPxcoi0geWPrxCuibtJJtv47
Ji/HBuxlQ1Q8NDAaYGiz0Y0ONFscIXe7q43UMYSR7xR1ODZsYBBcqE8ftrCBEVkWv/DBMMDPqkep
WtFQhD1sZmCmO/ESgSQvB5j/eopBbgOhISBu9+epspFsfavPVNlvs6ryjMENZU1GMEZX6sMbif/n
CqUFk0A6krkiBncJy+Ao1F4PHYPfakqkURsozy+O0gEnaWnfPFkOak61QSPXNNt7vkTfsfJYI52I
MfCHKYZS/8YHXa2wEoCOt9BMS9B/Vn6uUmfgG0hXj+iv+54RTCz/xVrRD4ELVRqLBWVoezw7i5NK
LVS5chMygj1OYPHMYQWIQMnU7aJYaE1UwYVIciq3T7bjZ+uVw2cvb/CHzpFqCDob8kqSyVj/Gknx
vxYyFff3JCYnYNfD9EA+wggilMM6pPvYQrnCs0x0HUnsCHFj9a29i7Exd6AgWtvbcqbrIGa86nyt
PHe0J42m/zOWZgBevJWis6zxzDvSpnaUq0ORvR3VkOIRKEtym7dNpAEa+Qz6eCQPSsh6otf2J3Gf
kHMMFgyNAX0hsctQGs0utygjg0W2
`protect end_protected
