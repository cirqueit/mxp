`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
2VGtM1DB936iBpafOSZ+W9JO1CU2ndTm2+FCYCWaYH98XW0eGiEIwyd+8lM0UgkxyCEiUhy9D1nV
D67fsr/dd1V/5Ca0niLu3m+xSr1UkHPoi+EsHsyFAlxezVNqJpROG5OMUcG2e0PlBoFgzxcDlr8d
eONT6G/qjbOqZ9jyVwvtbtxhwm2H6SlebGofyg9HqKAqKCU2WwM7tbXps7iakUlMpUJDiE8uOatS
Jj7txMG4fLemXdaqJxSUw/5KUKUK1N9jfeYZ3hmP1mTJltEmkdoaGEpQZ6uD63C/Xcn4RxJKiFb8
KJ/7BiZlyiHeONJ8C0SoscKJispjM0FBon3MQlkPRKmexWFLw9DQwpaRM1K8VD8yOYliDaPKEKxS
ub2IL2J9/AxxGzOeZ8H7qL1cC2k7fRHDZUMQQsFsYaO6OeBoZwTyZYYYnAqzj1YYKKNaPZQBEiFw
XwATIFRa91hq15OGVxNp1aRSpEiwkqYEh9L+AiUwfA60NCSUxggku1McYjw6Ztztu6ZCGkeOwjtI
DsrVABfQ1mcMscuQcZe4T8ApgBmVNwc4ODtQCiOOgKIsQNfmyT3IJuxWzIjtGXm7kx0UwF7Slqgh
K69ZkARL3WWKABjLZ65I8oz8kP5r4zwB3iUXbjaIV7aI/D7Qz+8nUob5ULJk2dsygxhjW6pD9hiP
MrGfDyUxv2WcO3Ngtb+F2VqoKzX6j658OkKPAy6UfVzd48PdnHPbz3WEcq2Txf9CsVfohZv0wGfO
e11aZzpC4viGsPxjSmFD6zthyOvKbiKUUd3ANxHt72hoW9uY4Hsr/HHuCaevipIbLI/faBHT09Q+
Sm0NEf3QsQoDoAC//M7OS2dgBh9IK52mogCTMsSKIglIi9WInxfkN3G+e5jsiiN4p3XMZQSA0729
gTIHTru3ynlHiCVWPvRurL3n1yoA6qh+yRcrBB8EldiF7rkv25gYWg4wWn8N5egExAiWLnDzFofQ
2jWrDfPGyn81iAkie4d1U0YA4opQfkVF6LeSeBfvJkqQ/G+stNKaa1XkE2pATXKUhTrfYvKErwfb
OnYpKiC+p6y4vlmfY9rKHPcV9Gtf9x3yhHs2/py0PIcwE2DokfDgPiM3EvQMPGQ68XsCF17zGSQx
7XGftkYJJve/hkEGnAWOZPV1F1WX3Zd0dvZAsXRGcM7K4sTUj20DTxIjE/4mv3g98AZkHH8GxUq0
VVk+eDUZnETJLz0Ynp6bxMJYdj4Z56fzpSA3rgxMG1lfDmYR7WSwDezdDXD3O3trrqs9jYsRf/Fp
lVN1At0SVeYC5poTT+7vCZB/81opnYUpRp2Jgz90T1EtTfWFYQddB5/2Db52XBwzbFoygwrRAuys
/Rgs8wqGt2pTNZYKcmqau+l9mC9rXEf8f5dSXVrpLUhvWa2RHjhjnsGLyPqp4S2OXFOPsfjAizcE
gYOrjJ0ReZtI84fpUf3DGSJCYIgiATW+m6a5dmsl4P2oFnejHZGjR5ciXtFFONTxl0spxRS7yi+c
fmzdCJSR+hzDJHA1sPwmV2qrN33oKpMRrL6raawfnJi2LfQjsc/fxC7aoStkbfMUML8BeT31pV5g
Eblsew6CKQgp3EkLavA4ElbTNFdrYuDdwANT6MGM5wLgl/ehbEqX982WCrM+C3izGIFQJDZvW3+W
RkltH0pz+auX63GTsaYndqp98WQEDDf+zAs3QfejaTy0G6zyeCwbt6F0MMwm6HSIhUA3iPCUnvy/
//0s8DNoPmW0j26goQ0/6nTJ9nqQ9VyP/1N+3ThmKqkmhKfLy62UHbIvK7pNzFOKoig76VBE+TOM
yVqnAhYHMbYV0bJzXRIJqw+XH6+9mNe+nRs8YO0TStV5LVqP6ENnyjyrmDPgMjKjo0ktavz5nWBH
6YdkpgueZ+7YWGX1JF5yDf8dh9zSgXOH1Mxe+QfgqaY1/X4QB+2rhui0jj1MIHlWmLYIMjPTo16c
VAgWZ8GlMt/6GVyRcIGm5uVa+tMBI3Y3JiVZxZlJbORRJYtwHaPSgM0+zZGcRnJfLIj479hcod0s
A1l1KvPGcwEKRqx+NcrtrTKl/yassacYJM1/u7lrdugA1uWk33PQvQ0c3SqLVB+nfETZdh20ZiN1
sNU44MDqSZ3HMPovi/3lS041vtPmrkmkry3PHqBE/6mQI5Dd5xw3mDGuNy5n9jdzMgTC+IhZcPyB
WxVLEflTJwrCaArJpVrVUIu0RHEoA/oAgGbP5NKgcVDurYQFGWz3suQZ38MUZR+SOmrb+CPV6oGt
2I118oY06HvZdKw+AbfQOLOk5TNLV+KW+/oGTb+YyIVn35FNgRkp8seKuauFqyZ6hnRJnmXp9Y9t
wcorsJMRAWz8gVEaHsqBAG1vSxsyKIj8KUFrHqmVcBo6D8q3+FJH+sCzQXMs7QBfOMaHpOJkLH4e
1qEOz3/JDiPBLup34NxQIyeLtanjjBOa3oY/k02DZqm5cblfFfs9WjgHhz/7snzvjRdW2tZosKlk
PMxv2ySMhD3333ueosPG3hjkFSS2svSJEXDDFey5ycIxxqFrRjQnlTS5R/CNUk8Fi3pCW6f4+u6W
Eg4I7W/0CPo0cz1pE0VYcEpxXhzvRGIcS4t5qpZi0Vrhfbq+jxZuKqDyV88OJlfLVa6Qg2qKbtTg
c/G1zj/vZYFt0UF2amRCnUOgKUKCmpB59K+UkMJb/teHWE7xPJaU7rt9whEV0Lik8cODQBXm8963
OZx8DVwflHWR+wM/EBQRtYmRiK+6RQdRh0KAKYveHn+blJcS4DIF5gQ7O5C2UExBpQ0n9ZyCz9Wt
TyJYiQu6b0mrgQvz253MFNtrs83322kynNwFWfG7In7emilGIYfGe4MTTa39959vVo3+
`protect end_protected
