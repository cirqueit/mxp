`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
6TUfLXDFyyT+JkEsdVgMdy9BzCR4cvjqLOZNMqXr+DJG3vbcDlo/8fwjVkKfOrVLX/F2L820OsPr
hUPXS9aePAYHErSSU7WmbAT2Nqyf60HSzV3SEbqJjDSxky4Xu1usyiFaf8fju7n0wwLACKLnkZ5G
RnxYmhHK27GV6QOzPgrRXd8tdi+X1x39NmAx8Mccs4CTy+MD1qIh2FrqN+exwnfdWPXGGJFB2DN3
3OU2zyx9LGSFMSfokkEJFjt7kwSlPwGaFSzTSwOFBgO69n94vQwMBvanlBXH/OM/QdBHG/N0NCaX
uyDk7LAxU06ie6xO/mwPjzoVsH5K3PKILfKSagwoaGo5tAyr14HgEAO8NRuqjEWye7DKoSr1SdDi
7QRmH559HyiOZCU2rsE5T3PE7YaOE7FJldEAb7MlGiJAQn8uqs/VMuxC8I9TvbstQq6mNsetHCVO
r+WPHP4xuHv9K5/PHjYf/zyuO5VDsBWG9QLhtA5pxO/nw5bTaQlXsk4nmJiu9GnZPbYtu6nKSRhv
i19ybwgK871hxvadSG9s1U9n0IHrECztMw96Gg+WVZ3eR8U9C3AW7nQimJLMyPjBhPqMk9E0bcd3
UQa4VTMo69mGOmlRdf81mCuK7HyCwxK5K8e5mRdKp5x01+Mq6l8NuFIzsMyk2u5PbHu6kicE7HMi
zrDk868iLBmGqXmgjhjjSBVl5+QjA47AVpWxjG9elCv4AfRv8YmDcQR2+OiQSz4Mwk6/Q5EDJmb4
Pca/cal84jCxTEOP/i2jt4d64S97upa4okL5bh9yKIVt3UH11stw93wOUGF8fwlcsoFDj8OArn0N
IdBZs0XTMqppLRfZ2W/KzbXu54QxnUGs2dycRWW4Vn3FIy7ggTZdmyKey9TaqcelkJBHPtP+7pxg
YoFWSSK00kqJPMSTnw3o1L4Sn/N2HPPM/2w4pkovG9PZXos4AvpvzAx1cGeTOv1Hx8MvQ7b3Q+1S
/7VpNxTr4bAsjbV8a8VQDlEqw17AnOjXm1giv6MJRU3Zycr4LoBFLyjvIWp8K9T2C29cpRyon8AL
nkaTLEVR4izT1TW72aJNYfRY9WZW8TSRu2VbUvT+pU/jkBxBxllcu6dNqR57GRXuNM21JDsypG/B
fZqB5tzWj+sneFQfJhYV+x3u4RPA7mKxXqiV5OlUKYJPzoq998siDvAGuKDdo0iUTYP6lcbHvTx6
kUuct7sqmfper9/5TqZpj1wsqt9vujn7MmK2gxKiG8HYtWtBND6Biw6DoV+2bQqfBreYCmMz2AlP
VJlVS82ClzTrOaf7aSe4Bwm7y74e2IVJ4M2IUhUiG1RfE58XUUe4we+7cGD4Bgv76MZ32fS4ahhu
4BpUNZIwhZsC9AzDF3sxX75p/Ay2XBduG5Fv1RqgCdK2RY6DPugH1s2Wvdq/lzFhchsdr5B6AwuS
In0utTpAmK/6vTrqR2KY8yDKOTERSJdzpBTpMbdeIiSqc6/I4jR3mGnlWGVZtShDoNUZamFofFBs
oDSH2sv2H9F8Ye7182otJd5TQlo9CNSa2cYzitlkwHmuL0BinKP+DASm4E9eaBVehXwSE/Ddegbn
04MFSQF5JPRniZm/2Ep3RAfsxukOSK3kadaQh9mbYnZglYiKpNaRcJhZXYlpftSUOx5VMo2Kv+Hm
am1vTn9Li2bChMv/dY6Y7YAKAEzeKQs/n/LjLOIZCmQY+eGqVH/c6n42sW7WkZKAspQkaNbw78xF
ZwnxfQaZsCf9WIv5pW71kRQO1CEgo4R3oWnczCKnVHtBfrUdhuAJsivtWvUdINjrhtZsAu/VM26o
sh9gnk8McFrQInp8eKpWJ4AjH530raDiniXa1Ao9qK/AB7w133rN5QHvIcdVO66x64SnNRsRV/pG
NaYra1u8yOqWQwLnZKWyfRS48hFB9DrC7ODqI15BdjjluSrtC+tpDutJRZzgT3wMHlb8ZjTAXT+Y
THm8yXEixYsNvvmAIRpqgBHg+xZ/GVkXrdMAMPu9GCy6xeb7vX3LIRpBqMdDVqMoqUhfJDYTDgr0
AXb+BHxsqO/uuoef0kekx687RKPWq+iDNCfdxD6TnCW7qVHoKROZfrOVzh5pYZCC/cYVV5V66kYv
NR72Pu8WXwA8zTMLeylSIHz4QdDbvmiaXvKeDpVu9bclH3mRA/v4+fpiOzXHGWLqBlXCX3oBIvuA
EKjTT5UgXZvSOmLj5/Y/3iz6ZxzQWQMEjR4mJ60n4TelIMECcSVZ0YFQaxdb4A5bWAdqWMgMWuNB
VrwFfOo30yys2nkACpiHUMBbii/RlTcl5uz8DVbMZXW4FJW5QVVLUUNMGwp6fbt/Rl05jlcLKsEy
i3S3XegwFMut7CgCRRcbzvH1Q/Xk1JXsV9Sf8ga7fzMGG178FGmqOF3FgjnRGt83hoxlt9Bd6AZS
kcKqvD+8U689eCA1ZEWCVS8vrYI5T7oTZhXGq8Z41SvHJur3KPDAvkRGcr6t7tu0S0m4bcKJ0mm+
eHK5q1ARvbFWznBtDZcIVQxYSEHGD3ahxJNKIXCTxpTlhRdt24H0UZn2xF46kKRNlfLXhmLE503D
BT3i/yF3XYNDbQpQ1/wAAxMMmnhtm1nwZ6W2KnL5UOuEoQ157ZBGlPk2eEjuVKy+vN6rk/Vbo/NB
hHEn1bKNUVN/QLL3llWdqUOb9+SP2OpNCKvXhZ2hJsH5Ly6Y3UM9G3XJDFSPvi1wmmzkirbKY0XL
9gII9Mv227qJMSwSUSt3du6F+DIVfAilQ92SGE8eooloS+ABqlzZdK0c7dO7C/YCVkdi6WL+6ZNz
SpkzygQRt9Hj6ssQd6Fnc8CuopPxqeJE9q3+Hz1NQzAKiQyrDHSrBAPpzN/Bkp0jbXoj1xU/d79t
8RV3zMqUDeDnI7dNyXMkynaRa6TWh5qoXfvylvLQ9xTstqSZxskFqTGLdP9jv3ZcLyOpHnLxCxyS
o0Ao31kRdal4KzdKzfIftRn9NsPJG/Jpk+042NL9aGbiQHSJWPK7YLLkKXKhpjKrh2A4uWt0ioYs
GAugk9azPJSFvZgtz8/3D19j+4aZ2AiF8FR3Kp6MDLTittF3kriaPEA8GHf1eP+pBxwGtpn8xXLT
uHDRTY3sBtuONA4OviElBdaM5AhJoox0h5G9894SekFXL2a9CHumps8L1nlfMye9NJCz3aoX0myg
xggwhSK82MetXyjUwBYwrhfehg+38RH+Hs5gYnS8blGZJR8vrA4Q18WJbZfWhR1Ic7FfEgQzxgFD
1ldQQiNn9jbuumkd63Xs07C8eLM/0xYqz+kVnJPkQcJqwYp4t89NcgRy8lNw2FNcuvANF9mNG+RN
3C7ylzJiBxxRpVmv/eY4CXQcmACE2gwLnBDeFeOHFTOWfAbOySyQT26rKpkipYocVvJfp09qX5ew
f1JquaBfcala3/IV4+lDgmupXfSWKMG8r6f9w8QQ4cOzSzV8iiTUaqSEGeoV+xJFWY0qL3qcEcXO
0ejQV2FENGdDOaXxv6I2A5XX0TfEiEtCV1i2DfOpw3nGW+Ku7vxJQov0KsNU0ozrkdCrjXt5Lmjf
a0hkA+X6UupPcpH9f9I+6+nAEtSLL/2G3xrvTiO7SBFmg7HHZwlYXOMTUb3oQaR1JIxw1jyETimU
sEDAYqrYIoym8Gd3eA0cTt/QFJkf1Nh8QSAwnBmTiqIYNHqx5peyu6zfHjOzS5YKQu8duoZGp6bU
ftnHPdcl7H1rSJOd1MNk4RkgxvKnF4n1ZS4J3Q3l7rN4rkYLsGNWVARI2gJbSQekklOGwsoC8Dxh
s5wHx+n2ALUzdpRlSkOioybJvDZ9k9pz41HZbIjRZ6Oa/GzL3Ho0YSClen8UkLrRT2/kOKyyOXYe
MKOQaVAwgwj6XJ18Z6TTsEurUJPeDHmp25Nza8sTybmDzggiGk8TCxgmuKYObICIDvzS3ZRE1B8a
LErJmZnrlsk5ZnrNrMqedaSzXaMbm2LoBg5fkZuaOsIcL5ODN/3Q3HA7uZ4gqz1hObNoDxQKdV6m
Xh8hAoei9h/9Kjht6vjg1Y9U0aq7o6vOqlM2KJSMj8KgQKmgwcAjQ3/rdkJi2rS876U1E2h9WijS
vAUMGb5cg8vAcADxWGLvelkhi1Kp0tX1qVlRDgz6Qj7ztfc0Of4LdAKN1HCkYqIkAwSPtphlrPa/
nIxL0FM0IlPVVngqMhUTXX/8QN1CAxDcb8AkSeWr/cPfWNzCPrXBI93tah5XWQIjsCqMmcc0ADxe
XZKPqkJh15JDPT/BezUl7cWuLot5bNl+rQDoY3rlx/WNv/sdyNJetGAaLPH5mnbl7WHERJAeoEVj
dF3Pn7o5qe1JM4i72f50iiWoiaF2TsaoOrBBAJxc1yptW7dXekTAC143dqgF1o9dtEElB/h8y7cC
DzPg8RgFBQLxwwC8H/P53erpwjNQvQNkaFu9rTlZFlla9n8Ci3sGI0T0Tpth4i2W6Pwne+CbTIPK
hJB3jYIVvMPv9+B4vkGm0rFnUbnMmoEqfCb8SqqeAf6VQNS3fZzAPwtZN1nSFgJa9zvqvYbJq/Zg
hp8/xI6VEuHektVYphmu8CNvfSG20llvlB423bni2rOMuy3bqjOBvaA3NY8zuGFXrc3opwpzzAhN
KwK/Y+szi1/Vk27T47VrAUC1smOXveOpb+GzvSd5aMJS8GZkuoFb+E2Libu7n7Lv2HxyWUSaErF9
nbTZLKz+5GvwtsaYq3Og31FpX7kQy3L15qxMraSkdJZw/+FE38+aeMuJykR8b+qGALiVl8sp4Opd
JMy8o/Rm8ZI2GozR2r4egq5ZSwOL7hYH/cLNVWg1tD5Ht3PQ2tkzKEg+fUK6Sl7C9QUVleopkKaX
Hu9WzM+tsC4P4zcq48Th7/8yJNhtfJiVKXaY5cSWMH2hdpHZglPdRvmRO0StUUPLpZDso+5P48jJ
gJSF1PvAIn0N77pZnFzj7nEgq4aH7A+w1S5B3M9qoYY8+z+xxrY2I2GipwgQiAP0nbIkhNkOCj7s
SyH2WtmAQoVPSqcdpGrNt3a8IaPLGb50saS8v/fHTKRAYB+lRvwh9oaCcpoflmQrERU7gMsqSqSk
HH+awSAVvoABxXI6PO3tor9BkCq1khQ2byxqs8Iw6+6GNJnmnP/PL1/voOfBpYgLZdHx9wuNxKM7
kYpHJLD31FE5TZwwHnkhduWhFl8jRfTP9q7DftWGBbyyScHd8t7fcZ8KwRz8Hu5m3n+drMySz4vz
hP5yTW0WERvAD8v2mqdf1seGlRokfXNHA5EA4Gr1WBR/csnFbafZ1xd3Fd0fymJMguYyxcO4uRBp
r3XqFfkTjUn6Rv1EKtGZhJ2m7cZC5MaHRfiEcGARGuQLd+0An62N646R8DdDllYXyirKaxDANBLE
U3pLeZVqfSBZaKKY2o0cy9vN2IahEXkvH8ZLDApAk4M/UvORZML3kqUkiuiYx80VBpz7IAWDXR1c
9XwbG4vjQienW14TATLU9q6ZrNgPaHFaWgTszif8HpSXr72SOZhm0bRLm6NzUksRTt2SMum8XhM0
3e3TnoMY1T+NYcLQbGdPb20tOnDsoE356ljTu+0XXibCa7rtSR0KcEoSlJX9OvFyedI93d54yfNR
cT4n14Wg6D2VAWB8Zl2PBNGCxGXrRYX74uxRjb0+PN9KPruhYpYaCfd3d/oVd+IHN9VyDDoBkK89
rYwwihDiDPQlIBy6THLddJvKIHbE13W7Y+U8KetE8gYKlIYVWEEqAqmaYAmWvDW/FkWDEwAxfF8n
hrauiNlK2Gh0azecvll/F1fB4R7MNc/imjM24M7yK60WqrLFnura5iyniTBdUeVpIRg2tFYyLYSZ
qqFJLRM7gNghLcveG78lmUrkSesyIzHq8TnAz1gG5zDODmaS19xEfanNtd8GBqSbBxsZfeWSlUt1
Xt/OCC69fqTuNpeHad95tHuHnYXRv+N5FOXzADyeZNB5X2jLeNKtc+C8kzYudWb7HR974QkJQmXe
oDgFsuV25Y36PNqL0FMs9Wz+V7uXIMHrBkgxF00/Xk+XzBIWmHgAIwbN7DYOkfxb+kHWZgnx5JEK
QnOfrvhL5HdhxgB9Cm9Cjpnx8i5dB897zlkz/z9QT/xxGIZgFuTWe7TET4vi2aVhgk0Oyy2/FBP8
Rfgb+EB7s9y2uJrcAGIvkY4jMsSAxNA99f9owfB7bwRrmg3WhlpTT1oHkOGQDB1Ru+avr6xAMc7Y
sl3f4bzxGDKvXz3srSAwwRDsAOxiornhzI8lOMrAWoj7iDHCEt3RaWIyd84WJ5edvFn6aYZw2UZ9
xKqAdnXxFsCkRo4Qr/rJUBi2dbq2gkawpNBEobTw7ELscYT1Sse5RS8jotJAQTT0Kycu+itWBTDX
6l88b4FxMfhtAg/kQATO84SLimLkyh5bjgNsq4NZkS8D2+g81hHud96v1K80O77ovuZA1+NC8MfQ
IQsa2h3rsksxw6CryQi3n95I7Om060dJyDMfaPXKb6jSE/Qk99LJgcbSZl08l5JgcjGErGswWUm2
jr+9tWiHToKp6dUKR5sWixy5lvYxUGTsBUXBQhZcAizVWDmOKCLojMgZLfvsKJQKYVteNc3Efm6M
GJYjyrvBydEPJ/1qoWu/0JC7zU0psPNQiIYMm6yYD1bGK2r9vYNhlIJG0p/3OPjSg1PXrSoyhDee
ht4WOdHfcIyoS00Q+IimZtrMyQ5xdt7x3UqN4jN59Cs2prM3KxtnTjvKUqIS0m1lORa2k27/1Vbr
pZYKemBA4MOHOwmcSxyao7NR1AwAwPdiZioAguZLSUlBZWm8hXZNPg/v34e5XUm67fOZcl03zJiZ
lCE6/5F2wr5yxtOQl9Uomks8SV4pz0KBSjTPIz4xrs1qF6mLhzTfAXubCVl6Z9pfsdgG5RiekSGn
ar25my3w8Og46GzWtQ1CekP8oahsLAH7ZYJxMpMLNQ60B1Goi5rWx9miklsAOQKX9y81iTfErI+y
qGTcbhlb7A7J0zM9XKNIXU7Nik72/oLmufC3ohFj1iMTqn8P5QtZGyBKCdqNOkJmK7K8DB/fku9X
CxdgQ7w0Giu3Dy+8u+gObdvP/Hgw7ZS9HVwVPjkMvd5tYfTo3JVVp8TPKFSWnpqI77CoXjTwDNtm
bCV4mNkY47huluKfc0mGivROTCT77gKWrEVjXjMYDm2AhxmddLgFcNi06kmQ6hgapMdVFmdqMXRJ
gozY7UknCN+5Ht4Q1PlD49IQL9PgtSdJx0JKmri6YWerFMfxMlqKtKynwOkTzf4u9FzeIEWTziwg
q1rbtVMdhcVgdURQZA3IHsQga0QATW7aQr3jS6ZtsT98biISQLV00I4g37vTgv+vkwVMBFHh4qH6
qmJcOC3sT+oyf6u/NTpWeuCmB6lnGuz6rdiHtScYEGUZDwHrbCsauRXlLIz2DDkTjGaZHrrmxhTe
2E+h4oPh5v5qprfeYT3kPJzkv1UynIiZNZ3bD3a95p4hVXY5QYjo8+dczsOEKdhv1oYG6RFt/zfq
D1H15vux2BRNSEXe1gfAZGr5OwImOG8ueuGbOnKw1t/1shin3Li71hg6vKcdzU1UTHJing5tb4FK
L2dGFNDFtbYIOhjZqTY82L2lcCfbwYxwTKBzyKe3mbQJCmAnRQ/N2Xb8AA9GIGrasqXCR6i4R9Ev
5p9aMtcc0/heWzDl+30ZRuLDTW8KHNpkVpTL/nhqzGDlToj7jnf/uJ1oox+CLqTX6jB9uaP62kZm
79Hn6xLO75pegnsKuvdaCFMefKLzJsDtM8/O7MBvSXZOZlItxGs/xCM3T9BrJ0wFbyN5jppDahdg
onqwiPn4OocLAs/wdryoIUMs37KM4I76cIjwv73QWRYGcBpDN8O8lmATQ7InvEC1f4LavWnp1G82
hjK71dM3uxFWXMzCxiv6GHLHMZfnk5o1IN5y4QiYtYTbQmTeEGLwicQH/qZpKedGAx+iqOmPsE2+
mzkKhIXKGbup62/l1BlKtLVaHlDpIGWP6gKPY6MEqKeOXM2r0IR7s8RQFrfzDUxZBTJHsyrfnlkd
Z5jRN1N0RGqaiaNBHNrUErgzRTwF8pj2OniLucSfJgcF2W4NA6Xq2LiG9nnSP9UeY00D+vfErIJh
LTYmX/3OveKuX3VNn0PxAhUPl8GBdVJC3ix7yw3esbh7IMp94i7WkjHJuZvdYtI2p4jxNFVZcL8a
PU8fpJ4v0FxWxSynb1KqmFcpgum4fROzyZxMsh5H/xSoGpWYk6emuAjhH4+J3BldMSGiEywQ1ASL
alFwI/bL076ecw461Iq/A6ucbIKTb6bd6gluW2ukUQ9P5RoeDzJjSiKsq7rFjsnWq8Rr3vYl1qPJ
hRExnXCdVSWmZwZLAvY2WRd6LFE2ZTuaYPqqtrKYsCcXPWQUpb89HlOC1sWU2iXnCoEhpxzK8QL5
5FRo9GE9hrikoGNg8DeojKPPPRg1MF/yzsplM9sWqLe7vqLv88NG+SocEPBGjEXnHAneH5AoLJTZ
xRS7d7ZCROuY1UQdW61kjw==
`protect end_protected
