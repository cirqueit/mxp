XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}#����NUe"j7��/�g�;Xռ�Q�(2/�r��m��9�O�ak
oN�{K��͋��K䞈�6p"8k�y�_h�|�1�X��������Đ����n�;Ӓ��V]�g3�������S~�U�[���?8�{���M_8l�͖c����^/r����	�x� ���~�O*5Ԁ��Z��Z7�Is���=�����A��Gy�g+Wa�Zt��u67vȑN�*^�s�2�ؠ+x
�_8۠��6ˀ�}�~�!�������mF>F�5𓏊8�L�{#�d'x��}Ɉ���
��2�-إ8���byX%����
��Xs�./��r�����Sͥ��cp����Ez#�xM�$�l/z���G�K�t!Sn��g8�bcy׀�)-����Ye�^�E�njM�:NHBބ����uV�Az�
�#����������<1���7��4��.<-�Ěbi-&�K�ŕ�������_�.�V�!��V�{	W}/�-�
�z|��X*�EVU��/{��;� ��~$�2�;�,u��S1y��˳�l�䧱�`�{f�e��At�ŖWa���_"(�Γ��;�Gd�9݉Џ��������䆂�|��gN=��ii��%u��a��)��Ͳ�N�5?����|D�*� (q����b�� T�����T�<f�+\ ��z�)V�0�� ڒ
/�Oż�[���r0��`ysSvw��'([.�x"I����.6��6�:����pf+��ن���f�z<&I�=�Bi���6�XlxVHYEB     400     190P<��Rξ���xIK��f�ho,�m_ePq_���N���C�j�؇�Ag@̢3v�JĿ��ʝ�������?��Z��[�+������7��{���jn�3�M ֦����'�A䗷l�y�����N߳Oٝ��Nh��%�#�y!�.�����ٲ���h��x�A�|��� �G0 ��w���C�J�g�闩��9�]#�E�����_ZQ,
��oKB�.�<��7}:!�(X#��9a�K/<�6c@4� 0�̒qfU����[��#� �����`bؘ8��(���9LUD��ej���E�+;t���̀����'�����F^� �q���"%<���=��'1#_��g{e䌀��l�M�4fP���v��.h�̿�XlxVHYEB     400     170&~�*�0]�����t�&5��&�W?!�J�5S�6����Hi�a�O]�K-u_���ƒ~�?�������w�+�k�eۙ9��c��j����1�zR� xw�?���|��:���:��;��!o�<WD,M,���e�e7:1 �P�����V�lbf���~Q��ON��cwݣ=�ouJ5`=+px�8�S��w~�e�㱕t�4)2���[�"Tj�{��,�63�ゥy�2����e&e���GN�.8�@M���)ߣ����NON�2��2��"Mx��M��9��ޅ�a[a,U���^u�úK��A��{�uu���DF��|�2q����aCA?��Y��P����W��ao�JXlxVHYEB     400     180��lz�� I9����;2�g0AS4�1����l~�ml����X_�v�Vz��W�$AW���:ǲ�=n) �m~���	X��|��Eg�q�S���7�W����W$���:�L|o����z��#'[�9�!q9g-��}�"P2q]>�� /��$||sL� i�.�:�3�PH��\�~�E��P�o���އ��!������A<!K�'��J�6E%b^��w��4bnD&՟���voT�V��
8{�B�9��]�Mܰ�0
Ǟ�MIʛ5�W�4�x��#��H��P�,~�{t��A=3��u�U�NBO�v�����S��-P����n$�$~�����r�9)a	m���n7nz������G�V��J��2�"XlxVHYEB     400     150�9��@���l� �;H�c�;����`f�`�rA �5���bg��ME�#-�Z �
�QS�0����
3襪�ޟ��c���Go����\Q�I��bq�9.��Bi�A3�\���`��W��Y"RGP<�Z�W}\C�,P���P��!j  ���ip�:�2k�k.M2��m�N\.&"d�lg��-���@���0�nO�����b�k^��O�����5�~S�vZ�`�Q�o�����2Q�|q�3Y,	������O[r�GO>���<���p�N��Z�D:Z�J{~�ף�w6E��h���}~�iЬ�Q.P��o���v"V��M;/\XlxVHYEB     400     170	�:`�����e:�ϟ}�gL�$%lS���8�T;��,P;ٸ]Ɇ+�M@9'ywqY��������J�)�p?m�
S
�С����Z��R�����1�"�Ա�L$i�95�y����@�yc��<�iŸ��#A����ZV�u�����cn���$#P띾��t�~��z��2`��n��q��@�i�EdkEFJe50�:�Y=Ƀ��.GCoTLi
`�\��;⦜ᝌZ	���|�^c�� W�4Wr�0�s������b,�r4J�[���c�h��?O
I���MwA��3�eTL3M��M�8)�D��|�h��s� 3��*�����9��#b����[E�@�=Y��}��[XlxVHYEB     400     1b0B0������o�KUe{dG�Sh>WK�˷��������(\0�L�{���LF�	��ΌQ��/s�BHҮa�a�Z���4��[��x�đ��ã��T�A�U� ���),?]n����C*�N�}�X��#����,B�0{\I��!à�ڳ�8: �P=�K���l@b0n�Y1�kM�k_�|^O��!P�P��ؽ� ��y$GN��*�:�d- Sq��/|���p����% �	��6��Ov���E��܊unS����TMZ3)�[��O������֜H��e^3�ɷz�B]� �%�^��x�Q҅3��bu�aE>���x�HԶvE(�F��� UKb�\�]>?ҳ:)?z2D!s�#i�)m�?r�~���],u��r�>3ep�ͱ�,�k!#X'�XlxVHYEB      e0      a0���1Χ$/8��0�u��i�K�UB��Np9?EE�H0 �=��xC-8��)j�2����u�r,Vjφ���2�ޒ۔Oj*Ow���V6+z�(�ej}��5��K�i���a�=ﾾ��a�|�ˑ%�I�d�vȬ�y��']Z�)fq���]��6�L��