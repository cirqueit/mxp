`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17984)
`protect data_block
NDXv5RyvFc83mN8b4HoFHZOgn1Osf7Yi/T8q00bTU6TI1GqMt6OPGm14RFbwbqUK64ZdYqaKBvMZ
7+zT6oj62PghdXaj/jVk+1KIq4KHUQOG/fmX6+43cA7XEKQHQUeeOfBCuqOCzR+Y5fmbgENb4QIS
BUN4HoyaLOqcklorT6JtXbNxPPc3e41jvG5TRuUWPXoD28XIHInyOBNEKRDii39qb3+fR2eUfJfP
jaJLsmS/FCX2JaFomJdwdm1uJANHUu3suSMlClNBSeKGWtQ9SksOgTuHFIHMI3KzNhS9zMIWGcB3
R1gwK5P4kmeZyUWDKUkq38aBimkoUNYS61QWuXRcUoTdQjvN3YlShEDckF0EvQJ2REUcnTU4E1DB
dbl6LH/F5qww+guPxQZBbVEyP/RF1Ao9UZcHYEHQFCEjTovKJEKFDdnBhgogR5ZcAhB/qMQhWA5V
cWMsgM0+BFfOSS0W+seirOv2lQ3x8DRvyiJR33LlZWslAwIWFmn4L0qipGvJ4qez9k0ERfE2Ddxh
/DOTI0eTktMz9b/R9yP+BslS9pM/nQjKzruEQVaGLWIw7FhRlAjuRfiO72C2472U5L4jF9N9aSMW
J1HElO1YPRGsxsQ8P2XDGKe3vGhtguk7ICd5NcB/XUMjIL9dqBMRNH0LGdqCwdsivrfnugkiOPpv
rICcxW3ZPoDtXojEdjNwpGRbPq3yi/6lxal6MxWP/IbW0Z2KNYrADGqVgrP5qPxExIWlaYfmyuQ3
SoFRrDl153DEtjLYzVPkz8F8IgDeRolIZ6ZYKWDVL5ovO1aJhA8M2kZongKG/W91bAh3Qxlf0zhb
PMx87jaPo78p3npb0cryNrssArxbdPhPUUcYZMhypQX3DuGZN0q3ogRLu/fMQ1w/KEU8XkSURbtb
IgnEd1Ra7gyJ+5iVJ84pz9+fHQ2mtWdu5WtuuMirE5f/HwMxCxpocTo6pZbohUuysi7OpIM0x8Su
9vL1gS0Api1lFGYZYdRfGJWr169pjxKt1lU+BBvz5Y1KbTnqyc+jQNsaxZu5oFZ7Zsn+dUG+Ekbg
Vb92nfX2aFYntRk+LKYh6IG+nbY3l2v1fp+93RdlQlXVFoo+OvVTl8szeHHdO+Ec+Pi5l2A5bp+j
yYUQ7rmjWaODflg2YRVohMfGOkXUv5bHkBN2LgJgHk0Y22dK4f7ymS2fcYzHztB26MnAp9O7NK/h
K1s93RGUN+IrAdWsCYAvk6n6/5AnA4Y42V4o3gyCuEUY2erhjkHJa8Q35UH7bef6kYbNn04cvT6v
XmckHtCGLUI8wWYnTccRBK/86++RYiL2PTwu4MV09Tqw1X6mITxb1hqEXwhnAgclxeF8cbfw0K2i
Lp82KQSNUepv4zT3BeMwnBS/XwBbtSt8hC8ZVDiCFyjYqKa2V0f96anajSxl7WcXQbJv9HUq29LI
MICkDNjWgqW+VNQN1qSM84oqQq3tt2N/bxsfJlxq2PgE3Yl8h4ABbgfkPOL9a8cRA+7AzfV8nN3T
fqdOIUkVHwVScLF3lx0mPzg/C7ysMoWomDfiKk/qRpb0P3tYA65f2+OwwFSAVwLpcSflt4sijk5a
diTmgqXryHXafV8GfqemfT13aP5XSawGsQBYEBAlaeXRSUbnT8zi1LaosebPODKAmEQb0pQCYgWn
4lSsklBlyMGZr/5KDmLHoG7ccOBxiOoIw873PU+1NKRNwxNXrQOm0hB3hSuK8qfhGLoKSO7cFOIM
XFH7rFi/e31baGWnFXe1rAWcH5YEkSWjNLHbwUVCydH1AxABDD98TGIeABXCCeapgFlcS+YNd026
CzF3ll6oA0ky4RIZeXNsaMdSqzdNuoQYdyGbF3XiSmf7F6NTQXB13UkIDswhXg5N8Er8GYxykZvt
rcbF+06XwaPi/3OJXGM2y5dtLpxHqlLFTOwNCp7plgD7hJDxTPWPAwMbhQv0AtpDCGvptV7snS7k
/jOi+9n/VRI8ZputP0umBSguHRwsMP3Q+I4ijZNMenPF1MRR8eAQ4PYQtG+ZrDeFtrsrgPFmDYjL
zefmdhcKXBqg28qoCESqs/8uG5QdBcbVAhE46/cUCT1qoStX3U14TCksQNio2ehInfMnZxOBcA0Y
m54LXa1VxsxYwNm5dYlifahhy2T4EYYoCXQxHVEmH/yFZt8mRTNbG+sRN0IGve7Yd1DU/+yxuXdY
jNrNTkzTMdQ6rEQl9IFQ91aT5EL8P9AXrylUBfvtQnzZOjS0EddYp9gBuVTZkdisiBdv7yRJr//Q
kkUOmqQFKaIxSRC+m4gwFBFUedM2qGhHEtRPjYxc227pQpNeB3iCNqgQfOhaZNREDIZXWkmzTv0H
8o6W19QvIQ28AjL/evNEHW2MZmgKVKhzELepTZgpLdPjyiaIBWAHS/GUDND2W0DF/+R+ipYwIqoB
o9KUzm9K9+xOaVOaqii5UIJ7ywzetfAkvvNUg60vVA7zRHIj5VR2Ag88NXikYfHa7u4ufy5gQ0tN
wzo6hYKnLip9LC2lJmJlF+vN8r1zmCZH45CBb9wPRut1SOuoDfHUhCR8X8d+xXwBZ5LCmX3opTJc
UVCnordp0TVipbDgey5FqQ47BcT9AFVvfhF87Bu8sF2FvFAblngUiwjsKn97lqFrxXTIOiaArXrd
17R3hQNf9H07ZEaJcAWsEvoz9B6WzsGCvd5k9eBUPFM2fmjFgSl7eJNl4X7qCElAiJkdkZgmLe1A
/pSLgr9N9b4wRwafIUcLTktoJpMVnyqlIGKO1tCV3dJbt6im5Ph1qoKcqfhfT/H+b3AtW7HY4f+N
q7CjY/4vBqlQVOvfNNRAx65ASMpvQ0z/FDAZNcJrzkDs7HwyppyhTVmTjUaRJcsLMEiCP82oMpO0
bIIWgq2Cs3om9Kky3SZQadG3E7jCOa3ac9RxlCFBKgSaySYe34irSWqNNjqPrfs19Ob3nPEhcFq4
vfYM39LPOpXhyApd7IQpP/p6Ee/HS1hKkv+2SUugn4j4jemodJDXkY425i1ukBeOn4HK70Am6nWR
7QPUm5XB+ARU6YGTmJuUE86DV3hu3upDuOhs9UEgBW1yFKbLbq2uWTZDKNNBWqT/d1Bo33fbebvm
WU1IMPW8Eycz5iSUtWM1WxGJgs/fiwccUhJDhvCEHCkIBxJCYSlTbRd3px7JxtPRd/rbEAymjYbf
0oUZ9gYscKQMcgQNVhWmwOmZ/jz3ycy2Aq+dkLR6Fm9S3Wh7Hne9ZZF2kB/mBTjIuAePAaFjpICq
FAT0KiH+P8Y0SeJV/ok0/uUHvtPfDG+QdJ/D5J8qyFqG0A3yQvE1jfJN0UysvFYCIyQR9Mqr7Ye/
eRZgsIApIXIrD/DDu6aa459DrX6NkMhg8GdXAAVmF3UYsB7wqwJVSEXaxDb59hTxwdiSpjVuncZx
9CSeFH8qQly5RoETevTwK9h1l2LYyHuSxgr4LDmkm6r6zQ6As7Y5U86prz94dtV4mJ7bLUSxQhhG
lHZGRORoh65apnEb64N9YjNSxlNSGP4N/0ILXUpKiO8xsM9DRfLGQ3+78k8QBJas4MRS/J7eEUwx
3wJkSvqOKU83t6YgHZGLuRY3Hi1pxGvayEQaLpEnNyVkd/ab2PYRXycpdQSEFN9Y+aBws7je81mk
JG/N7SP+BQlqS6DJHL+fRSE6eL1yyB+MLLe9o5b8IcjBQxqumSLSH6NSme40maIsaW0rl1Xiczzo
/7QVctm89INsx5Fv7BOa/nZnS/W+E4S0H2JQOl1j5wqR9OmPvF9Jhw/EgW0cU+/Y958T9nNoeqeE
AmriG6Q+52PXlZE/MRFIz/INKkUtQ3Y6vaw4B39I9zupdRShcNzkphE9BUbMTVfHgrEueX3/ROTE
IbbBFOTaJ+/lPz8LKWp7gSdWGiu3cjCoNeNpCI2wy6DAwZPZcGffCZdOBrHGcPffcq0hqTor49fS
ZTjsCznVWWeSqOzdYnSDKT5UJN/DSveYb0UShDg8Ub9zTMGyLCoporBm7qB1UjwyTGjWjZjcv8tG
h6jdy+TA0rO69s+Tx1qVhx5C6x9yfxZNhmmbVve0Ys5fzMhH6FlLaFyyeeBnj/PuPbbIGSNCZUA0
7CwBkRs31BjbZULtIZ3mVfhKyq82zErYK4AVenRAGX7KOIZnh5ZW76/p3y08w0JDpibPDjoofZhT
UMePFYqPeM1LjYJ7MXYyb7Oc9Gd/C8kWptfKR0lgueweecGV/dMwyQ9BbdqY/skZgMXGbhZ5ddk6
bh/Mh+JsRPK1nn+OU30sDhrq5XHQjDDFTayZIiP+wEpJXnmTrhuwLxRhGsTAVmnKu6CJdegZvyle
YQNMn+J4lJyYHuFn50NOhonwgJUo+y5plMjjq/1S/5px5YNvpE7gbp7a6Fll/Y8rKBE9vhKCOTer
qemjdTvVwZrXHw0UmggPjEiWwsL5pk51MU+fvKuxi7R2KFY3HLhRkRJFGhfgQd5Dsup+OgtLODqE
A6I39QtQYPfNYBHEPvF+GRZeUU8UYADNs4BN3vJPYvq8gQdkG0tnoi5wfx+VnAst/NANJq3WckzX
2ABhKJBMyIWq+axXpgfMgJmSsFbFZTB1s0KHTtgojjQCuMfEzNUMgkOHhC2TOfy4LcbTlak797iB
q+4pvKkK8e2AdHyWfKCHiYGi05Xf136vFQfoOfb13CSeK/4LXTgISiDiLtKnVd3BjzRtf/3Xj3YP
2zmS8wlJgPSo1wthMG9IKViiAvWB+DxzljvJX0YFzAUBaDTAgr0t9RbWYiS3omsZmJW0luOM+rTY
QylnYhXSDqOPQHyBQb2EvFGDZynqM3qLs1+ki360iDEP+QodYEh5u8dOrpQaoY5srHV6JgB/N/uL
+5iKqP6m4gUnAWYyM2C9iip9VMySD0FSdnvnHJjwJlxc4BAYTL4VvBWzVSnGZ7HFjEgn7I0VRGSF
VM+x42cJ5x0e2sjyg23NON2rhcLz56K4QH+w4wYSVloG5O6M+Uw2Be/5n+9BujlAajwCRQdmlYmt
DjHCUQHwgKzLcNfn0k6YIQL+em4IK16iZKWgp4eJ0aAeQrdRNn/SdANSz+bfiJ24jUFJLVZluxZD
PEnUgdF/l1DwrPhgPeUaPZPbET3jUmN97OzgBxiJGfVZ1VhqW60yw/bs02r3aZ4z3tEjWEW3P5uF
ZUhdrdchodji/EZJ6htdpjL92oPDZq6H4wJDQ5w2E1r1cE/IV00qq7yppZgzqqJG++Xnki9v3C+z
tqVqJDkz7aJFNiQLktWvVwvMntck9U4zk30WyeSkjkRxoDZ39h04cCuxMgYKmRiNwn6jxpl8nOEU
tGt+e9fQuP7eoMO8lY/skq/eD/+B5nhe0r9+SwR/t4d8EZCuNJQHfe7mMg0EUFmUc6Win3oj8TYE
Q4I75m/CJubORzrPYZDS3mN63xC0iAW9tEn3uL1vpx4d1hXmBBgdgFWRIcFCjd2A0qox57Ku2Yf6
bRDvcUm8OxsUQp4mTb1IBUwad8LjuEZa9FHOhryqIk0C3rIjXEbui5L63VThkxENE4BtIWrRctSa
SjMUCMjisHkwC6QwLuNDLpu1HWewMR62Kd4XasvY7Ajy3przv+ZIdRoIS4tGhYMVhkJE/VvMJEbP
hxZVQnE0tih6JN2OzlHbB1dCHQ6/Kj7+9p1ysl5p7XcmnI1p9BrmqcJnW27Fnf4t+k5xAC5lyKza
8iBbZdWaJ6GLXcOgXVBrkX6u1C0gv0LphOsPunyOUhfgBH/RGnZRtAn1SBFi1tdNk3KwvD89fy0O
LavGRE41nkiyKUrYq/p22mtbFTKCevlWRcdHD4mihKKJIKwr0lRe5oHO04ZjfgXPiKpgEGd6Oss9
q698Cx4uNqg49EP04b6AElcVuuuEsUw+c7WGcdPNwjPU+2YtmPS9C5OG4Hbls9t0YAB1o2XxM2MW
pvQfEgHUmdQBLqNXb2HcRLfCn2v90H5N6NXiFNexYW8cQopCnlXC28zvp4K+HshY8IxannUk23Ui
C5SECotsxQLyb4xRqPATjd/3ILH4zMp/PMVchytxE7SEMUAV/nTdH+BBU1tuZNEyG/sP3WUIbE2F
MXDAP5YTf0GxJxVrCz6LyGtcz8yGeTLwBo9VSKNal5yf11y7zG3i23zQP9wnDZrtT44Pl3bp2dLh
SUUxEG9pMCXii2kXPw1olgSuFHBLEvJEneFyFchOW5+f+GIofUtt+P9oNqoSYSMJCDHfpyc6mWLU
ZsKr2jTgqftapSpAMna/cSce2TKLAsYIY11BhF4/Ur33ZhM/n6fquPl/Y0OYZ1VHtcWlDNBlUSZu
s04qJ/Jkrpr/qUt5G3rCYsAL8wtD8E3mQp2ecZdYDxK9owqFCN591lg83ANlUlPyri+BK4YT7z1d
h2WblsGstCKtCN6/HPfEtblksV77Z9pHMqa/6vexygKEYYPKqV3wdi51Amr6Z0eLmVixKkjvKaif
fleOUVcWG6NNpsDu07hJ4lGE3MHJ2Ox3WtLq1cfxXj//Xzp9iiQ7fIjm7ClTv8DbDt4JDZ+jfLB+
Qy046UxI35vRvLTetaed1Byr0dA+mhqPg/TCAPGVPfg+o/qfOjWKsy7JyJRHlu0xMjnnnV04z5wR
9ecuZxsz5M2EXmFpn+JWnVDe2bbT62lKWYANwoAaKhtbZtKAooI0Pg1EXoxfH1pOtS2+80WXDtW+
xcVTW1LWjATvGx8H5qASWumvRohhJC4qiyH16Mi3m+bqAI3dVPS7bAzSw96cBFki3R0ZC1mDvdas
t6EvO2RqrfXO3igKv1tZBwzbxg3NcS+kOOT4Q7vrWmkgoWhIQUdT/3FW5iAZWAxwp+RajfQXnTKb
DZJlepwWU0zIy05sZ8mjKvXZO4l+QTx+hMbZI/O8pEqJtJzB/pd6V0XEhryrxKg17Q/ooO7Y/gy1
ysh/zzcSTz/Rq6xFFX8f6PAbgMBfJlDfDwNpfzn3pMUiQRF8hshNSMH/n354ng3lbr9uSRW7sUTl
BDPPtf9D4Rx+bhyYq07PmolhMz2LRNUj1j5KJVKVMqYrU371OzdFY4gnjgWw8qjPzFyMkjDkuXIA
46cNBbtr37TT3+BXOHKuLMNNLSQhl++WPc376k3sDyo+G0goao6n2tf4AJtxr7e6qMZtshbAVi9q
RAd9VX228CEg5JaMu7VkYHHNvR/Ruzdz32PoH1/TTzEXdU3ndIfpNrwJL4zdzy6rYUZGhacRZLuK
7qgVaB6/hmC4dEofkxZEwOx5C1SBKpx/F9zJH7xTQA1wPxHXC2ONsFy2mU6O56a6macp1fPPdIIz
AqkCLlW8O5RfTaEUHjgSsPhYOg5ZBrLHkDcgk5GkfYwkht1v7m+kvjEm5xpvIhRu9VEbby5irzis
4vQOuZAoEnb2TI1Q1Hz7wS4g6kkPyzZ+jKfAbGQ5dysZoNtjqrpxhxX/QR/zwxCKbXmzbd4MPit+
P5Htd0b3ERH8wIsJjlnWjJB4fAlmchb+jNwt/Evn5qTuYD/v5+qmmv9eDEkrIr2EBygTwkrgGl0v
I+J/Y0Dt4oWGpNbHhZf6xkV4ALkK6rpgsNEJHpp3BFIJoEO+E1ztLkQeSb04R99AIUQkWAq54NkM
+yIVkOpFHKbNjmrSLGhlU/S1rrnLyHb24fbRxeVo5jjnv/Is5WfMaYAQ5tMQksRR96foG9VekDjR
VH+fBnlMBzlB4y7I3lAVtu7iucn4HFQYf5LMTsV0NDcudGAxaqAhQrD7wKZQS6gBGtzaEJjCCs3B
KEWLDdCizBPEKi/F279b9Ci7mCiauT54tC1Dx/aSAkx/GIKHb2qXyhI5kECPk1T714KSu/TKNJ45
5q21uM6WFN9dywtCYR4OA8hB47OZFBZN+X1TB4poqO0uLw3bl/0tlcG94iKZqTVcQaVRaexQtBbZ
BfhAeaG2CoomPPDXeBTn1/ARq+yGE1zpFoo9J34WS0pxVjkQ2/r8AaCIQ1UdaBRJdl4SHBp4e6Xo
B9pOYf08Kv7//MtUYJAsMNwEJCv/niH95Fd+i1wQiuogxcb/8H6P2XgHeUwGVllIxQFDOoq/JYvc
QxXWXfApKDyv5pH+l7dWTJI7sESGLJ2bICyaUNvw70L6LVmPDmlhtc9HYWgrgQ0GRjCtpKppBjvj
OBit8M4ecGSvdbH3HnyK9seNCHvQ3FB5CU8i3O+rp6WFJ4zmvNMD/kUw+UDhmWWvn9ctgsW4GRAb
PqPz/YZ/4SVMtypWUCgsWMI2+LyI0yCq++hEpAHiu49jry7aFVnVR2OmBi3wazqojBo3VzVwNx0d
EcaLPVexcvFfATV5V4aXXM3yCu5VVCMh+nLZKgm/aMxNE01VrZ8FDMaftA6sa20UAz63zh0E+5Ix
4NtGC+qY2YFL5eRcjjTGXzABuKd/goSoA+S0OEjYnylAwGAXJazzCGDsSc2Vp1jzPHyufAVKLGc8
BbKdviJSgXziDFKP1gFhEaBoIV786iRwNytrxT7qy/cR1ZKnGW9A2o7F9AMCbCW/sGvR74YgAJPg
ddub3s6xMNNIGnxE/iyo6od+4OKYLNWrF/NGOYj1V/2auOTn1DDTS4GL+upgJKaYumy+YKSKQjv0
btU3+rKNVD61ledFy1mKJ97HgTjdH42K3xJPpITn6xFIV2KJu7b+TofjimGFv9W761oeWdcijjuN
o8c7p0omEU1lL6+Unt5oJa323c/0BDBjvo9kl2XJQGaxkRVUHwPT/uGSpvZjYqqhsSEbj/AVBEOj
StKL1QmxGRkNUi47hzV+UJnDoRyh83yhIhTZfi/cFI0OUDM9GPEy3vLaQA9abu3L+soajcTMpmcv
HZpviWUKrzPgiFxJpDAKcI8uS/7wZpHgrpRVVyV5mbMvWVbaNsOS7HAWCgBXM7g/V3dBlLlq37Z0
JKg7Nlnci8OZ3OOXlZxIRzRbi+/cEGTu8AIkwGWCqs+A4WrdqSRAM5fU8h5ibOLzegQPgjdFQEf+
o0jmc8cYz2HQregU+KyQDzIqvm2+jigSonwLbgxdiU2VPJ2ZVsrDWtwLq3haaInsSjYr2vloE/nn
cuIv/gLlUHc4MbneZMiv81nsvchCto07EwnAWGc596bcJaroym03xOTOQSkctnGLhc3mKaIHFPHK
ZCzAqAj//guDxPm7nLJU6p3k1RZQ7YxK7lPSMZVadQGXn1JGmUy8IxtSsyN6YrbILwqGShK5JW9x
k2DB1/z9Od2tUEmn8g+LWTJzx/inoyaAnhk4JxPjNX6PTaAXmaiXsheh1Z069rdUuRTFKKCm7AMj
PF8nf31CHVoiiAFa+x0nRpIxpXrmft4QMjRjv4fchTWjAUHtJQkZzTtJQAr9Eu/GWScQ/VixL9+l
r+s+Hk7+MjkbjSjiCtjGK2mOA+erFjcmmVKDFcSn4aonLeLGuw08xTMNwBRyngTmbH7sQ0S5wYZW
K7Vk2Qf7tM1mQjEO6lrZBoVamJyUpRmRWuBN30xFKEMZae7WarBVk9yXNQagtywCB9fOAGJ2ng1X
LhlL0l66p8shBNAq08yBndp6IM/xjQeUgRktXOeTM8OBbd/OvBvlFf9AXgPKNP8qH98ZLDWGcrcc
NWlZ6NDeZjmXjpIpAQOBDeFCLK+71C91g5CdEzCg9m7RTZCqF7dI7ic8bAQSYHU/h9dPJFRSCrcY
Y55qmvbuHgESWt3Jn0LWW3mBA2zPuNo8gyLuoRmHIKzrnOtgi+3Um90NyL1FntvpnawF98LWMXVJ
4chtnc9rCkyfzpwGmdjc494215+Hgyt54sPH0oUq3v4TAR+lqLU8T3JjdZixQlPIa4YPqjRvy1rj
r09Qby/U6TaSICy7C/cB4s7BmM0VTWr/nkDk5n0AzbY7/jhkt2OWvQBjZBfW1kijcLgcjtzkRZ2h
PuDL1Qe2sLaJ0g0CzA0+g7Z8olYfbw1P6zEvdY8P49oSb3lKuaUOKSmJYTDo/eS4YdSltFWu2sl6
ou4wmrJcT6Aqdz0AI3BxPLJYf2+I93dENvATr/9oc7dzz1QLzsc8oVV8vibE2yu5fpt2LM+Gocot
JoD4QfZkwJjfjX4TMtrXKeotHowf3FHXiVnQPR6OerxPq7GNNm+2r/0jwRXQAZRL8Y831nqtlXq7
uRzTU03iy3i8j14E+mJeF5bvGyJEHzsNDsEDDFcqCOjirzzTAxXduDJ8qe8XjSQeDYRMoP8Tk3nX
yks+A8Z9hbhhFiWSAOzDNn3BboZH/olZGdxilRAW2JbqGXYOKdPDThD8RN4bkbecpmdEvDRgCTdw
KcTTqCFNgQ136JWmuLG1tkJileAdujTD0MjtRvfPCMYJFI6HeTJ/lMm25kfURWH4DQtDc28FfehJ
oFLn0nMWOkdfKqFsz2+DSJcAhlp33YBcOL3mAOn79OKsDeZOzM0uiST/yrWGEkrsP8yGvv86SIOJ
oTt0HgeWhas38ARG09MvXo4qYebQgXgqxNATSJ2InO98Ydy7JVriAv+cFDHrSsBBzHO7s8q6/n5i
4QMbI4pr5yLtcCmHvGXTcWmvzBnhUdEH6wJyFuA3iU41BB22UIn/Q16ivmmlK9l2xg5kEEaIPZ83
3/um8s2GT9eyQrBL9AaSdlE1iEImgILriU0+cA247PolYMUxVAxLnMM9lrc4VAepTmGeMDVEeF2f
SMRs4agdvmzIGDzqVomTrenkxpXmG40EKA2knAqTNgWzol4P761Fmj2cXHMSjV1Txa7b7c4EpA/c
h646+6wAcULrUDzHI8M+j7S2JP3vAAJsgYbDmH+LGBdfvbnCVXv9QjZ0OBqCg4iPO0AZZ8f150gw
RFrC4jP6baPkj7jc74pkMW/Z3GxGf13n5urpy36kgPw1iyDSeiBqrHo3iZHRycHT86tKuiMADcFz
qFDeqCO5Qxbs9PBNAwdnmjdYmNXhYmiGluVZZAoX9cXQbpCxOfVSOQYS3Lw0nYSYPHZeQSGlwAcf
ETM6RiBTNmGkv0v4LDSiOI6T5+COw8WazJOZam/SjUD9vFGXrlACMen9Z7EMx6miGiIJj4dnNTYD
74trstvKGclAiav/j9R6R9fGUseW05PADGKh4P+CeJFtTM1Yc+YAgMdTyclyD/rE80OkqkR0m89r
M+Y1we3ufGwiBPlydpDF/5pK5okl3/mNOmzl9K6USlJDy3V8iF8ueBOArko+WIwhpCZDaBbOv0WH
Ww7IRkGxLmGMN6+kYdFeUDxjj4+X99jqc8Chhc6YXLyU0nufKHhoMr7BGg2xO2h6ee8zXKiHydcY
5paMGfb81apSHKtws5Rlo5O7wW0/VVk8ygveCIjSSpPNpjATESYprJopusDyKB6U9DFcXryVlR38
ZVtWvo9UktL+6SpsnPn1PrGDm6jDUIO/ZvxIZ3g4+dry6m6VYCJPTJe5WeoyTjFr9kC20f34ZqNe
s5VsmvOAzpzYAN+NuCsGcgHX2zqGttmIkJQ34lr9RamWbYDr2PtNyRyZZKYl2/jiCCHuTwIwFwR3
uwztR04SHQACQczqsFZ82g2QOak3+DVa79MqF0jgEYYSgi36Dwge58pfUdEeuJoMeDvqLA4QfyRV
KxK9/e0jVowm24fKT6xcHd9cgCOc/bhxaJ1wTQl/0TTtaVChecBzP4ZYrl4/l6KIF5hH1K5TIWS3
cucISCEv8HasMkRjyDxLrUFX6N8b9GVqAVjVzqrbdATOAGLQXvTx2jWC8fCnZca1wLhpGxLRVrzW
3O9lehQ82pLwUFHUdxVUSAy91AoODXDIjBBV1Y+Wu5X86/9j9RiV7fxITrCAFj68XJcIMyOdsvNf
Hg1ZI6PkIxclGli8isfS9guxyDGISbfb2cuq8t84H0FOLiEG0QT7LHh2VllgKNYEKPziaQnxTt3f
KDfrAFubn1ZAgfmYgmZiAd5633+qXYOvYYIjTF3TEi/g2VQ/SbUNWzzmiQcqpoPcc4nsQqzMMlGf
Fop5kVlmiBN/9OXhxFQPZA6hA5BXh4P60Mq9JkREEzt7sXpHXmqFrh4d0ZuHDlLAQbHQY3UNMU69
4w9Y6kOKxvUotos+ZJeJ/4jhRg/y3htL7CKyixnj+WfFQxBHnq7GfpbkTguUQ9T8uLxSDQMdSeRz
XMgGB/mOxPepbn3jgQlUfp1UNX2H50rafI44egRY2u89UwNzLxiElsPuH6unLLOdldTXOqE4zF17
sfQ9NPyfZtRaDJb8iJKqOhygR2Dumy7mRJKfial2F39zKmVn4nMkBgmnHeHJFOH41aA0AUWm1Cto
6xZjRDro5JPtylp1tV10xQZlGupx/DocAGYHCG3uh/OhVkmwCAYJ/WjYoeV4fN3j4NmMPdMA4eE9
Qys+1yViRfgGpku2SIAV6Th4wJMnlog5BBgUk80y1kZSN/WVifsOBOPIzXAIAPmPUMsEptzBWV0+
RD7OXPvZyaYxETT4j62w1yvgY424DkzGbd2mUqWjZVKf19w+nRQOSDH31dikeM+RD3692sOD2/t2
7VAxN8pYORCVyS+WOGNNPmmsBFgbjlcc08OuVloQHIrMc77BDsqz7I+/LBc3nHUigW2lk8QflJRQ
8I19sXq49MeYOTujFvFmn/feWbNUT6orbwhafI/kFjDvbq8A7+BxgmcTAjo5qthQqEdYBDDaGAuL
ajleK1qxhC8fjhFCpudju3oDddF5L/71uEVIhviVhdz7Cw6u8r+afnkbd6K/vuFhtj8o5VIN7hm1
d481o+l/Lc9AF0uwJ2UkNTEQhJl1HVbQG2AjbgJFmSBC56WtooCjVvKcXj9D0diRUWZleZ1PAmvn
5epw/KxQ6HD0d+G6PyhTupZ3n075tb1fyjKb9JTkmMpXVIWWwxPcwaTHOBLXlRMv8k329WDrNxMD
RmtZ+95PyK38ySDWzP1SLFrowXbL3gPI6jRoES6ydKpNn5pxQKjD7zQewdcRZFCxP/yunz0UmCmJ
WGSNeN1krVe3hBY66gNfRHuvLiGyuA7Hqx/I9biAxLlZnoG9sdlXMgB0GhXnZ0UHETyER7ARb5IG
cMmsRvudsnZcLpDcDQ1OECehxGZ6yWeyGVUKvHWLW5wNi2Hmy+BnpZMOYENRWmoYrSjhPG9Juyv2
44OCnNtOhG+z9KBjRQxHBVjJyFO9ZbDeY4l56TDEWWFMmdZvlQ2R40EpQDTmTYPRFGC/+hlinJdL
WMIgNJngbJxmKKP+1edMDC3E4/7aKFoFPGDC7nxe7r5RXERRHFPOjWNtRqdqmQbEvKM4pbmYJyO1
vD4IVlyDMvTWkXAoBd9M4BXZ+aDhrKr2L8pXGGRzvSwqSEBiW1vCRJdIONYgnHtafojhRe1dYDDS
vDAsPmtLnyhHsd9e8hHlPSWw5zKd/qoqsXLb/XrrehbVX8npDIYqJ/FaRnqWHshNAu8Bvz+UPpxV
dW3Lnb8zo+5yjRUGuLRi0Y6iZFK3q/8fZuCcYmfIlJ6wQb6Mc1MRCU4xfu6+lfQbq1fUeA/umryu
xgqYMvZg2r3U4SjHhgYJgqHYV12qaDtA3NMH814H9pvbsIAMCHt2QUoOiJ4fNEDjFmx+LGmeO8m7
ZfP4TEUeJn+W+EmdY0gosalTwIXYzVTs6wYLZ0Z6pl11rmxxmklqRvsYwpCWgKTBPBIhgxNxSTWx
aMC66BQq7meYaCXe1DkzYtNmI3pvWWW+/gH4xOZMUih5mj+euq1NixYHdWqIiT9MN0sD/BFFj2/Q
MUIgoxbkQQd+mr+xPAIAuwl1a6l5B+5af+WX3h9T42hLZ+zj/L5Qe3YdYGTmbIg1lrcbH0L/PSSW
9clj+dQzosZ6hbziqZiEMGn/Lf6SoJsIJ9086VHxt89JrD/QUvtH6rIoKx/xRjn8n6eSvqCnQP3S
ZytFjwl4vsHdOCe3qOId+x0fuh+06Kc7nMm4c5+llh0+IEBaDH9y1jSM8ySbIaOj7jdPVbr21fie
uqHKHjq92HwSBFU15ggJ2i5+jNTWP7GiwjXehem9SRBFb+9roHIfMz4m2nY/zHyBeSSA2gv/Q2Tm
+8w+UerEV2/FhIC6cTD1uVeN5xgPKIX7/Myd17su6aD/deY0JMO8iMoDh8qqFzG1qn30mrra40lf
7x8kXemImDAGRNp2khxxKBC/RIWrQrLK5A//V1Yk1eCBfbZuErutk/4ePSa7zhnUo+F8ndSHN5Qg
08IdGgWbT78BZZ6rbrQw8Nss1iXQhQ7Ntmw6FmosMI1CcxbEJCXVX5WdzC5fG/qjAtqUuADVKd0j
F3y/HTJrmTXAilu/sriBVnq/m9VbA26cuE7ztMNPmnTaECOvrzWK3q9zsk8uYPXucSod2bU9X7e+
UIm9l33xsfOh1SOnjgqpL8Od+rCO17/aqQkJQNJ4xdE2wDnwro1kzB1QRNIZAJWFtWc5mjxx+NRZ
+RrgcB6A4nAkQgcWlDWSdMTxRdaFa39biJ2h472djRwidaEiZ5dBDHu2ta/IkoMyuWkh7YYX2tTJ
xRA8yTpP46ZHUdt3lZHDe9FLV0l0zjZuBrpGdN4XNXLkIiilkGxf5Dj82n5A1yYl1W/6TANxtzKe
wJpQJ5SlphKk51FUovutfaKRdQWCdz6scFXVS76DZflbQbrq159r50lw1edYjojmPwsdRWXo5qUO
h2GsgFfKpeIKpu+n6p7azlcJSHTEWd/d9cVj6jempA803x/K6mV7nQyd4n0G5FlABcA8qD8o7iJ1
WBmgNwLKXzcM6CHMCXUv0Ew7FbpkAhHbCicaxFEs5+sRV5+oybJUSFbiTqV1c+afiahFgyn/AaIW
MelU7V/SPeGe0q7dghjtKmrQL9U0z0c2pGyMJ7DhFVsva5ex2GnBoz5hIr8dceY0mUsNhj41zis4
u1plqe36+vBoosJWeEpYi6gzgA6ef9StugjAEONIcJ0k6MQy1JAFf+Qmceav8Prkam1ou83AQZOa
O33R94UYtzs5QM+H36hhHe8nyqtIRAbKqCVpJqMUl5pUOtXwIrZKoRBlGMUiKvPGas9QWPXw52yu
AHQJSN+ZoLSwVQi9IfxIt+z+Wmz2QNxO5Av5qBSlyMOOQj2wWg53hqQVWX/X8C69jw5Raad253DN
lR+xUpDN4iXFGgxIvWLyvGcPHry1ZEGy4FbVg/QPcvOUzuSImnWN3p7NQDW4qghvhyJHnheCYV8t
Gv5urMttikYNBVUboijQ5GTuXur7ZrjQa4SZDDnfYEPz4hBG8OAGnwMhHBDUKupG7V8h+hpei1Wh
RDCIVlfYQ7pBtp5LqSZ58ME2tiA/GKSjNkllAg84WaPzm2pRRy5lMRAFMPrCHETP/FA8uGVU0oT/
SYxORTFBd44DGyUBAPLlOTG8NYRz1hjF18u5VEtTamqww6WDVmWATZngk/RM9DnUM9UXiKry6S4t
niFoX/XzjbvEsw+ouqhPqJSfS2htNfZuM5wfp+w+Pn/eKUvDFlp0j4eU95HBrWjz766dT7RI01X1
KhxWw8OqNxbyV+I+q8/mhOt6S8r43LEbPRE6iilQBwIMHCFFSpFDagICllNqb044aI2Cjr0eW561
D76QwWQjbJwccyZuDHq3K3fOCFvJSbqi1y9T/tIFA9iKl3GhyENGZBTbeaZp9IrUIrqQXIu4z2L0
22ESUZTn25j+BPup95TukoQjk1pCVLaW4SEH6S6pFrSF4Ux+OQ0EZ5a7a6+RdmHAL2BLTNAB0RGe
KVJwfIEeVI2ym0mQcaJU/gbpumzXWRtnmWx/FQW6fuio0Vy1qaDHjp489qCuAuQK32b/hszkkdR4
VEFz6FjEZzGVBh3Cdk6yQEzk675uLd8tOkbfclZ3sjW2pAIhXzKmL9LfA3UHOuZ/10QfoAl3R0F3
o7GtOqIDPPEEUZHFY++7Uy6RJlcIHK8FJ0PufHmfYlYZKop6+Cl0FltQXa2oRprcH8Awe+lIiGOg
TWAW6+bxqIH5BeX0guVjsPDT3bm1K+Xn6WO5GSfBjo83Lqx8yNPKrMiGW8Pwh0ra42X2zzUVVEIt
hclSZ+x3PtSIenl8QRVZBh3VcUsbK/qR0dpLFyr8o7nJfXLh8qY6gUoz9y4EGlXs6v/0b5URGU57
32n7YO8DyXHLZIN5l8799MkkLCEQhfPz9RwFH6d21EjAE1ogEazi4i7HtlY/jObt6xwJVaTcYbLL
ZRNVwRFDXfxPFvIABSRbLp3v57wvVlBMM+ZyE3SR5qtQ6kGfdkOXJNTIvR1f6Nls/bAEG1nv1Sdq
7zJVA6d+UqXk/sVrnpanuhbwB+6SKYZCiP+rXQ8mzj/ANOmHsqsj9XGJjm3Ki0P2HN7MLR1MucsR
IUKJb6/aGau2Mg/Vz9sjVhDfYDaWpIKxZ8FWk/P1nEvta7jnN6hWENMFURx7h7v6M9yDGHskSyJE
6JRxSjXkQUIlrMLxvRv2ApKWRoy2oEwyFqXQkXqPE6PHmMP96640qYHY9zEqN4mp15rIoeCeXYas
hQbcsQ32CPaWt4sXMEuTrpoSTiqE9RKzAf/UyAIF88J+Hv4nyOHGhMR3dNlOaH9j+9MbeMA9lg+r
mvT+2QnRvSa0ovjnknmgDC9tbbisLpjT54kgp+z6Pr/g5zAggSlf7bwS8th6roqo3M9B8gwuVSU7
YUUpFw3MBXtmzn+C8ykgAdsl1p02CMMg3qouN3DND+3IcLHLnGM/s/MYzb4cMAKHvITIivwFR0My
1crzgQ3nJcRehX6au1ImLwvz3/emlqlRjAA3Pvl+HNorSHJ3zPQ/hsxxIYZk1RVzPL348lYl/VF+
HpcXQkbvdlS4ygM2QCT4jOkUSH8hl31uygsT10e4Rq0OBico0xLr3PVXPhIuk5RYn0RsVMonhuJ9
UIMqvs1+Eh+Mf10TjaIF0WObSDy5150+VZ9aqTFYxVER7JcXSMqPBDXgJJXGS5QbQ33VL6w14Cqu
h/CNeyoFfd9ffpH4TszcmQNlzxDjx9R83v2l+ylD2SSHYCr3Obywk8t05afSd0eUYiqBDWQ9C1ad
4eCnhA+w9EMQ5qqAYNON9xCpj2R11H1bPv6lZjQ0bsyhhrmM/XN6gdfMB3l1zkDR9PTHVP12cr5M
6YhDtlXEATKaCuPaFbC9k33br3ld07teort7pQq/rQ+/j3jmS8GPKY+3pyckq2IireQwDjiaEC4Y
NyiTYc5o/lu9yY0NdVJTFKdhi+Nz/cbDWxVIkbs3r64Aj/A8j5ycG5x2UfKkaugrWaKL5UtzW14b
NhiAFWeo6gj5ikShjF8jo2f77N//27kun3ymDyTiQwfsTEZSxmkD9Af+YcPDWbJ2eRyr7edkM3U8
PTprE3gGOjb4lR209T3UXAOuW8ejlXkf7RbI4sIilxlcmTlWKJfgve8u63Edq6npn1PdpuMFrWAj
MkXdTlyh8jP8tUUUeH60pElqi27VUx6DFwELtWjSJcGDLZYWKRnvv8KvA8mZOIrBmU6xGExqaveo
YajzVJFqvfY3JKdjEsLI4+raOOUYebRPZ57Jbb3z+UiJ0geUE5sLXwyD/bgm5+LXubMnaWh4Pwg5
2qI2+H39zCLm9yzZ+kaMKXoCrPMQ2Xm1RcEqDfT3iU/aq5Etphh7YFGX2B3a0rYPDnTiflD8Y1m0
kfK7xnL5KM04PnVk4AJzMVO8GGrq92hQ+tcnOQMp/GgxaqC/mR7d+VmyZVycbglBSqW4qFp0TAPi
57SNnwswjoH3HR5x9w05mFEYprALk7bl032xcScdkS/mWCrpOz44zR7M0yirzMM50Wc/9r6bWOos
2bIuLJDtQg90o97UvjE8QKkTxDZrpD31tmCZ2S39u6Yu1c154lIoRvqz93/F+7DMOnvZUbuSTX/T
PEeH0oUjQ8Qd3hUar2wobfcOQb9G5s/ZStFSjMEZ9bS5IVEavOlSH3Nocc6yA+XAIz1262o7RnhE
gWMX2NTmwdt8EKTwtP8oEDknQ+EtyZ0A5qbYOJn8WnCDQap9Avm9UcXWYKitgbDGJ8CKRCnfBviT
vexZLtfEXl/EIKc61au1tdFs3UHVuE+gp73pppVatMRr/2cwJHFLuJuGImcdQH4uGdZ/TMzsdVe6
2tG4iQmMAs35qhS8l2gpyYIIoA5yVs+a981arIga5XxexaZEQVuAok6Kd++vL+FgH9xjaedfMTJD
bze2RlndKU+dvm5A/HxQuxmoiT0AHLPi6cfMONQm4BNe3UweXXWW0in3dNE+SylBJA1t8uNFbf62
R7A3TekyWW7Q5GJ/OBUjojd2lnV9qFqxWxnU8MbtoVsak59DazjF2ePx1dkDTvyz/qW0tSnwHM3S
BowsNKtRKA+vzt8f3W7XbSe9G9iAj0X4SCrNrJgkLoe1wdGg+L9uPZedkrfoxHJDJ0022ZwUqkTi
tL7ZWMqjdegVbd649UXrtT2TfGMYpjukFLLGvV2L95SVCKIya3QpLfrMuSbOXS9Nos5usciu+5lu
gIktyvQvMNYUNWPX2w4QcpfUzA8G9cUMnbyBs2Qxvv44hQGYj6y4WAqGd9sTTAV++pJ/M9K24l4P
2SlAOvwRd8/smwno9oOSgwQ+6192rqwHCqCzM26rozm/1f0qTdtQhHx21wwL1Ipbcc9xRoSZ+lRl
iCDA4/d4GSqrP0GMZDozeJ6iQLmLpk2reGHikYQen60o0WDUG8+vr3jCOhAJZ9Xhgta9Cml6Q0Ov
Z+KWXWrNTlBb60iUUMljxz+TdnQWIeM3JAS4KO65670ua6Vke+mRylSuF1FykkbbGTZDyZejU4QZ
fgmvbazK8o/ZW9mN624ldbZfH7+pRPUwxgIrqk+xw0wDDQAgvtKAByWpxlAY+e90ZUJ8YbBsMkZF
HtMOPBQ8kLLYb+LDKI4PZ7VxEbmfOeSA6XINtJ5LSQIO0IUnBJ4YSd7zEmiekQnioiiWlgq3xyR3
kQVh9DiFs4WUM+YFml5i6vWeKPMSwkLo1RxjDPUi7p80eKkA9+VZ30ZT2vPOazEA8qqN3zDjQB9i
rxITdvuraOqTH2oM6EtUHa/NR6NIsEPWiOYvJHOedYY/htmMC0hFqxZAPI+yLdieaZ+GHnMqPKbj
1OeJ0nNxVgM4d/xyIUEJ9OZGZ+JfxDhiQlmmoFbfJ9uaxCJpAGtnK+MNPqclTrZBIV107SCTwf3o
Gr6Eq4j6x08WsssoNKk+qt/8nPn+FRw6QLbL4cvdRMiHTXhjkRhpulcZjjlfiTxJ4x6P3w5/XHDC
YZa0M9dOtWZCW0j8JZEjWLaEtG+lfQ73jhYRGpTKqrVDvWl3fIy1Rw29dbK4jwjo7rVBc9103tnh
49CQiqxym+qPS6YJ3qm8SNvOawrbh4aGOy1kYAxogmolm3AgEtauS4xLcH8v9YN2KSf43Pjb8yEx
JFbdfDzF2vl9EDUrpXjMQVSto80Flq5nQk17dp+o9HttE/eZD1WyzQVoriPcEejZXVaalGKNMGMZ
NtfRYLsKgYw06UBb6OqIjDh0HWjQxQsbEkb7i+UO+75E94439hz7jjJsKpLdRSRwQW2siE92E78L
WMT85VC9Newfg2q8M2GqCnBrODm4OzTEjyMrl3cf/TrjWTFEb8hEaKcX3d4h/jycdxi8p133m/Ka
dmu6lNu+2KguUCiHQ4hTg8KUZtdYC6C0qfnp0ZBY6uybAALB10JoBIaLGSzEA4VT0BkzTizQKnhW
er1Q9wxy81Rxkw+2dE46J2BQDyBHDUYKsw3G69awKI7wf0kTz6axTIEwIHAe4q/RV+sjgOOOGIwj
s+SFjawBKM1JIxp4XjyHZwdPKUixvXmEZq38yMI6jTPkq6vyBGtYZ+lF1sdMAyuYxRN4vpjz2kku
IuBew6kVc3iCt0IJ3xOo9Aj8s5XxCyJmcUFXLq3mbZXvwQIFBh/cyq7wieRTcJCi4IVK6O1zKNb6
NtHm/Ip+N8sSO/ntLbLB16NVi/LTyMtkDM77EdpN4kTgR/NfLSi0jXFcGRI1iDVbawe5FdeZLo0v
CgzgvVS0wHv20aX4ihUlt/LHXYwYqXL2MtALopEz/nLTztbkr7+H2Ovug6adlfwq/Cuij772qJbR
VqkEBEFOxzEwHQ/V1jx8pLWON07Ru3XfWkWsuRJnhFLGm+/TVhAgj2+l/MwSL/WSzZ/ffRuMrpiJ
JIbLnHaxcOonTnKyROWm8LxAOLDywEbN5icO7QoaFqebwJxxdX2+bg3ENwc1P3/nhTHPDnpG2P4C
6NnOQx3A6isCsdBZplr+elr4pwLU+uC7RHqi7AXaVAyCZrkfUIfH0JVbWpA8lVfzG4P0sVIrr/MW
D8uMY1yfy6GwUSGcXWypWIVZDuMPe2RvTdxjHFPMW2G1ti+86Wsc791bSpZUhjVyw0sBqWAv5oPX
F4goLVi8WwxNZz7GIlPBkbne/JsQaGED8o6VDOpDLibAI0qv6Yy7aftZi5pMyfJgJxH7p9f8H7pb
MCye+KIaWNu1hpLSquRg7Xbc52puDJNi923IcxHUMGryuXNRbzcEhTL1+Y0UewtxUP9g5cKDv8/a
B5E6uxC3Q3aXGPd+zIhC6VC9+wemOq+lZQXmxoBzVz9lEZn9b+/xRw6OhJhu72VIDsYqB/5dVYcP
NQ08P6OPfFt6PnwWYilrsLinPp22sWB6E49r39ObQZvG1lmqjD29nb1Q4DIjaNenx0TTebHAHKqM
BB1PHKTOsDX7N+dcWH5Ptagm3r/eX6Pq+39AWQjOZ+AvjsRMkKrULkk4eIOMAP53Qqg0fzNBv+Sm
1i7HRFCCqpIrmJ1lQhdPJEeJVU41yTgiwvHPtvrfg0s+rYNh4PvAS6mlGQtIoG/IkPbNZjdX5afU
bmARz14lBGJlOLFkPWeBwbIyEuRlLdq7/7dTN8Nt3PoxYiyhbgDLR5qxUOQv+kg7b+gEd4z8j2Bp
LOSjEkCE+pT7HWjx3jO5OuSj6DHxZBtrWHPzxCgs/wfSZE0sHXJHSWCERkuYeC/lN7vs4wiIO2NI
uag8ZDSpNlZmbE2mHlRspEZsxIag5Q5T5pmErLz3njqmqUwgh7i7Jno73WfOe8aXVAG3gMCdPSpF
xkYcn1q5WqkqpoXfX60SbKatL7yl8ZQ5FS6vkjj7kSfmF6FPg971rX0DMFLlsPm08HF2bi9vvIMt
fh4R/Jq2ShVpwGsTATixG0Zj8DkGivOlEtezZMPjvccG+RoIsZR9s3DokPNppNpf46g1Eicba5rp
p+baj51SeS0wSHDDCO9yOWzUW/DghPqusWnrfTgXepiH6fFItikF2anaVUhQpl+J3TtAq3zk/TbU
/Ora2u75ITAFqDFTUrONrFHWqCn17k/zaspV4A2CyCIkRV9LQIAabwzdVeVMhQMhE/ZNiuPiwQ3R
ku3Q7EwE2/bFggecxOX/QjbCVer343mpX8yAPGnMvY/6tViTqeXashfv+IrtXzI/DQOPl5oI/fJ1
NnuD/GuZkota/qiztqHFZItvEg3oO+KupNdA3crzgAg5mFWKoQt9kx4Cy2+Y04U4Pz3fQd2d4mI5
Q4FPd45+ZXmE7noFBGlhkgIaDBwQpna4ovTKbbfb8VmK2JWQbp2vWNCh5mKlSGL6o5R5LRGXsVsH
VRBF1wL+cIgWomw7hYtfcv+R4zLRhGrmWhsVU5CZ7YJr0grQ3XBN4UKCjzWd+MaZK992m1ff5neD
gtUYfoVTeYG7WfheBim/Au9ifrTXHPWFOpJzWLpKqpSnS4l0vZzvQimw3gRL61zSPzwlRdlM1TJN
zioyEaCIBGX9DmiorTRWSf6KMUK3PNipLdnnB4LTV0AgCEIP7hdgV5bbKJOBk3sY0g68Sj2S+POf
TCS3dHtBg9nLrduzloh6SMjeIqlQyL14Q52tRfHpdrlmTq9jOU8dihqExq/L5Q0lotXSv3ncyhns
CFwa1h/u5rF/GdQbKayQTFy0yfzX94cjCCrRX50BeoVA+o9sDVefHfo0SfEIbrVMF8QdyVDXXXUr
/UInN+COOH6FwJDlV5W1PsV+/yvKfZK3cWA01aX5UxAh0hMX5YtBazVbyXnizO9Cob+GB6DjawoO
60eNdTVBWwylfKzKVPohnA0w7QjU11G+beR9xJXnAi4d0jKDTn/yNSRx+F6zgpc93ca6ybVmires
P2RIijQKc2Jnmypk6J8gYjDMfD5nSEEmNgfOd47075QHl363gAWh4ZjDb/VUINztSkC7du++TdBq
xYY13HQMaqcdHqFEedZUwwxz4UDGoDEKu/AZuwHsA7AJWXH0SZnQ/Lm7f10OR5VRjILZKwUl7qYi
DqsMJvMBvX3YmWsgveZ9DpjS41aKxwPTnjmPejA+vxbKtTeR2ZJjyU6oBTAEEs5GDjImpcE0q/LV
UMo6vo/XFog2gtvNejTVrJ8QU3GWcQaH/BrbnYhyuXU265AsI5aPojzpOMtnhj2dkM1n9XFrsBVv
JA3aVU8p5j+WeuayWtEfdIY3nO4OP6vRlA4a90N5nm3tbRtIbR4SF/SCGS9bYs7g6nhCoNqNFon/
8/2Iq5gj7/W70zvWoUiTIHKKbyEmyJQiQS7UU20BLesCi1Z2s4/Q/rrIG6fYQ0sg1Yby0PQdfDQj
S6tGF1INKdrpRvzLACJcFl+jf85wo/ixk/ctHVtddOJAmHZYEf6QiMmx5om2ddY5aVJfXOEtXpJt
GudDDXCW2FjqO16VoWFSYxdbbPl4w3rtbWwmY80Vtgbc+sM3o0N+KrT9a3xUELrA0dZp+HcjpqKp
1U6/G5FA29OBdubgdYC1mWsfHMhyIQEJcy0w4+Gz6XMG759pl3bdlbcJaV9duWziqNm3o/UdI+a0
uFY5ZYC6Kje8INdsQtym0PquxsWuasyS/MF2ULxdOjqhJAJs0x+YfZBe3UAbHxvDVrNkqEyNHFRk
g3vMeVEQXL9Crb/zVxtQ617qu6O8SFfNYlvWHN4mq7xMFwzvxVK+N3qsTg9mbdUQOSZZaNxqOqnU
cwfo+pTst0uCv0mNW6Hxcvmr+uFOHy45UX6DOOpl4xSNrIm6593pE4a++KVLE2qK2IOj7DykMzmw
+e8nSmC2ZsEMz1NDt+RzfWUKcgigZe7lf04JDDYxg2m8rT5fIrEP5ndKWvKEouIOoZPMe+e3rVRg
tDj9Aex/lGrivUKOebPDInMOh0BBxsFy/enttvqoyssTeIUbSC7m3qqce1Rre0VhMM8z6paL9xpJ
2nW7DP7yKKw2/L4kgfWUjvXVx2fCy0u1F+f0nEYdE2iSvoI13tTHs3k/hf9iwm5cLwje6l6ajpG6
UMq0P5iucZcMAah1Tj6TqyXL+yMQc6Qn5nuu8V7FVEHzdvGx5NOcKQ6XvUKsii65ggbTzf9aAf6F
HQ4dwwv1h0q/G97IMop30OKpfXKZ2lUEvIQPhd7sToAsx6f2GpLzi5o27C5Eu/hxPmnU6yOkfQf0
hAf+lq0EFz8bcUoMP1lW68E2wv/bEYGLSpgs99OwPgO4Z3ywGy9jEch16A11m9aVVc90BHAtQvLs
i7M4mYejjeJSUmBpvSmlluEpvWG8WJ+g+5zsqMbjhjwCOsyjUXlFhZ0GUq0HHhYrVKD01RA23NVL
h412RngLXdtk0nJniCvy8UxxUYpuo7kFfKtooZ411G2CIg7GszLf7psWXjJDCYY20qIxdm/Ge0fW
7hdUWhWmUPCYcpIg23swjdTaIk14r73MWVYHS/UbESXeuSuwr68DMQFhDQB2Z+d2rDV6svLEpasO
cyUX72HS+rPKJyWb+lNzm5gDfVulsOHCrnjspuA3hJqNNoggJ1ltqYPee8Kntny39ebgmFNNAwu3
HpQwqNpKMkjtY0GfwRUBwUwqogS5oALDFFUTPA4xzlwtNeFRhURkydevD0HXoSvo5U2oJMR7uKVq
nCgcx1FZNrga0YBNyNXy6M7XZGs+QXNQPCXOwYolMjfctqdFr0rcX+c+dcFmE/tTil0lnKXsgt2W
qtHgZTZ51K0RJQeUfeP0Su5Z/O9gyMHFz7sFS9xqmxz/cqThUvJP18hSNx2p67dF+xmTjMwPyyQM
Jl1HYSHMpgyoNLJL3jnI/H9EiOZJt5EopIGezQk=
`protect end_protected
