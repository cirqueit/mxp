��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���|�)�"��(��	��I�ؑW�=�#5��q4������(�	b�.�ȍjG�#^㭤eΛ���.sq�_X�^�rj�!�FQN(6N����j��4����͚rA��&�&��b�ϗx���bV���G��/�q��h�u/��,��b�{|ƖJ��^�����u��3?��K}p9-�:eN�ar�55��ԯ����f��լ�g��m�-*x����-�nә��\3c���*���rK��H-�j��X�}���/��p�2�`�`W��5�7�N�bRK/�nMs�L���'�� ��;��0u��;�B�.��WG������	
�`�񶓳[�I�{,L��G��o��@�H�u�z��9�@��&��&^��	�=g�)�f���,�~�\��&�?�W&`�^�#}nП���qڈ�U��7#s��l��K�U�婗��o�	zG�0�KJ`�k���x����]E��]�r<���4��y&���r&MfP��r��7wh�iM�v�U��:��c4�\פ��Ϭ�����鑴i���4/{��j�6߅|X`��.I�*��ܝ����<��Sc ^����p�(�#�M��^��:B�Ƞi���Ah�1��ouv6�3��H�0�E�c{��,�~�{#�z%RA
z�oʚdU��}+�ݦ�W����]~O$��o[؄���#p�7�"B&u�tx����,��8g��($iD�%��i��)���9m��r�ɲ�T?�F��ʛj
�	��f�?���
~xE�� J]���z�I���qS����뵜��A�4�i�|[3ҭU�B���p����R�{j٤��7r���KC��i/�P��?���͑Аx��v.ql}��H�(>��^��?� �B.���|�wm�X�> �a�@k 嶒x��)��i�%œ�a3�ճ���\:���H+<D({�g��&�hg�e*�KB^��0.=�amc5�m
��x���D� O�LO�Q>�,�b.�����հ��a��P9��N�����jE��%�F�n2�
аX� %8E&yu�gP��E��2v����F.z���d�~z�my*?w''��:���gs��|PWm��_SP�J�9(f
j��92����91��ԡu��~��tI5XRKR��xd�R���I��_��<KYXPS���[��,�9N6�-E�Læ���r|
����A�P �� Y��#�A��:�MI����@B�ذ�~�� �d��t۞�}�� #d��;-�z�&Q��,��]�ڇ�e3a
�%�Rt�,G F�zV{��`�"��K�k)У�1W�v�+�h}9��>����:��ʫ����FM�݃JR�D]jd1�c(?��)�].�w��{]OZ�$��aM����x�
-���,�D��A̑��9vB�a�1f���������V��˓�P��t�� �Б���&u|~���T1���b�`9WJr�d�1F���M�E�I��b�Ԛ����1fҩ\�9��\M�������c,������L)�����H��w1�l�/���8(�kW�YO������[�j�Wn�vjǤV��<�i��J�	�g�"O��e���g1�n��Nݾ���dĀ�{���/N�P\�3u���k���H����kE������&-]�.�����.�y=s��#3��Yk���S錭��&����k��-���g�=BH���0�î{��ג��2~��o��=��P"���w�|�f���EvK:���9�aΏ�TQ��4�@4�@=����;��8��gM�n(
���o~���[�\������ǜ޼7�>�T*a���%�3��#�R\K弗��gpZ�����ߓ��f�e�+-C�Q���m]��Ou?��U�<%�_	H��"f���u��!d�)�� �*a�N�c"�&_H���H�X>�����vC�R=�MA�D���*GH�Zo�.�eA�>j�=���Ex�����7���Y�zD�4AS��|�c�l��]\o�d��1嫗إ���s�Ҹt�!�EDs��`�	&�:˩a���b���ȶy��&S]d��O�/<��T~[�~�WW�$�|JGQXW�O�-��;;�y����m;_��w$է�0p�U���z��~�����G�q��G�N�@��4$ȸ���Ma�z�K��'�XJ�s(��o��2�W��kM�8��(�kU�ԟ�7�M�fP+�*n3�v�yl�^���BPCP�[�����L 0Q5lL	��}b���H\�(Z��Q�����ҿl�s���	/e����n;vm�!O����@#��PSw��*�86�=�Mӏ�)��Y�K�|$9��g���8��&���s�^dF�b_��OjԠe��RHE c�|��ʸo�\��
���y�{�LR�������h~լ�@;���a��豾"����hm9�..6ZP�Jla)���Hm��uWoF�%��,`"��)�X(ٚ�t�w�tn�RZ�����0e���wVO�������Z�؇��+�-�>�m���� �I&��S��{&&<s
W����D�,�� h�K����D��}���鎀mdBI�;R��z��96Rd|�d���x��l�?��\��*�,����gU�PQ��J�?@�{�U=W���]�D����x�ҩA�� �y(6b��)g��)$�C�d��G�5<�� ��I$����������z=�[��8�� t��O1�,~y�5F�d�=�`jDn�;���u7�Je@_�'��8�JU]]]_�'n�kW�Nl�Ni�%.��i�q_�*�Է��ŦU�����Fx3�	F,�T�IGD�f%J�J̟�bnBF�%i�:~���OE��:�h�70RRlp���q�n_϶�*5"��(�����S�y��;X@�'P���������花���&�u��̂� �� ߽�����~G2A���?�C���o�Z�:�BW@1롞���oi㩓�j'���W6ߧ�m�M Ҕ�����Xb��˸kB5p&Xq�W�uT /ݪ�z b�0a�z��a�|�,^5��|��QT)|��T_m�|�-����R���Dt���$�P���CZXh(�`��LL�)�r�IB���>DsMQ^r������i_��.<)R/b;��u����ߝO22�7�-N�Pe@���6#������:�c�ܠ�"�.#��u�T��kٳ���ƒ
�g`c�������>N�3��ȿ��9�8���>�=JL����!����5�X�T�g��uR[�|�_+�Qe���:71+��|�{��"�ۣAJ��2��i�l̛�}�^�|Ѷ���W�Ru�E����"�U����w�v��Ʌ=zP!�~�㹁S%��k�����+*X����+�R�
2嫗��~���
AeF7�bZjgY�
k��T�g}�S%!�$����xdsy:�����i�Wh�>J�UO��C"����~�+��~e��CɌ���唻��5@a����v�8�k ҽ��r��.���S����v�od����{Q��\h�j<ޥʛ��gXOU9$y�]v(f�h�z'W�~�9�V���S�g�c�J(��/�ͻϥ�l*�c(2h����Y�t�fa��ԿA�a�BΦ&�겅d��x!֒A�غG�Ek_}O<�w��dr\�����lS��Ax�g}�l<�p�d��y�R*�Q�e�N��
���s�8q�J�{L�]�����R���I4��K��C���?�gE~�;M�VqM���:�\����Bv��o�|�T��!��Z�kl�5�ro~8�N�SWV�B:+����Dt��$�f��&Q�gu&rv�v��o~�j(
����R����z�w�����l�G��2��`2҈���-��UM_���h@/@iM=A��l�Mʲ�ԭ��-���O�O�8Ta�z�������;V&�6Jw\E��* !����;�׸׮�Ğ�)n`{p��kO�G��ձ�(��1}3��o��� c��6  �7��t�|^#��3z쯝*��3�b�k�r]g�K�*���$��-��C�\~�����Nt��6I�!�G6�p��쁣��G��Tgpq���������ݫ'��H� ܣ�?�����>�)�^G`��ea��<;&�"�lе��V�w�L$�1,c��sn�� ~+%����:�j<�K���Nq��[��th4��E����L���v�BG|�,��ߨX���4T�6^QB�c��ʡ� sp��:��?k�<���\�vR��TRI�lm��k5f���f���ě^�$�C��}֎>q��]W^�rHL���j �J��E:+�Q$㈬��c�m�7�"P-��>zW��eK^��m�2�����W�>�怀t�3|7ﯡ��#�z�2�,�ҫ�XK�������3�"�5ƿ1ԁ�+�X�jق��2��N�f��r�/�G���P�o'u�����Ʈpj�`�<�N��Ω��[_� ��^��E���M�Bn�;i�����"���"���]�?X$r�71!��y��#�y>�cd ��.�����A��{ 6����l���mS����|�~�[����Y"��q<M���1RH���h"��0�:$���	L��N�0��4����� ��s�KÁ�^���aI/��f��u��r�gMPer+����n����o2�~���%�_�(����մ+���Jވ4Jz��j3"{���	����!��	���$`����-�\Lr_�P���䫲|��`Hj�W�r�Ql<��������v��<�`i��dS�T��]�ȫ�M�`lk9����D)��b��2��)?Nܤf����odNo�Y�=��C8!�{:&~�)̩�^�^6����\"���\&��$g���K2���G�F����V��=���ҦN�E"aL�v���fQ!�ҷ�`�	
#-��Ȧ�oː=�ZY��u݆�h���Z�J��pEt�+sw}n6F�>4e.�q�
�xC��`&
d�US]����г����^讆�x�@��I�#�S�a�/�=�z��dbK6J\��Q�
�.D���] �B��H���)%6�FK>Z�7�_�S�#����j���#\gu��yQ�� �rK��B��L ���$���oOL�$n�G�C����������$�)`�$���r� ����{'�����6��e��9:������`;��X
)�� ��� s�����b	ړ�ܷ�D
CG�E��-�/�\�μ��O��|Y� �3%���~A�X~��a�ؑ��a�;��&��,L�`Bj%OҭVm�-��F�h#
([�S�i'�zlZu�����s 0x	�J�����W!֡��;SZ�����y<w!��[�����k�gI�iY�h��WF�f�����Bsn�g�m��Lա��ᖟ����*�e�0������$��e���_��kZ���_y�w���c0U~�AF)@�0Xm�@�Φ� �-B%;��*��&;�SE��?6�)��n�.�����F�<�����~�����z��%�s�m�E�Oʺ2[˺�1�q�w����"��bS�U��n2���U��%�٠E�|;�w���١h�fd@���Tc�"u�Js������o˞�Q�Bᨣ�� ��ƌ�ofȦ���ן-�\~M[��X���M^IVH�%@�uZ��w�뭲 _s����}(?������?�� ��RXC�-������C�6�r"��U���e�9�]T��K��$�� �[�(2���4y���9��m���/��j:P*ZEO)ّTZ)��6A&���p�z��: y�
��ī �t0
��Ce�_�3���'��L3e޲(��شb�ȼd_����*)������W�Қ�����Ǧ��ɩ���f(AA|�Z,4O/[T�AJ@T~ߛ�J�����9#�E�	���S�m:����{@�A���t�̵KN/�z};ԉC|ܺ�R�}w�ݯ����Q�ȴ��-m<��Z����A�O2*�mǍ�i!b�8��K-�6�5{d��Z�:��� P����
�b�����)y_�*G?��!w��QΜT�����;5�a�bs6�r�O��
��|&P��R4�2�<�e�\?��.�tI����n�"�5����\��g����]j��~&N�'��y�QȲEW��Qr���P��.XP�-<���F���Cq�����#'�*I��N�i����j� %�ǘ�r��(�0Dp�T|��6����P�Eiܒia%e�X�J^l���+���f_�msD%eƿ�s�z���K���z�AH���֥��7��5��<E�QJ��s�I���\դ�ō?3Q�$U�Cp��<�6d��Ub�g_�KBB�Epԉ0�������&xp�� z��O�J�~�%���:��� B�U�����AT؀�#���x	Y+�s�㉿�ۤWFG?��$�y�:�8��l� W��>R[�3|�=��X���P�1����x�4g�� ��X3ƨ���6Cy�n��K�f�p����hզ��F=�kKJ�Jȧ# �sf�
.�-�䨅1v�n�#@٧e� �PP�e�{<�pSi���ꤢ�/)� -�H�Ǐ2��x[!�9O�@�`BD�)heIe[`��{��1Zx��%�����p������L����]�e�.{ag����.Ci���f��Ʊ[.�M	��%�J�|eA���.Ϭ	������I�r��tLk�aZ��%d��(�@؅L
Gq-Z�?�#�1�5Q����'^i/�Zo.w�;&'c���R����{��jM��*�G�$����m�cܞZ,��*���;���j�5�'T)p_��x��8�S-������<͍��eէ�2տ%.��m�B���Ia𘭫\A W[y�j8�8�Iea�ݒceap/	���9s#�hH'1���$�o�U�#J�'��(*Ȁ�����Ӟ�׎��!E�0�����*�S�zi�0Ih��3�sjC��i�|6�D��R�hs�ı�Ic�R��K1� �m_E�fT�ТT�@$�2��ٮ߮�8C�d�|�I~��Bֺ.�8�W�I�_{`��-�uiC�b�f}�iر�t�Bc�J��Q�yp�����?�X��=�f*��+��.N�vJ�Yٻ2��rZ��HJ\�!P�}���,�z�M[�Ju����݉FC����/�Y��{�f3�E��Q�SRYK���o ��������a0��Jt]-#�zuoQ��n�Ȁ��Y�����|/ɺhw\���m�d�TlX���=?���"�g"��;p��]>�Ήu�ۆ2뫭���)�g�/!p%[�8 ��Fe�8WR�LD���`������ !Б��#)}�Wh߹W���Toe"q�6ςz���4��6���5�O|C.1�������pT���Ɇ1`b���m�5P�DC��>�zc��;�!{oʴ$�ngບ�V��C��'��2�U{ �bC��L�-u��#Q�./P�	��"�ߔS5Hը�;�%�"�.�-��vcnlS��q��.����PdS����,��w=���m{c�o�F�5���P��$8�h��>��%X߮�����}
�zu+`\ �V�[r,�`2��y�Y]�������('��6ψ�����4�ڪ��k�'a�����$:{h�VqR�K1��m3�~�z�� �M:w���cdE�SyL�>1&	������(&2�SS9�����h,�<͡<��SĴ+�v-�������s���(�	�l��C�n���*Ҽ�GL[�������,1�}��꺊b�_��e�T�Vscr�s-%�_b� �Ε�r��x��&��n�gGXE��K����� ����=�I_��l�nnQ�Y���Pa�����j�rzG����®ǔO����"N�5[���<U+�=��h�D�?;d�����k��A;���4�4ej�5�T��$2yo.�!s��f�&������l=�@�[h�j[�|e���QLq4�=�U1�,��k�k��	��]е,◽�p	���3�~�D]�GA0wmǩ��4���% D��oSl&�
&�}�.�J���Kʆx� ـ}�6u!_��sZܦC��	�2q��c������V�ql�6Ӷ{��>��1�ھ�-��	�D�rV�$� !\k�>��(xt6�Ԙ�F�x?lk[dP�v�,Me�C��zz`���:%���i�NIzH�uT�G"� Hώ�#f*}鸦Tƪ���;���Xu%m�/�u���"��6`��C�U:�^;\������5��gH
�'�c�ʹo0�.���~S#���~��u�6e~.[ʖ���R3���ĿV��C/mr����g�M �{�Y��Q �(fD��7�9��W��N-C��w9i�9��$Ì���L(M$��lxZ��d��9o��x��g�r�`3��ts���V�����-�%QY��2+���NV?A�C�Cn��3�e�/�#i'9C�gj��W�����L^��L9gH.I���a���X��y�2�l%1d.a]g�~��ךЦ�=�:=���D���H|�le'<*���v�%]@��{=�٪f�JL�;K���^^�G�k D1![Z�Ԓ<z�2��n)>�W��o�
�1�T,ǫ�^�Sk� �$�&�?�[�"�眜���0��B�k;F�<��+U�KYύ�����!�u�Q����~@/`g{.���eN�F�bI�x~@	B����h�`��S���L5&[��ܙ�U�v�:�4����O���/y���T��Bl�d}��[O[:�`�{jR�
��,���%�ӢGy���ϐI}�	�8��3�%Ho�<��tK˒�U��)���)H�H.��7�3�K��9����I�W��Y�I�>�V��_�3�-_B����PmutiN��-����7��Í��^���c:uS]��dV���[��I�7 ��!�
]D�\f��֬Gq)�>p����� <�
P�����dǢ��*m3#��_҇�ʰE]8@��4v�ھ;�1%�a��6ڵ�/=���'�	���|TO%�]��*����� ��ۦ��Bѝ�~_�KC�Xm��/v�
DL IS6گ�Y{T
���[!By�d�_���]3���$���;��Q�i0��\]��5���� ڙO���<����/�2TY�Jc�t�H\(6c������m������#Ҹ)>�jf�B4���N����%S�ag���8d뎨zN�*R�xS���:��w����X"�I]Yl�:�3x}���ι�S�@�|QB��:a�&�j��s1ߊ��q߮�`�t��OLo���G0D{t���~�`�8�4E!^JL/���n
[s����L_O:1���J�� ��OG:���{[^�"%ƨ}误qs崵u��J�� �Nb7̘�?��	!�!���ժ�]�ŅK8����SC���d!7�#_��g��ɕ��GD�$ùu�o/��u|[�ĦKO�������Z%��/��FX蠎M�������L������r�2]Zi�cpU)P�e�s"E�d�z���
M[I��=9$)IҎp��܊��<�8M(����&�& >�/Ɨno�|T��^��b	�.Ce��T����Y�
�����v�׿�9ΐ�&$�@v�##2��K�Y�����(@���`3珉[s����
˸�;�a�yV�Y��U+��Ƀ��O���CC��*f�)S"���osI�J1�`�.�~$�AQ�"ٍ�?���A�$dz [�Me�D�>fZ;�z���ʯ��Q�B������D�������˼#�JCe��-�i��r1�ko�&}���C?I�_7���|>j�m���^�!��:�lO����Z��wМQS-�f�}���B�ڵ
�[_cĳT���6�����3��[CI��J�)����R����(\AͶ��8yy�EjyCJ�K� ����!*�f�˸lĽ�-�ā��8ٔ�Q���[����B��jwX��3ؐ6�7ZD��hH畽�] �������:����\�2�kR�/���
R>H#��]���ú�aY�̃d}���${,�UI�rG��J���;jǕ���Y4��:��ye�q��_7ʤ��y>M_��]߉��W5�K�:dw�q��9쒼ֿ�z.0��%�L(.�	4��FN�[�@���E�s�W B)���W���T�,[.�$�>U�ɕA����H�
;����u�=:���ms6*Ӂ�(%a0 T��d�8�Cc�T��[��+���[7g���1���f~aR����qf�*��~�iI2="���a��x[�8�kZOea�h���CE~a�Y'�.6�d��ܛ%-�ד
n9����>�Z������;�"=�`�3���7H:�t#�M����:�,A������es����9{���r�+�M�&�gJ�Q��}�툘 j��"�l�,�2�{�g�D��?�m��!؁{Pd�譻$��[�^�_���� t�l��7+ŨE!�	X��ne�v�ur<����Y��͗��;�I)�g��!��X�6)�>�x#ف�3 �Q�y�ރ���6X�k��,��;��S�`#��	!��Y-������s���i-Zd0	��v����S?KpO1�����s���#F/���f@�*�����7u:<V��z�9-�oQ�	��Sگ�-�`�qi� 3�5m4":�k�4���Zj=1��u���?#�������k.P_��3��	�o���eW��m�_����B�R�;��A�xR�|��N�ᶳ�B}�+�{����[�f�KA�Ր�����\3JL�+�KZH�׹�C��	�%Bl���X�%"WK?n��4��r������a��)�}}�5` �F��Fp֩��Xyhx|��%OP֨o��̜t+͘��z�Z�D��up��#�L�z����?`��?���iyJ����Ş�I2o2�j4JH�j�L_���ܠ�}��_077�n�7�Sn�a��q������x̎�4,z2IƬ�}�3�6��|��g �6Dh3@�P���e���=hV8��k���a~�\����~?�4Cz;p[���F��H=62�XT��9[�;R�F�@F~�*Lt̫���,5D|�1�v;�?d��m|ȵ�.��{{�2B��ܶ�q8|,����nH�R�@���0Y���3�{[sD�P�b��Yh5i%�`H�A�
���cgNW�SCG�e��A���˴nfzs�05����;IX(�g�h�ꧤWừ��@�\��~ֲ=X���a�O?$[L�$1�X{���p����W���#ǭgѰ�À�k���,}wt��V��m�8!����g�9�kؖp1�g �X�>�'�݊G�P�lL�<~�>i�ƚI߸=��3�H4HE��4��tl#��T�ɘf3�v�����!缀8�P&#'�}����������qN�6��34w��JU'@�@q�ЫҋC~Z�៻�OPDY��	�7:���L���;זރ�%�{�TI