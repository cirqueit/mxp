XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���:��J��4��B^d�l&��943Y���J�1:�hm����L`��s݄�J�p	^��oZ�M��3�����Du/� s�Fح��1P�Q'[	��s_p �=X�
F�[������&~�{�cc�a�U9����ǔ�g��V|��)m>MCie]���;�~e.�M�+\xzit���iicR�����(��Q%�D'�J�`�>g�@#��;C�K�4p��y���9V=i�Aj�u'��m���oA	~ Ň��gy�N�Ʌ�OyϾ���0��i#k��l�ӈ>��o�)��!u��*�B�����Ƙ��ƅ�6��Г��څ?�̗���˞��Q�5s�և� Z.�{�Jxnε)���T���
�	m3�e�`u�hc
r��ʋ'\Tȥ���jM��]חҪ�/nPO����㷄�tD����>&�J>}Ji�+I#�|���@G�"�?wm5�E�~��ɐ�D0�7��q�	,��:1\�U7+9Q�	N��a;h~��ȁ��S;����e����%��{.�/�X�%Y���aTh<�Oh�j��_�u�iy)q���՚ <���އ�Dy��.u������B���P)�$���8��#S�.�p�kb����_n'��W-Nf�-��g^�kz�A�ȱ�O���\���Q���.K�](�j�Ǵ4�d �:6u�:������oŀ�#���9K�$6����@�j1B�b�9�)D�7V�G���}�)|���k;�;���1��[�]XlxVHYEB     400     190��!�8��H�~L�T�"ްa�F�͸��t:�ˑ�M�g��
z�������J�z|�Mgᎎ��؟�/��Z�n�?Ȼ$����鈎;�뉜Y@⳨"�QG�g��[�3p2�ţi��"C��nY�S�#��A"Ș\�ەf�(B�(����(��D��i�K�WvŴC=��|����U��t��� �ɀ�WE>�^�;�����^_Vphѧ5r�O������9c�l;$� 7�䔣gk�*t]$Y��G�<
��-ݬ"+�Y�'�����[��y \�E�&�$�s+�azn]�ɺ���� �^����S�/��}���ۘ�h.�P��̿�H^�3*f٩�m|���x��֧E�;9��x�tP�v�_բ/�r@0Jͺonk��#�8XlxVHYEB     400     150��Y���R��"S��[���maL��$)�18��E"�L1�d�j?��ϼU��q�k��h�N�usN�T�*���	Lgs�u��MoT�%5!o���]�|��Uo6[�e}9�\W���]&A��dX��~Yb8����8+_Z����՘!��i5����%W�4$�����^C���T
Q���>z�[g7���0i>60���QFT�Y2n�Kw]6��l9/�!%Cj\���JxrB9{ ���ъ��� 
)+5�6�{�w->��� �V���ܣ�z�D�ϸ�4�q�������C3V�G1�k��|�W�c��F^XlxVHYEB     400     140��?&�� Nɺo$�G�+�>�5��e>	-�����ZS#I"�f_u��e��K˥�<������[Uoƾ/�4�6�:��@rR7/�VDFW��s��!tOA�EX=Cy%(��c��גP�5��1D��\#��`)Y D�qd죘u���स�RGz�x坴K���|�|9��2xS%�A���p�*fh�YT
�%�V��6�%��zӴ���3��^-~���v�����@ʠ��2F�[
v��}�j)tj�(�'�B�*�z��Iq��(_.�E�h���o���������,Ɂ��XlxVHYEB     400     180�|o�=�Q��HESti��6����w�'%��z���kUJס���t�C3��
>���VQ⢽ �D�寲mXְ:Q�Yy3��t��w�@���G���m>��Rf�~'�=a�M�1�c�d=��E�lJآ�(����b��0/�-��?PFrw� ��_{wV[?�["|��>�=���r1���쳢a8�����x�k�]��u�7�Y���V��f� ���W�{��k�Sp&5�,����)ז��x��ޕC���߷RFwiW�qu#�)hP�ѥ<���Jے.�ϧS�Pn���N�s�U.��g������� �*��bd���m�(5�:�WTS�H��4�.'�@�q(��8���}��0�tZ>{��|���݃�h�*XlxVHYEB     400      f0�VF#��Z �����Y�.��5v>��#��D�c6JF�.
k�n��r�����Ij_񋰚CuL���{ 	q7��$�"�y>�G�rNݩ��W�=%�_K�{. ���� ��������; #�6IpT�SLʾ��?��\{����6�
�gH�,�:���piVBzBn�ɾA9���J�_0c�Ⱦ��:��h���!�a��@�=U���6P��5!v������h+�"��XlxVHYEB     400     150k���v^���S ?Zku���_��k4d��8P�>8�@��TG4m_��'<xh�N�j?*Mm("�!���)%��//㧰יq�m��x��`+�?�Ո�@D�A�	_�0M��	N
x�t�kj���^���G��Ƅ�{���̒������ ��rhV���xn,�������_1��0��0��Z��P�tT3� �D9L��.o_0gvq��Z6��=�s�5l+q{PoJ[$��WJ'=�i�<��E[����eB14͙�XpU��9d���db"��-e�=�Ӏ9�}�qr�����9���۝nlv=VB�p����6�����;1M$X8H�XlxVHYEB     400     150�W�N�jb0�L��P�s��L�bH�ɉ�h��?uy��a���/+�%*]VE3N�۪`=� f�%p���'��������rt�}�#�;��6YDI�UI+m�A]�o���R�����C��;��D6>:A.�j�pIJ��Ԋ�z�@γ	B�������Q>���:��e\�����z��h�ї�.\������Z�TL�
���1���M�5R+��f�W�|HW����l�2W�uF-��1Å����r�d'�WtO���2�ӷ�+s����.��P�½e�*�7\�����x��o��)�u�S�7�F&|K{M1���(>o�~*�XlxVHYEB     400      e0�s"y*
��'�7㒞�z�:���,92���a��;���R�^�
Ps�u�,G����%�d�+B�T:��ո�0K��x�BB�w+�F��p��Ɗ:��Bt�m�X� ����˺V������� �̈́��-0	o�q;3���ʚ]Ug��n����aaϰ#���K��	�A�lH���ޤ6���
Akg��x�V�a-�Q;+F$o��M$<�RXlxVHYEB     400     180�m�н���Z|��KJ5�]���r�L㐚��n�L6�1�m���X���aQ���yZ�1U~9�4�cͅڌ	�}��)��D�<��[>�� ��;-E�)'C���m�v�z0�Vf�PPITdz�tU����:f�6�ϼ
/�Ƚ��넨LfǸ�C��1W���������(�%Qz����5 �ʤъ�
V���9-���p�%��,|!y/�%h�7��q=}ьۣh�
�4!*��N/�j�9�j�6����ZF�в[3㫖	ZX��o�(�蔑��대J,��:��Ǫ��>���8������c*qD�\~�ž5 w2�Ѡ��;��@�o� &Ȩ
�M�-O����V�E��4���O�����~\XlxVHYEB     2f4     1005�?�� �&��@�$�M��А)x�`�O�@v^�gs��&��]��ˋ�v�+��(��Y?���cd�����k��L���j����>���m�&��]R̘�V���6��������J� �(����?��
P�Gէ�]�r�Vd����i�����R1��_ڰm�|zRIG�+}۾P��A��x*�\5~��ʎ`y�h�*~����1�Ќ(�Je8]�'k7�߹<�>9�������}q��DJ�#��{