��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Лo K~��9�X��Ȉ^���ji)�z���C���j�U�8gqP5C���!KV���Z�ʀxz�p�qm��W����z���ף�^���*LiX��lӃD�j�}z{�X(��u/��rᥲ[ȠQ�/HǤ+�����k՜Ez֙�I��+�Bژ@��O�y����3w�IPp�+t[�c��*��j�$�V,yp��Iu޵R�{�l@v,==�΁�_�&K�ԫ6�LJm�R���!T%����V��J}�9eVH�
�e��fC�3���bD��&���V t����K�e�ܖy�F�b'"O�*yR��+
{@�' L6�!��pw�|T��:��0Z>�~�D�:�jB{�45�y���y�h�j
�<�:j2�}��<N(�U�j�G����d���ʲ<�(g��9��δI����;T"K�<�6'�H�u+�>���ٲ�������@vlEjz!���5���X�x%8]w�!���x�h{��B����`����-�z�_0��T���m��=� ���[K*�jb	���h�C���?$�#���՜q��ج�ߒ�]p����h���G��U�t����}f�Kf�v���8�*q����ߵ"������2>�����.��ў�/	A��-�����^��af�q8����Vc��L2�칂\a�����z�v�� Qs���M�A.��G��	fN_��f
{�~<83pUIMY�GiRѦ40Urn�&&�q2"��g�#��sTM�g�5<�=nk�X�����Cw�BAgN�E����;o�;#6J�]_����[�е i�o|DЇ�NGp���Ԗ*��2m�Ə���)8M�d��@���-5(-;nj�dvc�]ǵ��͑v*�-޺R���p��Kͨn�gЦ��}�f9��G{9"w���(�Z����H��P;{n�V1�98.����o�ԉss;�h��VKA4;�N�X������V��O��z��>�H�s�f�J]{+Cz|"0g�--U��E8ʪ+��y�H�oO�++>P#i��_Q΍���0`����9��E�y�`Vf���:cՇh��6ٔPݙ�(G^��5�O$�%��؉<^�K@?�N\�L�Uy� ��ߎ��_�o�$�f$ G��{jշ��j�����`�`�6�YZ����3��r=���Op��F�b���C�,��v����$kQ�p���/�XοI��/Xo9��y`�P�O ��/�=e	�*�B��\A�*�C��<^?�
���!��x�M�7�9��cy&'�Dj.h�#j�L�&_C�%��tW���qL|��ۛ�in
�I��'�L&�%�� �C��4��UE�P�UЧڡvH���X}����O�gP$�*��7�Ky��sx�f���"�4���H��N	%s���R���}�G�u���(E����ٵ`.�k�%�o��L�7�SjX��T�.�a�}`�Oq,Y#�BejHS���*���pssxwރ�_\���6�3�g���K-��	��p�E���F���J{��_9�Wi0,Wc��|��boiW^]���f��?��]������NY��$cٌw�ޢT��[p���_�&���/�� ����t��x�3�*���ٽ���'Na3�N��RbD�. �S�()�}�5r����ݑ��K��d��F]�3���,MQ%�,�nP#h��;6�N�^��hc�ޗ1��/n�ɽlh1b�NZ>:���u=�Z���a�C��Vu)^���8�r��H'�k�^5_oL�ފ�ʂE�N�X����ݿ�<��.�xox��X����5���{݂�o�^�G��ِžİm���+��E��9���wz~x}O:���&��)�\%�Ydw��`_g��#��-W�^
�)A�N�	��n�1�6�dd�h�hd5�� y*��h/8���s_b�JO�QbQ�k�p��Mc�F�P,9����߿����c�$����qt�u�{Gy���n�]3*	����'��N�.�>��҂pǇ�2��+����N���߆|��p�!t��J�(�+W��:�O;2<V1!������bŞ*�m{�|	�,���9��&?t�mفj���h���Ѩe�2}�r�DÍ9���8r8�v�J~�]�bM�;�]c����=f���o;CkB����l��fX`���u�	5r��j���� �UX�Պ��`��i�+��z���n�K�$
�=��-�<ӝ(&�w �D�z�����T�ٻm��@�6*��* �|��`��^�׋t(y���N����a��8o�������g^1ώ�1���";�����I�m�i:�_�ա�Wי�kQ��n�L�E�҂̹����ߴbqM˯���R�>�!b/iJ����e� ��7��M#w/?��.���{R��\x߅������ �8 	�w��T��;P%�(m���>L��g &�S	�w�9(����*¥���t,��-�w}��˨�Y�Ae�K���5Jas�a`熾�U/x�Z��ٛ�>o��ۻ�Ǭ�/�Q�g��W���Ω�qD��q� �#�e^X�M�nF�х�[��TC��ܑ��g���h�����p�GC��I~��!>(�P?�dFⲆ�|�Z��0�pTD"CTr�z�JV��
56CG��]2��'��-Z�����ZƂ�y<j.xoU�I)�2��_�����0�x�e+����w�B�{�Ғ<Z�S�w0�ɡ����ZuD9�Nc;�̌�7�^�ݧt���X��H��m�6)��;G'�M�C5�r�sU�����=k`Yh|:0e =�&�	�0>)1?�9����+q��W$&�u��%E���~V�$��L�p&�$aӕi��\:��A$�(�yI����tN�ȹ�r�	,hڅ�#�:�����\U�2P��)|[?	bl�g��|���<:71��[C�)=�(
�ɫo1뙪�����(*C�CUi�-���K:t���,���m<��߈R:m�݀l[��	�N���ъ��S�w�� ��Ȯ�<�߸8|�|�e��M����G�(�8YG@�LH����{����|ZO��m9�bqÎ�Bv���D�~CJ{�)�y29��yL�-F��>������U����O�F�b�����G����6��]������F���\�<�[mm_�zu�w�y@�şj5��(��{~�cʷѦ��U3�!��*���T9`̯��o��4�A���5�&`x���P�bz��F�y��N�ei�����q�ǰ�9�CM�R5�F`�m+������!|��5%�4TT�|�+�A�x��uν5�G����=�u��Ӱ�d&̹<N�c��t����@E�ͅ�|��3@2�Z��PzLx 	Z�De���m92M��ٴ,�Y��K���z�(�� b���1�����m
י�81?�,Irx�O�֗<ܜ��g���p��P�]��Z�6_��z���A�<b���\�}�X���O �*���9���b��D=�2μZ�[YE�q/|��m����̯#]��i��M��ט���������ʖ�/�Y�6( 26í��჻�w�+gީ�=�F�C4al�]���\% r�]ӆѺ^Rμ!~���UH/3�d���pm�0�-�/A��]Wٲ��/�9rF���P��&�-g1�<��m(xo�&.�m�n�P���$�&��!k��S\�(7ZYΠ�ue���.�8i�!e��-o�!g��mM�6�{ ��W�l��B�0	B���a���/gl�^� p�M^	',�.���|�꼹���eɑ1(�e]쁡�Y�Ga	1��()l��$��U4T�}����,�,V�u�9�P�r���������/4�ޠ~2Ul�qfp��ʷF�k���'5yc�W�Y���X�i��5^�p\o[Q@W�4rmBq��t��i���]0	ϵXfx��b+����� q�y�J8���_��u��7�|�U�<��t�q�(��	*A�v1�o�R��&��:w���%�鋷)����b�~+}I��$�n�W�,CUk��!)�7G�o����h�vu�1Vv��X@�v�^`}����p��D�[ ���M���n�����H��9!j��MzD1Xp�ʀc��@��u��נ����t�>4��/�������H!��'�pa%am!��u'>�����1�h۶��Ҩ)�rv%8N��a����w����-W�.~B�Pf�����#y��%f�*#��\�u4�����nKk�E��N�K�,�������6(fDpz5��	�)�z�`# 8#;�r_��ŰG�+A��[�Ç��5�I���]d)��"&������@y�*Ttzo���Z3Ӛ�6"��F$PWE���4�������2��I_[|�4[8X�d�����cLW�l<犓l�X������ο����dU���i1�7�q�j���`7H=�8�w1�%=�}$�-��7d@[�Ǝ�����rEm\��R;Ң�t�n�vt�����Q�{E�AY���~f]�|ħ��YS�G���?`6�k��3<������"-�c����X�]%sF(���Wb��b���x�z-��ѿS՘lӜa�E��P������ļ�l��6���"�\Z�A�%�Cin�*Ͷű���/�����6"�\�-Abu�,��r� ҺZyz�e��kH�5��+���H�!X0a��S0�&~��s�Ov����h��;h>�٪�t���x��g��@K�ˍoF��/09�!�En3��:��ń�7m����~`C߷}���T4��ջ�P�����NJV_q*j���^bo:�[�~#\�fgf�^V��,�(�X�v� ���-�_g�᧡�1����:�;�S[����7�^X)��ђ��a�>S�/;�,�n�	������;�\T�m� �`�>K��5?�s,s�������K���=�>a?#�;n!/,#E�iB�Ҁ�s���������fOR,(�[�V�v��`���&}��@鸤�lgqa��(bP�FM��,J�;�Aq�|eЌ?�Q5�[��/�{�uţ�!Mg�OBЙ^���k��Oѩ�*�I�(P[e���=�ؽ\�w.�����k>��d2Sk᧺)~�Vb��RᷢK�>zlu��f>��!^^~���\�I�w�a����J؀��)��g��^
+� ���tB��^�X\Y�1 �/��az�߬�^��DsD@ Ժ錢�O��a
���w��Nia:�z[)#+�G���Y˫%&�i[��[E!	�7�3�	6戅6$��7`��.n�ہRz<sq�k�Y�QF"_�z������b��H�A-Ϧ��E`º�n�\x�V��)�?�!���;䢍K�|n��/w�2��.����A�Ӌ��f���$R���ja�7������+4��:h�`1��`FV�H}��k�"!EΎ�_L���Y�LL뺧z�@�'��(�=9���������m�dm���F�"�����k̧���J~�v?�hz�.��a�bC���r�����T'���Ǝv��Z]�M�k��gD�-����v�f��	��N�J
�OAc�����CR�)��Es=�h�A�m���.�`b��ƽ؁�&�:�g>���6��=��˗�q�V�N(¼�O�ou5"�\@T/s5*����Sdc�7�-�KpJ	�X�%hݶT�o�W3��8_gУ����4=Y�_V~�e	��2�	�z�mWdݛ�sG��D�
F�!��7�$Qi1i{U��D��6��N�"ח�M�T���y��	�k� �a�up"&3����>��B��(/���.�yp� k���}K/:t�K�nT�j���&��w`�^`&~*��yl�-\����2�>��aÓ�;��V�{�ih4V3tPaJߖK��F���<�ϰ���U�~�e�q��w��Tyd?pr=�@:~�	`T�c`�v�ar�K[µ�^VY� S�h'/��]��-~��X���1�q�!=G�ZCP?͒ە����)ch��% [Z��H ���2�'�P{�`���O;e�����} ��"�(��
�#��q����OZv^7����aq�\���01'�}�^�T��⒬M �A�d�� %��.���e�R8����N袎l9\�����N�y:�n=��M� �/z��]�o��'�?p���@7�i�,�����+��y���
u�-�\6 ����?��:;�`�:<#�5�}�����h��Թ>�\��"h����0��s��o�X�@U��/qR�(7+8`���[�s��e�|h�?�$q��C�<�A���w��|}�ɑ����q�z�̸�=�>�ȆrUB
��F�^�b�W�X6Y;��i�?!Ii̙E�K��t���*,tl��ϱ��[�g&���t��=�11I��e��=�E�e�\/����a�?�� �r*X� �~t�|AI��nV�In�@rKI�2�f���ӭ�L��i�P�ĭ=ֿ7�.�ՃQ�Ym{���G�a��[`i1[V"�Z��d�s�Jq=Ŋ�� }٬ n���!DsӴ��0�0����nºՒae�q�'���W������%����PD�Wg�CY!�(yX8��>'2߰}xj+���Nӝ����Bf���BW��FΉ����z�{*x�LJ�v7ڵ����-5F�������JrM���W�Ae��F=Y��uf�'z"Uv6B7�m�-��i��)1�r��h�)�ܿ��u�ɔJD��5R�w�B���թ2�κ�?vIZtX6�lҵy%iH��qW;%�tb?��,W��$H ��P��EUd����@X~N�~&����]iN�d�<�\#��@�A��YS�]��C���!;{��'�y��-
S�x埝�8T4ԕ��u�#��M�S�����bW5�������c�D��1�IH8_�5��{���*/,���7���G�~x5�7�m@��L������q�P^:H�o1���]�nw�W0뤱N�]oֲ��C�Y�k���;�?�j�-<�bn�[�]�VJ�7X����%��"*߰wB�H��jf��Asb*�=��e�#L� 9������[CM��B��#��a����	,��U$�)�,)7 �$GF��_������ѡ������*��fN�jA��X��	�v�������V�p��R��?��8	8�d:��?�!6hfr�(e��}�����3�EZAi������	��21-/�qɵ�֮rY����lpGy��P3k7:EX�V/��L*�����k!��l��|�����<ll㖍X�Z5l�|AE@��ȗ@�}Xh�N ��H(��>��p�m]�G���&]o d	��-��z����/s�rvI�·֫#���R�����NbN�y;ؾ1���I��4#Tys�1.�Cm`��
3�O�U::�[�����-��o~n��ٲi\�帎�RH�>qZ܀j8�h����)O=B�M �E[?�[M�K�J�H����.��w�n���*�n��ו����k��i����[Q�Eٓ��"�(���G�B=x���`�(P���qc���؄L������ ���*���W�AO���eS^L=�y޸�؂�6��5v�~�ا@�A4H���]�Wb��a����|��'����30����MC����������t3k�]>,���urx�N�v[��d�	^������#�<	@���3#��u�H�� ��~����P� ��&�c,Tb��TS��i�;[�Ա�z.�*_�l|��k?�F�I7����d�z��ѺLۢ�����r�eL�|y���?��!5��������7���q_|��&� �Z��&]s�(�mKf�n��@�� w��K�.��b#h�{V(B|eI�g����U6?�	p�(�b"`�x �:��re�(��g	�b
�7c*��XolDw��r�!D�xYXM"^͎F�0�Od~�;��+����jX�d���OY%�n�c���aT���C�y��\Ĺ)����O��2"1WGj�.�A�N+p<�V�tgh�DX���B/�1������+�L���Y ƧF��|�>��t��v��0�rc���Z�w^j����A�$���A�/1��޸� &�W5GOhp\y�����f�t�'�$G���M��&�P?��Y�'�-so�r��CЉ�`��0�������[$g�א}�����C[�B`�F����o��b�3�������+�]��~������1Bq��'\0'�U�J��D�Xڈ_���!�W �gf�Z�c<��D�wI �Um9��wX����-��Q֤k������_��-�q��d��dF��!�g�'�:Ό������@&l�J�8|�ܗE-��(��ߚ;��KI�1d�g�y� �J�^=���l�b3
�����O�d
�W�s"��1W�)k�1{M����YSsҤ�DfkE��l�'�����iοso�1�M�Y�@�+��8M�y1]6=}i��P��K�>xJ����7������ezW��^�:�o�tgюV.�L�w:'�Χ���$O�yc]�xu�P2�ɀ/u�`����~T&���B�k���z�$�Y�f��q=K��|h�/� ��������v=H�2j�g����z�]��
�M��j-�J3���}�;��,����;3ӿ!7!_�U���\��� ���5���Vq��V����-�����RN�)�r���	_/�XO��6�ݖ&�=G
�\�w�#@|�,�ϐ��U��ކ�w|�a]��Of�� FAU�e�rd�+��f���7Tǥ�q�H��,7�h)�!=��ӂsC�C��6ya�s0.�KuU���[��O��W���`jF���~����r��⫳���;�yޓx\����Nh�0�3�`�^yDE"�Ǳ\;��d�.W��c
&#���6ې�A���k4���+?��I�	T��Oe��;���-�������aċ�g�[y2�l���N8%h��F R�J�(���ө�*��f�qu��:f,[E��Qǽ���َN̸�@���u�I��k}F�w:6�~�- 3ؘ���ȃ�x�����'|-�P��.��IvC�x��͒� 쿿���E83K��UT��:U.��,qʌ9o�N�!j��iZ�R��{���/V&����T�� {4S�E��-�oۧN[�zj������"H��1��4�÷�`"Fb�R�5��]+T	��~�S�u�"���i�y7�=c��|��L�G���M �j�]�:onZ a��� �h�h��$����2�W[QG����b)�-�ه �Q�P˿I����^ߨ�/�4[9|���_t�K<w�f����S�������`��&Z��E��*��D�5��-7DuNa�J1�v�F � v�=�0���'h��A#m���/d<J�6h� �)^���������r�DK�N5_ྷ4�w�<��������w�����m����2
!ɻ���4�@��6(?S>�m�!�56���*?vΑ����AN(���Ay\\����1tY0\�;���E�r�OI��
�J�]�P\�Tql�����PL���y�]aGV��<�إ	�C#wF��t�<���U��;��O���!�Q��r)4\p7!��2 ��"9	�|\��Q�B}Ks��m��6@%�N�1�l: ��My�2OVٖ���W0��e�������]ٔ����W�R9�%��Ȱ�r��~<�<��ోY�42!Y�Di�&�H8��q��eX