XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=I�DL	��`��w|�S4�$������������ԋ� �E~àh�6V����il�y��ta�A�1ͷ� �4EKȗivX�����|�{��0h�#��U��b+S�%������LF6�Ĝ����̠Sb¬$�:*⟦=�Y��Ӿ~v ?��/~�i��[�\d���k�m�����xɷl��hMN�c��� �2� ��#�����J�Y����!�
��1�����v}�o��YuiPO�H�q>ߔ��8��������6>O�d���A������u��j�瞗�s�d}F�dC���@1ض��@��!e�_�4	˶rDl�3���h�8��A��h�]��U�RY�pe.[����R�W:}�H_�/�K��n�N���,euJ�0/@+�>��� �(T����&�e�.7#�R�c{_�mcx�������,�Ђ�������ъ��M-���x��������,u;��abV	*N�Wf4	� x�9kF?&�r�h�(��l'����s��{�/�����~�U��g��O��!�>�=
*�ş<�(��#H�
)@��v[��%4#��OИ�*�tY�
��1�$��,NK,�-�e����ǒ2Vl�ki�����N�(Gp;S��ESf@70��n�"�O�]���L�PŬn�Y�I�3����0����?��[l�[@�G�H�] νOs���J�bK���~���g��b�R��bf���q�ZD����A �
Ui���X�K8y��XlxVHYEB     400     180R��(�fdrܝ9�2���(\#}�� 77�q�ư/�9!m'�css%oX��K��_��˧Hn��}�jB�xiF�!�i+qc�¬����H �~뎠ş���w�~��#{
`2l�p�!�:�W����n���ƶ�/�*�fb���'�ˆ�-�5v�.3uy@iSn"]��,�qȵ\�`���Y���?�딽$�/#��CN��vZ��O2��	8��� ��Nl�|cL}2�2&_���[N�nD"=�lp�I5�U��Q�$w��/_��hr^��1sO��^���+_fB�h�c��E�M1�Z�fe�������"��x�u���xH�  ��h6D�z�!�������YJ�&}�S	B�9�P.�;����<XlxVHYEB     400     160 �8�i����VG�rm?�t}�F1Q@s�4(ڢ��l�J��E��|��f�l��h�ktX%T�9|���Y��w�KV�oRW�/�Vt�iֽR���_�䬐Ѡ �徙�^�.8KZ��@!��b�^��<ԟkf�mbyE$*�D1�Y0D&'�e�E� J�VR�K-�����Ʃ��ԧ�w�yMb�A-]]CK1�זL)�(s)=ć��H���p~fPR�K8~40xu��!.lj��I�Lp:�ۃ�΃"w��H*�!����v9����/�O�L��<��V��1�T�����������9�)����2�RV*sg��f(�[�ָ��釸⺮��!N��XlxVHYEB     400      a0�R�5��Ѱ�/��[D�B�T��cYy���浂+;�"�r��&{�ULkO��:����lfD�6\Ŭ%�p~@��Wz�Ƒbd�i柆I�E	�3�+*���������n_CП�>(8��6T�3֥�X���}]��3�&���g�R-j��A2�XlxVHYEB     400     120!N�)�K�M�Y��ـ}پ��	��Vة+D.���\�5E��q����C33x����>��b��L�N/�
&�4�1�uY޻1�-��3"������Jnn`�>�z��cEY/�������k�t_~�)�'^���Q 	�mo�rW��P�c�e��������dZ�c=I���xf̮f��J�� �U�_	J�	(���HKB�'�5Tר�@�~u��ɠWN��w�E
@9��6{�
E��,Q7���ѾI��Y�QJ��y)�x�({�W�yHتG.�w�,tXlxVHYEB     400     110R���T��(o��O��6c��h~'6��8G�E������^�j=��
@�^����oHSX0��R�������͸מ�\m-�;��_���[�IF��o>EI�wȓ����Q
�7gq��pW�ޠ���V��P�j�Au�i`��B&��v�Y=�J���fn��˚�d�K�w��e��p.��AXs����;�j$Tp(&���m^#����C�~��=���pք-�%�����cm�L]��k� ��El>���j:�n�u�XlxVHYEB     400     130�#t�w��oc�g�Vt�o I�ߊ�8�����<����%AZ�ِ�m;v��	��j��#�e�;�+���"���G
��Ub*S�U�$3Z�#��n�o�G��؞��Ol��+`d�=�s3xƄ�|}�������뇗> �����_v��ܳ��+�a�"~Q���Qy��	�-Q�̻�k&J˯�..^�a��QdV��#�a��OiTouP������e���0@��Ư����y� X��nvx�z>t\jt��
v�z�&?���Q�݅����h�����Q6XlxVHYEB     400     130-���],�P�d�DE5��hXE~�Xu0	�iL�t��	���I�.�1�o��vq�,�Q]w����J6{���)pm�5��?�������xԜNW�����O࿿~���
��S�,�M�j����UAq�?Yg��z�����| C:5%���!F�j QH��
��sm����'��kT�޴��b���xS�jY�q⟼c�nuU
HlAV�zUR8h�:��������/��
�%�<�<�re�!Jc�L�}�R��A�v�h^ƚ��^r�z�.ƛ�wu7�E�����r���dJ�A}�`�o���XlxVHYEB     400     120���Ǭ［��R4l1@�+��윆�+0.�/����, dL� ����4׳�����.�zPr��a_�n�tc���fE{5���n[O�b�՗Y��p5�ݡs�4�s����j<�������b[6x��fK�2g�l��&ބi��]$#Q�����a8r�|�~������C��\K��dD��3���\��R}� �j��_�M
Lx�xմ��:s�RD	��G��1{�R��g\V2]�4�ALĮ0�B�b��B�&��U�M�('�Wv�5�<�J��S1Q&��XlxVHYEB     3a6     180�HU����H\Z�I�1h]����)��SD�2�r�J%�@*�gĚXJp3�V�i�M�b��4�Ql:#�,JL����rO���+K�>�=|c��N��ܮz[fE 𒯊�����0�-�1m]�������n����À��DηZ'���)nʴ&��i��x�ڢP��?.�����]���+c�܉!�™;��[շ%���uy�ҙ\N���&�#}�F}^჊��'i�z�T���}��t�ؿ�xM�7F} [D
��(T��oQe;���VY�e�;�խt�("%��'Ύ{�E!���4yOI@̀��+	rh���#������s?X�ҭ*r� O�j�Wv�_Ҳ��U�VX�˹��<d���s 