��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����i��9���KQ��n���02��ę8�&pB�q���wShCH���u�Xj|����1�N�vc$�v��Q1�4�����D- ҽt䍤4����-��-.����tT�DHׇ��@��䉋�r�`+tT"[:"��4z������F!��� ���tF��	zi���V��	���r3��E�D��G?<�+��`�O���s���~.��
��zI����5{��'[�@;�Y]���ifh�9�s1��(rJ�?|(I�|
�j�A�8s��w�+�ue$��4ށ�M�0��(�;����T���9W�",�P޹0���Yq�	w�}�QI�Ұy�J��躧��#Sj�z(���2���śI�B�g0Cn�9��oQH ��y�v��˰ƽ��y��Լ�&�T	�7��,�gx�X	'��*�=@�1� mehX^�r�߻�a��;��9�����e��Y''��G���/7μe�ji���;�)�L�'v�2��a,G����,�����  #�ο��i�]��ﺁ�q�k6 �"�YX񪽮*�!9y��Y��#r�Ƴ���K�q��e*�I���������=�"����R��˒C��b^׆�?�W�o��g
�N���>�AWg�%IO< E<N��KM�$$
�ď�/�I)��w�# ����A;񐻈��T���2,�N+8;
�fާ0�[@�<ϵW���>L|����ǌb�����D�A����Y�T���kL������e3��7z��ji.������pc�r�ܠ���Dh>�6�@ި׫8��i�Q�R
/��i��ExD�&7��z�����9jTH�]H���ja	���KS0��Y����nd�T+���h���Il.-��-Q��wH�a� _W�f�5�"�թ��^���צW�B�0�4?� X����T��֑�Y1`Uɵ��0*�ޏ�T�w�8���������'�����N���qi�vQ�~%�.u-[:Jnb]�2'���ݦ�xM%?�ȡ��%��~�����+$�|�F��͸����Zf�c��C16A�jw���kH�c�O�z�6S���Z�4�Kߕ��F_~���q�<�M�sq%Ja���G��E%*1P]�V�g��)�����䥙��Q]�z�Ɛ�=�.ă���<_6򉅳?3�e�UH�'j�4|r���iƹ��HH��"	��A�qL�U��v��R�3�Q�oc���ZB���]����&��s*]��h��9�gm�?�2�(��|�$=�~�jl�r�h���).=/�vv�RX�,� ҥ���s�V�w4�����_�b4��:F��,&�mM U%��kH�)}�H�fx��z�Ǻ��6���Q4T�LKz�LR|T� `q'd�� �
�\����ga���\F%�3�=���w��{rU}~���z��(!#���X(�m��
]�T�k�����w�ZȘ��(ch{%�I_��w	9ڎd�N�6sv�cᱹ�_�y��H�KQ
�
�ɑ�W�p����}�rnPu�g� ؓ�<]�i?�}������ߪ���=٘��;�����s����x��Q�݆0��!p0�2�m��WP]�2Me��\�O
��lK�^o����������-��e��A��1�1�֠h���w㚒s��-�&�[{��](�-_�8������q��x�w]@����ܓH�c�����1�4��*�=A�������\h���N'��H4���9b��;E}C1{9--Y�:�.�F�)�*���03�(l�k��JY�yL?�$Xi��۫��_�`�,�댦l@Q]Z����ٶC�g�<B4xdj+����q�PH�i����t��ݣ�BLtsf��LƜ(>I���(�I�V�YK�(%{B��ঘ��֑6���\9��B1�e�U�!]��b�C_ߞ�j���ư���M֗_(z��"P�>���0����2�2𩹊�sV��VՂ�ϒ H�I�&��DFkyP�f��v���M6��%�Zީ~�Kj�c�o�p�,Bg�̹˃��/C����/�v]�3E���d�{C/���ay��A�ߍJB���t
p����fe��|CP��!�����2!�ѻ�i^���b���<|%�*�d�e�x�pi%��W��Sw� t>�_تNt�!�;�N�Ah�������rxgˎ��ڱqb�`y�~���^��XR2,+�;�VY6��OT�ӨE�B��tH�e�2��*������ C ��f������ C�7]s���m[�1T�r�&��>�Zl�#:)��I�>{�Y�N� �%;���ET:�w#&�}����Q6��z��jN�URt�f]4�$2X�����MM��R�nQo���/�-x��X�y��X�7'���zWpɹBK�osٻ��DL�"E��<����<�&�G{���ƨ�R��Z3Op�3(�7���2�羌�76g�2��'`ѣ�����o^4�zJM`�P�x�1��3�|6欁�ZO���ᛡ?U�p,U��]	 �U�4�8��;�|�)�]��ff�U2�g�)�c0r�f2��ɜ���M,�Z</�\=].V���A�)�$�2b�%�6���-�j�Ca�R7m��^A4n�o2x�,�!G��SzE6��ĭ[J�T>$)�L��rY�������6�;!1\-:,�q@�*e��3KH!�6�����?��8 "6e�����.	���t�2"ʠ�b�����-��K�C;Bx�Qs��6)�qd:i )�S�{�ŔW<��r��NZ\8=p�9PB�(��mtn�ࡋ)���	@��Q��H���;y����͵@���>��ˇ4"�#Ի{VMíePWxuu�/.�j����D�e<��Z��Uz%��ߵ�ֱG�_Z�zVAK5�\�	��v��^[�R���d�7�.�������dl5�H�-|gr qha��_A�~|�����b�,����ύ�\��98���� 6�P��.n3!�!�V׊�joggI�	bI�N:�ŀ�-7�ݥ?���ywSD�K2����q��'�����P�`�&;��JM�v���F@M3zm��q=����%���,<��
#��z�X�����*�ϵ���|Y�q]̀�#��կ�(-|��|�U7A�ULȲ��~3Ube(t��z�	_!��-�pα�w{QT,j��P� �
8�v/�������D~O8�Wj�� ��J>�K�ǯdydA���M�0u�u��̑5��7�/��?3��q��ث�\hϐ��'��Ҍ�rS:�8����( 1�z>�=�&Oj�y�9�:�����7���o���4�Q�uH�y`Zk��H;�HV.bhU���7Um6��7��m%��j(;|�h
�����#,�\4;.�/怾<��%��5
� jbGΆO'ti�C��X5V+n7�QC-�o��A.d�� �b?��"ɺ�j1�7�G{O-�Wُ~�h�6�6[B����ߏmUR������0��W���t:uijaYy\�;�zͪ3��\b�<o��J�n�L�
��s�
=py��*�63!��q��՟�/^0#��m!��>��D���s�v ������\��.�y^;r�np���9ɄPqkυ}�%jfa|�X��g��Ko%I�x@�j�ŏ��h)m�4���&/Vj�9Ҭ�dr�8��6�c�ֶ�!�΀04����ɂJ��٫̹Ԯ�ma�U���b�J�����HǏ�P�}���Y`P��}�~��sf��J.���*=[ k�RColo�q�H\��P.�f�VV�얭�9�jI=I)��BQ�[�otf�S��\Tܢ��A�ߜ��P-#�� �yZ/�5$92�t������e���@/�u�Q[�$����,�g���,�OT+d}�J���k����{�.�?���8��+��^S��rG���1׆�۬ j�����J�z"∁x���h�[$,�8���G�����ՊJ��M�a�TFc</7g�c��yh��ha�8��t޺g�z��ٟ�b���ppSfz�.��6�wIKn��hZ�#�����@��Q�'d;�K�07��ժ'U�y8$�ĐNP1`2)a$ [0�
��[j��m�>���z����L���x~y�ԕf�݉iዷO��5c�*���;[����4��v|,P���,���ID��V�l����WTZ�Ŝ����ƞ�\ퟳ��1f�u|�h�  `��ig�(fgs�m��f@�%�(��y�MP�rb8�|WeHfb���_S��&Wv�u�P^V� �i�=/�!V!�Z�V�����]�SƌF2ds�$i<��~�#����َ�߱-)��9�,e/�qNAm������D�z3
<�f8_�ɓS�=�����E;��<_� �cQ(gbFzӲ�e���<"�."x�	��'
֕%8����\Zw`2r�wu(nN�5���r���O
e�wݥL7���ٵE�zB�J�#jX��̘ɀ	�U	Z١��9<�i�A�2�婠{~�I?�rFu_xȃ��*ܭC7���*�b�����jh�1�x�*$��J`E��ى�U䒖Z�U�Fa�����Qً���� �l~��,��#���"maFI�vO��G�6�o��&�j���Gfn�rs4���9.��3���A"�$����Ā'��]�@�jw�B�옎����q��0L�+�nqID��Ӗ��0������X"�D�I�a�/Ib��c��yyt�'[� ��r�A�M1]^��5k�Xa�嬺��>@{�N
>�z䇻 x{{�ԓ04n�-��&���f|UQ���ٶc1zkK�o�>�k$�X��g�)��G[8{i���\/�/i���A��]ZW}�_h��Z��I�oFa��SIG>�����`KD���cwH���J�b�݌��5f�]�����#R��%�hͦ�=��B��H�屠r���Q��|<�%��/w����ee�4w~�^�npP3"3���(1��M"��T�zU�4%iԱ�Mh]5B���~?����z3��F9��/���Ϛq�Q�y{#l�ݧׯC�}��8�`���}�wC��t"n�G~�g��K*	c���(��L׏�a�ԏ�GA�9�[^�,�����^�����:�֚����e����]�}R�l��q��TϠ�[�1���S��1�/�?
g�>�NhHc?���yRot4���T�6`�"'j��c!�_ �V� �LƆ.���/�6��ovn`��J��tQ���2t�UH���P��eYg���e��}�E �!ć�P��w���X���*c}ƪQ��F\]�.@e��w+mVc��7��}Qu܎�9O��z-K�=n]����ў�'c�+�;Vbj�����3 X,�O�c�����V���$7������H�������M�^+r}���sA�w�VA����e���U��<4��$ϭ�I�CV��Ax~�v���&ښ`xx��8u�8`�߲��X���D�k�J���#���X���?���kυ�_*�gs�j�Գ���ǭ��l�e�S�C>��\��L��n��'��@s�G$U�z�0F���sԘ�
��x��M�1c}݁����)�*n�q���ap�;6E*�`)�$[
��CCi�)�����M�E�`�P�t�|M�L��m�K��p̪��jlƪ��nqoMw="��༥�2��+%_���I��9k�ӝ�%rT���7H�K�Í���&������1�7L��R�:����w����F
����Dr��[�}�(DH؟$ =���o����9���h����wn9K��e-;�4�#����y���5Ҥ��lQpo5Qy`
�ǰ	��<�d����Px�@�(�!*��������ĥ8��t�G�7E��U� �Q_���5�F������o̲��rCX�6�1�yl��QV�����=㙛X� �'UA�& �9����$a��
� ,_��[��L��ƌxI`�(���ߝ�>��x��a_x�na4B{P����'BZ�P�R�9���u�8�����>!y5�T>�<�jM���1,#qC�
!��m���E�r��.��`���t�0�/�>����h�/��x�O
�b{~��a����