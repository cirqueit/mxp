XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����4�3;zb5Q����'�=\��&����׷419NZ�Cz�@W�97��l���E�t �Ǘa�P��ulh�G6���f�$���0K���ȴJ���2-�x2����l?Ǿ
F�Ѭ�����Q�����]��h7)��M�Xy*$�>����N���Z�԰���#kEz�}lX�3��i�� 's����q�Ja�[t2d(�ˠ�iev�دTc$�$����&IpH��U�
��>�d�zh��A3�I�ĕ��^��x���^x��^E{�K��zH��o�O~I����{荵���?^u��j�R+�}K\R�G��B�``24{Ҟ��tFn��R�������H1ʦL�(�o]K,����QJe�e_$��ԓ�X�6���l)����&k��� �(G��{�͇��s���J�i���5�:���X퍲�]����\S�7���7��]1�sQ�q�8L���wI�_^WI�]�1�=�Ԑ��C�P]��|6��*�&���H���u�e2�r__�E� ���0��'ty<*��Q!�%y��V�~sG���Ɠ֣Q�2\{�<طĩ�.d���奿�b-��)��jU����`�9e�+���M�����顃$t�ھ6IL7�-1��Ȋsc���x���l%���+b��]�ฤ+�0�no��N)���'F��;{����`%=f�&���rv=r�y�&;7��"{Vp�<Gj<�V��5g%����.��쏍�<��"���XlxVHYEB     400     150G<\B�8\��/F���Uܣ"fXW_/�S��9�Z!�ru�*����X�E�|��U�@��h���*)T�zCtA�t�U3�_�^W��V_��7�����ha#q��=x��z�u����m���m��H�XX� 6n���)w��.�p��|�(��9gJQ�wx${��jv�	��.�z[��vB��ջ,���PDt����|���#r\��+O���,?��e��:��QNrf6��*=P����t�d��;$S**.:f��#C 9L�H�=\��28&�൘u-�E_� ���_Q�!��:��3~4j���������l�D{�З��0�:ĩ�a\N�����XlxVHYEB     400     170A>pW���}rK;(f��S��G9�1
�`��у&Z��͊�$,R<�v��>'�����G� |$�xlH�)40��+���=�Wx�G~�;�O�� �Y>�6���;v.|n�Y8?��#�pz� +]�Җ�G��s� ��7�6�z�yӫaI 0z�JyxV�?�;�e�oB��^Q���G�MD*wI�O�	�5���\Ko����.�<�f�5F �c�hf����M��R��T)��Ȍ�e:���R���K)�u��p~�j<�WW� �ӥ!�{��U���#M��q�܋��ێl�9�K�`��:JQZSm7ɷS�z�i�~��hE���H@��S^���:m�Rk2���WW��N,�7C���x�jT�J1XlxVHYEB     400     130ͷ�;5�InH�Z���JS}���l�&ʁx�o���(Е�@��J� �L�g�rg<�$���Z���%����Z^�Y W�%R+]Dؐ������D�Rq��\bH��hE�ٸ�6��Ul�	X�1���l՚ɣ�>*�`�G�J�J��!�I�l{��bi�n�������W^���KHg���fӓ���`�|G4?��kh�g��w�~lE'�h��_~��v%W$1 ap��W(�}S(�@Py��"��OT�Eu8|g�2��
�����lՔ<���/(g0{#ߋuQy�Q,��T*M��ɍ�*XlxVHYEB     400     1005M����b]N/����j�,�h�Y�JpM]�b�v�Kc���������KC��]��<���$���РM2��Ȗ��R��bf�j��n�½��jG����^M�6��x���dǨ��f��*a��k�כ�|�L�k�3���c����EJ��UD.JI�����F�6N�� �E���?�C6`]�&9�Pb�u�TL������}xc �9^���l$g{��l��d�ޘ��@��E@ߴ���ӭ���XT�XlxVHYEB     400      e0�<t���%�vG�n�<��_ۇ���;�RdVB�'��Hb����X�����!Δb�#���b��O���G��~3q��Euj�BȬ�@��X�b*�+�����zdz�bd��%��}�A���̒ޞXʦ0"s&�$e)���Щ�y%�P��y���� ���g��RH���k�fh��/�ܬ/C��VQ�&|�2psWe;a�73����S^)�*�XlxVHYEB     400      d0V|�:W�.m\��d�[_@T�J��}��}8�}���h�!�i�׮j_UYf�,�4���������K�A���ڿZӢ��ꨋQ��t3yrN�)U�{�CB�`�H��|��zP�s����5bѡC�f5[Tk�?7�hI�z��ZE��NQ;�:k���_e�1�,0�}H�"ee
����㹺��K
��&Kר(�.�1���XlxVHYEB     400     120�W2�-~C*%<D<���⯗i��U��N.|���
�������ֶKQ�x���+h~܁$\�K��'�9��-N���� �x5Ö,ꫬ��Z��Q�R
C�/ro\�Rl$R�R����*��'!��/��dzp~�KS��_B�3�ũ�1�1���
_K�7Z�l�|��������@Joc�g	�O�*2�M��5�Z҅�Eӧ�oR�C
��#�_�%�p��a�(K���'.�/;��e*�g�?���}�u2eg���*�0&2{�q�Y�R�1��XlxVHYEB     400     180�����c� �9!6�0�S�@��o#�rCвC��>um�҉����x�V�vU��`�]���Cs���˄�w��~W]���*⦃�p"�09�)�N��Q�s�Ol��;�6�����������jB�7F<D9��n���ß��ˋYF�T��~@kiW����:���]SN��Kj۞�ZoW����8�a%�<Y�xz�AC^����������c�����X��yTe#I] ���X]9Y��[A⻸Y���m�B��]Ã�E}��ɽ��Nօ[���`�1��0kuי��-�af��л$�!%_X�S�&�
~�4�}.:�	�z�����pw��^����Þ�E�*LǺ,�^�k>C���3XlxVHYEB     400     140���r��t�|�
4�`�=����נA^�1Ę;��}ݦ��FjL��41(�u�ۙO<�r���H��)Rs�/n���f�����\:�m��'l[�)���v�?�0����f)qni?�pDG�XsǗr�Y.�b��^*�yj���r��T5D1�zj��ȃ��<;���^��M �äN��>���<8T�c�8\iCK.�8�H��a�������BCk�h����4�ToҜ%X9�b�צN歰���Ι����/H֔^���`�	[PКe�f��3]���H/�9�(���p�&�1�5��*��XlxVHYEB     400     170�N���/�|,1�V`Ga�VL�}B�2�E�A]^q?�c�b0ו;��"�d����L[�� ��y������sf��=d�ݼ>�5�q��L��*Ȃ���@ �l��d�$���Wm.(�K�?Z�+���"����D-�����"MwC������r]X�������d"�0�n#���`�meM����3Oݲ4��$@G(������E=^����KRR�:Si>}�!���nT��w y>=��:�*`2��*yH@��+~�L!J� �v��t�]�b$�M�Qe����kD���7��G�cϊB6�'���2J>�y������o����t�d3�g瞡W}��Am�
XlxVHYEB     170      d0�����ް��P�%���QX��t�MU�s��5|�� �>\K�X#����0O1->�r�;hp��T�TCqQ���V�aS�P�sG�,r�{�R�&�E5�tB�-��T{gYh��~V讙JHF���Q�{c[1ujm��	��E]���<�C��h>���lj�L3�mM4���`��BY���D�_���L3r<1c��