XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���C��R�lX�6V���G��^������V��*�?Z4�y�>�f,��Q޼�,+rм�N�C��Q���n%�٠ڋ�K�2���X7�3+%3��&Z&R�!��_v[bJ�F��Y=;g��^���%"P�*��'n[b꤅�u����(�+���K���]����}�y,��i�UL�r#Q�|a� ƥ����qݏ�B�l��QvB�j�c�D��l��8C<��^��mxvd�f�5nx.©u��Fd+���Ja؋����QC�K�D�Kb�g�)	3����X�9�D�ZEH��?��F������c@I3�F|���*�w��5���:�%����_��*z�|�|���`7����g����S3[��1w������R��4�Y��C\�
I�B���	E��D�<����L����V[�m�Ѫ��k��+uu1�;*����޴�7�{������Z�V�G��<м�)2����kj�?zc���L����ۤ�E�\hĭ��"1?¶h90\f�/���G�lqx߆�C���p��"U�-0��n�F>��`ŕ�[zʝ-���Ÿ=�<0لV #�<�W���ǋX�+*�/�"�PT�,L�����ٰ��]�@�asK��&�U�@��	���'!�k�6Z2�%����*9��Z��n�P/i����d����	��N�z�SY�����=�Mh�aƴp�&W��O$#:rc�e���Ԅ�e�u��a�v~O��?Z��ұ0
��=켁XlxVHYEB     400     190?��"n0��'f�\���H\b��n��Eb�*I]��ӟ��f��
��M7$�Șg�����_���Ҁ4�/�����_
+`��!�f���͊�jI[�*w0F}6��9����})�\lL��Y`A,�.5��=F^/���ex��o������J�cN�K@���q��-�=�������0_'S	����9Z�+�������;d2	b{������}��۲UY�ټ(H���mz��h��q�4��XTY����am�yz�f4��8�2�y|Yz=f�V��F�̚9�2ڄ�,0��x�Y�ǱW9��.˹vψ~��
�-���(Z�2	]qs/�|n�k�����
H{�N 7�����}';�u 0C����ݐ�2��˽%��	=�z7XlxVHYEB     400     170�M*-y댳�EJK����pԌ&�f������[�.ӓ$i��L�[3��1��5J�����!��F���-����6�km�-�#��WU�f��� �	�G+z�T �6(fT�C��E��Q�F}���2Š�)�dCX�X�H�o��ǚ	��4���@�x��ґ�+a�����Ѻɜ�M�ec^$�q�f�����2�K0Ӥ)���U\��T��@T���#���&؃�2岜p��"�b���q���(�s�`��
�ULI���ъp8Vb���Mn9�����W+����/g��)����{��Z>��f%��{ų��{��+�(0C�9��9�@/��*�����f4�-�E�t|�PXlxVHYEB     400     180S�v[xe��Pr>�z���@&?������9�&3i栫>�R:^*`�.�Y��⮉~oGZv�ˉ �TA�O��03�BheL���������'�|�5"�aܚ�-�W*�vt�:ӊ�f�:�.i���qk�Ǚ��0�hl��m���ͤr���1�L��Q z���� q�H�m�W�fh]��gۆw�Ʉc=Õ�318��_원f�הxA+AD On�D��e�H
p�a�ŝ_�Y��aH���/��t��(}�lAv�¼��[�k��qN�C	D�%$GL���Ȍ�I�Gχ�HݸA~.P��J�WO��V�`q��z�W�����7�cަ�av~!	�<��6�������$�m�	f�C���o�����C��~շ0��u�@XlxVHYEB     400     150%~�N$���GA�"���B2�_t�,J{�1�z�`���=���8P��D���AQ�熋%b��}0�̮���eD�;�VvȆL0�~}��g�K]4_C;�����W	�H`�&5���[���"*�ڬ6����~B�}Wtx����?��bQ~"�1G�Е�� � ۗ�� �C�˗%�M��՚Kc"K���5#�PQ�h�lA�Lg:@�7��YG��;����cN�ٗ����[�ⲡA�P��i���xb���g�̓�MWܺ�@�įo��LÌ�%S�!�����w�a�6����`�va�����\i�h"}��E����XlxVHYEB     400     170��\�C^���T+Ō	�
��*��:5/�y@������*��Eh�b�u眯ek��iO�
�L_5�]��VZ�J�������
��쮣m4~Yd[�ܱ8�IV��d��U�U�O�5+��1��0�3/��+-�������c���Y��Hz�W�y��Ɵx�����Y�D�wN<ӥ%%C�h'�������jGQs��?��`x�ͥ���u{:=�e��������d�Ԯ�g�u��L�5s���-��#�A�Ҭ�3�V�T�c�,���c�5՞Μ�A{��˷a,�^�����Vn\��`�g���~�?����n�Z�t�X�/hF��Z���KkB��y{7���-h��y�7&�XlxVHYEB     400     1b0�Aŗ~�ɑ��3�? |�v���p��/�����	��b��Ӧ���H��Qf��3��O(Z�F��06B��x|�C���>uD�ߏx&�Д� !��	Q��]�����<@*��:Q�ѓF&2���f���u>B��S~_7�����u�}���G�K�Ӛ�}^T�%1qO�.�efQV?U�q�|ҥ�z�KΟ���'�C='0��om�xxk@�ϲŨ���o��ڝ�o����c
أ�\T`�9F�m������i)1lSEn�,��K;�A��LP�=��Zf[���cPǒ�ZvqU�P�h�5��2jƽg=�g�l7A���y,��Ȩr��t��v͡vÉ_6R�c�<��9e��	��Ź��DJ�&y�-)/X�B������-�S���B�dd�#cn% ���,�`��5����XlxVHYEB      e0      a0�?������on?��oRڨt�JZw�v���-�l��9�t_$�H��R�1��Z�K����oit� ���;���$T������ɛ�^��n�(L�ZTy�g���P��gX>1p�#�M�RQ��yN��<�g�aZ��"�jS�M鎪�a������ 