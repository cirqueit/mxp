`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
5lXszTI14XBynzbIZW3H4xUHCG2ACYeFl8Pf/bvPVvnPRfnGykh/BMCuFp1lMiu0lNENQbOdg1Pg
FnmLKZvsdRKFOJcCd89JJHSZaqDDqG8M+dMcDSBsR7yvq0fksNQmIm+SW6Yr6asiyU99uatEvtNu
v5gnGnZSzxGBwQ4rP4d0qQhkcPHntfoB3SIUfYoPWk9BFlI0XlX6Fle4eBOsddhI+QeKD7B/rgrh
V2SuOpdSRvogaazvOtJOwsY/6rQhtFJiRJGKoPo6XjumEgcPj6xSqjq02aVXQuptZbN6ouioeVet
IVix5nvm+AqSLKVTMJNwgh2FHRmwOTQKO/jRm56iRhydLxDne3iVtvb4Nag27jCiVi0YNFcbbHXs
hz0pBqB0Rjox5Zi1Jv4gTQgBClTsSXNgnl9+u9ZWzD1iwii0hT8i/0u0EJL3N3+keSruH8cIUw63
XUm0QtAzfMijFz6c+h7CzWNRRnNyMLDvTiiZ93yeVPIbs2g54fPSP5YshcUgmjgh56THOZGQpYzi
P1p7ojgBMUo+kjc6jxEGRG1X4Qt+utKijloLqS026OY4bBrTruGxkKEYySDs+R/HCMw5aZ//083t
+n0DvJQb5pHFhQF5jyul63Um6N6h1lu2T1OsVLAlkVYX1jKU8B4ShYRbBz26BaBDXhnAoT4+AQR7
HW7BncTMJz+NQNjRhr9ZWxvCsNRx997pjqYxPi0x3rSUoR82mJgUQqIOzdu6VHBblgljpwLmJYhU
LRycveG+NfW5ne2DdCP3Yjy2a2+KlMPZ3RWA3715dYhT//2WmGpJNuGfPwMkBW7i2ruBJNOXaSdq
UQlOnb0BISemuj0eoXXkrabJjnUPQpM0YtV6jyQDEZSPIex7Xnp61+IrjqCCgcsQBkBLzh0zJwx0
Ywf5KvVYDSGBt4zbcuiMKSyqH8ttI8Z/KHiXVXgICy4wMZ95cLtIKFbnOcwNr7nhujcNuuhcI8S6
S6WdloGLTUC4VOyg2aa2y1A76OmvlPm47WGDsuH/C2Oax40NCFAX5AZ03Lbr/fCafmErG+FTc+di
RyuLM86xtGly6R2d+o5UpYooEB1ef6DSK1Cb9/EoW6aicB1akbuJkRv/iMGTve49EIqnx40tDCoq
eyuYOSi9esIP3+J1qvwxqf/mBuNfKG6SaFt7oiAeFYchAaRsEsGxu8bZaSubmpRuhmG/guBySnTA
PrPXJzSUNlRnFNTP8aaXDg==
`protect end_protected
