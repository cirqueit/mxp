��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����¦`���IU�e�Yb���PJ�����N��V�A}"1!�w�)�Yxx��?f�2YEV�V+��I�K'+�lOB�xWѷ��/�'E���#~~��F%���jlO[�m���׿��JM�(�o�.6�|{	t�&��T"'@����v^��B/�6��W�Z!M��\s�az!�6����g�������m	���?!|3��nc�W�
���R_��`A��tb3��y��3�1]0}�F�G�ғq>E�����c���D�j��ش԰h�*=����6t�Fz�8�G��"_J�=����ӨM��QV�Om�����[�՟���B�>~�n2ԕf��F����ȱ���$�A�nw���6g;]���10-*�L&��[N���o���|K�+ݡ���-2��z�=5W������ܳ)q	{�靋�PQ�5-b�*r�G��U�3�����T�,�^�pϫ1Ά�D؉mH4W�i�� p��@�5$|��<�*��Ҧ�<A۹!H[]%4	��?s_z�S
�!�H��pw}���0�m_>�P����i!��
�Y�{n)3�T������~�1���R����XC�0�3y�ѓ�.B� "P���7�dϷNK'-�8 jO���$��S�>j"ǦZս��嘉��/�V	��?I ����N��Q�)Aݸ@/F����d�q��-�cǘ�Q��!W>�I=���EL�f��b��40�|=~�4�'l�!�KT�ʾ3UzC�mK�	��Q���&�Nƒ>D�v��|a�P2���~�o�;�:#V�����<*L�$�$E�ΰ����6�����~w1���E&zi�tڌ��4���y����N�$�J��9���BA�Ġ�/Q�F�̅]e�"w7���_o:��p�L���#��zi*�Ș�Q iF��k����*tx>��><P.�ܰD^�;:н>=0����=�#lV?g�=��h�WG/��>�5��.�	��L���t�By�3�қji��'��w�i��A�*Q�N��|E2�ߵv������ij֫����ʔ������>�!��n��H��Y���A�8Uf���c��A��uG��6,�s��]�Ǟ��yK�v9�G^i�~�nn��6w�V��a&��y�T�MB>�3��)�j���+�m~1�9\A0�C����j�r
}J��ΈEk���x��wt� �+=����'y��k���k�e������O���ݥ���J�ψ�sk�x�,%
e^Ӈ����a������N+���� W�AS���H�d ���-��T�j��*��N8�>�ۻB�!�nC L>�j��jO����b��x�<X��\S�G$HŽ-l)Q��t�jۊU�,T�L�x$�������/�	%X��/�W���9e8ʕ���Ӕvt�#�,Da�=r��s�`r�g�t6B
�O��oK�Ғ�������!R(��Ⱦv�Sn����=S0˵����'��5����
𞏜C�P���hEY8a��|gt�w�����L9��i31uHcУ,�@[�H��������5�%��-�%��}՞[�HRp���g�ɑ߼�T��v;,�a��yz��sBGeF�b���y�ja��ӆ�0�d�{����w�1�/�c@^��!ۛ���I5Os��L��e���v$8O�hK� �f���df���?*wjS9��46m ��ah�i}���bv�E�@�\�3�'�3Ÿ���b< ��ƣ�ߞs87���٩,s\h`Ф~�i��IϞT%F��!���'"G�r��������c�nxCA)�CG(�Y���?�\�����p��*�J������qѨ1R�vSD_���K��R買�[�U�;!�{�P̗D�YH֌��(����d��@ky���8x�lrh�.�Ňb<B%��8���;��<ڦ�)D�A֞�������07�t1m,����H�p�H�g���2��5t����'�IZ������r�1F�\��Ck�5/)����e�a9�����Њ������2��ƈ�5L���K4UQ
&�bǛwր)�yt{2,���m�QZqrk$�Qb�tJxˬ�m@+X�[/JQ$fz\���[q��ڌe�<P`t�bnu ���C�e�p�ڑHn[��[4���ͯ��&�}�P�=���p��'�c��IN���\-r�	��eF�k!�7���� �K�}��R�������Li/u&��^V��pi
��PK|��O�lk'V.૩��h�$�i�s��&Z_ixW��}{3�&Ӭ���K\�%�����	�növ�[(����I��9"ے�8��$�v��v�_!>>�"2��P�3e�#�-"�^u�±G���8Xu��
��AB9���<��� "=�V��I�l�ԑ����d�*2*c!�8Z�c,�lUbM�����/m{�"�E8��������\c��4 {��W�s{v�B\%�������·T��T=m}e�`XÌvݐ����r������X�
-���e f����̗�yX��Y��u��!���=&��@U"|�K��r5�ǃ�슣��� Di���M��d�i>{�ݸ�n��p�ڬH�w��>`oU�jH���o��	�;Cx�S�,;˴���t�SEx�e72��1N�5�����'2��L�YF�� 43�'�M|��ʈJ�e�mil��jc�����ql3�j�Mb#����a����~bs�E�Q5�SY%��1P���3-���?Mڭy�a��!Oa�{Ӽ���u3Q�?��N���Et�oZ-ap9�]���zj��`�*�
}���#���8�빌�l�b�e�2N�!��pHw�	7�3���J�a$���Ӕ�$lB5��'��⨻���A+ӬM.H�~Z{)��j�L#=�"��~���X��0����t��I����*@W/�sC�=�[��%���)v�XT?�Da���'�	Jf��j%~e� λ���._F��2�@�Q�h���@�5O������}��*�8s:õ���G1�
�N�G�Ħ���ʓ��Y�Hz�&�k�A���f��htWMd���D4��Czm0�9�W�Wp��Ń�F�ڏ���C��g8>P�+�n�aoѝGs4���m�׸�KBt�	�l���$f��N�����^�� �+ۃH�'�$�,Uq�m�4�Ks�A˨����=*�UZCoCl�����XJ`�[G�M8��/[�S��nL�E�_[FG,�f_⋈�����`,�"�#��d�l���
 eI���.�LOj��4�;�Q��D�Ļ��6�F��ʍE�ѭF�ȫ�8�ۻ{U#�����˾�c� IƧ2����uڭC�h�����z���}�h�Q7A��]���&�/�
l�ڣ��ٗQ�9U3�=�.)s� 梊R�Ka?(�k�Ay$�F�V`Ԟ:�\�@A�<��K�}"�Ǚ+y�.�kQ"��\��� C8 �!�E�~�8F�,+���ZС��5�I5��M�]D�nt�O�G�z����B��6�r��Du.Z �B��vV~�4��TQ��=�E��E{�P��
���=W��xq�����؎��bs;����a�����.Y�h�SXE��%(yK�������|���³[�ڋ!~_���0���)��^����6�d�P�*M���6���i���V��L�G	f�����Q�Z���R��Of�yC�#�N�*�iNUU��l�2=Yv���B����]ǎK6 _�k��U9G��~_|�jK�nj#�� D��Q�����Z�ƩcN�|u/�'T9�i��4`�x H�hn��^O��4��g�a�'�נgP�߀�`"4�%����ЎO���}�떚����~h*iXU �@ ke��3� ~����:O�� �a8�1~�F��M?��ą�?���G$"��5[��� ����2`�sGkЉ "�DI� Hz%�ǈg�4���T1���2@���E��K�y�̸M���. �i�ϗ\@�+,��Ի�k ��9��t5*:\����a���~�qi�E)��˷��`c����J��P<^P�NQ�����Ƀv��a�چ-	�w	c����.s�7�עr},Q�>�"�ǆv��)=4;�f�`7�nBi��	ᝁx݅u)�m�S9�s�	��x��$��_�C?��`�{�rvZI�
lB��i�=���:�xP�~��`p��;��ߩ�ء}�3�Z���#䁶���iIy!ks��2z�V��,`!�W#�����t��5�5db\}�v�Rb��>��5�?*�]�,�	�<��Y�*(D+�lB�jB�P��+τ�&����x�Y+�9C�Cys�]��r��K���M2�%�(o��(�rum��[|�d����L7�Mr7��\�)N��n����PM�V���Xj;v�Y���	�YJ,�Fᇓ�x�B�j'����.K�ߏ`��MRM���H5�`��C��qp��;����콖��7+�nY��yLe�
��SI⍪ܯж�T�G�@<�e|�omE����fW�)L��&6OXĶ�`��{s��I���^����(ч���-�F>q��Z� L
�]p`��ҵ��\�W��VLŹ/t^�����os#&�o���v�����T�S.8ȇ36��Rɰ�EX���w�a�O�Yzt���3�`y��9C���n��k"�@q�v꒧�{����dN)��m�c�m��#�W�k��J����{�+Ӗ�hĄO�g^M�-v��O�R�أ�>g�^���XG�u�>���yv�?�'���5e�S��]�$7�zj~tVWi�^4�Z7��|H�-�}p�1��b:��@!U{S|-�� ����9�Q��a�UJ^�Y�ճ�:��׍ c�`Б�n�t��k ���n��ѭ�zi`Tp����f�K�h�륮r϶���K���������~QPIk�Sj�;�˳x\v x8�uNmd�Ӡy�~�o��w�T�0�Dԧo����fK���ukv�wa֢�!��αn��ð�
?�~�ȸ�j�݋�Ԓʓ'�_��f>U���h�Fi~���90�	 j}vϝ�ʕ&:VN �5��l�-ǟ�����O�¤��p������@�4Nj�
Wc�1G�:��d;"*|l���^��$�}Bm��`r��Z��k�4��d?vxL��:����'Z���*$�pK��-�8L��!��Q��O�>`�Y�H�@L>�=��@,R��́���L��f �>��n�mG���Ь'�
vz� �YڰJr����H��<�u�Ӫ���q������ރ�Ϟt;j��v<'q��ȝA��Z
Qx��H���V�'����(�0����s��u�Vp�V}���t2��no�92�tIӒߢ+��U�TNP��o� ��a�x��I+��ew�O��F.	��Ÿ��4s����v��9W�9�E {_�S��o5�>1rtG�y)>K�,��]�$�(g5����^�T-9:h�&����٩I�C�M52<�O;�
� ���#�ȔXF�Ef��3	^%Fm	g�A��Lj�%P@#G���a0ӂI9'F X�2��s�c�#M�	��Ys|�8�$��l��;G5́��,��gY��
F�ޛJ?����4&ª|�~T�~��\�<��G���Z�y��
6���v%�3[��;��;(]u֏&Wf6x����lS� :����s�o��*��[��Q}^'k�����wU�&�ꂅʽ)
�V��Ӄ�(@F��潊�N��qUV�x����պ��*���`���Y?�Le#tE]A���|�_8��Z`d��i	�q�·�,�Vx�=r|�qį�70��I.�v6��Ҋ��R�x@���O��f��܁��-��`n�:K��P�H���H�(\�!G��x3���x�W -=�����>8�nʬB,_#'U��4�������Ew�I���t�#��%�A?m=��ݢ�V�L0��s��tM��X2�%@���*��)J3�F&������؝�#��b8#%�탘g�Z�M�MS>�
�aV�����\f%iGSG��rk������t�U��'��N[�z��ܫP�INӓ�աX�!Ue�v���xe`��I5P�ܱ�"����ery�����{�lq��@`�|?��\W�c����i�&0�pnI���Ӯ��5��,���[����H <�Fb�SC�@&�sj�>��,��}|C�<���v\���������5��R��TF������������[�,��*�$���P��n�+5��غl�����s���<B�I�SvK�$z��pYV�w����h����;�.9cFU�ۈ:;@$�����O�0��s��_�4\ Q�A8����^�]��5���F�2�>$>Ό�u�?V:6"=w�����G>yg"k	��x�4��?˨���������\�*���)x���wc�V#5�(�6����3U��̑�>����Į�g�Kp������+N�%��f�Kb~�m���"�MR=W��ة�I�P�aY��'>��Q)xʤ;l�4�	�p'܁.�4äW rw�qm_^RfDG�y,����-��}�J��ڏ����u�[���0�+�?��b�3@����3C����u�����*fm5���>fhO�;��h���������]<�&7�P�����0'Q�^8
Ɛ��5���c�v�bY��_��x$r$u���
5���9'�۹�Ns=Є�w�Q���uQn�;3K6��>��o]^1���3Iif�e{�e�����|ڮ`~'L{?�z�� �����5w�y�<�۪����r�V[�m��-��~B���R��
��gH1캎�0�Ud� �e)D�f��S��s �+�v	����j9� g�у�����FK���_��Q��Ežסٔ�1�VA2����{+P�)tjl�T�d�*GV���	"� �XL͎W���Aqe��w�����A�z#P���K�����5c�qA��ꘒl@x�7��zη�9�Z1�o��:��bM���J�O���g�#����d��kPm{ku�9�C���'hC�\߮]m�ZF鞽��O�^ܵ ٛ�Ac���y��z�#��ӅE�I
�t���� 6��ڬјx���WD$O;��þ�ȡ�4dK�%U5��(��.����T�6����1���N��fh�{��܅�-U����6�A�S�|�<�����!��K�Q���{�n�� 7�"�,�d��T�F�GY�a�.��O40ui���A��o�m�t$6Y���|>�#���3>ɘ��L���˅ L ���K���νh�J�2c��,cx���D!ށŧ� +"U�$��W2�(ÌD}�(�<����M�d)d�VX��4�u��2�C!}�k-]gxS3_��M�V�lt��d�X��7�GMR9)O�ы��h�����b�W��&O��.�� ��.h4Iߤ����,��g�X����V�
br��"ee��V���˪żwv]��W���U�����Mj�İz�c�mD�N��?�H�T�?r�b�a2p"�G��\�5���;"�I?�M��樜/�}ɜ�JO�PomN�c�t���`Nc�w�W�9�7;��1у�n6���F�b�r_6��)�LGM��P���/ aM��
HC���� o�x���C�VÒ�dJ��aX	[yc�z�[�"!��y�{^�a�1'q�	�Uxb�^+O�+У].�b$��W~�.~�^w���I� ���_�<`����!4��Y��c��H�G<��KOq��[�k+�#�:�zmf]�Ɛ�t���ࢱ'�s+��sx=�kgb-Q��HYO��G^�Po'�-�u��./֐�m������}c��ƙK�u;�C%�u�� eIw]V��hCr�X�
�iCk4�����(@?i�G��?D�7��������>� �����,�Ak-�/J�q��hh���O�=/� >������I����F��4y�Ð(2.�w6�.���1f�����B3�P}�G����b@p��;�k�"�{��/���k����?s�����BN�1��
%‸������JX\?5��Z F�I]�� �k��M���^g�ղ\S�H*��=����*n^�E�N-ؚ��_~�C%y�2I�2�:�&���{�N#f3+������y��,��>�@Z�Fv8ѩhoQt]�� ڒАt�A�ݚ_s2a� �����xnQEZ�	7�{���^ !��:�h���[դ;���\�5����!2���4b�s��O�O-���u�O�?܊���x��nN"$�i�	FA��%����v�+��L�[��`����3ޑ���o�Т
��hegW��{�,�)Q�k9��������<3�Yt-�q���k��! �
)�1X�5���G�aΥ��/,�N���s�}%Ѕ�or����P�{6Dc a���i����1�-��ss�:uL�=�<~�&��6��p�y�z' +|�[z�CEK=F��`�5�(y�����m((�P]$^��1"(D��v�OL����M}�<��Q�<�
d��x ����f#�Z����&ޤ[�CV�愂�BU2�x^�9xM�+�_2E�	sx<�͐�(��peyV���<]�h�� �r��,��m-S]�.b�9���Pk�DR~�j�S�-���ʛL�P"�Q�w �����j����_)űM�k����=Uk�0sh�i?��)������>/����"_z�y�������3q�3���8�	��M��OD**81�I�S��������@o�E"����ނ�n�j��/�R�3���M��v�r#�nW
����@-u*K�x;�����K�V�9X�q�y�#�F¯`�us�b.!����_�  �u[sϗv�]Ĺe���[ƶ.�x L��hS`��l⎟-ϐ�h�=��ڱ�<�Ҍ?���v!����}ȶZ��I0�c�{�уR*�*6v��d��G��v�%*;b�q�������eByE7�����o.c��E�Đ���w��В���c|B1JX��w��*�}�f)P �:0�����q>Īw�0�d�ܜV��5�k���|,]r�ԡ?!zB2���;�#�n6[�#�J\|�#ΰ�0`�UXD�t�h��X�Մ%�A@%�H�h�b�9�1(�I�����bs���Tv�w�#��jb��b��E�]e�h$⽓��#Q2��ã��瞨�̜�}(H!-��$��`	>F_wbGu���D�m�Sa#����/��Q�ja��(x��:H�u��XPZ#�7�%lmp�����;�5	3��y)�͹#d����腷g*h3x�0�]b����}�1L6��U�OU�:����o��n#a�ѷ��yjȪ�KR�����e�c��S�Jy��U6` I�+�P�l\�/���<���J9̙jI�j�aKzp��\W�az:�3�c<�xj]�
S�\ls�P���7wL�����,Q������Q��������<�(�8}� �ثQh�}7�	V}бuo�O������D��e�K���n�����h����=���cP����'HHE�� @�s�5�0�\I�_����i,:e���D�A��[����QO�q�ה���nZ�4�Ni�(��q��D��)��D��wC@��\~7�{������4�0vr��	�p�=C�;�s������5dדtw��d���@x\�A����n	*��%�4�ÑnZ���i�ٱ;�ђ�>�܉��kW̻@� zgy�I����ՄS��o�7���L���E��qfS%Z�РE؉�4'Y��Yq����?�0�HXH9`��3�9̒�}Y�����n	��}wAŪP��""�sO�NY�^/Շk� ��3h���"*G��bvT�0��_(ؚ&p��'��s��������9���-I��C�y�������yA6�~�t�p�~���+�U�\Y=r0Ce�V�A��������pՋ�$�ѣs��	��		���6�y05%�����kMF�W|�d!لaF$��i�Ϊ(��
\Y�7=:i���}�Xgҟf]X��H��\��w�"&��ݡ�����L$ƦE��������ٰ�d\tF��*-�]���
z���oe��޴���<t�S�~��Z�O ̭�DH����2Źc03-$��������	�a�/�v�������{�6��T��z�aX1��{��~ǣ�t��OG�G?���>M~���x8ѿ����5N%�Q�|n.5�O."�4d@�����@�r(��\��<���O�����e����/��T��!^��y�g��u۽�%��f�7�QQ/y�L� �xC� ��J����o��D�S>m����*_'�f�7���o�?��0���L�݊J���;����	��ٻ���P<eBu��5�� �������9[���G���"�Fn�Ψ�=����&����l`j\�:pir$+?���.�F��4�E�qY��ޭ����^gp���dP�:p���e�F��9��+��Ӊw�S$A��$��[H��s&4��"&�{:ڧr����ѭ�����M��k(��#��<e�;�;���
�buލ���b>u�k�P�a���O`�2�h��>�j�� -�Ҏa]��F�O�Gs���&o��v[�m��zi@s��B���%�d~�ЋC�]+p�ix=Bdn/"��Ldu+� �M��F�G:�AmG�le��pϏW�@�iר����#N(nB�i��مs-���g���?��^V0�}�u�?%z�7�ɺ6�lB�����m�@�S����Bm-̈�_��UˣU�kZ��� -���.�����P;�tZIF�E<s� A|�f���f@��v�>9@^CQ�|f���"-w�P���؜Yt�|�E��=/�p�x�-]���bY�@�>;����	��7j���9Ǐ�gc��O���gFu�vK{S��$dGS�m�3�C��R�hX�n��
����#YZZNm�����q5[+�t��=WOZ���E��[p2h8Z�؋Z|=x�ÚPv�T8WP�t�K�R ���ǒ	�^�� &�џ�b��妙񍡦m���g�!�4@'w@�gZT��d��
�VaWDgtػ�2��m��
��7X�AkwG�v}C|L�8� V.z%a��5΢�B�O8%U}��� �l�T�+��5�z�� xdz@f���H�@�7n��䛍J12&\{�P���F!�M�	`n|�L!��;��AҀ�BT5��L28pԡ$櫊@Z�*�
1�$�ݿ�ǣ� l�H��x�&���dP�Gq�
b@}P�7vDUEX:N>�T��� �7����D�S9�O���_�����*� �g�!�u��B��ׂ��w���'��<��=<��H��/����p��#���=]����n �j��p�[�\*�t��rc�6�����7�h,���ѓ��M[rG(�\���u��������q뽏��H��RW�c�@�«i��	�B	l1[���d1i��0o��G�����.`��߱�s�;�/��2�u=l��Z�U�U��y��	��?�
�I��& +V"s��l�~�{N=jȯ'd_���-S>��6TP�>ɬ�hrl�)�A'�
�o.>1��t�ª��$2�eT�b�
�P@0�/ɛ�� -��~�����&!4����t�e=7��7�����:�2	�xU���?�y.��b��X��TH{P-��ϗ{��r�YM_�W��
8���N����=PK,���J�ũU-�IZj���W���b�l���1��L�A�k[\2V��*�f����>�gi�we,�@��=��|Cc9�AUo�,0�I@���z��5��x���(�rY���L~YI��"��蝏��	C̛$��6��Q3"Ѱ�
��
���FҴ<���l�mX_������&������CH�#���}��/��-^G	�Y����W��~��U��͢��|"�t��p�+�$IÇ��%�$Y2�����	�Q���x�r*��y�s���.�{J���X�[���CW0�\/�g}m��z*4��Te6i�a�(WL.�B}��`�,�%�KZ�ܤ�8�3�1M��b'u�C�Ͷu�B��N�k�׷ӵZ��|w�NcI���ؠ䪦a�.ہ��5%�u<�*H�kC���&����l��#�4����~	�S���^!���4T��{���;#<?��gŒ��!"1��״	8��Y�� 9h+%�`�a�>&�x흹!N�� �A���F���ٵ:_q��Ӎ�c�1��Q��[ǣ={3�3
�$��ZX�a��jԼ/c�9|D�Y�G���
e��%)y����	ӻ\���q���x�*boOx/N��{���l�آ=��Cxf�?��Q��*�g�B�M�	��Y���/�_�p:%V�~[�,�/h���<�qn���JE�����ozZ�6%�뭮���3<�?��+����Tw&�Ә�Y�E��U9�Q���Z:+!�J���ן&֩y����$��^ΐ�D9+��il��e�fJ<��ʜ�rX_�	2�UXm9^�BvAp�`�`���韂�~u�3����Ǻ-���m���Q����.��̩_�l����06�� ���4�����s�&o�ȫ2��+�)!�#���o��2�y,���p�
bDoa��"F�0��+m������Xţ_�l�r��L�+�廔i������J?��3ő��Ν��8:�ӑj�zCʩwP��4&��'�c�HBM.]MN�"�e��zV݆�'r42˥!dEU�0�V4؛�E88;;�Ò������]��m	ױ!��2F����/F�`'ꬸB|�m��k@o$�v�ש������fL+ӹ�s�pn�ۖ�6e$�=��tT��?��5���󃎹����sL��T��!1�]�rl��eF�ix')���'t)c��ܘ��e�&)��T�ۺ�Gq>��51�Jn:�-�j��/̗��f9gK�	Y�q�}�&�;9S�hNx�~������țް��Y��=����X�(���g�e!r#1ݧ���!1@^��jsg���}����d0�c��P)Ix�g
2����LfvUcRf��t�GG_i��Q�賴]�5��B�O7� ���Y�v�;��o������OIl�kn�iW�8�,)͔�����Q��p����;�C���c+�Ò���hNS�p���-�~�6��^8����<$��
�
v��rU�e�G��c�}LnE�V_�^'��ձ��s��7��݈p���y4?P���tq�Z�|I��ݖ3ӋR����`#������/n���{m

'^c����p� g xM��P#T�ۢI��� ó��;<�@"ѝ��d�#�Pok��E���9�����n$�k�LүL�~N���q���F��ǘ�B;[$X۵�x�Dc��6i��n��ֈl���i
��E�= ���Q���c�8�D�'/Eq�[�5�&'Ȳ!�$K ��z�cV��q4:��$uR�WN3���3cy@>��7١���q� i��8EC+v?���2���0�P�Jҧ�	�a�\�d���;8ݷ��T�w0Ǝ���g	�]��b���<&����_Y��]Xgs�$M��}Z������2г�n���w�P��c�������+�,k�=�]����y��w�L啋�QL�Ά��A�z��<걚l���v���%ړX�Q0��I+Β|�ES���Y�|Ń�*h���= �.j�Q�jA���9k[��;��5DU1�\2�v!)r�����0i�j!�m\R��QIc�v�?t�P�X��pu�jň�P��q�>5�Np�����,���}΃���Ǐ~�à��81����a�e�f��3�m󣧉�.�	�C�s�@߽�D� �On �#�ُ�Y�_4�wY��W5�?T6q�H�����)*v��!�m���>2T�Y~�Θ7���n�W���`��-��<�?��'�j��]����"���o�B-�D������c�D�A����%�7����6��"R� =�����\�T�S��;���������+c�c�r���0ٻE���D(՝(�u�j�W�#��G�]1��\�WN��'3�p(x�K�!ʹ�F���Z�S��`.��cĝ���W���wsl^5A���B���v���_ǁ}��z\���ֲ��aac�GΪ)�#�C~ӎ5�]3�{��Vqn�0�0.s<�;��Z�Iw�����Vu�N:<W��L��w���`�U����9���G����[�Y_Iȍdt$�]T��e0,Æ
��x�.lq����k
R���Wp�����	��x=ű�ԌŎA����P�?VQ�K��c�Dl�n�ۨ�.��?��?�RU�d�?�9h�����S�������/z��J=��AJ��L��Os�����5��+������2���Ph�Q��gª�����o�l!�I$�6?�D��T�J"Z�D�3��(BVh�:��%�G�-�Ӽ�r�v�B���e*p��׃�>)�9��j��oU��`Xd���<(=7;�Y���Q��+����g�<;����iӕ�)g�y��Y�NmA��^C�A�Zb-ʋ���}�5z��<ԯ���b�d�'�A�|(��#���������ԛ՛��y�5�<+�Ǎ��q2����6��H�`��D�j��3l>���D����b�(�m���\jn��|��8����?���p��5�����ߛ��'�I�'�
N����7�btZ��z�_�Y����I,6蛨X��;� ���<"�hN5F������V)$��Z�A�KK���|�EMY���(�����3��gh�E����r���Y XLyF�����rݠ(}��m���4����ʑ�#J>~id"��A�KB���(�yn+f���?�b�d��n���z�^�L����<Q;��2!�Vn�s�NpQ��3�6�~�Ϥc��%��/h���ں�Bޏ߃o��I����'/rދ?�p�������o���ZڴN*�f��()�m�#��m��O1S��û#vu?Do��������e����	�t�b[�Ȕ฽_�aPJ| 2�\�g)�X�\���fb�m�n�T�==?�.����n�Ϡ�۷�+�0�]+ϵi�1`�vI�YUϒA�����F�sM�SU̺����9�BjM��1�X.+>�̊�(���5H�KSμc�N^45����]n��6�an�A���@J��u���,�H��� ���M&Li���)4��j
��^�?Ti�u�P�bp�/a��([�;��\�v�=�f�v�.��Sr <�)A`饲�?��>#��,�7�l��0XX�q^7��>�UhPC��4���E��Z�I�B�L�u�%0��UB��WoG�����/��|�XA:�n�z��G��6���!d'��W�@���y�1�};ߘ�M��g紘���	��Va>�~L	G�#�f���ʝ:��1��[m7��[&��w`�T�/�i$��/�Æ�[�+��T�M�o4$����I��ߕ�]�Q�ހ����:ԝ_�l�c��7fe�3��b������ͱl��-d��gg��R�bB��lHˢH��Be��4YQ�*4�q�\�kG]
��NawV
Dk���(����>��_�!+�U�b�gu�r�H(}��	f�3�"n\��::�G��ь���?�[�bTST�~�ك8�.��������/טv1�t`so���̪�^�L���9C��]Ɯu'����S,��y��z�Xۯ��?K~��,@��B�9=�5��Q�����}�<�VPĚ.��'�5�B���R��H�yA���O�:���;�<��Ə�F�F��GWv�O%�:k�
��J�t+�M��2���7��/��
����wS��i	p�	���c�>*_�}k��b�8��r���!�lD+�,=��!���w�3
�ů�$�,	50��:��?t(U�Mb=���;�G����sv��p���7���y )֖|����}G_q�w�1���0W��``-��P�^e����D�zG���cm�z1�y�RB�ǼIA�✄׹ȊtC�5��;�b�{�}U�����U�ֲ��fW"���?�,.nB���5��o�֢���NBh����hAH��w }����Z��\'7t;qed��s�#�������yEK�[_&]��5�<��7�z1��䗆��x����g�+�?<�e;�<֐o�ioR�2��H��>v#� ��9��]��a�E4�&=��*��ۍ���4�.� s�}�\��uZQh���P�M��Y���'!�$�C5P(�;@Cc��%����u��ЂV���/9��)��)�]�:r	�N���/�Y(��F��}��ɚS���U��jp��q�&!�~s�al!=�0H	�6�q.��z_��8����S�I����I��ӲzT�&C����xѭ]	f�_�XN�k���E�Q�h*V� ��S��TH������~=
�<���{Ė���|{����iɰE��E%Bj�`���x���|��gU�6	Hb�:}����'�0w�9���,V�J���8�ݵ=w���ps93�w~"߃����l�%���0���)�2C�Z���� y]�\�>��x�z
n"�Y��]d1ؖ�����C��oA롌©���:_����Y|�yπKs�3��V�h/ÇЅ�k~���:��77"S?2�j�T3���Q <G��ϊD�e��359|U��#0a�x��dra�b��'�"�j�L��.-�4������W�f@o��6��?�Dվ�1iB�֬��QmĔ�1R�>�@�ֻs?���%���%uS�o�Lk����g��8��t��U/R�n�%��2%���΢�"���_��'��i೑*8�~?���b��ӆ�=�I�Q9�ɳsᑢ6���	��W�9F(On�d��Ŗ�� _�5�|Ѽj�� '��T�k�%ˣ�����:�3Y�T��>�[W�"5M.;�x����P&z�O�cN]�TV^�-�A�
;oۜ�`OO��]��w��E�������9�O��!&�[#�Q���h�7M,�j�;Jo� ]>_'.Vд'Y�m��َz�T���pF����.��)��x�t��MZ����heuF��f�P�Q�����r +��*�U���fA��ǁ�"9��O8�h��X'+C�1ԙp^��gګ����3��g���zly��=�J�D��8鐷�Y�_gi>��4�z�0�Q�޵Qkس�Zh_���4�@aD,��C6��ʪկ�Y���,ܘ�u��ogw�s�< �%�߮a���AMƴ�*`�H�
�G��
�#2�o	$�rHޏ�,��
��*�U)d`4�^A~�����L����G$%����]:���`X?�f���X����Z>��'���id%i=�9eV��k��Eg��6�l��յ4 ��Y�Aq�		��!�	u� �i)];���{�h�9�K�\�-���=�`�e���O?�\sMw<����ֱ��U�>(�6F�H"l_������\p��zQ>R0�h���f����vb��c"/��?,R  r����Ox�C���Qƕ�4��to�na�J~��aF�-\J��NK��(E-c�iq:�{`��x��+��)�t�8��܆��5�匉��ۮt��`�a�\b��3��Se��rJ�$\4L4����Ϻo�i��C���e���Z��h��k�(�o5y�+G���m{��/�S6��]�Q <�@ZY��$E��uJ�+��
�O��;v�P�k I�6�<�$7�h�=-s�.��R�m�Oeq�Z�wHM�Hp:�M�l��$V
��c��}�7�:llZQ�U����R`����>���2z��	£��s+��wӞ,���=bg'`��~�:Y��=�̖P���(|Ƭ���e��(����N�ռU���D==��uk1%�%#��W��>�R�"���,Sl%��V>��#y��<F|M�E��m�u�=�#���gپ�X<��[�S��W�BŻ��X�I��uNWrE���
ߧ6�w7<F�H�v%�y| Iw@��j��1��IV�[��h�V;훫�KG��7&�z�%�+p���%�.�ᴮBQ�y�Z����뇥��>�l�{V����+�&j&F�\n��m�vȀ��!��-1�{��o� �͡�o�)��f����+I���}�b	$�����k�E�>��]�QL��^����R�_���R��B����r.v�|#e{�.�M�����7��\ �w�O�=,�~�H����Ί|�������+Ɉf��S0�ix0)wZ�޶�FzZд�A���{?f}�B�=f̞j��gɹ[���C�[��b��Պw%��3���KA�`�h�Q�N�!�ti�d!]�����]☯�a*E%p�s]c�L	D��M��z*
���l=����K�����i���2Y��=�n���98�c��v�P�h�<�J�I��ky�;Ŕ�@8�� �4h���b0$�s�uq�޵|�D[3��Ѿ�-��Р�jn؂��̓4 {{�p�gPz��ѿ�r`:�c]N��<P�U�Ő��(A��6���4��u��y�3j�� ��a֠e��8V��.2Ww����N�<��fP1c��*��Ee�b�A&sv�ap�*��u��!tXY�H��{�<{9��%X\��Q�촣���/+��`&}|\|��E_[z��O`��!�3�� qds%��R���}���)��ܤ���b>6���$5zƦ"\�'���D�*>����QQ�<ޥ<�n���[��J4J�E\��c
�YV�MM絨+5oKF�;L�;�Q��sN=�=Lƽ�H�O]���gҪJ��= ������z��8g�����Xo������:�/	S"G˭��l�!�ҋ��s��$.8��1��yEw�lŧ������s�X�Vu��*� �|�%zx���X��ƫ&hX=�	���,Ex�~���P�������ҶL���3<�&Ky@�8�0e�im���I��P���|*8�zcG�;^؝��}��oGr���U׏� ��\�縲}}��P9:�05;-(Ƃ](r���ҡ�j�nmږF�HH�Ҝ?p���l�o�@�(�|�D4"h5�E�]�o�R��	�o@���-�̖�l�P0��e"G��k|�~���A��V��|�5��H���4/�a�GDش�;\�^�2&�Hw=��E��0�BJ״�7�Ms	5F)��σ�w�k�!���ҁӾ��2'�S��%u����<�?r��g~�.fNc�3��ʦ#�O�H�U��@����j�\%
�Ќ��\����Zt��1�A �(�C� 
�f\;��Q�Q����D�]�C�� ���v;����M6�0�}�������A�w���L���8٨H�ؐʼ���O�f��z{)�Z��W?<P��ǰ�(��
���D�`�y��rk�el�Zl]jj|���6�r�	��d����fR��g���0���@*^��;�2�]>�_�<A����K憖���?��	��A�s�)r�<�������II�o�]�Iw�j�8�~Q�(;��ï�j�T�|C��x�U���얃���4�\�5����Y2�eEԊڑ����&����@���R�o������Q�d��c9��-MO�m�����%�;c4��!�jS�ƿ見ø�F�"�Z��>��I7.Z�徱K��{b�H5f��޴���}f�D��U:�9���zb�m�<&���u��"��h���2:a�	Zs�&kE���)��3Ͱ�2��  ��E�l��	�'�/A`+J�RS�q�����[�+��@ ��X��3�b��O�q�o�c_�B����JJ�7a�H���w� F%����庄�0+����t~�/�^ѫb�*��w���FT�^KT��?|�1ѱy�$\�i��ߋ���u����DU}�r��i}(-tݘ�'����������=L�Fw1'"�ɠ�tQ��2B�B���54 Z;1���*�G ��Õ �]��!�gPQ�ϼ�a�щ��� _S���5{���;�ٰ�k�k�T�g����p�X&�����9b�_�n���b�D�x]�����/c����+A	_塆Ի:�Ǩvz/���1oA�2Ф�F,��g/���C7�~�EꝂ�"�1(y��{,`TP;'�:���m�#J����W�֕�`���A��(k�HR]��K\0�no�\Lę�FT��:*��\�SÇ���b�A���O@�`hZ���ø�~�N !ɛ����g�]�l�~����B�o���r���G�\�n�&��& �m+&j�kl���|�ڼ��,�U�>KJ#I͖���{��sm?xp�9�>�#�R4)MM���m�=�1ؽI�e���N%���wk7'J勱�/��K��h��[���l;�$��Bݟ��LvkbǴ���餒Q�r��C�]0��O�V��+�5s�M�gť���������y����O�ƚ��i�t��r��{�L�Cst����kef��-�k���5��+�P&#q�
+��1��x�:b[,#�"�57��C���/��g
R}�~�I��� �����\Q�#z��.��z6U�"���=�Q��Nپ^���C��ހ"[^SŪhS���o����Uf�A7P��0ղC�*��3��_��lÝ$�T;�ƕ�Ə�[n�8��9Ʌ����zJ�<'���fEm�7q5	襜d@Q����{/�d�1rֻ�y3�jk0�&U��F���׀%V/o��5�
�w@4���?*�����0Qn��T���'�ةAv.�N<�`�d���(��w_�_,k�v'ZH�d��s�%�=gr#_�ޡE�R�P��[�-F�F(�md�������o�4�-8�֘q ��YE3��Y$5ˢ��9T����bFfS��-�iL��R}e,4e� V�d"* ���v�^%�*�]��	��{��Zc�lN���D~��@1"���C������S6�Kv<�/O�1�T�5��S$�+�cS��;C�3�$�U��5�q���Z�դ�=>{�H�[} `5��\z�5V`ۏ�̝���`���*(b�n�R$�"�8�[:������M-Y��^�1�����yrt���t5���0Ϣ�эC�^7�U��+��Z��+�I�j7�=���y��O@��Uw
�b�D��7=�p��2C|Ύ��_pN]��LdS�@�,���uF(��c��^�^�>!H)�*&�!i7��q���U�9H��g���3�{���3d�pf�r�ק>�v�U��we-w�\|P�e@��?��[ɯf�>�� �G��'Uy���t�~��CA�d�f�)� �Q��sj������v-7�kZǌ�s�!���&N�:Gx�`D��݈In�\
�Q���G��\�M��D
�� �2�ԀE2i^��si�������~H)�⟠�3䙾�S�0�I��]S�>h�6������{�kE�[�m[t�݆�ӑź��o�\�b��o|��`t�Y�`�������F}�$@L���1m̓Ni�d�9�hY 3�Σ�Qh���� ��GlE�����&����;�H�C��L���4�� <����<�(���5��������d�h�J��^�[�uA����U	�!��v�����Y��# ��w�� +�xPyP�Q�)Kyf$a��&�.,>�t�,XWs�m�-b8P@��'~��M�ɓc<֚��7������G"�����=�N��>��1
f���x��P�u&��v������eM�XM_`���gM��PV���H	�H��3�j����O��FlA��9yjV0��U��XE�����[��Sen(��`Gq�w>��r+���M3m��$\���t�ξ�,���h�;�˅}�|Km��~-�(�ʊ��{�Y�眿�s� �H.̞T�� ��,u��^�'�l�iDxU�s��Ǘ���1�,�)�s�� �ь�|���5_άl�0_��C����u��<�E�`Ո��	s��TQ�<e�����QA���Ҁ�)�`��.��� 9qƗ�.jQ��`��f��
��ǣ��^q�cu��T�����Z�`�1V=��	�y��~n���RQ��"�e��ӘeBw1���*�46�NZRz��'�S��G[Y|�^r�e���aǒW�y%��DF$��W��(�t�?1)�xVw�oE1on!9F�*�/�yH3�6�1�۩��P%��9�5�#2J[E���V�Y&NfA�0jOQ�)̴P�	@��3�U�t�����
��ָ�O;��C��$�S�Ca����[������ۛx��_Ƙ+�*�S�Z:Wp�Vve/�o�k̝B���������C��|Oǫl����Z�l����x+����z��bYVhU��6���h����M�P���˚�ZD��0ٿ��3o��_�G�m[:D��$���p҆�����p��N�QCN�R.N��G��M�DU�眼	HP*`}�.3R֋8�mߍ(ԅb�]���(X�w�w"=�s�#mY	xkE{�"ϡ�*
�:`���o2�̾�ݹѐl���V�9}Y[O��-���Y���%V�3l~P��r?�S�d���лΘ��dΤ��U�5_l�������";Q��&T�j*�DJ���'��E��v�=�ހ~������ڄ��{1310{�0F��0h����Y���Q#X3�m7���/�B�T�R5Sљ>+�� �U�*R��c�ɚ�B��<0�L(����q���|D�Yߟ% ��G�Jd�����'Q�������#����^���<Ԯ��a��	�*�$|�ɂN�W3���e܂��r%�Fq��.��O����6�����j3j���DQ��9���c��J:B/�M��g��/�5�����
�8j���8ُ�1M����b����BX�L��-��_OH^���9y����K���cA�~��� Ō���AV	�z� ��t���!�p�Y���F�#��	������� 6#���"ە=���jz9��i����:�F	�o�����G���C��Yg�S n@�mԊ�o��f
0�1j�xÀH��å��	!4��
�	A��}���`"��uq0�$1`Q�N����4��N����sI�������}ƺ�d|����М���e9ꂯs��P.@����st&K��(�-`ͩA���p�k�,-n� �Q�C݊�t��af� _��<�I��?�4� 3S�7��P��<��؟��^�\vwD��׈�j/b4��vh��eL�KR�>D�� o�e������>Bx0�]{!��0tt�$�1�U�d5U��T�yq��Rm�~�:l1h�/�̒L��ޭ���rKV���ܑ]�W�ܱzv�4SYk��dd�j��Es1L�Z�O� Nh�}t���`�|Jѐ;���.gk??V�U���0b�	LM�G�*���Ye��.��k�z��\���S��'Y'�@��#oZ������Ϙߜ(mT�0��(�	S�P�a�=*v�f`P?/\K�JC(2'*8�?����O���q<e�NW>ryQIb��㧫-�,�.�CM�+bC�s����M�c�I5B�x)MYc-�HT/�J��ou��[�n�>q�l�J��аv����9Fw"x�D!cㄼ��r����z!��c�(2�g ��
����uV3��|���+�#�8�2��w�k��B"�,���%��Xf�Oȡ\�1�>�ې�h�N.0�fl�bf��.1�������I��o ����9�c�,�I?���Њ��$�R�*;iMdWЍ��	<���:���X%��.n�v+)F�[7����XlJ�آJϴ���C��A}�.E��<;��O���(�n�w�lrUa`��<��o@?>�!��?�X<с�:�9�+fI�cE"�ϰc-�'QѺ��R�;B���9~4���߯T�������|+;�Se�J�r��\���e�c�k��Ԛ[��⣵�o�]J�{�2p��X
;���}�_?��d!*�͝:|Xrī&nf=r�ޘ�&�!�6�@�2��1p�|x��)u����}��\RW���}��8�虍g�����L���h�L�gxoP�@7�SZ�E��*��t{#�]�Q���q����9��1��#T�Ǌ����jgL��c��q�|Wz�I�!�Cޞ�(2[�}Ua���U٩����� �w�^�,���1kkb�O�"���h�K�ԫ ��(����"=d��f��Dؑ��6�95�F* ƋY�����k�\�1����Ə++ }ℇ�@`�a�Ó7^�/+)���~[��0Z�