`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
yGbQnXt3Pc9RB8X2wlk1OBBfENPdEyHijdErEwI2SJezdgQJOFaEjyecAi/9jY5GscA2MadCf5sz
o/GRYL4y3XTkzhcTege20SSIJKVm033qv3uosmlGEy0pueqE1TQt77SVw8FFigRclTwL3bV+UKge
c+rhtIxM6amEr1+E1DUhXmJh7RhFQNL2ajmhJrbqIt5B8SMDuMGQWSjUtCpv6LDW3qjBjwurx3Nt
26+B+jV4xLTlOVNdIvrZQQQu0Ocb4lheMbYmpYv3mxgZXpk5bFA4cM3tOAoStr400b6FmYDXi+kF
wmW6jn4Yk3417ZlRXvNNA9lXUIGGEXCMZyrjiq0vGOYf5N64rLQBTB119HPXNXq38IPAnrPge/Xb
OvGkZyx5ph9MLmRP7bGfbdGSCsa30RAyZLF8OGHu+BblGHEwqSQZ18R33+ThvyetDzQHPNuJ3D2G
PRp7dWGt/v2JxCthrcfF8AXBIG/wG/3x2WJu3+vwh+1xOqLA6o54Wjf+LpX8cRNwQ+npm0YQz7Q6
bX7phONIruaIax+MRiTxLaQ0YC4E2KFfDUbRY56IcJxEzdoXRBXlkO3A+6AdvWDKnwUdJuIHwDYg
YcyMlRR3O5M/LvsoJz+CA08u2FRNl2w5LjH7qnr5Ml1ws7H9Y15aZienqqEdqlrtkaJdy3lQjqgk
gmw5x8o7pODuz8jYjsjqJlarfvnu+X4O043keQdylgMk3Wszm4Ew2hNtkBPK/X+F9I6VLmlYVMDD
GvPMRjtCpGKV6suUfhGEeYpLYBQnopmQSacb0vbZ8ZPtkyVK+x/Mr9AhLRj7k2mlTxGo7/KgzTGC
uLEO0qiaNK1TX+qMiTb1+N7JhHFG5D+W7hiTbuBE6cNAGfw/UVPZLeyRLD4HYtHivZEmqBAzVla5
SPm+RgWFF7g/Q9/zEs/kufM5S/C3J5UJRfqPD15+lkXnAvDrvHM2843nontggUE5371hgQqI4kVx
Vq5n+PLXE/g7CUalBbJV2q+JKw2i+P0Jh4oDoSrVnQrc++ERHrZ0E92JJThmsFEoNAzjHiCUWNfe
iWvUQHdWIa/XjmYqE+xlI6TZP4oXCairftxJEUL7JEJ1k2SH32vAn8KEdXeD4ZyW3aTxbuoD/GZT
TL+Db3RJFPY/wecH95E/DMkQiY/xVD3trxyRyOqOToIcgRGQiFbPcAxKC5lZywrTWw4kM8Nk2nUR
3ZHBZ18zGcFi5SGOnRotvpAxjRonMk8qvmdtsb6rZwuFAvrFZB+JobJ++8FcnDpXi+IQ58Q1P+sX
s8J83KnMRy3+UJ/NzVNCV0kyQBzytM9DNOFlDVd0LCiXi1SLi5DxNJLcNNyuVL+hDveXffqetQxZ
d9KPmZ1ZBSmSyPlYgBThpz1hsMTdZbIJc5pkbCHKmS01FuNiR51iA257CZruSqkEam9R3YuMXztI
beoo2dt4RjmnAl9VL2Qts3LKcvUN/0u1t/pAQ3fphACt8VqLfgSIG4fEC6uKLFhjG0xxPZ4E581/
3KdQwX0yFCOllAuJkRZ9zCowe+EwxftrhJH9tC8DqqMNo2uQq6liOut+bd4fqQXREjekrfUEWr+j
4YvOau46fYOtE8S34lpVrOLmxaLQCuLw6Y9DApwUAozBllLaML6DuqV2LH7BARSEpFzddAQKY4m2
FqWrZ0t9qvTNNbXdfX6xJqrU39ZmTVLLkKIGLWVdtimysLtNM8KVLyktfn5q34jAndZU0FwkMnAH
6UW5A3Ifs2eA1TAupNX2SI0/JuMCHs8O6jjqEByj+ANeUblqiWdCzz7BxAJswURT2hUrwtCyxfXq
SHL93L8PiSCxzAkLhvWMfa4LjjyKX7c1j2KGvurmGJCMvL2Sb0mKFlFpHdJYRpoa+Qv2l1bq8mIH
E3n6G10/CGwFdwA+aBBgmGaVkfFwL44PHV+bTpkXBtKPFsoFGYDERlkF1FXbbzHpwg7Sly5cCkou
/rB+u9Sm+/mqM/dmBQUKTFc7sGqxj8pc7a2Wzbe0Ls2uj65MpHqugQgJ6GSg4XCxt5jJliIb6cVj
nSNP6pqQJUlvnOQ5JmZlWrg7w1MPVMINSazFNAww9VlllrJmz9/+3tptrASNlHqolNP02ZRpsTh7
SQlg5clYOHpOpk6zGnyRsrrwZP8NAmdJXbkcUitzGX4hB0LB4gydbwvXSveNb4PM1pzVyhm6Edbe
s2obE+9h0UC8etrIcgmm/DZC6DvVYo1M/qtFXnOdnEsYSU5fgwOd831BjId2G9rljtAprUQEk7Be
Le13osxmzhXY8gZEqYLG/ZY9llq4ZeHdMgUyMsbgyG+aoPWrg+6bCVEJ6x1ZS88gxXXLsc4bWKyB
ASBuMDn8IY9+KrIJVd9zyUQPgp202Ee+jvBRIPNnigOEOCndurgcvzbN79ZBrDRbJEyq/n9/CFls
d55F1BT7OHP8fH7eXg18ANUxcSjqnF5bn7kkvzSsvQgB4tH/Cw1ipgIha2+xcy0SnQ9lt0LItex5
1KNZchSG9++CjLAMDcJlF43s18OdBvrkxWuvFxoafN8Erd1Ti5EYbHdeP7ySAd4jME6f3UnMOqxU
mpEoJaqZ+8L0C2ibKNRfnOq+4LP2rmiRyp/OdxX77Iw942Yr6CS0HzIyixaVLW0OW6w6bc3f5brh
wUdkqVQ2S+iSlpZR/7Yr3mGuzpgMt9va7CKoPcW++endub4/peNz4T1XBbt6TkbpWi8Op+xYxiJo
V8Rncu9/f3Sbc9pqeDsw3QTgPHIfmDFPFMSt/KZtGllq32P8GeLvVbjDOweRsOr21z2NUv92O/So
46o4qvD3k8efNV0IglUBEhO+o5uvqoZOmD2DE4S5P+ubqIdKU3rLqSclpRChhtbQ1oKXPgfyQ34N
nybVf3ayvw38+rTVFoxAnYBN1IS9jrw8SikelTZPrIugHvs7ysiTev9iospuDS7ExCo3xoNWlc8c
1v7uNc7HkOinucrm5rQ2Qywn8YVksnZ/L9e9Pmzvu739956isoNkNBjOgZEtuWCm/y+6GZk6VkeZ
zWZf0acFNDt3ywGFQPsdc7lpqqQ0wSDx1WS4IsXd9qoeFlz2VPw+QVsinWiTYTZUmrxPvt4czL4A
o1sB89tyDBJ5c5C4w5kw9PcIEumGjSL79z/a2gxD912XSCYDvi58RqphEfpbscJkgBGPxthqEUi+
yBu2rsXxkRL3QiXH+Eg5Xb2S+eiwSft6m+YnebDmCcvQ7Erc1yZIYCSzfdz2crLT4uonQOdNOD5V
WZsCpNuyQ6ujqvzvqoBB+64/PUqhWbW3YV9rwfdu45yKj3B+r5nROtvgmIrTggiBu5IQgkG3TaOv
tVrpC/fN7GxYWacH/SPR+bMoQRpCb2Xlkbt2p4AKbHKsQWVojgSCCHMFC6DOBRX7MzVVP7Qao6Gc
DGl1BHj92SICoQEJradtx6AJsjowlc6hc0CmzOKx8LQOhh5qYUuwKTVLKhyzAY4kuhC2KO8Kb4vQ
rC1u+jtxr6K119UeAQorK4XoDHnT0fBssD+7njIYFYtXrgvaROrmVzoOzAiMPZhIi3jvpxdxEscz
fJLu1xd3ZlQwQf+euZ2SN7Ri9gshtz/8VkzENKBh4mBOJItLFgJdW1SgGzKfnxk48upHhzo3eBbo
gTNaIJqjlNXagrEm577ohT8aDnY36Lj0OqK4wSykwq2jqKhBOIBm4cvOeINWyT9QcVxWmLUHQIeM
A76RKVAHoCxG2IZAw8frkv94Zi95fmH+4A3d45j6imqLbsTfDWxpC6fMTUm16ApmWoYOj9WoMl+h
Wv0S+6BB53BC0E8QZJ3Riq0nPZ6C+xE6oJkUrwdepuoxgvYtO3icGpneXTirFKZP0WD5mfjV5CbQ
mFyXG2iPUp/IUuVcSg6iDtPsuo+eAycuZSni65yxb+s+uIzE1/JPse3dPI7pZtPETqbQwY64ERlX
ym1kMBe66jLen5GBUC78vGj8aA0XZfkdVdsdrzJKWRWI1h6Mgo6XY1QVSchLiVlS4faQuJAeRkgD
/OucnPpxN4oV689sK6lbqWmgUxbjfWp7OTZBbIOnSdEuiLxqZFvrIfy1M1q2ObOHIKAZXz3ivoax
isqRFcDNoFq9bsog3HVtLM5KAY/stfqHYW95j9KmN1NlkSoyyGdy3yu8edBUjwH9BMtlotvhv4F5
Xn87kPFH/zdHB4dNGp1ljqYMqFple0YU0+N0aIozRVTCM0U67iovnHMGR9xknBg+ht7yGzNATZFk
8uLhlGoLtsfDi2VLuLiRS31cZjyESg5oyesVATX2zF9mHlFkQQqTb6RvbJvqt5SLPnVTDOu/OOi3
NMEd2AnMVG4hIq9dYMTNPbpkN7LeL4TZpNb1eSz1gKcXmQFVQvThwo0tZH/46ehEZTFJ+p9m48vZ
8vvMz5iWhYTKaQebhntEu6h7h6KMh01S47cRTgSLiR4PC/iuGsssiKYZoFrQrwNPu+h9Bj5I2e8X
3vKIXxLx1JAU29PwjwovCBG0LqYchxEba8fCNAkrDufR6fKalpnkZh5VSUq3fv6QwFYfp0OehMse
CiXrMF7mCZtZR/ttEHkf9LPBG7IDgAqfJYT3F8lzcxQUfCWr2DS2UgA0CvY7YLPpanmJgj1KAaZ9
A0qN06V2jFBaS4tvpEhn6HqolQUsIHaAcByIdfJIzmzyB5uwP6RYaQMgqx+aa1JoDIlQ0dFELZWO
bO62ckklyJqcUGKaN+sLgoxOA/OMFtTMs0ipgAFnZa9A95VMEULJ9OthfX3rTqOkZq2kZCZ3ygPS
38zcl5lh6cw7Fih5W7mXY8DwkGkQAhDtkss8ND7SxNATP4cmiPohPIaJ5M6Mpsmz6VfMR+XoTyuD
fmeZAoMNjxFf5VJ0a/W6Tkh2jjBIfGjgOOkjDqE22zH8Un0YXGFVdfX6jHeKJtNTC+QTxzT+vuws
TFstJNG+ZuoyGrqlOZgB0SYGKujQurvf24sANFmC+Tub56+bZVluXDw2BIq13EQD5sHQ8Tu/htsT
1vsNukrOuFlTT+ybrDQJmMWQv/xahfhfi2/cTrFMYG38fg8GG0q6zzYzglV9SkZpzzEBhF1d5tq1
6ChdFzYwMYfGL1lfPCKZgnndqcjVdL/lKCrMwKJ542G6R2mBVBGNNNwl+SqeFKlbC75cj3clEiP9
cspll+MVyPJYCJXW9pIrmwFWVEr2Y7qJQylyuAlo+5M2skZvaS0vKm/zxbUYVP2P5/gdKmZQe5CH
nYuOXLwqKMubFlnMrhDni4EzJpD/aasnUZfkP+3MM9CjSM0BczAVp/kmQZvB02UpkFYwCmkDa5MW
rtAgnylJRasR0OvV4w2FPSQVhCb7vQz2bVBqX1SFo2qFvScA4gfSFZ43BnM+tPmYcLrvJJ1cAgj2
DdBUI+vqEnIYO631WX0WYWV6D0FUsEt/3PCGMK6FMfIwyDndY+zXcYpmXAV8fSq7BpY2DNqpY6gd
eWjnZWSDDDgdSiANRDM5CtoHQRrIt5lfiGDqqXb1tLpi+E503ozqaXROAkPy+a+oyqIeLp6zchMY
uTpKXfj4F1Y64OLcyIs0MyoVCvZ+JexLJZ+ePYli7WM9XZMiXuLXVMoQ8SP9Q3wJpAEKtDqvxdfL
SHFIEMfAaw6qxjZbZzKCZ4mSlaz+zecIxSx+oTQEWbkhvey0K52+VA1C1ElVZg7MV9/QawncYz59
/ECb3ezbJ1cZZRAvyL+eeRl5I4zPuPtC++P2pr8eBnXRWjn6ZM7VEILyxLrNO/OnP+558y2MOweo
Bobt43GolV58JsIYdHj5bNdm3GLdVgdwHorgO/yA1n4HsJ6SN0oVOtcKSnMxVPanP3HPIlzHhDut
gxHZGBEj1d7rvF7fT+hPNeiGJLH/RIANvWuX4Pkf//8edgy98uy3HlBtXfZq9fiJZImIK/Dmbqt/
1D9X6652jF+zO8ak5A4Bo0o4JHbZEDEqQTFgUrZE7xOH/VzB1ju9KiZJzeh8egf35DjlBXAse53N
nvCWEt5ihYftyYrSe8uk6vnYwZN1UrpovtVG79E7uuQJ9ibVER057R/GGUvfU2q7wb+xFSlB9etP
uiiJbL0yY65dt34RiLFlXBQijRSbDHE14S0/0ZI1Q1VVhEWm4f6FqB1ErXKikhKgISqMMuP33zCc
15YrGRaKaspuM8IBcvCcT73FWaJcVPZcmZBij3Dm3m4O2ASrtbgXJO9IZDMYV3hIDiMv+mhWvYt7
pragsS3lJ9eAJKr6pix1NBLCRjWoPkF+OzdaLnjCK6oWAW4J7FKbGAnlmWD++DP4R8CMW5wxiGnk
z5snlzxNVi2oXbpDTKyXjkaq40we4Xe4KZLtrQ/mJ/1+OZF0RhC4sVVJyk58NcPxt55xjzdtY7vx
rbwNLLrmvnarRspFgwQ1el1fuI0JwpBprVmdKnDfQqLQZ9zC8sr3k4sQdHkD/sdRE2TBIji8EjGM
I2gcXZXzdmKmIP9kL/9AR1SP4JEx6hdud2AtgHvh0EnsaHShv/ZBUpftnbSl7yvUccNLErkOYKk6
uKGYfcLY4Ht8r4fYoOulHFj7ej9ghlcPFPOuv1G5j9pKyGQ/Y5reDezy0mxZWgfACTUZV00PJJII
EItZummPXRM/KlHQ0fygc2Yy9jCm0qksCByVa7S3hBw/gkav6uXp+m18S98Hmc//VaMS7Wf5M+ED
i8ASD//OE/fRB2dEwVPkUjNVT45OrfNo/1dpUOe/AUzYll6NGt//LR31DLTYMpa3SKxsc36Gho1Z
Tm84KLar1x+dpnLXjw030RU9+5FzbG18SItrVGmU3zowse6P2soWLSFjWrf6KzchWCJYTNMwpFd0
IuM3Yghqx85gBrSjBkZzWBjDiLOCa0Bw1HkWmGxw41U4yK15ODJzXb21X0kcV59CIteSjVtoVL1Y
lLLui/bb1ugQZbEGxemLepw7NGllCrZ8QBoLaPJea05WZBJMDETd5JraV6GFkGLyHTqhi2PirTFn
ciQXDZvuk9eifPECU72NMovi8e6DQxedfS2by1Jpc1JW/+SQPypB4uvjnDNTdDJ8jA3u4vjCxhux
Ur4nsh45HqVM6HzFoROe/LU4BBd1IPp6TJEQfVN1C1b7QEVvVhDAUit9DBUJlqq21lHR0qDj8ZXU
malnty1372VYoydabDf3sESpqE5mfNpYSWrKekerqYXNYcIhnCyTdCw+hup1GfHYl/P8Z0WuIH6Z
lORUJ1zdrfHSYimRGJT4o2ifO8SRCF0eMBP+bniTdFkj9ev/Men3if0A0zrvb4dcDW0QYxbFapU3
eiC3THvdQvD1rPXZ62qzFl4Lo5CdMWdlV/nnhhOrU19lnNGPYd7Sncds7tStLGVqbJ0/5QY2fxUL
ZsyTERyHjoz/PD4TA4eohH1nQwH6Avd8DGPN1dX9F3cYjy0sQKU4GLEDeLPXLY65L/fOXAOSQO38
I6l200yQ/bZccDgo9SLiuvItEKxRnifx+mVUIosfuOXgzbWbKQTPj4FvZp/uruCO0LRCaxbioU2s
ngebhJVDHeQSurT18PlDpZcLmircF2LjcPJhgMqI1iGAPGGTSjp5LOl3abzx7thY4UOqLTZhFP2w
dxOeXo0n3yMlDPixPlwVdpJX4pLNzwwpZfq00jEKgTwbIQjd9OW/Nb1crpGW39Qmk5EgmiECPx+N
ahhgdxFOgEAbRPCGA4gWrF1UaEoFGp71mWghrVyJHjfLK/hNKD6p1mo4/qoJRN1aiPUxBVDZMbfn
evtL8/BpMWIvm1QMqVBWRhcDUQn1/i+r1W2kmaD1HtFm+v3g76OoY6RI0BN+62f8Q530KJbDuA+a
0eezldnmwlSX25Ry5AUcTz+hXHeDyZ+SnHyNm/dh77yNFlQgNf/qNO5847p3mxvaKVXwwze6YP+9
cp2g4Oeux+mBO87S76VJdIBq9XF0qDAF1l7axk+b96dg9BeV4mGPsrttIOHdvyz35bnZGCK4FfZ+
k01xL+QbRlsAMq8XVGvnZAb76cHEyFm1VvR23z8pUwd4ogbAx6q/bnntxJQfQCZNNkqFgwnL4m3l
ArVb+G1Qz4Uy4tFW216bCEjGpR/ghLeRw+2gij4yyguiZcJGgmh21d+uDFbS2aUwJIiZIlAnifNN
M3O5465VcrFCYvrM1MZVNS+XAo5qgBzLncHSdmobwSSPhTWxA/W1PsN5yFRDwT28YPtVMSMH3EKe
2o+N6OjGnAz7jjuoz3JVn6xQRJ1IKfSFY3PyqKNN3PlSfXalb0vIxY64w2LNHzJJIHyT8H3xXlm3
IVfm3BViY1xarnc7kthju0cwE8qRCWskDGBTaM+HZZJsohr0l4MW2nlvrV0/JppM5MkxLI40H6lX
HMlJlGbHPiF/iyrnkUxUkD2Y0pA7Ezt6SafXvGrCffy2tkMqPprLrfNOS28Jaxbhsz/P92+FInNz
b6Ar6aEZN8GiR3f2t74gj1X/vsYCIIvrWrRTaItZ+uwDYfnfZY0ok0fzf/5+0aLKAqFrxe1gQ/lq
pueXnGVlx2m0R3jkTEySiieYMh2xxN2Ar8FjIiFuyBDIR388JMJJXA1wx8937PqRhdr6BRSJcWqE
+ODjkLzdSCCFg/zHc1J6zuLBO7PZ4giQjHd+Ocz3AkT+4X9e7FnWAabvZQGOaKgXxO9JQXbyt09O
74DQ6JU/wBS/pRj7eg38Oqz5c2IohDVFVjyXhJ2QQlMhcd79kt5Gujth6MS1DWeeDTyu0j8enU/u
6Xnd2KTo3tKch1fNE1b8ZMIwCEtrrv0xP+wV9+yM6FZc2Q+ymh9NtNpM6ynh5YRtL3QwGnpraNEC
r4BSpp0AYhyPC29AbjuT3ixpJnPDR6k86jHIVhAIynoj17F8xUFEyIjH4+9YJB1NDcl7EUH3efN3
vtWyA8gFoMMU+lxpQFAJcquMmNucHN+zzbenwFg4avPx8RME6sn6NqxE1lAjcfuXmAZkRkGeMqA6
0mXCtCkteK3wJ0NGsUpiwpbygA0+HUA4fzfmvHfFrRmstRIlimahy10w5t5V7mkB/7JpOUAAmngV
77VnhEdmmMgxSFPFlV6HRmC0szcU6cGRzAWVcaRb2zTyt4c0tTTT1YxG/2CQBt+eSzwW8nh0vqoa
GgPn9bw95+Vg2QygQN3iDuButzZa1GccpWmnBUWO0COODyui0EHkm5ol1Hk2cVv9+73ZrBOcoK/S
sFqXChpwPIpM8GThd+Jqi3sUBpWx3LqEZJk3d1aG4xb/YdBUtskECBV1hn+PU5o+sAJAIAtLEcHb
Funy1u8+16XQVrsfUxHKmE1f1kKqmZHdosQXFgifbE8q/j53Q5v1j+3qE8HYz6BpeUZ9MosT8xBZ
+34TVY/JQuGgHvYoss0la8QivFk8AwkI6y1ok3mcLkDBrn1lgGXn4xZvQ0/4MYETN2c+SHXa5MBY
ap8FDB8kA+P6vRl5mzEmeSvE+tgztG+c1EGE8RxUIqZ2Z8rcKiTHRRciStF586fckgm44oXjE/Ae
FIGYBMkI2UE0UcRq8NRK8Jbih/ogdn2BoM5M+ZjQXRJJzjrbyF1N3wT9rZltfH2MEbFBgUGZWSGq
svrauHcKfwDlP2CwoZBwG+N1Z8+becWQo1uAfwvssWWjDp23O6HMTrm+VpyMSdzF3ID9IpS2wAhP
WUcRwwBaZMjAT7L3L14LIAtV3Wm+PRXSXOSr+7khMc1WhbjwTjINRhSXUZRNv2tiv9JlQ3RtNcUu
4F2LsWwRJpbGhXC5injR/jcHNV6ToJp4va5Plo7PlG/o6HqSM1gDpgIA5Em2+hnWJeFmktbub96g
9XpyYsVJqgoGJPdX8Fu7rp4XH5TzPPAabVwvXtCK6ZmEh8w5igUUKFpAsKK5m3pmCmAeb7LTBAlE
mbrpKC1GBPF6mkSRdhSVECMtYF8DOK8agEBi2EsfhmrG3sGoR9BgERvUOZvzTqk+l+5ruk01VYRE
6ypmJjsKus2fs5ijMttMA55Wv7ToZBX5EaD2A8lEJkV+u3yAiXiFAXB0rdVt+2JpZyYthKTIqQYJ
QrB7YxeSdEhZeXqb+msocKE9Y0UTDw73Jg3z5ju+Ww4tjMwbHXbQOCtDPZXuFJxv1E8idJuf+v+S
tw5o2HrVRyQnhlEKXGZJMCfwfQeNGK6P48YKXsR4VTRh8A6I2UqJAHb86nI0OoUl64//PlCdlXk0
edHAyVHLVWCYZWNVPtEVTOBRCZUWJnV5BkUO7nlEx6AebCorY8a1GKdC4xvnr4K4//3ejQrLVh62
VxQtG2xwAfJmu2g9YiA8bRElZN26mzqsIunj5MZ/FKZxo5zjc54KNvHbRFHSFYhX7Xq6jAbDaSIy
BYuyF3b31tlJhYKOSfoQ4qEYp6Z67F4EO+8gwA7zbJBMbvrYSsYeYzrZbHIKyDa6uySPtAQw5qpM
fYjag36Sa8csHJirB2N7x9uMR8LWAlJZZBqBMPHXbM0k1/2OQKf8EIIWAhOiukVo6LkRM7tPyism
y3K6e22+vDsdJoIz4DRoUOMzXA0jlBqnqwFO7aLppaV/4ynxR1wLxF0IZrghBkbCCcD1oeJLywZd
VhUC9p9bpR+YHb5umFQmE4MlabXvCyorJSfrTUXtJo/11JGvYqVzOM49hwR+UVhblTN2hiXhatIM
IuHsPpXOY/bbQc6ph9YX4OuBJqo8z9nrRVt9m/9VPhxtnMErjMcmRUKt2B9AbfSIq3Yy0ipQ/d4t
PciSR4OY+LbBZ+TS79RBRk7Lh+4F6tg0/fowX7YVRejVnSxf4mVLv8tvbuvf9D2NzNoHVVzLt9OZ
FGdFa8nBkA/fEqrpGuxoofrGBtNtV636ZyjBH8UHRaxMwnRojcYiPl9+ufU6sWSZuoxpaMv5QWKs
cKpkzbob4NkIDX1FBNq2OUMBJMIjaVNQLZPcswQQMx2xojBKxxzw467ZSHPoORr82L71WxWWdpf/
t6DrXj2L+ZFCyJytgob97B4GeSzGtOPW67RHuhCFvfA0SAy/uNmhLWJW8xVnFcixO6UtNayFuL9b
wOMm2CHyfDidimQb3gk6PG7Pxs/lB5sXrdE++xm5MFHNlPFoUmJbq2zTXnwfaD3/6PcUkddZVhmx
j4v1vZwdNaB7nH6E+CasyeBiS6fJ/lsxpzDUuYc2iylAdR7G4eBZNsf8n6rPyfDTYz8IdP1HGko+
3EyzVxDMmTKZ/fMCSCpXL7ayH0sGUNzMjYdEpGA9KBUC9iCfqc6GwXFPzqkPzHPFZnOJQxQzWUf0
R54jU4r7C7qoF6zhYPn4y9Mp7TY9bDU+7boqMyL0hjMP4sjdHBJFg38dlwNxfSQKYSQZKZ6PPQHC
Vu41BwnUMy8I90SAeG1JY6LY4XnpZZM5KAoTRLKQ5Emykx0euK45cRDSG4pWk+xXgz9xDGlL+Gg3
x68DDZRuFM4vQjVCf8Sfv1JqPoa5v+lUJDJgH8r1DOsM53KC0U6j+FnQC/20cP67XZGRiuLKuqtL
+Mrecnz8ul/42qcdi4bmpBOvs/DFHFTArXahdkqpm46MRCIHnFNKBBCFn7GMbWmUSjmqGjl8qBoq
VLwEez3KgTDCFfZOB8bqjgpdSWczhhvbXDJsqtwb0eYAQQQDYUaJOG18Hfqds0Bbk0mwb1SOIRX1
QAUrtFbvOJlF10hMrhfHJHITyfQVLBUt+CoJYrH8SYKmEwuV4ef/GQq/9XnD2AzY5HrEGHcB32WA
kXuxT4Cx/KmWWHI+Wmc7Q8Yv+78qCLpwX3z0dS8iSuvcLnzZtxNt4cbi8pFx1dol+GKJCabvJZ5N
TDQs7v92yNGZFjHIL1rX5ahaPa9pqqYOi5LioevGWHtH0p5kq0QfmrsTXRk8cmbBpUG52S6o4Qxt
iMalzw3aFArPmalKUlZCq/fvJt3sXaA1Fz60Xty1PpZLKWJ38zTUJe9FE6BH9JLML/4VnCJbPadd
YMMQmTEV9qgr0nVefdRpvZWC59KHouLkT0VHxNc2IkKcNAJq30d4QBY9s/AKmgyJUbCpkHFLc+5y
SPz+58SSuzja6c/3JClLFhyff4jfVgVPwGZzRiePLH/HV8ynFWOuyE3NCJGzyH4bs1MpiZ0KmqPj
R66Ty+4YGtZbYxHPZ++g0Gxje5TA/196eS9010b0S/Rf+FLuoxuoYaN/6At4Ge7/RNJXHGNJeFNb
wrHjghjmmwj7GtMAms7oCTskvWzr3wm8+OlFoLdiTqkLfLx3/pl0SIQQr3KQ6FpRtyHy68NVfJK1
uWh7EJ+iubKeaF+7cTLX/rEyI0YWmBCr/B6+01Vh5waFIzRU/bQlmDdD3FcT6occidpSadOyAA62
t4hlS37q2p3QKuM3R8bPYEeloPzSUPKhIPmBsg7umgQeQylWaZ+v5SCMbd4782B/BK+eEQVdbkZH
fDY9PF1NdAunBTQmR781Y0PXa1C0qyUIR0mNpFZ41Mx+vGRa9fbWEyj98ZLmQMEc2vfFfWgdxYPH
Tc5dkUmwq22rJExP5YnrKZugSfvnp56M3YZscBwv/MlGZ6htdt8wcpTqAHAZwVq+vQagFLNx22K8
Hnl/1EYJv1ovNuJEUg1QuFruI1HEy3WI96Ee61OOEdRGwciYVCWjqkV5M45eNlKcTQXlsRoRTkuO
jzJlDWodvnXmqucsMIHRnsoKbp3EU+MCiDcdJ+kwg/V4zWrYRpOVVAdueq0sqJUczwCSmBc/Dgl3
th8iXy1LF+z2EPDbpQvLEo6P5JcBbfhF1JyPg6gJldEH1qe2xf1ROw+neqQ/aV7kUnKvqI1dp0+9
etOCPrLzGFULR8R/5Gw9b9P+iwkYjxaB8BXc2jzgCLe5UBN68GgPCY5Y9kKYF1n5fcjtfWvfLsSv
vVQ4CbSYL+ezI1cuSfCvRzWtMYfCrJ3qYBC7rpIbwRszv7/Ifh5dClt7iFLz2Trxz/eG0cizeNxt
08NC/hKs6xo6LHs3TfbDbWh8/uBIYmtFkUbl55IUwg8ootgwqAslIGd5oXci1wZihFXl15neWg97
hI/nxJdRAWIXCAiXvxipvEqxFMsOEpzDyXNCMVymMrSbEAgbySkJFbEJyDx5Ay/v9AuvEEj8zVTm
Ru2NFaDttMnrs7+SORBSaku9pfJIKoGu4H4ylHTcnnqM+NLca6/AFM43MYEIOw6E3N6uR5YAzlkD
oKm4MXCzvSTrwjvGM06UCYZPi4F6Pei1NwGWY11ZDvICycsju/jTnX6z4UL7Ef9w6hI/lz/H5XqK
WjipQudlGNHee5PAX3ARhmMXot6LCKM+QisMd5XD758+olhQpWKgrcVwrKk39XHmU9PzHi82SWa2
M3/kEuAnKn80n1NDcQjqx0Y6PgOHNcmTvbLEwx8eC586qHseOt2EB2DmnlXeRx1wRr0Vlz0Hr9fj
DAQ92+0HUyfjfpv7sSwUlH3v3lEoo4YBGcUOjpQMEN2HqeDXykV6LdXiv0JzArSTBHRpckPP0pH2
lK2jDVNR8kotho2d3fWSz3pjnB+zTCdjgNrHx3HEChuSzmA6AauT2L1gH4kGvsYoGZzE+ZR7i6jP
55qXNFDhaW6AcUUHPVnPc/+xkNa9J0l99brddlr371r637T+opz4guntEjiGZZHvdNtb6NAmPpRi
C6IcX//tPez63GprvUPwwPYWkd0tUNwcuKdVlGfdlZEoHUSkj1kCwx0WRfwqCPR8uZR/MycOJaLs
oDCmD/aGnpuqqpCJqendiE58hLWelaD4tJvxOwB9wVVgVtBbrBg/9je9VAU2uVouVWwkGGr/fwse
/2+atJEMntf4xO2uQ1QOqIXjDboR3FhP5mV57BFhv60CVcPJO/vA+WQc5PLRxz0Jv3Hcr659ohBW
Sm/Rse63i8qI4iPZHds79MonZXTGUc4MEED7BQsX0jL2zk96mIsiCy3oqzNiSe8MPoKVxDL9I6bO
gsSfICLXqCrktDo1/uThUnz2D/r/ZQLGJP7LvG65MxSKz7frvDtOMM5ehhnjc9gMTSg4mjliA7MJ
p62AoVTZZPTroJcpLNiU/LNlsJSz9IJWUndsbmXy9gzr3oGiOCwDLW+laiAgY1LAQPOTe3yeUYOL
4Busc7f00KDwEVKIWmawoyIIutf0xwTax2fNAAFFzixKn3sowq1WvGQv6UaNY9p2HXUWILEoJxmb
xIv+6AuebAfyvelyg2kXx99HEWWP0Ftvr38YOdkaw1cmVpNKPBzX1Kq7AMUrHvdTEnChoEKbX2UV
dpkt8Oy3IJjjcR/UPmD3Yw6QyR6PfMoKBpXQkEbCv2HsCpBXM3HxZKtPYZRymrRpapB6l+MOJ1WH
5rKueQtet2R1Jf4VNeXRZEDopLPK94Dj8AgPhKXcN2l7As0gIwEvyvgjOoGngP7AuxzdF5lL7s3i
l3J2DD1RaLWZfCFv+GAbQWc5pgw7VHHzduLfCMyvAoJT5mn7o7AYc7bJ/VCz29v2PsGFDYtpPeRD
TcU5miPUoZkYbgJLW150p90ohIoyDDSU8JH5NrgzdObsNQIZkNR2waTGE2afwt5Wz/8vS04AI0Sz
fE6wuwdC92wEQLcqNrOlE/ISve69s31sPLYuz/iqp49vcxe+TN3h8SsejS6RN1n0rWg+vul3weQ2
qLMCIx1laWjj7T70FokYjF+V1xzKoa01XTf3myfhBAytyWXeNA0X+R2xlYiYnelcM+bYNMlN4cMq
7hADKmJtURq8gXNAHq7WzOO0rXYdv0NlvAjlYsa4G2MmvF0VfoS+ISxhf/5u8109OaM4f8QJ1gHF
RNtuRwbIk0n6iEc1KZUDxJ2hrmHLzCwN1sQlYNdDc1d2glhqx0NgIXV323wtjrlMyvm9H3g5Of7Q
JeJibEoxVqY+0HSCO0j7oomsE7r9ZZ+tKm2C873WMei9QyiXmJUU0o1RpGLArZhQ/oFzt1eezhlW
zFWcTH27CWHio/KOkdu3qffT2wofVAYF/hkaH4hOQ5oDhbpyIFTP4lVQmCVCcq77WAqaxKBvcHRq
0n2gGTjSNAXicPpVybzfRyv/21Rq4yUd6m/LGwuj7c61DnJxCF6wtR3TmwBFA5rwVbT04OX1OyTK
VVMvoxUGZz+e6CAZCJ9T4ecEV3jsIFEW6fmosVRtx0pc/3iyqoiKZAzjr93mHHmPinY4XIry1bdi
PVDfLCn+Mv3VPJa/CLyq/ItH0HrMu8lOtRcPHz/OFTlkQcvrnXvM1wKaaNuhdXGLqgF3edHW8wJe
gWYplaldtUG9le4CY59OuwxAVAPbAzrtJi994lrjfIsvtn1DZo+rUwg2XQWMESKcLUka5AZ+hnxZ
rz5wxy8lgkpita+j+fAMfzFGI2PoBKrxJ89TvstRIJdNKXmDLf8r4mVIU3Y3OSx3IsVqOZTQWMrk
23uyNQCkJgDoE2Ytzh0yATQypxX+moI7rbfLioFHB8xsq9FL3tElUYZ/Z1SoLrxYh/raJP4iZuD+
Z8slP8e8U8PIt1PJvJJzB68cEtKYUt0BmBuYWo8X5dCPoHdGGS3WtMzHk8ZsDIiVFKJyvKmKjMGO
Wp1VJeeW6Mz423yEut4snUC4z8jr/KsMCY+kPeGxHKGXBIsfhv27b1ZnntUpiSiBamuA61RoSByU
M2FTP6Kq005RnfQOnrPf3KnjISKUdDO13eCGzw9XcVv10bjbSa2a5rWcusBNvOjvupPZmDMSDils
5OQdt8WAVnVtEnzq4FTjqlQCL0NEkpovaVxHq+4mdlboGIDPmbZmHe71JFqFQiiAolegjOBLyZfy
kCpcx8l0IxOqgp2F7Ek/13Y0uk+Gz1CGgXmLtAMbg0aBYslt6SnM9+g64t4+rc1t3tw3IgksOOTH
rKHgDzq1Y89o1wkgcWEGkElcLqXo8UCLOHa7rbP2PMGz5Kph8mnP8ETWPXF6u3vAwRKLRGmj7LCx
IJz/GghS91SM/lzTNgq6L5QKkGPolt8XUN3PIO2taFeN8ZpQuWLEZNL8Hsa1BhcAWDhN5ZGTeYAc
RNXQ9XoWxbVZVe12m1Y9iVYQRDsZcOYYeZwC5IBHKFIeksGobRf824/UX33rLV3huG0luwiiWYEI
mK+nwZES15Tih3Qph3iFYUS1rXmlGXoZuPCP8e6LMGBw6SP5YDDxbYitkTw/b08kqd7W8jTx9zo/
tRZo5N4zLCgbPOLYLrVtqS/UuSCECeBin2QJYTWYNa3WqnHd9xvBk5YjvoJ79TjWeouxDZgBH2gP
fIeBHRZ+conbXw1TtHFgWIS5LSJOJu580lVNU/ylIBp9p/idzSGVqW5Mv67oD8tNIgIzLEVhiZjt
MAG7pzuuTxnqzO+NchfWR9juOW1FR1Os9RVSaJPv5Xtpt/60ESSa4Dn7d4yNmg0GeAcJfbPDnwlb
2R/2EcrcBdrmU5XzvF/YrUz2Vr2JC8B6aYFJ2S473iOuhh/nC8F++pLwwcMjPWhwv8sByuxJIDkZ
8kDobZcoZ92dzkdD5zRsZBNn/kNhJIvTnPnLSm9KCDIdLwIN9/sF9Co8g5WKkfOKbyP/FNGHfPxJ
ReO0p/KBvIqpJYN033oLHlTO3iG5XOGc9MwIoZJDU4jbQEEgJiAlyuqJfV29ntDe53x6y7zByOk3
pRKc+qeYrKqNogZJRUYK9qrt3R+omrIc7DiKW7q9Fw+9GE4OCup9o82XEdqJokjFz5BBxR+lgehs
4Kxt/g3Eyf+oWada5VvDfVdjDLwOKtCGYLU+b19ZXQOWgyRS6MvKgbqShZbU3tiAqbvhL/8WQKB9
cds6Fwyz1QhQAkTyoTnoWnxmux/Ih7rjndezQ/skQ/3e165XIykq55CuK3S1Tp3wiyqc8T+e94bR
8JY5xC7xlkjStu9FcM4qBsJwrOkBblF5dShQ87zyDoyMYzUDWRL4GZTMCD6/vDBqFI1RNJVBGa2V
6WK926QCi2lOW/MuHLCgDIN/rpZFToMoKOQTPhXzIrHh+6Rad/HtYVxMCNO94xgE5Z6ZgodqARyW
WUWy8D9wP18OZU/Qx4U3a3Nkgv+ir341i48Nu3snO/X8yJ3IT3Q6SwtDHa1cp9WJA7EvM0sCMCxa
NSewOaKAXU6DpCPaRpRIVOSa55lh+gfXxAxaPTijZa735cWNV+Y3COIf+HWESI+egATW7uLJA57l
/zEiZ/5ho0nmbGe3a1k88JGikc8GNNP1y6HzSZX4cesjAAeERqKB5KuVMZG6SuwQ2GegLm/ttF6a
BGMs+/hEP3JUhyDUCpiQ3COFQ3limZ08rkz95akUVQtM0XYvTJzTxmTth3Qw1L1JTlb2mFP4L5J0
4Zvj73436e9vt1MnLba+QDngFC4mEXNXa4sUlfzjuiraKfstjCB1vqQ5827/1Bj4Z22ds1nsPSr2
Usce71pDDi8MORs+YQ/62CMg3RVUD16ASWF2eNpRPbiavMs4j2in/iApyFmSnooSBqujDe7fQSaQ
0YKZuZnMQQgdxTVvHoMyfpLmcVRdBMrAMJ9ehzpGmGoGbmsPAcwSGHvpPrvsGvWNT5YnlRTtoraK
ble0EeHU1OgHPiz4jP+cHmIEUCk5KKL2YeB4zPZuQkU6GS3IGJU/wctOuPMdXvo7WkENhJ//c2ML
oNQuUQKm5J6wOS7N60CoZusAao8dL9oYCK+Fx0TK65KwhYIL+zZ00HAks2Kkrr/eOFAix5Xd5JXr
FVnlqqWIRPn0p3omoYY8DpnX7hIF3uG+fN1zSYcxL16EceURzePHEIdeUPCoBFkCTZUiRCgAU0ff
Rs6GY/oeF7w2OXN+pw16xgjiofYZq7oLXP4cvJbCFfgOZyUhKVAjDNi24n8FliwFn9Yn4Vdfv8Ry
rQ9gLTeo8fYruK0ZUNkaOksdZcjTz34h3/R+O6+OpCDQ6g1RDgv4kfY48EZNUNYf4ghmqClFFOKR
im/AzSI3ghXV1CEAiis2z+l/jjNE2HVdK20V7RT+KRPYNpcIKkx1SXgaWLCn0EzwBRmidJRQlUap
YWiS8q0RcVlOjae+tZEZb5g/K77Op7PsYlXlzUEUeoi6rfPA+IFlcNKW9yOMeaWhUHxcEQ2AVNCG
ULEXn8kPLrlAwQlJFtpVLNbe20w41hgVmLwyHkA267y/xwijigcGqe2fTcdaH6jOpuvH3G7E3GMM
J52EdxoFtiC0pozfNT3S2dyj1MlOf5It8cHNxPoHuWbqosYWmvX1Xh9dVnXPrCqfI66hvBXtoNZF
4Pde8EFu1pWOs2oeBkm2mZtAbpkLifCgt3xtswoPpAeO9eRJKPsDjb9SqOwhQ1+pi/PWgdBM59nh
v+X4Jtn2CwwjRDdSOjDQVpMdmOBMBtmnum/UuCe70F5hqNBWeDyPgJrlP8Z6m4r+viINimdsEiVZ
A682mj/6wkonxVpiEo8ORlL4lya4A8hFOgjueQgmsTUXGHfRKzzK/lMuPq8wrfHkGyKWgWjQ+I6C
SzvZsriEVj2jQgRSMsfWGmDAjm2IQG+IkpQpaGLzL+bj/8oZtWVR2rbMTAXk8G04DWFJbZDJb7q8
rEO8zH2QiZCYQj3ADiF23uPsCXCl5LOI2nmz7EjZeL5E42CRvhHu4C5ZrQ5B6UzlX5M8+zVPlUpw
kv0jbcPj1+JQ81P3yawSRLnrCi+7UMmZfmzhP0Udu78tnCaHlq/m1ZJSMTpGxCzcLuJYH5wedpnK
aJGe/SFuwUOFFEyMxHv+0VMWC7z2TNysybuGU2Lpc05rD8q96zrjXi/DHgvBbyj8k3/LddLjAmWy
3CLl9EScZENPVyeoaRyIK35dgN3t1utzfvJE9YB8nonYkwp4P1iaA1GxTxhHlx9kWgyS5VmPmiHj
+X4243XYvfOXA8nlUDELHGx5QigdTUm/yycCNTqIxkONbQwg3KFYuR2sPwrn6vPax9wVOO0Sc64t
1Wi/yKJ5Bem3scuC8b35SVw5ifizyRJN9UQF61ARoj8t0Z+LLHFplcyC1QCIS5jGjVAyhIlWF9W9
4b2d6MQiIKTOdp7jFMrMKooVdqKqK9E8YWngJhV5Fm28xm4hf+Ea/p0mIdk5c5ww4e8or9NUWHS6
qulg3Ly5JtUj+6WY56zrHdwji2APq4dTazCAyxgI9X98vZlSqCl5crEszQ2m+Vwy9OESLSVpx9G2
ksXDbLkvIVFOnIy25ukB0qrWjcFcXemkRxxEOZQGAaNLWKoYMSKwtcCo8mXeEKq2wcQxWteciAUp
P6R4L3bT0HNaTKWn7JzZHAMzP4E6gyPcRMJ0WwSb2yRflOS/ZHF2u1pISKv2W04BOFLdlkIkvgn0
yEHHKzFGck4rsIxss7dmImC9+1L3DwTqjLU4nPOsGIWWy3+SjailwhBEsovLYKQm/u/vlzU58j+n
I5vIImK7KjpxLaoc3uTPvMsxEkF5dtj/rrHYo0lwyrUDq6QOZjXJtUEd0ZV2QHPFs66RIUoYdhJf
0wdmkUin6Ij7LEActRITwYSiPmQx9RFcgG7aXaZzxg4+xzOhTuscASgs5C8KZkUMfIOVlJmkI8LA
MlmWS8yZ9/TbStKo+pyH6PPDLEgd8RYZFUWxevUun+6KnM0CCMiHwNjzqg9JgvHiaRcSgVCAiLnZ
APnwafymZEoqPf94UUD/kBl6EpndMXZyxAFKHDAlBdbIO48BQFj4AB75+5vvgxgNfqDzgHvIZ267
oEOk38jCr8GAMefNTiGH2fvayPYIQOqoaOMLhaIknPOT62at2pDoOsvi4yesLkSdHTxSI83VEBRY
DIGv5TePAnbeFv7qQRUVKQwGS4IfOoWoo8r0iSVjLNURh1re9ser4D/Bsc/zvbI9UZWDew2xxlTV
fxxqhSRThH3MN/QrD3w6WIki0paELpjNSPg4Do+sO0EH/NgttD/rdD04xPe3itokjwVEoeAeNN9W
SiNa8AWdEVADfZLHHue0OAxVwkAlYzQckz/UR5VBJPoU4C/oObWDV8KJoxIm4aD3VPprJV8G+mRD
3STtGWtidDQZ2ZAt75HGadXOakjZgyw3wP9zOlJLOVjzDEJyl4hQeMJ1CqPCvEosEYi3j8r+fS0v
l1IAjfbs/IR0hHLKXj13cm9F+V3pWup50ym4yu/r0hr6Xc3lqEyaHrOUCOmTymb814iWuatQUR8A
17SIkx3jesxuKzneX+clv8p+MmSaMz8KSGELDbhV6Aq5OYjKjmy0xhIPETuLgLCEdOCv9rZhuLHs
iGb4Iuz/eXn5DXwj8V6f1VNfgSQ9hN7HKDmYSYoHpY0bJLbti9ESZtsZQO1rbID/3lMKyf9dzkX4
TRtpaC3WXgD9nmnyqcyiI3iTIGT0f47Gmhp1svB9czsL21f4vGcWk+qPz5ndKshLzCYBZXM64/6h
3zKJacrW8snA3LL2Snx3uHIP3tjwVkpatSJUKpf6gXt6ZxnJCrITGIuMXFThqP6j8GaMHRDU1Y11
q9N4XeT+JKvRdw66lZQuKzi3hbjsT32p4jjA3LtqZ8ncvD6ttRm5lcEwkzJM6LNtsZ34x1DH51an
+tmOr4KrEBniPgrb9VRv75Y9kyKmV3ZUVZbjWinWIch5jOFkCRLc8NuKgaChUTUTvvjtE6PGi2fG
9CQ5IUhB0CmSjQID+5fuVBDRvO4bdFe/7s4s2SkxWi9Pr/jMGBKvwqoLUMh0KVo1e5oG0trZyKmJ
o8pvwddMatxFPKjpHZWJZgMcoN4yAFEsBSVqbQGpKnmEvV0XJQ77oRUUuqtqx1p2cXfIGiLemowT
o07GYs73Z6qxR8SJwRbHjP6qt6llYaIdo4upsLJtqXNBs/1Yf7Pdn0SHUBgvLhPEBQjXjl28WoU7
ctfrLccfhOrwc2u0GmQcCY1kgwkjinvvjBtltbtkevV+v03J2KsYOdfTRAqL7qRc/5i7J4SA/qDo
5q+eZzfbCfrqXBZe3EK40sRT4aXkRFzR0Zvyt6LukRlKR10IFTTorMZ2+KPZ1jROaHncG/XLx/63
rmfdKjgTfjxsfXv56lLR73SXZ322CLjvCjH+lVdFOBBmTQQcagMvXtkaF7nsL4AiisLUMSaGhdj1
S3jRNmmZRUhKYmZ3G2qPmUAIuMXE+A8bx3j4Aa+2dEq3HA22Uh3SiQd0FlRbNZYJzF3qKyUvPsNr
eSxCGXWjtedVZDF2T7zvUQTQg5N/uCYQC2GQN5TXbSlJd5QLFDXX41X93BhMOgSAPeo09LD02LDd
0Xge5C/MoYkMu1ZqD3AJumdGfQvTuLfLCCgK0zel/0Cqx9ShxrufrQck5rqJmaxiCQF8JS8c7EDH
LNOeYy9hcSTpJHmd+EnwrrKmg9BRzyMB+oAoSj6RlNzlhVqijovkSJ/2aGvDKh57vNTGPrYylBK5
pkRcabQhZ8ZcM2ZcweccLTlYdtIEThbKtUxq7E8/EXj2Y6k37S6hx6aus4jlevPkqjFgMaEUXMt5
mnxcZwDZi9OhZksj8cPO93Koa9JlePt7EAu7mWyzX1qDCG9gOdfsTCrzvZhvnPpcb9Adf1aRcXrX
/YfkrP0Y3/cB+0J3SKj2zlPoNu5Otp+myfzqWpJTcI1ceA3ziZVunibxSni4T/ClRkT6ocBhoEYV
suT4lefKccbj/LyXXhvKjmW68l+EqLPJOjJL/7o9xniC2npoMMzz4Nl0JhYp7LgmL+8Au/ivSLhE
MaxoxCHY9srjYefvbXYCIltdhwDTiHLYBp/frPQ2MZi6RaJ3JglvwcasGPVGLWQe2D3hDghYjvTX
itbeBj/l+t55+J+JgQ5DsMPO5G7ViMe1fflU9L+ZzPklYDeA2+RGjgramDkEERAEROXX4Dd7wwDL
aArWBIw0iPTue7TcaPXtnCydkc+pUXlotN3NaMummZfF891xPbT240Rd+P+imYFAgXqPMgDqve5L
WztY36Dj9+76ED73tD883hSNcaWrUUup4emb2im51bzFGlyACZT2wZA7lgP9A8w77pbXcMMe8VVO
IRUsab9p2Ld4HE0Hqn9KiZOlHDSwx1RMzJbbJctgGVMgKl5YssDBWh0Dumj+xMtQ32mC40Z2H7yH
IJmPNrpuRsrjQzXiFi/J4a86O8npnzt7/FYYV5hFF864PDo3NmMryh4N6j3xJUH4ErRLqwq1t1Xa
XREkci1XSSxKhzvD1p6EXH4J1beK660ibCSXLlmAVen0dB0Uu/mvGq8ov+NRgAhlET2DV70AYCIb
w6/EXtH7YoI6pZpvE4/bUtpP66/pifuIbiOcevPw3Dx4YS6e9FmK7TuHdqUGGCgXO5mjT6Mk7vNH
oa1oiP1K2saCxMxMvAnmz7Dh0pivbTsrRzF/KIrIQ1I/FI64yZloUqz4rG8JvlZ0FXxaIwDpRQSx
SiJwoGdrWp2Xjj2h7Eg5yo3cUR/HPpsXPQIDYaPsIT19Vc6gjXTUk3dWnZLS3QTv8jIOuLr+7sD7
xEGvDXXXWwOxwRd7nUgLomgYa6xrg2RwwoUy3ljOswbL0cqGKSvrUYKUix1Y86AMcJG9jpHtmuYI
oRXSKYc4w63o426Iupi95C2k0kMasLj8kRfdYS9r47VtR9DDxDyMKhhS++Hl7TPgzlwcs2osHOPQ
y4IPkHbykk9LyzMjRzZ3MWJCsD9CTsHw3liUfImZiOiUQyyEq7CQQYl8I+/5cD8yq4QdEKt2HOBt
PuaqMrhiffnDbT4OAN3gRmADRa/nWXzySyCcM9FyDjVevnQSZzj7bJLQh/OWT8d8vuAt1SAcY0Iz
88hWlKzuzWPBS2F3w6tVJwiNbhI7dufeZu8W3ocadZmKnNolfEf3LbW8oD2JenlOqSraKMedeSZL
3e59RxW3ZJ+Ey7uL5cDYDU+DyLJ5DPTBUW6AzYHKt6XwrkikEaTxKp3ctDy5zXJ2GWZiqXSBCqye
UJveJ6G1fCTnQ+K+wLfp2FoAvbNNzbK4VFKPR+sp16Bmfwc3NgaD8qMrMZsbmHYwPFUYAYGlO7JS
915iUbZFVEWbpbsjVIZDvz4lRm2Ur+RdO1k9pYXssy8+RD/K6n7Hc2o3xCNUDaSnXS+hsuEI2Jnx
UXd7QtcU68VTyVV4MAhllYNeZe12RAaiLkXXqJHlsq7cKYYBplyr4BjWuzmKC6FYwosvCjxklK/P
IneYwMmScn9s9WGhkfBhooASlgfaibSaT6Sgprr2RKZyFKqBvmKKDB0cy9pozQGGoYlIolqzRiIg
sYJ1hAV9zRVIU8uqEvV4ayR34ZPTrGIApwUgsnG4eWnRLvdfvVEgJncDroDuFBM8r2D8XKB+G3Vg
8/dNfKGKTj0SOJx87gRLp8JSSyMUHXo8I7JzVcDuIprbWc8uFy65AxxIzQqAODwdyOGm+7E0XdU/
1pzaxTWtQ3+jIsTMEjrRHFCEkbtxzM/iK6qrxlorcPgfj4vLRaWe2hcScS4EKVnc9j/sBGrxMI0q
NBfdWqPuFftVbCTqf2XVxj2IJ20IKjEZA2DuUVl186MDltx1TytNR/OWvmnuL0LjfFCWXAT+Lsny
TTpcic/hAd2vla/8o/cLE3QhQnYUNX6PeCaoenjzMPEr1O5XVA0Bx5c8sRfgMCWhE2h765StCYLl
cjxeaTI53Pqydf1kUl3SwEhDslOHJNz1QioQzMUbuNKP8gdZNzfvnyXuF05WPebi4r1iHJAO8MtE
tHvY75h95tewjrxFMPYSgBMA9lPcUrrnSUywSx+xmh3Taj7ct8E1S5D7I8UAqkM7xfuIkaQmvbgW
RcNPZCa/QA/nFz7/dIYpewprH2wxutV9kmPA3nanUQi5wjBX3o0o6sgg+0kjDZXdWtDjnUp1MELx
CNkX+1Wl1UQn3KOWkpgEwiGs3W7Co9jYpebdPI2IVlKAEABM+elFdA4CFTKpQ5ZqosszXU4UBPoO
uRhQSlXdHiCagdxjR5/6crwdzfVmv7c/dWDrpVp819b9aURf0sVbHV+XZOZDme8p2Rhe9IuJ33Xb
9uviTKvMN7P9KALIqcr85qQAeYeC5fid+J3t0qsSegyWrXdiXeFK5dCg7zIt6PKNjBpnKT7J4UdN
oN2GV4PFwf5hI8AL7sFaAcIsUxzP4Taj9Ggi3GCah0+HYVrQNOK8pIUKv9e+Hjm+xgjpl2W1lVMf
aBfsC8To/hCN/94hZuaklH8ZpX2zBtwZEBwAyaKe2flOtWtINSNKugjXmmZozCfl17q6BoGyjSb/
f1QvLDgRWZg2SQChxiog0FyhMHAMdpAVxaPXAt1oWwyGFza2/D0ow3QlOf1vhAtxj2x21xjuS2A6
q42i3Fd2G4D2Ztfk7OIodx4CVLPTKklrwuCgIoIM1hwon6z5WsffRPty7hQ03tjofi0gd8J4g8UW
8wAEVngD1ljheWcJJv/3eM6oOhX+g/2xFtRvN/GFya1Y6hnJcbLYVKQS9p92lLk/snzYBSZVhojT
UkPrOhiyql/1XseyPM9Sc0CvO9VJovOk0+tqWwP9Cgde7qevAKgTU7QeJfG8mY/EUmnzex9i4hPP
4mxMcSrZ5N2GbStp9C8nEKGPdw4LeOYDMmiLEe9uvNQyr1JvU3+MRQXTeuQDujN/8xgx1lYWiZ6q
x7kNnzSnrZl3cr8oPWCefoUZDVYXMxIUkwi7abew4jh3OpacUY77xrgoNL5k14tzV0kRd2zLdS0e
VTq4jKof8fb86M5mGEOwtKvy8BIXaexHjSaUnhXy9LwM/4kS1mQCM7BpsGnv3/UM88nViXkN59uU
0NFM0kc8wwOem5qlr/zPt52Uq+lxhPieeq32seQjl0/MZXOccZ4b35o1ibH7CpbduxShriiGfOoi
jNwWdRgYUaAMjs+bUY6u3r39Izqgn+nDuWq91fQ2BEng+ed0XtRi4j5FJiCSrqjiZjLAshiqLLkL
7elJ6WtFVsSHW9tlPZQzwzPz+lnwfjDBJxVPHyZRxmKHKYnpwFB4tiGIWVlNBUZmh66yxSktKaWC
AxaSidORjVIn9HyM0JHGtiNkpvsPreR2Ru0zpyBlsNCRXf3uJ7ui2cY1YO+Sd7yDUzq/Cluj0Wtk
FaGCxFoJhKl0GbO/NfR4D++odIr8RmUK/Jsy61YOoZ8t8943uzs3FJLVdAUTnGer9kBFZYLGxAIZ
4B2ooLRphV3OY+YR0g+40UNknz2B25YCj9EGhczwTiPdSoRvFLNXeI557wXHdHCmbB+nNtObGSVw
XD1wOn7Gy3kXRFhQ/uVMbI1kdrvoH7MJcuPnuuiOYsnxH9RDrFVqPU1qZwjMzzHcfLo03lApQWZk
Ja2+o9SWGBNUCYqQy3iCUW55oGabzrD45x3Dv/8SVjuGv/gvDkOxtiR+qWy5nahRRF423k2rX3+F
3vpebucbG7PH1eXg2YJj59oJjKS/6zaTNEKvxfQNPbZTTVRECGT+gbqX43mcHvlcZcWEZguLYQLc
Ac0Z0LKvQfQB/6Oh+Pya0tzMOehIbMAvVPLsDpQ7FeTJZW10fZuEaYCq29g7rIJke/XNEa5uSsyn
S+sgMZOQbFfFT+jcvh5CjMD59nrVhY0EYfKYta9w2G+Z9DQap4s0ckbJahQVudbQkVLmX6YhSX+4
NfR5DD5eJKV2Pxowcbs1A5eatt5FGLFDsUVPl9cKVvYRQlRS7ZPjWjnkvYgp+fIT10ZVafIKz6ob
90pq9oFluLkbjOT87eXvVqSr33fESfDm7JkYR5TYInAecHOOoj+Y2cDmQc9x0yaWgVSr8kfyAw28
KGfngYiJvJy0ZjPmXse4MY/5F7XyBkDabrIAQ1nsejyptCUAweIajCRvfdLoIQY3kYtXIEEd80La
jGNUKodn+UrqiorA2dlLbGmjCrhsK6XStOjn8i01hEsRUsF2+PdsfuvMuORuer2uP9Q3ckXiN0RL
YkT7Q+sFwam0yWn3R2Ntrummsnneoh9P8wq3uaQhKZGtaud/IqT1oTJwlShxCsIa/PR6HTiVo/S8
CCAiXsAz9SW/JA7GWTTl0ND5mg3yHR+iPY/MIKW3csPhlcGgnR6XstirmAFgwk7r85gMtLXJQl9/
ucKBTtzDMcCXExuPrvQ4goRpbOpsEc+kAor5nmm1KGHyD+vRNZvKtULEFQrMX6ZRJwhWBhXMwXOV
DdeSQzm5JEbxOcnEa62SNjZ7BTdSnNPHrosaL5+ayvdVRvlEPXIkNtjd9HCu0lW9FH8MxjjrXcUX
tTbTNrt75s+6OIOjUPFr/MRHUtJNTnm/eTPiAJPLdBimbjBKtXaUK9Ja1f7s0YwBLpPUXvATspuq
htH0qwd1YDgYGX0/AGTiagZxKti6Z9SbnFKvbEHI5HGw9din7ZIA8wk7YLoUjjAHjF1g1kO3xmEE
CSchhQUgfpiq0iz107f6UP0joWXQtzcaAfB6pRuOLbIkf2LQSxUd/Uk3z2W6cegl1hiWJlBSk5Dd
9uNzJQArKoutk5i/j+icIS1hxIXBtGEMHHXLqsjtCGjoOos9edjhetBgwVsxYPpBgAaKrxO8kLvs
Rxo85kS59lM6JaCUrgB6/WydNJr6fXMkHCs1p3ay+MFTKPd1AmfoDFj9kWDG9eOb+SULtTLXWtKQ
OfhlSL9ZzJWQ2F3HJeqglGuOUTpPNi8xweWdkk5fsHNuZeYH3dDQFadGjVG0oT3+nPhBZEeIUmMi
iVff6hPRTFI3P5uzX6xP7dB7vB0DAQC7vjjRdKHv/ta4xy8I0k+9mDYCSXGmE/e1SLeBqa7eFZBZ
rMiYCUOFNjrF3G/JMchjcP1MXZbig9R5WyMiKW2Wf6JzdpXuXAAsZE43L9zJ0ZujQy9914iKKZRq
LV9m6UpytaiwTDyQaRbWnEUZsMiSqhSns2CwPNeUus2EOHUtfB2U8rax/mHLGMJjblPTXaK16vgL
Q703jXT5Un4r0yhfFOpZO6rLmDjsa8nAOAzlfKV3H7kj1OvQ9kv4NhfCfCXCrJ6AX9UHDLz6sk1W
wppKCAl9SWV/T3aCe1KC90bdu/KJqfPPG0sXJd0cE+km1mt44274FWnKZ54rNNwmHCcxn355SQHM
bLjowFMpEA9LNQm1CenrQVB8BowBMmB/yUoqSf5Qnl64iFdqQgzndkvL+CKamgkEha3gRkRZ/8Ur
wc5z1lvHsjSKAXuS2xLETAprw3y0mx90riAmYz779yS2/IZgBj+RrAYam83Nd+axBuWuwxho6FOa
M0qvE6UciBr072jP7to5m/4ELj7zfVr0AUCkR6zpd3tvD6R80BDuRXDTGb1VE6SQcxoR7BmIE/3v
cuYxFLapsFDMy5BMWXHX15zX2Gvf9VTemn3jntSIBguGetNTjHbLLRFI004UejB3QnMdTT9lT5SK
slpq3Ahl2BVUGIdIk759iV94JdnjWJkePFA3IIA2J1cYRKJthNQ4wGA8CI8U0IizFYt33FBMTU4n
mAv7YrRgPWusdoGxaIC1DIXnQj6777mnxYsh75b8WsmWxrCgVEiSo6r8Qzd1KQIq0F7tDSA/8Oog
xYGk9HQsL7GIcUubFI6vN6wnEJdG0w2M8/rGDFIe+gfXoqdWfyZ/tONPPfBgSxWssP6p28nKZPKU
Hmw1ud5PG84kdj6KCXZ29w8xdq1/jR63oMDtaNRA3fBZGxsoZ2Vby13eD1hH6A7TDY/Au8QQb6Ar
37vLEfom+iQcIEnNKMPJZREbXAecWLOgI6rTByB1+CVF/rcEwaQtuwezmD1k9Nf/hDzf9tCkN5Vj
mWLHJjipwDRiABOX11yXaGcPFfEmf0sL+vJ7MXJCq4yIUPR+OcsOQB0BhfZfPgQvptAvBlRNRx4c
pDxTIYwWwERQhRD2mLwhxSuXEHV9IC2RtQQ7AVQM/nW8wVIVjE23l/6Ugh/u7xaJc2LkYLV7ekOp
6xkoj/G6ZnaGP0VPLdvgL8QDwBf+5HXzvsTfd+31v2ECycqKtezLaHHgVtx9KAOUBNWMffPAv90L
0upDCHxGSLA9tznA8Aq4TgxP+BXR9zotGfWtRnPlKWpu4AN2GYGCZcoAHCDsXDnrovxgbktZHstV
m/QpkaKDzlQvrAoqL5fOnee3/sbDMgjT4gt3xqNejG4oGZSuUjMYChWZ3nUFyFUXc/5DBLpnqdHF
nB9CdVfI5K2hEaL+zAL5kerSwxj3FH3FpcsABaf1Pqd1b0yG1hIaFQdEHmWccl00ZKu4TH4CMwuD
mu3bKZzvei41YP745AhuPQWzUsyHR7AZQYNFdJw5qzXsWsh3sX9WQvzS57lcscM88dqIdTb21huu
ReBhGW/9CZKKblc/aZv3cuYcpQuZa9+7DkjMt1YcefTI4N2EcvwKmsP1JGIE7ho/3r28ITNxCk/4
Sj687joK7IOCZDmai3/GtbIhDTNn46kkHTOM8jIAgEn9z0rsJ8EK+KalEzr+PqC0pR0YUxyxepIG
rXjXBPtIQkVkHAi2JtcTfQFZTHKLIwpJaExT5itfXMayBr7aQgbrmqWFiOcUB7QLWPWx1aFHBXLI
EwM6aiKmJ9KPPrZJtnQFZRG95JE6ImcVRBscJaCrL2tNL2KjQgRvGtXgLTgGEIffRRyyNj3/Gfas
BKXgWEjqTVHxdOlHjQw3pLijOuoIO8sgiq5+kPXwRM7BPeNWsN75VIRO3bHqkxWHai3818Y6nUD6
wBAVUTMXcLg3BnbUvTojlHlWc02dII+hnmgUJPQGVoacVTfAl0U3ldyEcw3RjNUMphFf73pF0ELA
VueLC4tTkLLT7baj1O7JgJQo2KDaUPVhLARGIxOlUttauXM1ZyFL1TVgLRwt534ShGK+4QrDhH8B
3milUZIeeZCO+qQg6vZ09Y5IPgm82wMMnjKb3jqpQ/jrUBcz95QLyzkss7fb1zr9vYZNY+fKU3Vz
WQvrx5V3ZKrWyZBft6iqJibce014kF5o1T/WsFQNcj9ZPcWhjkdmyHUcIrBzFdTs4OUdrbs2qIV7
nn+AbNa2KIXpgZ1WucCoezroCBaD77Uml11qSK5fLfowKzDXwYTXCiR0LYUg+4WbpN+kltaAZY8S
CZ0fq2kB0ZVOy/EDBQyLdBlchY0vp0GhdNVpS8TWAvqc4JvvmjuY8Mp7iDv3r7pBe2+7ZLwjCT6c
rNOZ9ZPH/s67mJgH00kO8+AB3yoGYaODkFrAXa0W3czcRgLUIcLTNo/R3DpoUGyz5gc+Jvf5U/Ox
uBtbHEb65pZRPRjWkQ2dewtctVsC/DQQl/reG1/URg/VjZ5Fa5AqWLVwIo25QUYF+frV5wBGFkgl
CGwHvUb9WCoAOAp7yMFf4EiID+txY8CJiMBhp/bCXBzY9Z4dWFrvO4b80Sewl2eAcPzDS2cN9s/m
KXUHYO5u2ZlECTWevyAH735x0sgY0TKvRQPfxQ1rNWQG0lrp6Brfo2T7nrOimo1W09XXJ4w6/kaO
IU9FOoTGTjARSUQfCUMKEq/iZBVbdpDLq/0eDKsJ0zAuH3JnHS8nwqKMNSIG9vOnguqBIgXffdRU
CHcxoE4gG7ODp/VHiUpwxF6Z/tnGeFy+lG0hzUQpkKRoJ+FFLua79ltYSoN8yoVLSSorjoG+F6Li
mMvL6zMYFbiQZlbaMR0IXTbzFEa27LSGBxReIpDEEYnueP+5seHlCfJwisVJmrtJ4lRnzWJ+7T8x
NBTiMoKSMS78jISCdbbcY42qAOzJxEBBH+0AVYOgAmUnhyoanjElICO9D7Jxk26YP35M99GzCu0A
yoFBFatjL0nXSljDqmardD5hAQyH5bTWpOonYuiGDggYwDDaJU1x+e0dGoaSTxWhmKGIhYGdERnI
NayX4+9NjaitwyjXxaNOxBTbjy6YE9eFL4V6StfnWIvyjJo1AqBrV8oWH3fQQPen5ei7hCcmbku4
cPrFK9K37rE7lu4gN2QmkbLvC2eNrYPBb4A17LFkKt5c/A6xSLl1/anSQu2N1j6iPSX4c5p/a0s0
8uX5+12/EpnJqfqTFVSGK/i3/E0xIkT+tWuQfEImcnASNEWH8XxXgZ3Nv8cjJ4JNBeoAqfF71dtC
Cbj0oFJxbBhe4T8YU57LBMtQK9tGeqXvnJgTCsVO3FHEvK/2pC35SBZdcF3qJJ2zWZIE8sQDQXCG
bkw4bh8tsHABjB1q9o+ukl+Yaf96kRI5gEKU7xJ4JDCBVv9wySUf7Ju8ZD71dq+ijK+VOYtRJ7cj
VJT9FF7ePYT9j54CjdQJvmA8u+9dH+LGif1av1DnxGvBuHMwS9V6RXrM1QZeeCMyT4tLdL3EwhWE
/Lla80XM3S2MCD/fINBCzvrv3fMAxkSElzMJEqI2hUa717J6xhp1XFgMjqhxLAd6ktEmvamM8pxd
ITz6A99qiKV8hUZGFUFUz8zjy7emapeq2kZ0ytITRgLDmGm8cwEU/X++Bmp4fBEdB4OKFkI5DCBJ
WBPT42E3aXJkHFz5X2v244tOVkuQmDeOOS42jgfr1OaFW9S4OU5BbHGoExcaRkoIbAkiS4hNvAmT
VDSFucoSoHHOmhMjOFtlfgHd/a4iaAi5/mZyRySLb+i9PJnmRExi5JqQNjEz6cIUA0dN44ab/XQY
yWFyqaM1lrEcmBuXrHGZL5OeKFF3puF/NABVqbCJ6FIvUngMSbonwYIyhb5KAaCBnbGTmqiK04HP
FUZiBdzz/qqVcdzN6LbnFzJe1CZDDwVBJoQLNDk4+6j1vwATwtC+Km5/xyDyAf3/L72xbkIjGhnm
WFS/cACZOLAo5vMzOTtRH0gdOxPoZo0ufKJJvToK4kXXfPE5hITI+ps/koadnJ/9xYR7pfK6MGaD
z3SDxAUMj1DNwhb0K1qrQw3MjX3AtZuAjI/BljmX2KrfpCB7M0eFi4XMPFR2+v622UUhBeFsDhAW
KyGhFyRHv7lngHhKJzF6QyrNIyoFaikN2IBufREECFmTSz4IUE7M3L7J5AxzZVuIBkcNjklVo1y1
1mv57TKRQdMbsqA9y0xE7zB8p/ehi5Sh7WiSOO8yMBnosffG8qUgXqkvFvbiuzjGU9lSBgr+2bG8
gvmMtvJHQ8LOBRmHt/WSny/XpFPl5QmgHSlqFiMdbl6cISW6OQSG9Xevok3TmUP73cexvH1qOFkF
Lw0ZbmWeOiA7iYQneeehvXof05hmx4wLZUttZbjhokKfiVIWt5dj4MWNkqqpSjO/9rCER1mA0FDG
nHIZf2GBx7qqpyjuOEsMfcHKE/P0+z4fl7nrlJTXa2Ib7uuTUOcaulhOj113OtSiKParAAVnDmUq
3nyyrS8XMHBNrt2RjiU5OQoRk3MzB4hA8/cSl5tpfRMKNY7jQM+YNW0ljtik51MyhviMgc2aa+eX
lZX6h46IJJq0vwmEzCbljhJYekqIHxcaOku2CB5r+vfgTDMtsWhYgXgawhHFUomzEt1JdF6RCwUH
64tB80vHto9MfYI9t/exqLwbU0vnmWWJkQslE00zs5n2SdwYu+rlXjLYTlWTXk1A4ZbqWXnFkqMz
IvCD34Jc2VoMWA/OACLSTDYkduyWt3WMqH5y4RkQiufPSmnUF+hkhRnka8SbD7L7fdlIPhElBKa+
XHT2F+jOq5El6xRcFuHmVL254offdqEvc87myXzXQj6tynGO2UfeHi3JucI3vZhNjuvvhO6j7DKD
xMxY/pd5szoe4/R+GTonIgWAxbkUMu7yQMJA/Umkr1V5Zv7R4QaHIdf1bxgdolQ1ufCeMW8Q9hoN
hBP7JXEHWgyKLs779q4gFTIlT/glTJwk3Qi76dPT4QpKz9MnaRSIsf+07yw43SDB89oqV2evN8l4
jLsv9s0mAnLqD+gVIc3p3V+TZakb3YkfG5FRiTNxUZn+0gIkJbwiSRcWDvyI/4vqJhqDJu5P4VZI
7sd+z3GT408JybujTCPxyz33j7ktFaCAOmlMS0PrWqn2Sb5vcpWwhdTlHGpCLunB41JDVI3nLz43
SjYhBXLMMxB0Q36EqYZAeFGMzap+Hr6eHrv5V50YbxsaUPm4wgXHfxaMUWf/KuQEmlzbhZpJuwiC
QnMGBiUZ0bPxY3KVozA3mnIWEWnT6hj+X30abckLfKK6h2Asnq+ydQgM54gwybCi1MoXgC8n0JST
gGekUWJU3JmgTyxsBP/VQfBdaTsKwmZwV6xL3YjYYPLGy741WjSn8nhKBr/dbxKvk5klQ46eWN1/
VvhFTgWjclCpxZz0aaSalMjyw/7dZ1gaBzqWbJ93XIzCDypX08UdgTn3tmPyrw+Otot49h4rrX1Y
B3lQ7E3Jfa9lFLNnLf9i/l/sGLfum+9LzpAEoCB8Fg70GYIkSlvbfUNLp3CvA87OZcTuBBJ059nQ
DGwuiAAhvL/9N1+/+z+yZBC+PLsQMIHrQW9nodyvDo3uezcX3eIhU8UNEE1ZeyH0ASldGLzuLkmx
Z33UC9mpu2OunuyL7rR6bZUdNXnioKwYf43w04sbS7DP4F0Jg1x7dMNDEGHhEoqfrMefTqczx+w+
xOPSotTjHFoyI316MROwbxB9KMpoCNiCEyY40AYXAr4bWPEEb9IG2Oa6LjvHPsMcn6M4wefD4owo
0/QK8Ae5EmUZL+dOueaxMZkl0jD7WijN2i/hs1OpLEjcQxh+0E/QyX4lQ+AXfdSEmAKIrWkyGyZI
437uPoikh/P2K2ntFEheG6+c9X1zSvf1HoM+ejmA5HLs3WM0cPsb0rv6icUmHfwVpEn3OOdC0NHH
xegZcUgglFcDKUfJj4eA5BJw/3gV2enRMhEX4xsGITAo7vSNMb7HohLhwj+J5IFWcd/ZAZiAkN1u
Sta4BdRL8UVrlPAknBRFONJW2pg8tE00oYdhrMHSn4oCa61yVvWVLOsxuh10SSXGvyDrAaejAAoE
3zxTYTTGNhF83lIfdRrg9/KpaBx5BtPyCdCT9pvPR/5XwP7ENhgnO1cGCf7iWQSHkGSi45u4GKlE
e4ZzeDZqQp+/1E9Vevyn2tscdR0mizFYkAEGUknUyeqn7o0UXkveJizrVk/XHPPfUPmHtmryrBNS
c9GwNZ6VFDLLXpzZXyW74tKVtzJMlu0qCiEBxMKVFdhbcpi/5Hcqu8D13QXCa01WY1Uk2LzqFhf8
ymgEQ/Qf4cDBnVwtkAzV1wv59MACDPYXAU9Vbaack4FtJ5Fr8eGWOZboQqipCgqFbt3EJCzw4x07
SFfhofaTUpS69nP8b558jmE5MnuzIUokqn3kNsaM75qD15jr3LYckPoaqnh9/kehMesWlofq9FSt
0t4AeDNL6aLwdP4A6wK8fHLdXQyTcQ47A/32Woipmyw3lwPSTV7o2kL3cvDs341lrT9ylPwW6Qc1
E2JE6KXatbrT2kft85r3qiI3YaSpTBZZGBJgoK7M+gTr0fcCLRolMh+zIz2HjuMe1bxcVONywVm0
wFv1vrcSNZpJsKjDdw6ZXaC7xGP+Id7O+dsu99PAukMvzFM37SBef9IjzZPHhQJ/bBOcoGtwU7ul
pasV72lVf3htojMRVwHISfHZcmyBYuHeni8HJXhUA1F4IfD6i7hB7A690hlCvrHZepi3Hc1MxAA5
yolwp9YzeqHmpXW7m6yY1RztKfhPgQ4rA63ObMSrpAdF5qcl22wxWVlpx2f/9MK1s/r8FZT7pjet
X7hx+eNH1EjlKiHgnKV/s3buPCsU3dpcVP2HuYekal+zAxv5lOSPSqR3Ekdde+lhcehqLgLN+liU
1NioXSc70miMlWAu9f5VIq6TMIImeEAO1mPrUhYJl+QmsEgy0jElYSu285IWmZH90oO9w2J+I9kM
ctj6rCHyABlqx5ApYuVF3O4VF5Zo04TS0stiu97OryX/yBrC/l4w0TrBorrC+uF7KftUhWO9IN+w
UPYjJ5+KaqCnR3EcE/a97EOvZuKZHVwBuZJzyd3H56EijceybYVQPM/pPInu3t2l5F/VsvPvXHOV
Sl8NA59lJ6+NvJHU7JPVCmDUXH8kkaRf66oKBbKEjeJ8eCATc7RBeHOmMA53Ao/ofSmeguOhxVfw
u+qGk2y6tnBDiywsKlSVnRM+aZLp1/FRXheg7pt+3A8IZjLDqdC6jrMVRT7mM+/bWVJ3cUNKGg/p
abryJg0EUuz9el/1QXmFFvxPNWy9yFh7Uqc9w7jQp8LtPYb1nt3fd6PqIT7RZFX3DgL2SxQDCULp
6zv9KBhYxwjNablm5D7DVspSMXGNR3TvrrDS3VLCOoFN1M8yAmqi6R1uE3vpoCi4LEoeY3JpOfkm
wKWS3ifFJSUZ98d3d/6pW5vztQFYWjes3WVrZq46mkZPz6XlanaoxKvaJudWw348NBWw69HSeN72
fvJDa3KHIgVxSDIxGAWPCEBcDXwF8x7AvMHteTHpTEac4srl9cJFS1CLSJi66M2MgI1xWsorPZxa
z8um7GYZ8RqqqwO7LQ1wNgXbFXe/koz7Cp4aO6WxT/5tS+3gHze/JkwA1s/O2e48fsioS9fkbwnh
PzuO5SJ0TQLlUR8zOIzYbJFNn/PHkns9gEWsX8rVljtgENzlC4s2HH+nQOt20yrPe3CnVvYVN4Cr
RNfJz7kB5Jfea+I8IUntRIEsNRkV4IsNiWaUsr3JAkLCoT4EelLRFdu6pesvNITBceA74zJ64wVU
hlM1LvQVaJEmR6C2C31ZToJzVhLi/Unp3GohSpGXYuwTnxqN+3OxsoREu3hWlYK/m8rXGL/dhSMI
oo91J7kMG1BCB6zJOZGMP1d1hMOv1tezUuCXwnChibSUuI3ZujkyS6MBojweR7HkJNQaBbpsGAEQ
Jkw7WxbTN/iTW9m3XGg3lyoo6fsYukxQ15SLPOuEk+jd+4qi2vnkFhRe5KotHx5556A9DpzXpfdU
WIOloW5RWfImnCJ1U3pwTVVMZCzyU3FtpTPEVCMd792TmndXna6n+JQzmgGYWejCNkwIcLX0cW9y
LsebxN8YPuKtyBOePojF+WMvKrLBJLRCSaFe8UUBPBk3CkqqThly2o6v8yWcGf2WSZ7zoBdo0PDs
aG3rUafY488J6XEqvD5LOfCC6M//UncxE80Eg1FP8797MeHu++3irYFoP5+5/hFyjom+mgIuOYYb
rGeD8EfeM5gYzs6EtrTpp/DlKUwMfafMW9G+vEs3I43RBQbN0AddYyzN6yo9fAhHO/Vg1fmkpgEa
kIFpamGToS5hBi0gJxFlk2vigPSwJtg1OUq4WultXJYYwQheftEX8zLO1lIrcRjTtiN5dOStL7qC
D8Rp2VJyY4uIhCXV9LZ9OwX3Gda2nH1x2g3NUe/nLVVgXrZe4oC+KhUjv6sqisz0uVAYS2I1/Fyn
d4GVTTHDR/3qDVVVj6lYKcX2h9sjikaOZwhnBzUEZhu8Cry1OAB/dOmP9Y7ben2MD7Cb3XYCtJrQ
SQh8jT/m2/WKLzcwgH9nfE5KTXZeYWjGZXbPFmb8XygIjlHTUWsXiflCOA/UxF75P/R8gvcNFxTP
0vqmJ7GQ23uOq76per4j2TpUTn2ibmvdi9YabFYqzDuaR741ZFKB1byfCgWNiNuC2/vYiGjKk42f
3XSPtSq5L34b8LBkHp6k1fihrVix2r+t714gju2TT+hOtvHM+eE/OA9UwpqlNkfzwsMLeDnent7l
UDDVbSfIun/FP3Y4bZ6OMZRd2ETcwuaq57ljosOI0bTE/nE3FsrDdD1UFzATc/qzaIAb7LAoahPZ
vQJxZrDgtOsGdbGXd80Aeh6KjA3ERh19LgWJJjZamX1XoOJvtNeVAco6onz1QhbT+GiKQvBVXwRh
70D8pZM4pvQ5exXW0nZUiKJc+ul0iU3qz5CJT168wcg6PCfw/UC2r+8twNoKIINJidoYk4SbOPxO
5ubZWFx14reyb6xRWa5mIV2/NIIghLmsj68AWrM1v8o6V3203HYi9Y+eARyzc8Vsp7l9n5ynxJMT
Co0TFjUm5vwlZXMWffo/+gvGskCPrRbR4igJlK66KAxI8x4Nt335bmcVcQWQsAi/wXxZyc0X1r2U
7wIVISOO8EL3Tt++J2jCCJhhGLd6Reo83YJx02uFCOKfhFAp3RMVaphC4iumqRD/BM6xZNdHD3Ej
fQvoQ075TLQGOkjRMdFRCLqT08tsHSdTjXKV8SaTH5g72jvMyW/Le7XYbCN2smRm8HpVrwsse8I2
LPlKH9oq6godTSLShMNcfEA+bgbS2EEEeXwCBT9IKzBWlhjl1Eunh3FNg4g3XS3u75Fbbb8WCmmR
2uK4qgSpUwtCjd6hMrzCKx+mHRsl3aQJFiDBq3yLgUGlTPz5DTJAXfv3+fqP5mxt9Ju827GU/nIP
dWz28icu3q0hknR7JwohX2Gh0y00EP6CvfcURW3i6TI15Sea2Eqgm39GAXYusJpc5S1/DJwodr69
yM0nuSKO5PUVeTkGgm1EeGDCDXLOFMN+XKxKq/pXeFc9mBukZuoceqGEX+4MBEv7FZseGejE0+JL
zMsZj6XDWhyMbORr0XDsAqCrPRPowiIUUSKqW1CodncMtDBql8d5ZVItrm4Q7ImqtDTKaKxVUwAg
k+SbOOAxGuWpiLrqrz8G7pF6mxJyk8vQGi8+jS4GZdw0RacYFKF19+uxtUbM/8U2Ou3JluJfr8Tw
zMAsFw7hWUuze8WJhXRXOs7cgrOkXuLr//AJawwJSqm9a3hgNUXfkXJrHJEt9cQJAYgxpDgkp4sw
JJdfUNP+HxVM6WJh/K8WPwC6XgrVTdbS72+ahIpAgwCOPIMGuSAJv04U/CKNK7/w/mXpISWnYP8r
ccfARxu1qw9MVszgU0g2xFflKbJOT/XzAIBJhUEn3hQlluZsKwAnoDdDQNWGYTe1yfQIbRDjH/Uf
0B3DthxzxYlpAIJbH4Q2trYYXehdLjCAJenMlbOca84iswofWM3B65LNJLDyoGfSRaLq2sqclftC
yfCM0rX0tmQUxD/uYhqjZ8YsB1EtuVrKdSA3WUSmyhfoXRZhcKnVmjID57h0dbBPKIihZ4dwSutP
gI5LjJztR6ZpPRLvfBwODY5Ho6c8XDCy3glGENRgIDRLehNfkz5RfYx7kH2I2OuAmBAWmlmlxy+2
o5fo8d4PgTeEmlgPt0YffxFmFbXlmZvTUM8biEWDUOWOIy55/jaRT/uugzaNWnJNY3qYdjYqJjJA
MkQGNoZcDYyJW832kVri0iTuIVnaMGlv/iW3BrXNN6iclftTJ5DHaK6bSOi6/Qfzk6DkH3BOxl9z
/4K5B7+GygGzYiQuE3MGs8m7HHZj4R5zWtDGAolKcoC3iFHlzk5UBBksz/zI/ZD3pkP8Xf5MYKQW
dP4O0s3UXutMzJdrm3KvoxX2np9Msqhc40Y+ckoWnC1YYZqVZ3BEy8q+f1y6fRA/IMCadUrC6z+k
LJUyaC/u4Lcnkz42e56AIIqaPB5Lpe22GP9GLXRgfbksnBh6eqCAej21Re2J6spwnIFSZLtT1n30
j8W2JJV4M30z6aIdT8/G+jNprsMGPbeUroCc/0wQSPU02+w0u3E7XmKIse+IH9jgbtZdFQ27D5r6
V9x50p0OTnzSbCfbfUgX+fQ3DyJbYQhdOpB425Bcy/BCfTZ2qHHartLGvNscdK0eU1JCynphMfs2
bkqYEeQrz0Xq73Tg7KWEis4niQWPwqxYxHrA7jLrIuAK5LdLRVVDBVSHASE+5hH5gVVovVixvviz
p9c/ItxtCgiepdGJTPC/HiBW1KVPo8pbYxkuJ1jd/UeuXlkjlZAd1Od9iVQrWW0L/QOtw3R4pbjL
a+MuDPhsWFxNsyQJn44T0x6LLdQVtVn+8ZxBEWG7lBqvxOotqcP8/HtVESTrKBXV6Xn+EFYrghyE
SdxVU+BepZ5TlpdyhDiv/Ashn2QGOUtQ97uJa4eCbuCEfQEydzATiWueRexZKivoiqzSadLBmMn6
b+8apFHyl+g8ISLvaaRSwzrCs/JIdUGe7S6QZFwd1JAKpGMqyVioWTYt1to0GMvaWJGrhnatlqsi
s5aeNM52X/+gxz1qnG1qAF2hlr3a4BYt/p6qriaAOU1NY32SkBRLLJpkWduKmq3JpfDlM72s4lkW
PO26zB3CAftACEJxwB2WHwUGo/R42h5VavN+kWK4pKTio0EwSWoGHax+PSLmt4i95LKBwtrZjC5Z
cjz5AGsncSzXsl2mDErLvMnR1uai77iz/x8+0x7HehZbmUYkc22kxFlRm5LSU5l8Zmpv29UNmNfs
cQqRwlZNjEYru/5fXMRlfNlFwEVNf62DSKx42aRrvtCDiKBfLoBQEY0uw/lrfCzxuUl0QlIiHyQK
rF2y3DNcjtNaI5e1TQvYogjxyXbiOZCNac9bJE+pmjccggxWnGhCDlTqQolhTMejMUSL+SDYQWHC
D94uDxj4lUz+WxRThDtSj/4jxzQqp3jhl3BhZkzZamZM/9Yilcq/Ynw+iDAJz3E3gbd+n+7546qG
m/Cd2JIaklcijuYq+N/PpdrGZYUidXtfvpm036+wAF1vGxag0yM/didv9z/IGjlGpo9loetDGEXh
h5VBfUfTRoGEk7AuJDCqPm7ObGA9lY9GshtTFb/AsgvaCQY+ZS1PEQqrasD0bCZFouQGyoReSsn9
6O3YVTKVWhFnozmHF0vJSDx+/bty4JZf3Obv0eL2NhcdsbX3CyoiSBtiAyUz/7QE3UgoSWLwYOKO
4zmi5iyJZ9MZNwCCsQ93zbIR5q0kY/POrGVYd0+sznkBYjX5Ax889PgxiAPWg0ZA0I7V+rJP6bHj
YMZGc/uywO1QUiEuVKDibr9phrGUgn5JgQtzN0JpEvC+AUGh9EoUrPDqqnTxIXIbVl12kYirqtSq
GuGxlCgNqfeF7ARZ14ZJ0WT33o3WC+/YTPM4ucXRayVjleO41kCGaLUX4fCzH5IlTnEAOZ3MJhZe
grRAiW8s2N/lsfwhMXMN+egOyhBn2H4zDiBktGn4/xMMpvjjdDdRfo+WlZAGd9mMeLD+n6gPHcDd
smYqPkVhYR5vBFaxV8GytM/pKZFG2WmFzgutzo9hNwcuh0xRTQF3/OyoqlBySMuC+eERPpQAoj+h
7+sZe6xA6YImuMOsiRMINQs6cvd+rh9IKyKZGmGgLohtmTJC2Ns618IAmyo3wmvN8FunTB0vLjc+
vzO24hOGmN6GUI7IRiAGh6Jzjoy6w+KEZa0QsmSBYBoI0bgEDo20SmQoWjxCRsDEM9Y+uS+RZ3zG
SP0mHgU1Jm5zpE5dYeNbyXqcJSEMKOKx4TNx9Qq9R1+vwEQ7itJIGyTTNGvYUvoxcp2haUkqDgFb
+wCkGPntLuEH6op5Uve/mMV/4L3B3iuajGclI+1QQF2d1yurMhQ7CRvO6sgjUE+NJyApaSqLV81N
XbefTIWCQ4xRvsv5f5VIomUDhEuvVeOnKFaoswWyFaoxxbOVs6VkVd8PJhJgdQXfVK0MzWrv+vuJ
enFQyYA5AmQMbuNzD+MVaVVrwQQDFPcbaffOFTo1su0/mLr31iJPLb7duoMzQ/mAU3Kw4RqJTxnS
uKVgDY8Sdh4E14A+/VVksjLnDxzU0CDn8g5DUoNVCU36K2SpfY6fofXzbTQkTAP0MMyzpjvT7Ghm
iX0TsoINsbQV0wY3PFEohsorrf1JOEWSPwt948+H9eENtt0WYYsl8e6pE1IogIspnWHA738uUhZC
uMSUm9dZ20mtPOdNAKgfUogeYzCfXMKaGwijta5iaPzdQ633BFoAg3XWnGvoTp+OwQUMNyb6UUho
Q7v0DMSBzJ/YirM2qpwv/Lx7s86mMxuzLkOZ6lZRDhyuyOQDoBv3o5Vmo2NDd5GIfnpewxs3gz4H
F6o30lKF5i11CMs53PCfYHEQwBMk1YDoBWxnI/1VUxn1e8GpbDJlUryYzsAxOJznYJp60mYDbSvh
GRNy+oU0B+NnkKvA9INwV2jfloTvIn3XoQWtK0aTcQylJxvMc9jbAO5+s1CJBg9stMX7U6qot5O2
Q3RK59zInzfaWvjVyt2+TiAIhkkSC4ZII9j+en/kWzYGpHALyWLDUt1tmKHvfbpvMDb8c++heX+v
4YbiKKMpQWdsQpEuIjeucEFGpkCuigPAIbRrlG30uacUMlFsw6VRaaEKd6S3pCdF4z5LiMGvkcE0
XC1wfGSU8GhfK14fTR0xwX9V3gfOcyGwndG1q+lhD4cRy/Bo5XA/hzgyrbMXFVCoQYJTPIM9QVws
VEsJ/SiPps3w/dsBJsE1cfzVw7WjQwJg34lP9o3ioWrO8+phWtN7ujHeGiwCt0nB5neit+ATCv2o
+Q6booTgk0LyacAWTdn2cSmjUJBHFjH5Tl779WLhVoKcZQ3BULgS1DzsDaIHKE0RVYsXVlVl1nK7
evig/2tAn0pOYaZXFDNviVqVU0wO+hD2VFSiVgvekCIvtB3/txRoucaCkwZbrOqLe0OMujMXTZrb
93QXEbsyIScsbMrc7n5TAMBX8u7cv/BmSy6NEF1ljoogQaGYK2lABwnW/IKFpKCsDerPgtSgUtjr
fvwwBG1qZwFI6m4rXv7quj54UsdYoXJ9IqEMVbTSeXv02eGTUJctfnA4OwevGNnQFsXvN+FD7Tze
SKSkVXDOJ2u9XE+bHdh9TpqQLKURI5gKaOi58Vxx2WwGBmX7AmWBzgQCoI4VeaYgEHEVtawq8lhb
JxgelgyplFAxCC3TxfCm8IU6x+DEMqVofFqZeS02/l1BtnqKYklCLCHpVH4me7XP4MHP4E2Cw27O
n4JHrKFa/ZL2JJZTkD2EhVW9ZINWXdVGAaPJDQRnlb0ZAiAx1o8UnncO1OUaQghM5kNbg2oRO7Z8
sHhJZgNI9DjaMN1YouNt2/igFBzHfD9IIt5/gJ/IZJZRHnN+3u4YPjOwWPkoTJSO9damxIjmd+hT
/2X2+zIW4qDyOPXisaQBWHY/af1tlEBCPDQvIGCRHeotDrS2ds+2ofdackT9gacgmEck7UWlNCcR
/msN6zBK3swElIH0uD+VRd7xLEfNutj8GiItUhO5kkZO5TospOJtq/dIPgwPImh9me31YrxHm8x5
yYj0RK9GZ5WV+yunh+VLKWBWlZeoVqgM6uqUw3LtKQEWTuPFj45gXq8JhyUq20KEsovIlB3m9/Z2
yQOCoigFceYGi9sTW7pqDSExnMfAXLbRM848Ci1c2dGiLHWp0Md6c0Tedj3xzvLxZt4cH4YZRUUj
rA1ybv4gg7hyJWQ+8oweZE9PdARw/rpAXGkElGyx+M4vCONrImP2WRhhLaQWNL3Z3xDLaKZnc9EV
OeHOyxEK3SVmczJF3qzJ8K+WdukeUl895GytQGFwlUKNihlQShqvo/S+gY8I2Dw6hVVO9xxvSdj9
wPPGDkl0BNBv40pdUiajyc7ylu7YdwcmxiiPbncckem38JTFD4x7hnqPa79TZUm9YEs873i7OEeP
aeO6kTvCGYuoat3YYDVEhizctMpMKsse0q+8s0vOMMJGnuyb35RcSdlDdwgxPHt9CnUY5IPAFdm9
3s1dWtSBXujJZUtpfXJm86YQUEXUsDo5kQCTSrV0ZJSyQu2e6no+i6n8lhIpk+Hqg9J1R0/+E7yw
iADBe1wOr1v68aA9ZPB7tOCmHo4FfxcI2hEt6i/5LwG00wSiMM2gW9kSK5ulE/55k9UEcY+zR3ll
R7R2f1dzMOqglGKWMpJBdGCFi+nFKLCWKZKhGuc2/dulJ8AnTS4YQDd/yCdhO4CsbYferff25JBa
ZJAYZOhWIMllEJtRJ3wgMtHx/P30I+yCPtb0aTgNyu9dSAgQs2PIQsGPVLOTW53EJnjrS26QspWW
yF3xmfrTSk11pAtrvujm835Ll+3rCNS7OhLcoxghyadq2PcBFbrzCfv8HuBs4OkAmJLSDrExbSyc
3NJeghqljMo2CbPTo1MjMS7fE5/09eyPmXm3sjmgHGeLIzFKrGWbOpG2nURCQt2Jju7CDj1xsX0q
yQTUf+0cMwoVtUXapXX8Et9c2iZidkzAkCmpb99VDL6e5axBEiBlvThm8COXVNUk9uDiiLFEmL2o
yXaNhJLYO4xRTkAHGlrK8GN+NHshMxep0XqXPUX/CiKqPKg5wQWzkfPnCxxdnAe+JefUmcPV+jwp
gKbHfp7PDtq1TCbNKVY3xMJ9oAIROo1VQXQKGeVb3RL7cQ3yZ8Yb4jjLCbf+G0Gf2OdC3kGtlx2z
ib/mr6MenHbEZDi/R7FWGKlQfcEOa8ocaeDcNvcjxlptbmS2rBiI9z3mSpAxTItVX33a3Djs6iyC
DpYFZuacgXSHOAE9p9qGT5Qvl9XM5Tum8qpBj9IJcG0EpRBvE8QskqYBtDvG/fyzByiF7NiE32K7
5+lhW23ZfMNbDKACRO0AXhykMOlo91oFko6pd+Ft3v28xLRULeKHFocaPTwO+bLoqYJXhHE68bqW
JAxlXHSj3q0e4/6croZQORTiw7UUWtc4kzT0f59gD5TEOj27TgkNclVpSPJ8/1Dd8lYSDXBnX4SE
eC0Chj9F6bhoZcEeaclcqXodVnyqH1geI6l2oCP0OjJuJnhkQDj/pVZGqe/+6Hou6nm4czF9o9Fx
/eHOJQ8WQZx+fGerrgF4V0hg+sBV+PvL+hsPjLPnhTbi7MPRaw/Ho6j1N1l6XdJPWwzOP3kDNKj/
YmDxHouAMxDVivD6YUcquNbr/li4DR0uQPv/3FIugfYHTwNAEFO10YQpkaO60aNYHQ495SywrukL
zDnBoOqzhQt6anZWDipc2thNzvezw1m/8cNBCEEEAs6+Y9gvw8yA93yqg1s7bCdQDXdbDsEI3o9I
zq0gthdclNvImmUMsKQTborTuPuoviEuGm07E1Cof3jlP+I0cC8ZCx6tjstV2j+/6shyng9awCI8
Q/RhsOJ/6OUIcwUYJFzJPMkRF2Ju+05YjMR2fv5NYld+hFrWp3+8V2CV396iOTmQVc74D5KR4XwC
3x+4gZYeilm7g58/PStd5djMz3uS2fmfmFhwVN8sy8pPSvOqFUTtC+9R0i0BZZCgx610EJHSB420
L4P6JBYiwFz0v24zhXpuh30lBJZlHtD6lVmG0AQZBLct6mTGdNKvvyCi5sZVDTViHvE7JzQX9SX2
0pN4AJVFNHRDtlAUJjct+hGU1yCzqXQZHrFChpawIbYc7oVKxYBtO0WfaX4M5KrlBua+kp/sB9+P
pL5u9qKbeKEHtcRQXlwZv/2/KY+CdKCspSEDamXTuLcKvyylINJ+PxBDQJRS7y8X9SV/rEdyz+n4
5/QXqtDSAimqBd2dk0OZKy/NAu6LJKg7IrHGZhJ1c+ofCu0W+Zn2Atp9LPHTRYn8sBz2QO0+eYDy
DbIoim3pflKacoVjpJ2XuIbn0uOBCR1b5tsaPkJ14NuHAJj42FnMbfT9zn2IWGI9gjOoO4m9kz+F
tWmx7LoFpO2Tu7EeApGgEiPGk3XdJYA8S7kenGv198pXIh24PCNJixA300OHu06Cg5O9HXu8cvII
uPQmfvdSyJ3Hmy8QIJkZSC++Nn2s2OrLdu2PYu05vXsKdNOcvmamf5JitKRZBIIZsvf+GC69SpXY
oDYmTkL4vDd+rA8LEGauJ/hOY8XN8KxuRaxJTvAB/aZqVHCUpnQ8OyIxmMRI0Yf2k1xA2f1xx94k
hKevilAlfSTrG6SzWxJCWg1EJwk7BrzB/KXfM1b+O7XQx++KMdnPsajQcYgDGDT7HRK1QYyo34AO
TGn5+JBIIHs1O74ESUr7muMx7jRa2R1O0jx7n72GW8en2jo4R9C7vuh43j3vEyMEF3CLJzBMKylc
Xh/a9PqgbtGGEgmrtDsrZstcOg80SW62vCEsMBEswG84swIWhmImglYGmFqHwNeDBcVJRmFZoPFc
RE8BLeKrubLqQyo2Bq2McYquh/dJ0wFedRDVNUJDkPKazn6iuAbA0Kc4YwmoARQCbG3ZtlQDHTEM
5ogVbsrw+TfkEOTyJHFq4QwaA7/ZkNcIKe0tydUQJKqM7lroecZAro+cXc/gH4mgcnqmfpNrc/LB
0UENgRJmTCMRxY3cp9jTKn+9hb/6UdW1AMfywexSNYHpzSxsREDYo1WuME9RoVo+aGBqcfDwf+eg
crQwJxYEZwSmiXNowDBErJUltyQ5KhP1d1N8EdhE4hWxjVhCajQV+ZbqugW4gJa1QZwnH3kt9y46
EXgITa2z4eZ6ws/2/Z+dpuxzbBIVvrD+MzVgFPDBO3lXvDyJZVRM8FNEfCa+VFvFQwszqGq+M9kd
QeXhkzyt5Lzt+9tbHEgFeyiwo8XcUkAnmOXVcsToyyFM/yDMpj0OQlaTWyA7DmLY980Sh1EQbyKG
veWWtyx3GCsOOGzBeb9g7jP1wSoKpYFsnnAS4DXGZNC6WfGzqnOx4yhn1Fv4s0YxQEbJmZMZubdY
XFutsP8ZtCTMUaDnGsY9W3BeX0a55pUQj6rfpVuA4EhRnf02LlE+hkLCsenjvzuAIEyluB8VxkO8
w6kKI2BlzZOmHgt+zs4ybbz7qE5av6J/5Abm6dWOsoAO5SIYRU5jwJm18shkGacoY+ZHms4IJRV4
MB12ZNETTSzP56z8DexUL7FVKbp083t0qaCWh+sTeCzySEzkzqNDrgCI+awqBfRP11Kn9Ta+dOJL
5n5IJTywywm167dEzqP7rvJP4Bd1MIBUt7uUwUCBoF094miHRNfu9ph6bYMVsjAOjbt8WKQvL9vW
fSHfnxmmfNP5yuisEcJeqL7DDV0QjEApAZNszWRsfxTdLjbPwuGo/i89DpCeiRmZWdhDwd67ZyRT
Hskig8LFtWo4W0KNRRe/t++eQZY5YZvs4jMRPLTsDslpqc0sBifH6GDj3MV7UPj50VcQQXsmHys6
98IcR57io08LMDnfDU4PApVCOkRhNo+Yi+V7JKaI1rqFUaaVyTsCfMio5FDGbziZy9LhYg9suqTm
CJ50UMNdCt//Cww6SkFn3nM3qJD+GTjWi4+lADNAjG0RNwAWjB0O9ZiEUkEnUdyGNZA6U+pwa/Ik
KgAAX+rdWfrNTWeX8vZuIJ+E4sEBcV8kMEZMR3/nsQ/b0R8aUiJcSSCCNDUj7lxepc1x7lOV1X2j
L9aQleQUG8HD33rAaQ/12OayFtPo/uXP2GRBx1H3rgURnu+EW7C9OtW7WEYBhN84gg2MJP+/wq+o
AIHFcy+rbPkc7QJaGukCoiuQ/FR/C2ZOGyfpGzC/VsF9SsmC+9cL1Wz8ZQvq8sZ1WgsCJZhTJLlX
0K5J4aC69J/AqIK3z/jBJMrC1uxyv7ausWRpwVL/8qxtB/WO2v+ZJOGhqlzZEGSnEEVPojtmUSEU
eF79vI7GtM3dbRsat3Y4UNegb70p1FQtvDyUG/VjdOpg5XpVd1/86dZXKLjhGIaRf7MdRfc84nyx
kMxzL9551p4ymCmdu4+UeS1aHmBTrdBqRs1di1gKjkWYVuhuX4watEjAAulPLppMmtUEMClxn6U2
ufRdmxNZhdaWgJNYU5tqh3AIjqz+Fh4u5hdvhTxPn1KWJLak+K+hjwkIbOl+Uop8sHaO+WVSs7mN
+CbGrU0yxBd6tnh2UBcZQS+petF1/StO8CxoPS2tuOxfIHaMWWXEFdfF5r3fof1pN9kdGmDexP5t
DU/3tzfLpOxDYNcTV5fr4qHWtH1NWw2jF7zuW16BvJ3b12ZQTQmFYgmWpGNYdyNxKZ5qH5bc7ylx
N8lTHmhCpB9lWzJ8MUQbadQ8ALDWTI4TFHRsDH3VPGD6Ea/tFAb0VTXSLPVyaXqjJpZNkZiWx5kg
sO6YgV4u0lXuhOdH8lh4FcxB7EqsfwHpBTVjYK1i4XHarxn1Gz80OlZaEn5cjfZkXf9P8/+89uGd
yxBhz474NHX3jSa5ZiseQGreBPG19G0tBZ6bZTfiN6FhMoKo5DVVtk5L+g7IEQWvyYZ6dq4/op9g
Bcmtt7ThdXhzhYcwXW54AfOwn+amCYvMcLVHuJ0CZQ2uv7Y/D9QDauD2aQCHn2Tyj5zUp/92K0d+
jxhF+KO0u96ZRGT3akksew6XiG5YPDGTP/Ha67jQfR2MtjyI5vqDazpf8iDO22gZjZyIvXv7RgXy
qrzDanm5IPJaYA575dZhNJwVZhgq/Dg7JQDfHlChVNMPJO8kL/5CveyEFjfSNspDUSlYfz+9diUQ
lDo3jCHzbLd9NIwXiSG226d76Dl/VGL5254ZJWOUW634wpsiVqag3xCGE9Ub/4goZm5+fLgq6Xai
oBXNFnDhZVZYNiNEu4fpGGGxJ8zGXy9DD9ygi/9jAHWi23NrE1CVxjMJ7MQVyDoSE3A5LPNehHQj
SBsXh0KbBf1qJQQDPg+OnWixB1+FKpv44TKwtU/w3yomny0tGNnqcEtn/GtuZqm40JBT0xwgDLBm
4g+UhTnghiB7KkK5yjAHVT3Jt4ukbtTDphbzPsiF+jE/aKLratkTKZEiDR9rnYrCfUZnet1g6TBy
TjBbh7ESjyjR0z/fZU2kz52tL6rkgGwBqOAOc7mFSkKlpGxtxoVXG2cuyap/pgmRG2+DxVg1NW//
nZQA0Ztn+21GNY+qwVxfjq9SweYCRLRO5EOA1YUG3aSBKxQVA/XLbEwigjiSJ9O71LQpPZznTxQn
sZESvMFbRTcWcNErvtT0AIYtAHsxDqgokJp8kJ4uCtqtQZkCSfzymQUv7EUf1R+j0uEwrUsr6J5x
yE4BWqD7eqsMHw2O02S69pjWfdFJTbPXOCL722pVXDUHmIzWUWOvRSmdqtX+4oZFwiQ7xtDuc9Kd
5uSMvBVQ75eCQuFwf3e706o+ZrTTTfYEzuXceo3fF6qhPrH+MelEureiuDgIaTLQ7HCSvm1K7Hgf
pkSHWwqAP3F8z0Q4Mzm70Lv47APKSWqjCSj0sUXHi0wJvcP3UN+JZCxyiq6ZU9hz/hZiIfstdrei
/39ZpRwxHorkLOIevla9pov2b1vgmz1UVIFo0yTBTEWhTBndqwr/siO4RsEXxpm9d1KZX4lc0b0/
k3G8T39xGiPg+e568JY30s+m+7ZAtGQ6p/PZI9QSp7vuFL4rTaSQPyzlFEFrukrKU9MbQMrQDPIb
u8F7uqB2F6LTW5AVyT0fi5ZsEKIR3SMk62HHvFR5KSuoW2KzqMANfVUCQqq64uZdtnSQv2lp8CLM
w79yvH6FJkQuMC2qKdiAiFxOXlvHHsMF2x60QuAkpsZXfS+jIk0jrxrMcCCBF0Rel14bptCjJPnr
7i0rBsFfTcIjBV5d2gY6jGXSS/O+b2odj3VIYZFnpEsB123FTMPKvarF9rmXlf+wjZrQSY5oAEkD
RTXUaNsubfi2EKHOysdizepA0ME04MpmoVBG0qvGt4mYGieRcKQdz8SWVwY222FOtTmGv87f63a4
A6cm+gp3EK0NV09sXwwRPeNdDgBGuUy5H50HFsNLG/BlaEBkVvIyd6TEpzOE+gw5cmT2MIsl5pdh
8OpUnG6Ck8iAghegjMMIbiPRJatpg2SyXQCf5pDVg/RwZ5ahp7qUGYBEAZGf4fBZZdh2Fah/8ekz
OXfQV2yDbuuCZ5ZqCJ94UE/st7d/p4RTtS3W9HEPETSe6zjR6z+7K7KEQo/c3zF/Q/D3toCgEvyy
7GBfaqAmYBd3l0JxSiC7nuSBF0zsoMA8MDkrtOHaIH1KAkv2MCfnsezbvUFBy/qeOgnHEC5CEi4P
dpZeNjktikMS7Aws2oPKzUOtX8KurRaGwModf85ycxX5ZBKm+sncAqCtZYyg3v917PEa/dIGd7y5
OyjRyAsJzebBjiKpqncq/o8HvWA7UAEG/NaTJgqcWTQ4TN3QILU8UMHHBxv7QdFyr1lxLIkde3zl
YUIGeonnMj6L+ZlLGDuwRj++LjAx8d9dakkcL1/t08pgcHdL2zW1aHBNjR+NRjAPQI+Bd48nw5I4
FHdg4s+8dRF2qXsfoBAUqLgQ5McUcBqPUD44J/vVOiOnc4OiUiZzB0iw1NGUzHvealS0e0cLU68L
9TJvJ4hq+mgDeiYgXdoAaxtTUYGXM+Cgf9ELIYjiG8eRKJgZxPhauL2RXNxT7JQXysVOu6bOJ2nb
rdMWYHQDTI11CX2tlP+NAesY6Ne0ArnLmvbjNnuTb1S0sSeS/JQCmWaMAL68r2gQ+SdGPZelCxcW
JlwTOEQ68+m0O6pmqVJIIj1MsoGOEZSD7CSDfJyM1WEYBO91T6d5jFms1Zu5RpBZAp/rLb9aiwmZ
dBmmmTGSkF8mrmzHIPgoX5zomwPQdt2olkV+O74b3EYX5v389EomVQAxnm4VnDq6wMEiZHZWue3D
hf+sV0kuafuEUZel9OzA7l77UQY6vVYGs5tOzu4xCcgDYPxOkB0wjKn6W7xulLw9FcjRP7q23Bhl
Imvko2uVHuQNnplJHOLX2+FOj2ywirhXWdq5p/JEzLObeZvh+lxOAhpKK8kNrdjo/btk7oYtQT5q
CP2xmjcbURfkPqwuXUFQtT1gAmBegkBPjgmDxt6isBXV5HHrFVB4mhVKtDl6D4njY6/1f5xrQj35
SDQJrZJCsnyXO7z9EVUtzBKH4B0UXEAIb9P5YOCVAwf2nAe7ObKk8Ss1wY6E3wBIHMa4lAEemYqP
L5jIM59PNU/G7OH48l5Kohd15hTu9HMltZ34vg1GvCAtdSn2GkfFzX7aybLmnUuQeOpxMpmVZoOe
X9N0dGkI+/gsnFsZg2aAoXAR81taxvr7SMgiIbiWX4ieZKkbHrDqMLUuNCIiwbEwwX8bwu6z7ru6
HxBgctLTkF6r+tZob6tkJgGMIAsB2qN4vlPnYKa+k6b6hi7Rozs4FWAVT6XY1CfYKnUFvbvuzmZo
fls2ZOBk7768/ALwdI6zjfslwlWv82iXIr16T4P74uSRXpB2gYU50/V2H/fmsvQZVV07QHgEve5o
r9vl5mQ3LM49hRB4+pyb42aUfOFiB005DpfPXoYVqhizKu4CMvpNE7XC6Jo0GYMhCJZZGNuTL3zG
4GWhZbHo9A8c9QiNRrnlA227AK3Y0pQZRYuaeK0UM2DTQaUJYg4I7gE7e02IJB00ri8ZSEa+CfI6
5mY4ix28YWRyQH+qf8RbKNjx/iLLTgJ6mNENGGViKZIpvOKLDG8BfPg5+izdgTjiE2ncG4Fu+ao8
C+2SYm2DAOtzVwyl2hDe+aXR+P940FMTdWwst6UKvjOvcIKlaatVWJnJJN9m+lHY/3++k+6Iyj7/
PPND8GZ2tEGYa4FjK0evgfhUNd26qluDacUhqXhc2xi/huqnzPvEcPzOWIyYWbMP3pyv/qbXJK+N
gM92fNjlZ0B3cygvGGeAyMrmgUB/kXz6VofVot6V1+sxyza/dOhuvLe5SFcSoekjcG1C1rvGbLRz
0q7hS09Fx/VFwIexH+p/beAZ6HgyBZ0SFpSBnS5nJIyBNnUuu/21vpkhegR++Mwn3xNFdDPtmMNF
Nz80GDxIAyZBW2J/6QpQIcnzQvKI53+eVwO3BnjFHoLWjBbrA4vU0Rl5DD52u5E3hSPvgUbHRP42
4mSTtEO0qiyWjWppL5wfv2+YPdQEa6De2VtlRNshYLo1LEwbw2/+UHO8lKBd0HCMMbG2wDhfoGOg
SRZyVPpAcnwVK6PlxDVd9L7yJDdFonJkOQioJa4mC1f1Uk0M5uhRNItuLkMV+1CpuuN1bAxQB20f
Ud97xEMsxPlZcnv6YAfQvAqZ1loBWElXXsuaAAQd3pTzWjaoZOkwkk95dS0Vk8dA0L6ef6Ja+h1p
o/qhV/Vz9gHP//plIlBeLXZuzt6fDXCP9VkCrX/98brQkd9sZj1fk/zDRfhsZI2PqTCyJ7YkoQfd
kRXHQziPdGeX4SNE2ZaAu8iMwA9UcFfflo6nJRJevVdJj/r7nFPsfbiH3MiTuh5G8JzQSbrQwizL
sdA6Lm/dMGAkO6bdinkTJOurl64MxfuYN/8P8P9RAYCk/66mDQ3fcRsFCRrGyjWGw1b1F0sg7Szg
V/sBvSEhpaSjBryCckE8omVXiZXc1wqCcz1uYFAKSBJnTcRT9qZKOVEgA/tmp3+TSnZULKkObU55
aDgEasyQd/94WqddlUmdMnH77+GggZulzS84VR4PMO0ilZMs8n7goD3vWuWbUmU0Ix6OK6+BGm5w
7ph1UJYuL/YEX2V2ghsf7vaorJ76rLq3Ocn66bIESdxKNC+MSMCyc/FYOJvdwDDw1DZPC2PTvEFS
T/fe/9QzqyTQaY6F1+70kZWiJ0mSreI5UMem5SSiL0rVVf0z5kGRGlvjFue2a3+RI1NM3GS8xZOI
L5w6NtaAoUYOyniAWZdBxCadv9vdQp+3JjgHkgYvFMUiN42sBO+vJThPEMxf9a5Yovw6o6Pi4o3l
7pAwhwo4XTTj6fyA34QQrLDpukpsfgJWG9I6MDvN+F8oO6B5xBjXkuUEKoJC/ZRaoSUMYRtjdFeD
sUWiTEB4jV5rACLUiQF9xcuN+e1bEEgq94x4YO/urGy1z1k9KBqxljQ71HCHLpAc4R/4Ta41wd9z
A5kcW9wrqdspgN46AccT43DSH/IaQec+tdajShc9OoapINedO+QujG6E7kmJZ1AKex6c7kH+gR+0
EWYqhqsmhHUrx90KaHkSZv20ayosStrK3weyTNDuhnLzm4tpsTe3q7TIGQ61pUXhLsGmJd/GOWop
JetUdmZ9/3eIEh32d3laRY3L7+fGPONFaZlTOBErNHqMGBcabHUi+BBq4xanv6yUINlCaHcIVW5G
ON2VuRd5GVJRusZ7MITp4p75EX/m2fJtqsomCWhtZofpx9cm/vXx5qcGBJPCTGg/GzdgDW/HklMR
S4clGr5jzrcd9Fc6WRjCSj8s+60QkmZncgGJRxa0KzzMtcLlNsxPrkRsbL+Wykv4bVEwl/49PkjP
zPeBg7CZE1uzEMfpSeI6Ba+oTwBOO4dYJXoBX43xZ453egDPokF6gI1EialBdJmEg6zftMxNcRDm
1GDMa7oGJag6SrVLEQqwpfSS3JpBBzTpHB1YyIipuI55Bkge5CHYrb1btTBHfwUTuxmT0VgvdbDK
wt1YNSHUyWnaxe05TTTvEwsSa7yzHdfOM8T+kv9IZS8jmETmUAatRlZhKgg/W0Dwht/J1JUQ8b0H
J99wROcD4bmDoxYvIaacGv7UOX3GxigbLvKfc+3GG0cM66ghzOLRezdjYVpj8bnfYSr3MXWzRGI+
LZS2pq3ry4QECC8JWGZET4mM8OrSpB+ZZu8Wei0jAuaEezP5D3aHVHQzYbuccmcaiZLIMUkPCbml
/BoX5QO/HHspCGcGTjitSJ+Z7PZwKvwBvpZAFMKI0lpHjaD2KDhtAWbfMZx/+2+B9anDILQGfFZU
muMB4tfDqegi+etWwqUWG4TthUePXpB9Ims2bNhhJjZEg/u5PgQ6yxj/GBGgAQBeE2BHBuXP0/g8
GHvhQDyfHPDqk0+m1qe/7iF+/DpIXbfLhjkB5VL0keqUqFXCTZ/9Ou2pvUwh5WUVHJj8wIk2t615
uJOzlqNZWoGTHxY7afvFdkBfWI2xoxM6dn6BOBFPTbLiEPXQ1gd5yMu/Oi0c4QKzT+NJUCK/3jUt
d8Sk4FOTJyWgD5wnHAnyiZcm/9azxNg7F7N9HAoiXS5gYmvhIVrlLQqBIl5G9eLcxRu/g7NeaXje
ZEhfA+xrKtp/B12yILWpLksEOaLrl84P3e26dhk3NZMjch+WSZ7XZ+H7jreehMV4hsW23YvgLSZp
VKY8CNDObMYG56p0mvXyWYIrbQ0KmQaTrc5dsWfoo3c3bKDUuVLdSfwbWdTXi3Swg4Mx+4BQTmPV
mtzxR40DvtzQWTVeo6qUAYu3qiW4oQEtfPjs3qQPhUCp9LT0Mz48hIzA/n2bLC157nRtroSMzGGJ
QCy1zkYnQXjgrZJAY42ImOKoxAmfOAz2aC1kjt5QKUN6VsEMdSKY6gsaH85juWe8K0vOW8IaXuUW
jj5V2tCihdsfJls9Ofu18huxmYkC2t+N2yl1POCcDiSVKdsFIEdqwPrSxpXy0kw3qQFUewIuVkWD
CqPpEJ9PY6sX3lSAwSaJtNmTW5R0AdiwHB/RocuezOBYLK94EmoUgDZtm0H59yKlm+WNu1qRKxF9
yaictwxyJyrV5Y/l+3r13DIs9jJwsF+9+LSMIQr6mDdWfi1tmW3fNg7YyRwyUk7h2C5xEfpmM0yu
4mrEKwgc7EJlv3V01fqWMnb5Tme1g3KtSRoyj8Vu3Z3rdnTLi/nJVC2ZGMVFaOLAvzfSnZ0XuEsG
DljKVIW/4z0yrweV7v+HQrOvNZnGogcz9D/kfZv7w5FF33TTcb7ccgQtA0w0ejN678tSIbuABoly
KlZQvK/l0zjtTkFl9xTglv9lST2o+MkIlzvJHz5LEOC3+NtMtuwvnYC0wyEjpFb1ZU9ZYo7WjOQk
0BGclDirRubNTIQO7ketlMu+reiqHiuM1Xep7c8tY6EjOjNV7GkKirhqcZxAWKQgZUDZjUpKpp3x
7oAnBtvf0Hr+Y+lm1ANq+2hiCCJ4gR4ARJhsHmzlp1GGLD7xUuZkYtyjKSBAKgfa0+scOGkHq9/V
8mk4OXK9h4Y+m3h7Qx1AAYqBLrSrREBY4OCEzLSw+4jLXYdE0u8LLN/qbPNb6WoD/ul22VpeIjrL
ngatpRExGf7MNnmhNvNB2cS0jcwFQDkuDyg9JBV5LqnDZpzmLd18DSpNeUWmgoaHV6ejjpqBzlP+
0IZkUconhtxQzideTqbAPD5gHsjJ6nqayxL+h+OT+LVgGmJevEtIXmUvkAvOiyO8Jy4HuqULm1YK
Xqe4T0W/BfFF7fh+FzL2ixokvum5ISmDW5ydSXTreaj+v+9vYrv+wleqgbQKQ4DOBGn6FwtpD4gC
C/P/M5oCNsI7HlSAsgGTlc8dDEKZNLa06lfUnY2DO2ktl2Jf/iNhMZy3K6p3kZ+ygQD2c4074ovv
5myM6/gKDlTWmoNoVaI4C9/DaHVP4IkmfnGDQbSH1vSVDSruVk/3QipqxIvN5Zu3O55q6kCG15Ux
3h1mzcZDpieEYde4PvX8/VoTlhHEmG8TY8Yg4ISwPn7YhKTeK2W0ZP2XbHRJelT7boDFO0Qq9q/F
oixeL7174c7sE6XV93/WFeSfxU68Te2oMIP9XWR6/xXp4K9HtaESzAnBWf48Sh2/PI9j4aStOG0z
3ej97SGyTu3/v0JDkye9wUD3rJdo4UJm3O+j8tLQh+kAY8N4lXJoKrBcWDG8Nb7xJkMjZHq45xou
DRzFIB7/h2K+3Ep2YLMG+rnGZRwfJQcQe79Yax4oKnOmsN4sW/c29JhBrN1c7nqmLY55NxW75fsQ
6DH22Ll0sC/pA9jy/blDpV6JdgNih+YyWdtMV001JfdDqnoKFJkBKPsz+jv48ymGlDRVsJoztaQM
D3zIO5WCNO1JOmMqhjawFibym8jghQ79OrHU2d+jiKh9eEtqEofKRtkRtUnsW6Gv49F7zFRXkfxP
SLBo/6vkyoKEKypmaTJJrVmh3e4irlC0KlzAJ2OxAO0pgXMMwetyKf/NvUoYE6d8NMCEWH2fVk0D
PGS5K/9SkuI+Y1toLGxpEwWcpqZxrsYsYcKepfkX3eH81bX7qabr08lWukb/B1Y/A2wp0xINWTpO
5sDJCajehSQCFwY6VraLGOw5CvNLRGNW0pEwOW0ImqzSN0CN4Amf5+npdF5eifyUDoDPeaZo7BoC
qfuM+GBpxgzGZCg+hiicw8uZPnFlMswEvG+ag/u5lbduyLbrqkgoRRSVmZEbXyJXggQYJnO9qyn1
ta2Blw0K3m1rNWQwLHnDSsDrirV3nVwCo7/mkA3gnJh8TZJLCKW+CJN/43K7kS7eAlXFkc9tFd9N
Gxtch/hU+bT/Bd71OpOIFszTpD9UWXiz1mcAy6P6nZyMRmZA0fxgirQTcTjaCOl6bNNK1rwnbGJS
Xr1EVV6iL/aR9HU+NSIxUxHrOA84NwZw+5vBBIKr8ykbc/AE+zYwIkRioc1gTbPVU3uhH0yQvPxG
BQT/bhLP8bOFSg9HZcUl+wtzOCHz7AiyemNiYNcrNVOXGCU2i3z2f2KUchCQ9jdvea0+THeuV9sI
0hrpqvUk3wJkk5Yoh+NeO1Tsw28MLqHMGd/B9Mg01U0PRPVs2IZZO9bxeT9VX3PbnCAYcwMPZC/k
O2w0w/N7v+En+/4+zU1VPX4CSe60yTCm1NPN2/Lw+rgQo2VW3oL3G67ITQXcUbPjiTqgSQUOxPFw
tj0wggss3xYRqV6Hjq1YYcpxOJzbpK+MloFJV+g+TkSDC6jWPrqAFjtcHjVhTIZ4swQZ3zgI7wXZ
XmLNvDyLcOnK9qMefxWVcWA6a7fwUdgOF8se6mN9pPPHsHm2PJ2XxDYAr4e1o95fpia72mxDmUNC
wOceCm9XBPkm2MBGMHzkJLPLmrrGDJcquXQCZ9n5auzssADOkbOzikMMsyIl8VULc4K0LnE9Rl+t
YPkXe6D/fXXImHbUE+2iuB9ARWROjasrPtn07mhc8pO/MNuqSLbPP/vxdOZiizVn+coEnZJH+UzE
A89i14unui07r/vCqh6D/+x/cjtUbQOMZklmdc5/cvHcfdm1SW1rosu9HYjQFBSSvTOlVVVgm7fE
ixfOnUOwbEeVF6kpl+fqGKE3CBaXqON4M2tp+2RLbtP903rQ16dmFlUhN471Gca+BZdBm0hd1aOX
G3SZPaS44hHUcsEAlwpG5rf2dbv86k4cPNXHjhNzCSuvx1ISLcKF5mEpUkP5+XR8aeMghIDyL1/X
wDJ3OYmyPKwUCywjQSRwQZ3eXApKCb8iKDE67pukzgjKRG6nA+pB/XHOzGzBbQpcAhoaqk1AiYM6
jiokpZC1Vx5PlXzAEIqbhnVI4jvlNekeppjtXyBiV38BwEjIbS7Hc7sy4zu8HpMeXTBFO+jrm/2q
oeQtmjYjUgKTNaScHTF14ydRsc10HHGftfB6Ldegyd6KYZThyPp12NFqv14v/gLjN5G7ERDbpYAi
qJJiQdsJOw6UkjwAQVQozEvIu1WohqaVxmzCqBhK7OoputAZXd5VqZwUl5rCZNaACxScI3TsDbRM
OIErrrRA5OMISng3nTCPgCEmxNTA2WVemvTi0CLr488FoRruagAjruxcjYN7GBPLjX6MhoAPtoTn
VJ3HPD9CltzfbgKWh6JqRWHaB5hGvecBDPBMPqFgjdYidhySxhtZlZezY8eVvvrvEd84mqt0/BnZ
0JCzsDhRhnUzt5kgGfgi+CDKSiKpMEUtj8+PsGW9K3E9zAxfDuSSJD4X9sqFYao1wta3tlo+pLgO
hU7whbp+eymy3Wfm7gS37XFoBCqizVELrvE1e2AtPEsqfVe7wMLonSoOKtDcIOXL1RdQj3kwpRAI
CSSnR2e3FVkfVsdvQWb6WUWANSpkSzMJ/zerqy/JyFZ5wraB8mnxLlB6zqZV0QeuUvlubAoVuVnm
2HBczq/qPzp5VOpX3b5TEYPRpdS7BlmZicNUPfj2UWQeW+6hs7OdsL9Z5XS24dpj5XQ5sdz0s0/Q
lpqF2Fb+8C6E5rg569W47e4rKk/2iXwclOxwvDagVudIVVA3oYEqZAzlA+2tDf6/Yfrc/yPM4517
sO6URJZ+5nBYZ7/rCVvzQENcK/Uqf4ZXhvzSxDg9ifANJAZyQGM9hNCZrUDzJmNUmY26GYkAjtvR
POBDV/iWNa/Vr6U3pgZdhIPdbzBr+mgTWZ5MuWz0qirILvZj4oL3MLx5TghPsPzJ0Ou9fdpgSJH1
yxlQw4MRznSwbjIfbY6e7ZWzK9QT8LRcOtLsQio/Zv28vcB17iwbQuYHMjl+fVDXCFx4msvAj4r9
ZmGcZK0g2MotJ6laeu+T6gHbesJZqzeH5e1EVI3ZwPYsoFc76eBwPqJBVgQ3SkY55nIu2RKgHDMT
SwYBggFRwe3FMtAz5HP/wnoXSHqb2FuSfrG18WzBGO357s7tdUQHg2jje3nePWn9rC2WvI/kxDRN
LTmIKcAfLza1dUJLkx+3G1w9MNomuEm0YUmE1ok0jRzIk1rosCk0EbA19Bo4zf+L/1IJgL1ZhmhE
QU8NHHKjkcK1yh2Nk3PZ9XZ+P41gpTSlaRxx3NRRgEYodcYnefHcv+IX3iF1+FAnz2BMCoeVu+dS
t3+jAYF8KEgk8Cavn2VoRqjtIla5FMm7KPYkQCxlKeHaKCM+RhXW7OM5qgaKBzJ07J7d0fggDmn0
Sq1l02WaoEKmkRyJkUvfjGvaevuDzjmHU3H0yODfDWmQdvbN3Xu4vsXkSuDcoP8SBKKdQF/F9WZh
6Qd5vUlwyibAY5iCAjs8Fx/0COwKaPEoXw6bG//ZacowPKrBUXIthOLGX2HNdhXGJSbebTgTQM8o
j6K3JNyzGU0A9gTGisjhtX+ULdqCcVaBjzjaJO1fkvUZ+rMJ558e5brZpt+5ZrSANkNHaOXLSGFy
E0/VP+BfpZ7lAyo0ira7yLZpLHLOjCnbztTkHzph7UmvHTuQc7GeE8quOgmk7m/fR5wDOukRS42o
wdBO/GxibxT16Kym2bylp22Z0iMklfezhK4zwIOuM7y/m/nPV8tMjVmiugTtsAQGpGdt2FN659E3
mlQppQYUdQvEOVWH1HyzoGpPsPsJQHbuCqq5sfNoXq9l8HQd5a7ZwfMjdoEWVCA8eRP66vM9aJTB
ZLIhZdKDnCjKdDEznaiU2S8pTHGhwI038XWLlcC3FnX/woB421TkxYMc2dLjafAVfp5IkVIILduu
EzWlI3TvfSAyv5H+HAY5OubizM2ryQVDeWS+mymEBdCnhygOt8j+70QZiZPadyVH2B2vvhb/6lkk
VKjGpNdfsiLy3Eot+KBrxiiY9kmiVRnfPCP2szxk+TcnXx74hRWFp8UvR8+m7cKDyz66ROHh3yCU
r+C8dabmd6ZKQBfvzpncRdWNl+0lphPo1de4fZtiBZ5f33dwXCSrc2X+6xGYfR6hYTsTmOpT8jV5
77Sy9I0XuGdrNEW2AgYGmEHfS/tnDUKwgvKH9v2y615FSx9Wr2geF8n1uB4vZheRyB2MNJAc+mgi
ybBoVMJSmeHo6jRLCtdDLDn6kqdPHh+lyNFJP6rpMQSqScWr2vsGLX36k0hBn49Otly8iUMagu3Q
P0lEd+T1ju6fHG4lewpNJM9QVwRTKNz6cXfdgYgfeUrD5iRR8jPKvMvFLf2U9vJ2MYkQv7Hen/X1
HM5Eq1frZUshVrlFZvAeDTlPsRV4wvIf13xjYhhNrUqB/lEZxEy25OZgpJn6GtkWHp9iHmXst4xG
QRsiLLhqPQ63YbwNASh2OUswQPqyv3i+3u9mrq2qirh6GOPoRA5pbp2hykhnwztXH2X9R0sR+ydz
N0vbMGFCSVt6/Z6gHrZpWjuepHiZDh+XUytV4kEenYhVnLP1DQ4Ybj7x0f51SLYd9zK/eWilYx3D
P+y3L3Kf/qT4WXOJ8cYU0nRJbeSyAzzrl2VoVLl+AJlgXt8w7U9DMQxMrOjnie/oM/Z8fNB7ND6k
wbdjZardlUUnq6IJkVmrYfNZ3bMV4h8uljrFQeQ3uBJWEPTbEGxxWVfjHbrH/nGjPHvKTAYUdBkt
TcNSe39BLJJlosV3/s88kr9Qg8wv7yM9gZL1bKfHMQrdlD+TS7UT92pJ8K+eqJTCooJkAZ81Fwkb
35tOnHHvAAcq+x3r7RGzQJE/jGJwAHRx7ocXoXsAdV7UnFUXxfv9PELhU5O3q6f9cotfZVnx4OJ8
QBkRewjwrFzrsOcvckdXQBA0rirG8tdXhyYpQPwJAaiA5h5mDSVVjEVzJ3jgJmLMeSeipJD9xsuI
9ezHmdw+WX0//Tyrowx+uxzq5HbkMaZWnvK52pwWoDyouhXs9KvLf2BXcpNZFMShD/+mh5RExaEH
H4RuRDr1bpQbF+JhUtWVnVAZeR/y473hh+4i/tO7DqSEmHTPAJsqTCpHYCVVDjtubVA8kEWL1jc9
F5q5bc/8j6wID7JqcOs9eG3F29ywGnd0i/0EWzISMLqQMqdKRCIUOsx/8GMbE7eTbYRYSjR0u5Tl
2sbZKq7gkjn3rPXRPYW/gkAGnUXARRLozypSbfqcKONrd+Q1e1lWhwGTgAJItTVmpk3CoUf6K4/c
1amOrXKhcyIIYyw8wYJYEmEqoQ+9BrQemf0c593FBC+ms0QNShy1+rHLURXcothnHP5zAEYvARZS
LRwmOkoT3axJ9LELmM//iwBz7ZDKFFR6cO4njlrRB7LciQiVZrwzdE0mxJGRO8yYZHD5iG7++4s2
xgHSUEP+7A3lf0bY5KZJ9RpltjfcabL5kUo8cj1PtZr03tP70jnrnsxQW/PfndqqmuG0JBSqlAos
1M912NLZ9uGlU3/YckQ3q+nOfEjnjaK23YKkT/3uUPrYaaYN29zm0JYXOGOmGLroHSvT8d8dMq38
iGw6RJD/osG2isngcVAXv9ue9sxhwpZzkPxwPp6p9e2OOcHl22P/FMBSVnuMk09Tmwu36y6i4bE4
v5ZmltcaBG1ncsb1b+XoAuSvszYSX2zdQs3+codHiM1G0j+UUppVgrsYI9M5DmIEP5oybpWPdD0V
jAFlwrye5SMbCLotGpgb/kCrf2n/r1FoUmIMhJOV2dNCT8sdDbRUAfvcO0xeeMtZzdZaJhOE1DGs
tXDoet1/qjNgRH679os5ELujqZHOa8FwNOPbaKoV8tnwVrInUW6C2VmnGtoUhazHiLzQB/GLkIFZ
1QnkPjYInUgfziOPSv30FL4vrAYSqkysuuKn1wclhlfWhPAYFWSqqBJjFY11g/pMpbn91blHjtma
4r5xdS+zpYQE030bxmhPCb3fcyuO7p5zjng1jD+vxv4aLS0BZQ7UoFM1IWfNf4hk7FxmYoanDRa/
Aj/FIZrxvRaPmysTJDG/6fAW46I9buU3cOuppijgQ5OBp8kWfGbUnTDhrKTzsZoIzER2RpBMovc/
ddJhYejsRiTOzTs88OWCHFX4AsmzSsVOZQjG+1DmsEyvxDVPhb7DuRM4HQMYg07X4XlseSy4TDoB
PXQnHB5oB2dSjjWsZtx60ESpJiq+RoBJvDBmYUenr+DWZPL+e/1dJkOY43RILHxlCrUrLTJxfLm6
JZj3pGTSbFvdf0wvaQ8Y+KWF9ReeTKlvWJdejPZpU0Y61J6n8gfBdVMYhy3JhYjFzcj5yec3JKdh
yv5eoes/RXLSoojsPK7/O6bw8+urreN3fhbCMcZiRFNDY8BYqLUI2+FGZNuMxSmIIGZpab3apNQI
ywsqt2pvJQmSx4HzUY9DytQiE2zcLkhmc6h4a8ZThq67c3MJCm7jCVNzhWHyYC3crcJcfoXnRKg7
zu6RELf00KV4hULX6i8jj7Pz4U8dENvLsxmj6/ezsAHnPqbH84VKNCWPjw7dgWQCUxsGabob19QK
h/ybC97cZCtjbAsYLm6vuf7M4yNcKaKCMODMx/NJXGi9MjXgguEv0x+IitTGvfDN/Th1+z9AwJEG
WAP02OSDYKoe4nRtfq1uZ8tRpXkhKwvWGdC13zklQevf657o3IUQlIRPqp8IXK9N8Cv71hRirL1G
2JRr+HgHP0l+4C4u6xeinvkHPSNBeMNTuIUoY1byK/TvBL1PnjbX4Yr9lv2//EWTxQT6LcNmHLXp
0pV/oQCsddjI7De25FoCSW15Rwfl+Nrs/wIFYpafiuBCcHjE2TXBRYK/L/GZvQDEjo0f7Zpio/1k
wXRHweNEwW3fDFRZkvFcAzGxZAiSg+WFqQAh1F/gtSP2Cv4a/EV9L2zuQuJQSDy0AZz5li4hN2Qa
q1ilbeb3kSUGb9KRPg8pUAXSZ3VzLflFJ+MFAalr79YRZGb5uU8BGPKs0RJGZ3dE4YLYcMHHtpEE
5sEWijYtHntYLpuCX/R0vE60EROlEhlGnSH9b1PEjmU5pgJM+XzEjWhw+uqmNN6LoRGrSDrfz0zc
FwgfyD84F+3jvtlKzT1w2tG28cgQ25Bod58Q+GsJNsujlzIPyEPM95O4OvpXRfY0rTjE/y3k6Xk9
Khf5t7nwMzPLX3U/09YnMinoxPv344hs5f8bICkdBKqcnzyq0e/hOV50SRHlkZSSY75gSg1gBp/K
bfju+8NuL5V25s8bbwNVubY0nQ/Qsw6xsLh61avKMzc+XRoqzS9tSojIuQqIDBoPckcPV533BDCe
MwNn0gk6AlViR03WtpGMknN4XqNm+Gruzgs/Wi4IpzRI6wW9KYzUkRb2pd1mPsz227T61tru3Z1A
HrjH6d+q3s6uC5YU//WSIk4UzXnLwrRL89mszFqZ45YhcaanewD05e3rY+7nzPritGOmxUuXVPWg
t2RyohuS3JnrSujP6xLcD74+cwGjY11wRHKFemZZlvUtRCnQlxLGDwyK8d5ryZ1wFb1RiT55DMJO
YCxXMFZ6d+P+eEubx6G6uzNBsqhteBc714tSCecTuoU7JpJMi+X2WUfzx8mpRyMpgy24J2FJeGqm
nfKQvv3BXmgym1RZN3HqFghOkk/gMfQs7kbL5AIsfZsu+TvXhTgRIT5Tt8pjIFQyj6TNZDwLLflq
Wpx5DifraoWoaT+y78TPwCKraPLB4f9Ru69UyavQQvd/8bZX8ezVEdOeRCcIAgjxP8L1ocuCDL34
nQQOBJcRGytDTLN8ABY+Y6o04p9ofscwwbX4YJlLtaRT9PSA1OdByxfYcGRvvNUXQDeJAMXGGemJ
Bd92Cp0W9XnZCC7H/5rGB+RPCSX0jSkTN9P7F1AltYPv74+Mn8kGFm0MiAqi72dYwGc2JEwBQAuq
s0Pt5BYsw4KZZwRgeGJVOnWTjp4d3esuUCDKfH3J0prGaSA8TdyUj8vD3gD2i2SgTbkUjVUbmUuW
GLZ6+UmC52/FC5OBDkT+SWJEIXqkX1iK5x5OiL5UHR8JjWS3eOt2iljcpjCutmeuUENHFghY6jPM
WHH8vtdsXiR3WHo5iYrQ0RPaTIDXAjsMjaD4whkKPpbC6Mfuvgbei/2jYAxpoIQ8+XI+70brrBU1
yzuVNUpWO3MS4oC4bhx/AUbU3guZ0TRdTRU6FF71OV705qujN5t+TeG/A9GAqnI/DT8AS49B+D/L
4R6LZyZ413CRzI+t7M0v2ZQCxv92oecqSh4rnmXKq/NKi8tWIK3XW0jLkPL9uinX03gVc3P2Ctkj
9mLC0x/UDBDBVNQKvnoN85drC1WQlSIj5iU60eL6SOzPEvrmTXDvIxCTyHTlY+oZUw2HbgX3u8ZH
Zh/xjGx9kGOFr3fUGqOU3zBTHORHMMYylsXmKktQATrU5eGTcqWP6DjMA8BwPXrrQW12C4R1QyP0
a8CGPgSOGDwNcGWYqnSY/zAbc/lTEIV1bXd3rMFVEPlzrYNTTq4Z/o9OBl3jtByUEUnFhFOEJ2eJ
VB6/Sr0PAhYM9uc//FmYhdvGpnE8vfx+neCzYRg68W+9xsqrqw6ta7ss9RLpteFW5ZBaPWug36zP
+M27AhKbBtXMFxcrj21NpP024isKDNZgtJtTM+u8UJgWtJXajXOGeWXJWb4KLgZDP8/Wv1BCvMyx
gq3EAUmksdeKmjuAQAdlH9SYpUbUJ5gL2PG7nqrDub9MnB7UcYC9JVCRUM2iie6+7YHUywKm+O6D
/6duKwFv6O0H+zH0gPgkXW4wRLJ+UumIjvFN8lMyXw0uftUjd9DJzGlkluifdESNj4EQ6Yp4jiuT
pNlAHengoxgLRzoz7OUtG6uD9dfFk8JvFmYRbX5k5NT5GX+JCIRXwM8aaKV1+r9d3dTIrylxvY9G
vqtw5ldD0iLi3l/aTCWnK2RgSch/bCwsyBixO56aZIVGVkJ/rTidXHsOCzKUzg4XISL5fRBdIUP0
J//glU6lam8fiupe+kycRb4hDIcAOfO0hA3+f+EpHwGyhKUS7QP55yK2flpnjgYLpTVTnlS+IBsD
A4eMLV19oXf81AHCynQwZpuGscP/4aLC2Q4NtfX80Pz7pMTrKX62RLjcNi2wqIKhiEPGFDVqDOd0
pYq9lpD7rzTEZtaVqYHboUjl44CKrgjBGaBasW9IemHNxH63uhrh6DCKkZRVxhL0Xt0MG17xHgwT
DMSJXdMu2Ab5HE9S1DCdAJ+TZcrmCBmwgVSxxBKiRtyWx44HOcHiPgc/PqLy0/iMXb535V9biE8v
Q5VYLxKpe6KAvqNh8CN2ZzE+mdb8QJjbs/xu+R+7MVuKGFYzqsuR7fMjeNGNMv68RhZVGBS9Xhcm
pjjb1L8Rx4F4pYWB/zp1uJcfIgon6G9tfLf5sJdHy85Kr6Hx6yBHdpcJeLXJaHxuhXcf+IolbAPl
/tp9VtsU3M/XT309wJv8GeeM4R5fjVoTAEOxIY1/uBnJNlxUKdDU/rvDUKuvabFBCwm0TkhAdmR5
EbAzGWhtZsY2/2TEu5QowJ12A66X1nL9JGrpQ0tbcbY5ik7FgDHsuIHB5Fy7kZRxjUUKl3JWZeVA
r4fDHs/U4W7wYhqwCRd5eyKFaBaAfNA42N9cSHhp9ilYqa5dIscQ2kcHTFSQmBB+3htYZXgnrCm6
G5KyblgmAv3PUMyRGAEu2ek7BoaA7cx79gQSqhBnNk0mtA6J/dRX7NJILzKwOpK6NytbRBju96BX
DObOSxSWKRWaCabCxEg24TENj5LhwJZh8mlkCfMJdLudpsE05ixk01qLJMrZrXfRqlnkNtV37YdP
xjoyl+PdXZzXR/1mdgXH40gOiZzM3/2bz/+o3G+cc5MaHfTq13oq0Ejowj1WIj8P2uC4dRhmCXnb
HQ4L8uONNxkweNgevrr9FB972nqG+Az81djXgPOxGzGpReaZOXgucKBYcZa0rswuDOfgEfLOAlP9
ApZ25FARWS2If9lDHSBooksKo4JFMTwRjC1/oiYgxjJlCiTT5mMyae92kiBBoOTqqtu7J3vPkWXh
4nYS25lDxKojAbu+E23IzH7JHDlBBrnfAydIBZnaTSdDsRUCgRM8ifzUHkVq1VJzdympc0bUEWXF
YNOmUa2XkbPG830Ps8qH0YlXM+pUs8evuRVDK5qihme6Oc8KkZlQOKun0PPpSZSMIeuukRhrdHDf
lyI/SywmClMpymd7SxxXEUgz8tE9lyS/ZNBHKhTu5y1hPXWOGWLgUKCHBxVXOD1Oss53so7DKUxg
w+Wx8z86eCxrZgDI1GaGPHI+LkvG4qLLhN3FTelOjUb4gSVcmPmSeJ0go2UjldFFrGHAw48KQtXR
TSBJTZOKLDByYIaJFRJsKhOawySFAZwXb84O4inI36oPviEwE4oj456Mhe4Se1c7y7S+rVtBz1Vj
TvdEWuW8eX+XWyzNe6nwNIXwMznsC35R2qW/eIXvTKhSDS+Calg4M3KgimcEbtKaYuAhuV/aCnzh
cCFwecRkce4E6XLog3WnqB4BFrIwKdhQ98qaU5gBtb7ZrfRpKTuV6XxW7IE3HF5K67f9vcmzwWa7
pOlsF6AKM5TEwoIhnFfNsbfzbmQP10FcD7Eme6lk1VrzjMk9vR5cNQQ2KCcyhAnJINDvE82Mo2hY
Su7uNq+1PbsZUoYBCK73TbZXvkX0VTnd1Hh2GKuWa6K8UiJzhFt1z+36hTfYkNkjwRcHogN1ZEiU
S3FpQsIS/ZqK2XAh/hxROxVhDQEmyTa7kCdy0Lq4+AHuxahIzVwvrnjgkJTvIB1mJ6gJl70wMvO3
iGSRnMZmFbm0kkQ0g8ba2oY8DBk05kEoVu0dHRFGdJVLxTZzbxL7C9YC/bTfikIh+6R66s7rqF55
fM31Dzdd3jv68AwsQVPQ0c2YQYY1fdwqqRR4uraSZOVKedmPL5yd7pIEMk8tSWbnyq+acxb1KgZG
FbikrvwsMw10mcz8PgJ54G0xL35JlZ7e+vBWLqJXPKmKw49RzyyozkNKY0bro8OHkZyhuwCE1/tX
8Z6YgnY9SbmO/eFxEIwnQZmFuhtkvz95Jx+2GAodWXhcYoq1dwexjhQL5UhpvDWIafBrcf/AD8g4
BN7/y+4MHyhbazNZDOmMp4H+IolA8+hK9GFf8nY3XZ2k4D1/Q8qtfhpA6I6Hf5YLVmGVOZyC/C3A
uPrchk6LwE4s4C6OcNbR+LtBsrXovLO0AhBScPn8kKFNXMva/MlFv3lO+cBOozHl5LBSbUrJ/q4Q
Ab6vRhBlSqkDUZ6W3yPAFY9bFqZuoEb0ulrV9VIMn3iMtBLznhOFK+vwWo6vC18QDQWUd6loew7b
pIK15Dwfw4+TB2pB1b5M5UoA0PtbXaUKsCozR1PiP12HJpWImC/PGwnZauIkQHs/FLjyGT3VmYTr
NqOmZIxP8kfdoY7ATXHarYvEbHbCRJ3LK8PlqCtEm1kX16LLefVOvwOB8ukajf9GcVOovbZmcrMd
D2x/JKhMfpbmhLDy30qU4Pjo+AwAx1/T1kJaZ1ZcBCkZmEtticgukv42To5DITQkvvAg9l7RRF3e
wIMi3p+mms/+px3Vcr4aA5sSywNkWbhqYQhHVvYUJlAoYJBE3mFt00wqaj82hHI7DxMrtjj5gTM+
J0fAWV8SPuX2V3+3Fv84IgosF8EOi4M+boAPcQUXrrx6bICGX35937uQd+cxg4KKHXRJvqUyBGDU
hdWDzr9Qz3JPWjcC0bx+NwuMuof8/D/d8wp9bW9aBk+Z8PbHcxPFdr29QjKXcJXXqN1wynWuutxg
Y9Xq/DO4Nx+J/Ks5J93uyq99klIzUn1qnDXiAseAgE1R+oKFrZi8beYFgaYHSHslbVimPPhr90q4
vwKC6a3JJXDCc3Cdk+jlHd/mOo8/4UUTM/pZGVhrxSyWnA56RRoECBsspBWK5JalPyxR/2G7/p1V
7m7LbNZHVpIZXH64xxlSHSuL4iEz+7QES3huck6RYb1xEWXzMCbJWa/6DBA4/jFW5x/LjNQZPLQZ
QMaBYS/LX09MEEvHZvZO0/BXY/746CCxZIGCOp3k37dvlnzu0LA4eUvNHmXk+BZqa8kBTA+sXkRg
0vlYPaho3Zpu2T1RY42KNoo7jyXHmRgwOCJG8MOFKHTo5sVywdCD9i1nwFgvsOVkA44r+rl+uu/V
A2htkVYZwQo2ekrYxiaW296KLQSRQOoE35SkeDd+v117HI6ZaX5t9d2Ebe31knDs5w3bbFlBIaRp
/fep2grmFjOM5chjTTPUC6pHFry7S5ve3EcPvVp+KTageVoe3enUb3a+jK5fvpTXuGjO7DsLbSxj
d8cbszwEXhmICK3vVYaNW5+QMMcxKCxG32Wvr6BX4dCsbUR3amhqe42y/WrvB1BXVbd9dqzPXVzQ
+ZewOLIMq26LWInqO9cIK30CkKGqUZb9kTyFCAivgApNzF3gTZH/RSeJi60WseEtTMs+VDziWWQS
pBDU3WzjFkfMdbnlkoaPtRYuIMXuaNSXsKUImAz9NuryIk/9gVL+lto9qMy88Xf1SnITDyIcuVtZ
tEjjJCJkCNP6Ja0pdhWzgpvp44JCnm7Q4M/c4yvGCIvp0H6CToDlEkUDkf62XQTFnWPyZPUriDQ4
Q5oWmAnyQuvwGjedOeCle5mW9xBhp90ERLnTL01qIIzJufa98D7EAXz4waPdYqVN5q7NX/ufq5N/
Yj/xQWWqq2YJb6Ev3mXegPNmA/NhaRsg7U0EcPmCH3K7McMP/gPpKS7ZeQGxl1VO+3LFpoytUuBa
WfhLmkp7ZbI866WqQ7RIurSoaZ2XE4MH/uwZ7EKrQw+3fEPoxtD9yU5gYJr+hdMxtOGWt9alVUSK
2tLONrbGpkLcGsgWQbQUmIQngWAgSIddrIHcHTPBL4fJkxffmwv/Ag1s7Xl+S4659HioO66pJ54j
fRlb7Mb1pJB8AMPTihzQNWZkWk+zSM5HWS933HARE3xHgnILZzK+zsI6elqbIqw58MPYyRRvlHTW
L6Em9fAmL649pC6H4fHGPmnGacvAz6O7Bq9rRAHTEPniQ/lsOULFH+V5128T/CpKeDD7MtKOwwqX
X9TxSXVBCbAjJRQRB7cilcIYqcfCx0zMrOGxnZBpRjPpVZwfZP6W7txfYGsrpmJdLxNOqEu0vX7h
uMsOcn5N0DdBlClZLdiKoL0Hamd19alK4WHzkUlGJRAdPfFGZziUCMIiaqPpV/QebiJw3S4TduIK
yFHkd1/FJVP9UB4Azd4Vd7Ys/M1pDXDsXysH+p3Xbkva9lFI3wkoUhevlbkAONfV25M4GVT8Exz9
29hSrwhQAAXaEJ5U3PbjZAJvyPIS2WIeBIcTSSOJJdCBTMhT0jaVP0iCPotAP96S/N+65cNlJLZl
h2GFrYc90kfuomRdWCrZdwNoFWDciXA6N5SlaxIOXLqjKPmkTcbZZUQoCM/dqqE7QxmPVu87Ijgs
3ZANR4aYFd75niGUiZuNHHX2w75SJJakjzWU0j+lt9soZDxgjN86XV4Fngjqu61MJNnBRUqTXjua
GrBn5ta08shceelo9XzF8zYlwfvb1SAq+FlSHL7MJXFdVw8B3sd0EzoJNAoVYrIQbYEciX5MIzIf
U+363lurgR37LniUgrdnD4lgKtx8K6pXABN4ohxuvUqmnC5qSDWqUB0sKWO8ucgv8ker+oPLRP7j
iFeG9vImE2/ll9ym4etfTl/LaG3SAy62NQ7GR5KikynNZ3fo7+t0bd27ToezPEHyUkGcp4/mSvBU
zCVHH7zriotMj0m0IYRnot4elmVcB3Z5hytM3yOoaP/NYyEF4hJwIAwxonCtu1WIriOS12Xdzd9s
OiL+LQCm2DZO/ZhLFUNiG2ZxoPR8MSYPbpjJVR8jPD8byhU/P1fEbvUYDmi/uIao4Bfw1P965Em5
gIl0XnzdAyqjlsyky02xUqewg+eUyclVnEPP+BeSNYKtPg0br7UK0UJ+87J81Ii4LA3e24mHCCU3
PfQWHhgUOMJz3PpQAFLyWXE/AglDsuY1gBFqdAr7hzbSvnGH5iflSHAAqh4YXy40G9Pzy/6ixdHZ
OixKIL+lBQU7II0gK3bffMLlf3wLGPupbE2ZiJvMCqnnLLlSgrQm//0UYlkaAUxwLNBZSdonK0eH
wtUYdOlicP5esMoYyLejYGllC1aCMsRUGuIR3TA7niqJ+2vmji5e7ZDOeTIKMBwO0UOMnfia0GPZ
GMxhiq1ZerYG7w0I8AatRorVGJ7h5tMp/4Sj8d9TEXWJybNg/i4JbCtoUzOFAtg/mVVWoJgMgiLe
+qOrf1i1U6LnSp5nTCHNb+1bsnRrOwFDlAcf4+0J6GnwRMfRIpjIvIBXwLcTaX1eInZ7MoBY5z+9
ZcQ+rbkTzyX5+f5hxOqg9Ywn7gswADKCHeGaxnOclQKvB4q4+yBTpsxf4GQV5ozsC5NR2FjXg/kU
CYAL2uMeqz+nckE4DuKDuhY8AhHpnFIRO+Ny5azjJDtWDA17iBvFzcI3GKmKEA8ihzOuBFMhhvJ2
osY64uQ0g2mXOu/v/+X3vfbpQPVD3wLojU1kfOa1VbOu5BulrAj1POjPD2HBMmeEa4rE8BYw/IZg
YCqULkneSQchzDYpbbVwEbJ1mIKpyaVV8VOKSBkf17oZqUxcZ3iM7wVj67AAPCoj9C/SgAdpEMWu
c++Qur7VKUROzKxohYY8Cd2W+OBaWkXKhEHBX4x5R2JTtPQoIW1cC1VMO01YGCHsPBjOAbtfMBtD
Pt8gNsOzfLwlkJK2BRn9BrGAee4DSUxqHShUK4uSAnVvmd0jR+MSl/zvIulMsagHDmpFMZSnAFeh
50Ye/bo0gCcSDbjZ8zI+2nvbmv8gArL7z0n9t7ytqZoWm9sybRLklLV7FVPfmQwSSebbQsg1Fq6t
zVLPVdnelledh0nk5Muo/8wr3JRY8d5NKrjLuo5HJFt1yv0oC2GsJ7YD4/Xt+BJ6VqgqTsI1wShb
Cn/3w6nG7V+Pz95Gwv1RGesHJAGAfxP1AUaEpQ6hPm7iyhhTaon8AxuYAnCuAVxaMxWh79SC3WzP
niIfFaA9chP6wq6VH/GQPK85Hy9CKc0VjRD2Yx2GLbXRcNk+wRqjdSHFGDo+SBmIT69OkBavtjSn
claNTT54CYAkWpUS1ZmM9R7Be57UXjpBoRbYFn4VZV2UcMXxdX274Jk+VchDUfIOG2EAtUMw/Io3
PADGzVwh2RoiCs/nEtYLFWThkzMSqQG3OwBcCyB1xIlZMDz9YEmW6tC19J4tU7nmFxj3e2uooIZ6
1G008dySdyVbR0FWesn/J/TYcUgi5VzQuRQTGBU7pS2OB2FdZWiQ3j/nkxcc46GBkj84818HQC4r
/sEq8AHG2Zdp4HK6m8pWKWLLD7+041kdXU9CeeIdFUCS4FCIV5cg0FNSUUUwogLEUGW+G7S87JAp
ONZxaH9Ug4mpYDLUKUWq+EKuh9SCOO/jGn3/PSt4TuA2zRhSassoev9JkX4/K2a878s7AtoDymOS
RjGc7B1HnJL7+7w2830WTz6gAvotUXS801GzypJ/Wjl+5Vm4Io72NGn4LlGos4LAY1LU0Pc8/WYX
B6IXkAC9gTedY2QHhPaRK9YAtIT75vAsnlHXrWUMBI23cNkseV0AlOBDypt8LN9Wm4ZyqhY6YFvV
ukW5y+FY3ReDW4ZilpTxWoQW2mWObKyuWif9pHBcBGL61n/HAuq9qH2jSa3kSGT1TwvZO07xHDij
EiwdVrsPJjKrxuUITGlCjgvnRP6WNFJzPs78tQAbLxwMhA/FOSCqfiHrNcyM1ZAzHLZSzh5yPBtv
flW1v+XiV64z9Xf2seij92tU+e2HlnQKkDjDzPaIKKSZYGvbZPoiq8cNctZyxk5XC7tkMtL7l0te
pRbsDwCm2IYeS39sJGSCQohrCwUVsau1E1e2xmrnWdkRwjt162LXU8Y+7o2tCoouvsI2+zguN1WV
PBSc7vYaqmkJap1vo+FoZWc8979IEYf8mQMkU4M3PLbrYCjDLrRBxNq6pTQ+aKk2L/ehr3Pp3Hnu
KRHWhNRZTy4EZWIHgACcVvwMMQx8ULyPAy6Seu4jMV95dOf/GooY4wgRCh/RGNQEMrzql15C+gZK
eOdsPf56tWloeRibHHfzlbi10REsBfhGL/2Ajof86FP9/4TYJS8l5xQEtCrqBk4O5v9Y7Ci4z3GG
l9FwmpZBtSqyp+Fm4slXEDDCiXydv3by7gSUQO49Fp+soQUjgG6dREH4+rjWKNwW5jvJcShEiCaC
ICkS4ZmdntGaRJbAhcqYbmN7NP6Rw4HJMSYUM3FdGPlaoBVu14+Y1FAuYNmO5XMTuhyZpcrawxTG
acw8kLKIuVjh/y7UUYnN/1C1fMBqESPJ/OgyM5yVpXQkhzLwxpMNN0BEyrAxo5Ze04USI8P8I8rF
/zJQ893zpgLugo+cpfu0cD9wjRCaO9otonIUXET/L0vx5DsjwwoU5qw679xgjFnAy3LnmZDkY/dG
uQrojCrv6ePiaqEeLL8rWaVVTGH6wpvGkNst0JKvKee6EVw8TOzzG9Clkd3sKN8gzvZ3WRA+RPds
N3wnBD8kixvukGsBeFpOVuhjuDLnc+EWrGAbnBNVCfNjOvrcnS3gYl43K4sNqI82F7kJnOzGTFac
NUg8fkvPWiFNJYkVJgLhH2XgwQ0Wsh4HLXLpT7I2zPgt7XJXzQhKZ1x8wKBT6iWIemsMiAtAn+dJ
U71ywDbmEyj/VwUU/8FSQE4EtNBgW70htQ94YUuFrXCTTdK4DJmKs+5KkxGz8d0q56CnXyJprvyh
FCQs8dJBcU9EmEuGy3tW/dFSEdDM90fTX/dTZWGIaM2UrNWZT5TaRYe+9tmHTYiypRWpvfM65Y9+
6NI5HMrDIYznt87T8kEvggGTW/c8TQKq1hy+cYCaP3kilBcB3tx1ErkNS3SxTVkrw7xhoss5T+Vc
ejI1AxeBs09AUJ+JtGJ6uB2Gj+U/4fH8FkU0+ZHvOHvMZVKYBDdh14tjjF4RqOMnKqSYnUHqnKCL
1IbZ6PKrZLGC/NK/LPLaDs+t63uH4Yjuay8HRMZXLFa3co6LJx8Z7cVOpB41l84NusJvs2/SHu6r
es4iKbkr57fdTvolWAHMlpYguBfz2TXjs7E5QFKSXYL37HQ0K3sYZr/e4IXHapwvWPLzT8GH0H2P
7Lvn+WkM82sC0xhc64dEAe0aUkjf2KuioDhewin5+O8GdY3gTSEI1sWBZjENU6T8rg2IL7DVzQQl
DWFB6WxinMFrgLwxcVCbtNKDE9/UUjNX7p38in+zemeC5cF5s6Scu/HLPlV2DWzBF3kbF3L7VnzH
TnUP2zIkBoAkLRlJFuFzj53qU45Q0ERuPGecLUHFZdTAQCRcjy0gB1tbKpNDNroGPu7z/xdqCcqR
Y1plzvbeVZdxC4mjwiaDK5vKqxNdI17YfX7heANjj1vPLGn7EOFB0oauyui+Vg+2Lr4srD+s7E0F
MQ/vxZw23VcNC2h638prdr8UkTAs8OeUNW3jdabLvedngVgj7uSQj2ZmMsAxzEhIGWRGu//lPA4H
fRGuzVTXT8FRvk7PUKFam/gAYQxbIU9oC+9FRqAW22lhu7+RNZr+MCriEWWBp8PGoDk/zqrRZVH4
+moNSGKL6jgtKJEqA6i7fKwNxCFdC8Aau06j+Yx5Oa/EZRiuGc3V8yDkHLAK+MkjlTaceRSMlT1M
ad3PqbZGcbqLGGWMpA9OfC/w+WmeeoY1QJqeU/uV2U6TWeBgCEdDeW+xmTmsEtgf9S67+LxJmjmH
Vy08zt7WtHUgGa9iUrmQTJ1+mBMpI7QiSWtMfwy4XGA6MvELUX0VszBBSRmgTYfyPSnbGrv0tfBy
KXDJI8sMxacTSTZmbsM+dVgeTlFOxtzMwH26nS2eONh4f3O0jQoBtucQeerZ46MRZY/YxduhuUIY
oLY1jw0q8tigmYI3w6vvxut3pAVkj4JQIJxy5h5LcBUj1Hm9xbyLskLRUOENl5kXf5NLXTzg0TZU
XzDtb/U5pCkk7LbalIx2t5aWyB2UvyRBbJZ8PTHA8g3aurbylj6ppQePzdWqqAx0ouH966VR9WO9
JMaMTdb91SvuHwuejafWlVPh1u0vjK55HcxhddGlhK/VuQnyRnCBtx39XzWKVUt1QkugJNM+6bSL
haYWEGey85vJqIhW5iQJHZ9KjfHvjN9bnRpsELbO3erLHmgB/4rXx9G8qxfm+g+sYkACV0m4YaGK
ZymZTgQn3hlRqYl1RDg2G26fUqEB0+A6UUsuGb/y6jdmdKlh9hfXXmoT/jwo6/wf86q4dB2hSQJ2
WECaLpPPyxG4FKcwkRYfGX5vgdJhtw0rZGkZqVRUHDn3pJxLI9rNUmk8XcAHZAh8qw4oFv2bQhEr
OQMTcBMcpXjO0rb+cQLYK1I3TLbIAZCXYWYgAeJtlIj973SB7R8B762O3yeCshUejDYEXP9sqViy
ZLfua1RM2z01wv/QF9aDUe19ZDmOf5HreWzoS7dwhi987RKy0Kt6WMtKFwrJaz7z4jPfC+gx4yjn
VJI5O7IiUCjyGsLZj7TZIfZ+0pAjbVM8Vh8TIzYYgh2ErSHcj27sSe9d3N0cAcvBJK+6Hnz2Izor
Z7AZ2b0OeRR6SiYtgJQL4rdUmBXk/aKnYJSwN04956dUy+/WlQwOymm81CtTNanrxk3aqMO8OYqZ
tFmvnzRmSY7IG/pR98AcoZbKoP0MOxdvpEWzqHKr7p46pPDJplrqiVHTgXCf4OFQggtU+Qf9cauk
ssBnHDaYZw8yUvztE/S6hYTrJYH+xfFIhUXvYGmIPEwP7MpsBjG0tS3Kk1mALESYZr4qa2t+REb8
dd+H74BzgpMPfbtIs0nas/MSRAeCfWzYkaighVjN+VuQxrg1MNJhmiHiQnpgH+vkAka66UIGUrxa
3tkdgEoAYDttxCjQOBzSGyGC9DsdWwPBjWzFXEiHPF504I/ppdnJCgFngPppmSy6tUYe+rSd/bm7
duIM4AJKCwAnTkTp1BK9c+AoA6C4oBhMycX4U4/WiMNNoQzlaYEBzDoEddh6kygcvVJGvwQBS8g3
4zdp2QSEU6VP/UOksetFHFJv+LuF+eGd8gxf+mBXXGpiICXlEXi8XCZ1GQYMALkAhGoUccFxdlKu
ZfcO+p3qr/jtKtGeATpaqdBBeYT7vOIIMT0aBmvRWPhbRsfKwkxWJQiKNmrnZA18j4JdSSdW+2a/
ZTJA5SNXVC78a1RGzEOEQDk4VaNR6lfvHoNd8U6udxK72QR7ZloxPEYB8b+L/0Hqg1gmW3t1cILZ
8PtFevW58/bW+ZiYy7vcxvwztK5JxHvxv/qeZJxesUoBeYOY4qdDx4iJY1XEMlzwaBExUr0J9gRA
b0lBivlNqwv5dZ9ufl0lRjUh/1c9i2yaiG9kQM8qJqyG5tnGovL3SVgG+ImYbJfBfwpaz9ky30LG
yA9jfnWXHPYcfB2rlbhPVnkQvExmFRfwcVxAA1KKfxFMFG77PhCVvKWuQC8FioCLsj6YnLadXnhq
av3rtD8nT/FvBKaF3Wan06l9PuujAh4yWP6XjkzjvpUnX+NyhmPvIfQ4cO+XpHp2G5qMLxxp0JGD
Uoqb/Jjdi29NG6RQiLcfNhP5U6oJ7JSE8bmuGhTED76EDYGcLNpySUdBy7F8rmNrVleUnw+OhsIi
f4HhCkHYsw32MfQ+quEAo90RMVprRRb7JXVEYnA5k5HsQuE4jJk3d/v6AxII9xN+8qNsGTvJhOmt
z8oTI9XQ+0F9q6eXIgZbEUvHlFiY+zUF5B0MmmXpl2FMU2ZZxm0+Gt9XwRvMSV+vHtmkCWNf3sEI
zom4SAqivCAWPRSff5KJjKX7tbaHY5eMFock9emTlX12OKIyxPNkXW4QE00K5gm2eP/my8+hBCFN
bBz+9fMTht3aQeZSOmEPv3XSUJ0CYkqAa0k5hLHIK3UYJAV+SJidPrcncTi97yIKZr/w/xrf/qA6
0CSCce4F6mbkvfo9GjiRu1gXTfVKMJtWKJdkYm/6kiAsaCR3F7ZFxM4TmbgKVGiktmoUz4axZn5R
mDoUHp8u1rC0LBYy+NfdWmm7p0C7wshuK5SE94AnYsdNnZ8miOiEOTBkqFCu5sljXlosOXKUSnvf
S8NMKz8cojQRSHfwKJ+7kDgz6dpCQIgL1QOr+QdLOy9ESvKswBCUK9KwH3tW8h7M2j3RcxABF2ZC
iiIOB7/4+CvbYXfk4KxvGptUzAAPx+7AN0Y1BO2WEcGq6vlg9xAJeukc2W9+RsDQuISAy/F6raGn
ZKDSfy4tGjbhf+PqpW2QmfwOzhh5jr7l7mBnrHigMv9MloUd4S7zrfTl/jKMmiUys/WGNuVdwK++
QaBx+VNgKtiIU7HNxyMJIszVCuS5HuikRjDsQ4e39TnA+TR3GNb0NrrlPlHzT0Q4SFxZ7oCLYtom
2RrDrJ/0MVdOrUeuR2gfQR8Slkk7W9PCcqrfZaZ6DqTOHl+GhzzYhy+AfC0PiZiP0aIW1/Z0e6sP
dvFfsPMzUKvAwa0jbhWfL9z79l7PNTRm9meNH/fwI8VeD7qxXKJ+WeV4skfwDbrDbdfxi9cLLMyB
ssIG3UBzihAsI5VxG6Ny+4moVmm/I03a/s9xXlFFPxAkWZplx9oYhwp9fVJNPFaC7sI/v67hyUz1
HNwGdOc9rtqWf6FyFa/O0M02jFoesP3GDrQFPdWJ6MmulmgsajkoUwgasfjMJhjqDyNzmJlAgd/L
BvPOKnwDWfHMCmREOoY4/Ua612np+x3p40PLzr2o6lfiI75D54NvCGdU0VRm7cJtUg+cg2Cwz3EE
BtkraJqmdHEf6dUvYNganuMz53r3jSf9heh4P8RMCtBHafnr8hAPOKNYTGiyg04fGVVa3CYt6b+L
roCv0ANV12amzXTxqSx7XDSRfSX/SEtCPygTpYPmhbX0/a1XdclZCTJlLv8B54JgYX308041nWzT
09WVHEWCzHQmEIoWwzPI4sCHGfvhQFPk9nZzMqGPyznWvPhH6Z4Qi+KjndQrl0Pungec309+R9oI
yOFQbCmVAgGlvoVWlGqNUGmXI/YWAXaP78XGgqkpexrWFs0nB61mI8Z3o3YLw0Ri9BuVWmsQbAiJ
i9g24l4IHcJRPw7dDF7vLp3cAKFszTsg7MDgMv6uLZGbO4EGGZD9nG7qLJwbA3+0TM7dOhl3aP9J
zQCBpPa4X4XT/91CgfTbuseezTKyYPe/husdOVS4xzGEN9wLCvl/BTYIKOkZ8FKubwdEdM+TLjcr
kRGXZdRc1Bd/dBPn7YSYIa9LnaATvS3psUwm3nUElI3S3eAh2tEHs+jxrEFOOv1nVZ4bdU1uhKeB
h8njxa5Qq57uXilKRNL5NChigK0g2pYfHk6ijdCYSABV5WZX+mpi95oVb9gW1nQVZcxgGSBFeSAz
piT4FlnG5wGVo1ShtZDZfgnm5VogwVtgPal1zVNMy25ox/QGvEwSWGJbOW8mo+LKIZ/3e7Q/wI+R
p/q401Zusbx8aaMIInYtOMFX7WM5KLfBR8Mmk66tcRKVy+TsuM+ijl6MNq4UoR9Z1ZaU0wLB2APU
bpbwMizYRdipNqST1Z0ezk5HnJQCjPMo9DKdnnvyUqcizVsm0ig5SIebovwOqpaJeESTmTkfKccN
S0SnnAwWdAz/O/etTwpVo5ReKtyJ3IbJrq6TzQ0XdQ/UsoWOteY4RmTSmljhm0AJ9hfVBVyUtBow
b5EEzel/ppWWBKNzoibuy2I3yamEWbximJ8EQK5jOz0Xqha5faUCzAJr+XA70HIs/PzxOFo0DsGX
0CeF0puQA3syM38lFAjB5zsLlb5VAir64SS1ATsBPkHolK1a0EoWMephLtrB2aq9uzC0znNoxH9Z
ibOUJi9GWsaPmrMmvXOhMY1aziZZh4i2nzaTNF1jKjLWqO3b2o7w/Mw3/HKqdwVfrDkQ6h+Oj8nT
WSuDU+5+U0y4yS1loU0D5aci96MvIarUXAVMh6TT8iGImISUSEnIRhxneD29OMuM+tJu0yYKNJZj
b8hPVV4EHeYzMjhO/JOsJOF+/+EmLaJrxwW0nf/3YOIiFkRPuNynZiYb903fFrrpVhTH0DSyEtR0
30PUOuHnVUM5jRLxjy85FpcyQmbfT6GT+nLnGnIi7GmMJJ9z0+sWDSecRoy2HNBzEXW8o+JCRhbE
dFj/qqxnM/EIlFiw+HoIQfmn+Yth4NcvK520EQiAqTihQdYXkId7qhkRufLx6Z3N3cuE8uCownIi
21dqdpPplvTyrczP/S4VF1jYSft71q4pVLzWl8kjY5eHfy9ddHw6UsUnCNABC+mfcgU2MXVzHzjC
toChRpUvLU0quVoDu0Hp4gNqbCvOWUpc1Tuc+Brq3a35tjL0yfQ27noSVaMP7phd4fBSsBbn85T7
2QZ7pLWS+4QU1blVF55pulRYI6mIhTcI+jcN2eSa7wiv0cB1b/nV9LzUo21qFBvGq43EHrncAq6A
n3GBOCX52z5DUbZn3yNFPBeAjBkWK764eJ/Trjq5VCS0ds8H4dHaAxA6m0FBCDsMIeq3EzD6ae04
a3MgNkpKpda6HyEDFOSlUFB9A2tfKkd0ba2Hky0LaViJ+Q18Q4eew7c2yMCoxuM+w9c+j3B49usQ
wV41HhgC1+ams+WJx4HFmTaK2FC+c/hulQKGCBz4n7h4N1FokHt9rrXlCUMRxmsZympEKxrmSYVR
P7acxMgU1qAJDvKiUeegzvm30Lp/7i1HC6uM9tuD1QTXnbBq0e+iSOBw0LDIZEwA1rUJLMHBxLqn
60c/kMTc5AdwAQqSnXgLWmuNWggQYgUEHIE2q++PFoLFnK+UzbdfxaA85MXcsneyYDOxGx+PdgFg
nLOjdY1wceYCWKGWlYsY4NhiRlv7HjxZySj6YVSTeuOeQReejKfTf+YmTv4iTZ8b+v2eNoUAfBEs
q0LtZZZTkAZJWwHX0U/dIefjWP50J/LHKOy8bTOsnJY/MvH38UlolZCeWQznW2tljBAMvq5JgfVX
nrJrgZ2+Ykfabs+eMnKeC0TNphvRuiiB5h7KNGf47fC4K3jAEBCa+1y02hQIq6/cZnaubL3+jVWO
BN05EmOPPMuTa0gMPi08TdzcAItcj8dJ1FhtB1tTM7B8LR00EmmfA7imIuKp0PBRU704xpwL3GsX
v/jBjYAJc8UcmbWei0xE71ZpwpI16+qCCdWBscHbLBix/0IpmJZrO+DyAGnohbCnjYjKE0ulkdCy
o1brKTRFgLh7bGKG4sbcnMOvUYxbTeISoLNA6bafkkTzoJNEgpc4DWnPnVXqjY0KjxDAPgfVxlfT
gTs1C6IDqt0whTtdMQ39ANrVkorppoF9VXQpyk7FLxcjOA6U2I8XsjSG7oCJdffX3a6PDYdRRwKM
vDsELg71vhGfnW5KjOs9/uRMycENwfztgoYZHGfC1yasAQSp4/nACbyWbm+wM/urEzlcT+bLKvGs
wM3XoOhV/AF8L5IAzgnzcaDwxSXWzowNGBFPEfAq2zwcOju71LnMyZgdf4GOXTLjPT+BxlMk9EAw
5n3f9iq6lAhXiegqIQq8F7d+ydnT0+SMD4uZNqnOknVIQ7pJguoHdJrvxSReosFrRBLq1Hf804lG
fkLbrEb3ym4XnIUGOFTWKpzpae6OeG5iFL/urgPE7EU/dCIRrs6sE1CHMcNHeGPFPvTyuFH7YntX
soKZ8Bc7zp0mfyDdiamo5UdrIJQwdruJ0bhgiBieiCSMeAK2PtHofKDvZhQmd9ScIkVUqyT5P6vb
SbFC3474cX/4iJgNdO7DECHRDXPdFtkoqqNzoFJUXG8DQrXj9fRw0pr6SCQK1VJqRYPu3WcH8XR5
vGmh7n+lSCPxsG5SrjYhPaRZp1mZMqmctHRhRZxheTAIICwD3b5vsdDWLy4W76jUONXNeFLuBza6
HxWQXoAMBhsvwH6fJCqbhL7LTjDkRjH3hL4ONNjQACKUyYGN/QT7L79yiZh3GLFLZYc4alu9kA6U
kC9EQ/iwMKEPDA8bBLe5dIqfcPDAUHSQ0i1EhAQg0y9Q36xfVPJ87W5mnWQCoxZPczP1iEV8HnuC
8FrmCmSwRY5n6F2HmGkg1+Dvvf7qDub6jrBmuUwt1r8nUXB82zG3dFm6mXeqvceHcUP0oxyvzWNy
9Q3TcjttN7EvuXUo9VXpBKuu4vY2mb8ZzG1A/Vw6mF71OQKnowg7kl0GJklhoeyoOnuyYqOI+Qqz
Ts1x/+nrtJk0mhCjsAHeH+aay2/NzaFz/lNvJN2GoqO8dYBiHscvslgJ5l5BcvkR8JFpsnMNRJ4E
h6BjRnDCuGeQ7iDLhjrQGhseeIYEqz/JAqD+/OO4IBc4yMtBIX9QODE1MXBOYbTQbTP5oc4vRC3r
TP0AgRYx6I62+l+VSFXb/EhaXR7fsVMlMSz9PRuKPH1ejqWhy7uuktBgWYz4/XFNC6yBhkrv/7B4
87d01J8sydivsGpJIQC71F5uuwKEgweN7cYlhOOroLj6JJv6hHpSk5gh7OfjyaHXaXtL99tqXkdc
zXbEIuYjPDGhUwFOXv+OtSlBEGEFRfNIIHJg6cvmzN2/6imJO6y6pTz0ZUzr4P+cMoGVcA/AP+KV
4oNjNLbaemnkEY3rWUU1/YxFrl24raW+1YKvwp5/yFzMOWNX1CPRCqwR0QopYqdzkzJ0yrF4PeAn
YaB18KRJ2jibVXsskkHcgsIypeoEkB9K+MWvd6OUFec/xCHzygtHWK9HPuWWlmi2/KMAZmnj7rBH
8AjwRlxdDjPb/RXfLFNst5hg2OdgpyFRdLRjEaWFxyP59MP+lmKAdfzvsJuE7ntuXEi3r5bAL2jK
rbKTW7w9jHcRHw5Qa/8B1se4XX77UApub1V0BEyHLvNldCCQLyeJgFaRZYIe4gSvlPZtLUdVf5V3
eR669vwmQ7G5uIkichwos1QgjW/oBpr1GMOc/SLz3gv7M8xCa7eSJWJoL9ErtoiSJ9wd6olKjfW3
Z+pCe55uyAuMD0R9iE58zYjO8SpDykw/PQc7ZXfeTequYGlhjczdycw2HaKe2jG9Sk76Ilnwz/gV
NqCRQUlUqdC0nMu+G9cEvc0hAUy+20W3SDQggN91/w8gz4oG/MDqPnL6CcxFAFKqW4fHetzfjhM3
OSJC7Ux7T1vdHnGfay7m9i4N/Crmfv4AOKkiYRmgk4Qsf5p9/rRZgLYsS5AHwdvAn14kXO9NwLpr
yu6iimqLsXzHpnYEOefyeWC3OWzBHBwc5V4JjW/lxLgogEe1xJwpo2UMHBjqPoIpHnnXWBwpENwE
YFf7idu2u4uS+uWWPruh5noj3CsYMKAbzKcP/8VzDykC5AliaP3G2kG5MSG5Vwhz3hLqSRgB6v4K
Wi5GBiFpUki4W3byX3h9nBvpOHFRT4vxs5WuceDOy12lt+4D6W7pbqmY266z5m+Pa4PpFfqo6goc
cfGtcUNsdu2R+Rn6oTJZHONk/HMsefSuL6IW0bytyIXbFRfRPaRrpSHCO2AJW+ydOQ9Zz13iX9n9
Cdhwr9G8YIYgpfN9ZtNjQ3zLFvrW0PPX8aS9ZIkRz1IzXpAUaUvcg4ZlBMloqseMxaeQhmiX4m7W
NI28i/XGhdfcBFdYFhJcig/FFjarv96NO9PW+m9BcTjwJ6j0Jxha9kFzW0UelDbODKgW6fRO94Y3
Ewyuygu9M6+UEui4LrbMUnOxggfXVmKsfKSreDU8OFmVFyUv36g6Hw/kXbL8v1yvXgJg7SaPXS+f
2oXU04OXrV+PybkHQURrQuhDiUQu6vtHLjEJbfZmwn4V5MT7JbB3iyp6j8+tuuz3fr6ycMgdArMZ
LhXsgbU/JLdM4qsAtv1tglChRafk/VnS4UMZB3K5IfWXjrVSylaOkyxBFTWgfPzvTr36+QPrmXoV
+w86Ijo+An1ehDNZknQVhrjX3P/nIzEZt1QmCm6f61l0y8VZyNLcKq2nLle2/sHrAO9DGyp7Gxm3
aYbeahS7s34ulS4ecoufePyrUbM4lwGpHW19oSmKUETZZbaXF/42Vcxx24OOBmkfise3vvSipOcy
5Yl20mQF01Xh7UE4h478C8hlBTG086Vc9sOhFRHlKYsMckSUHnS6g2ZwXeePbi4A3xkY82qyrhGC
U2Yy46ppbnbfJCNibYoj4Uom8/uMMef3DUPVI5hJwnjYXjt0O+urYMYcRLIdY7B0VjlwE6trHimf
hddgwCk80FRUAZhgHxtXJt9aiCPXg+BJ7Oxor8HyTA6WsuBVAiNhtbZh/rn3LwR7LjnuJyjR+gQB
vGafmbmrYjmq6lkPYjWYGRRV790bREtRTkfc/rE7pMb4YLidwyLHUURH8oqtQTS1pEvWprWLT4+7
KaWrU/8QWq8CZ4iyMXACSn+AnFYkSJ/qT1JEjejc6E0GrOYaHUZQFxV+9mRT2GJELRHjstEUrfZy
FerVMjx14E88DubHv1ne1Bj1cVyeLOjFFv4vVG4yvPQjfb+pVzvUtybtxTotHArOIRrVNFhs6f24
s2gXXq3PtfGSxlA+2rkpjXu8U8nCk/0pr3HvcPXr9r5wNdISwoniTJhZ3GYXeGEJ6mwzb+MRs6PW
dQfq3NCoJpCCQ/FLp2AccXln/kOzOMf0nmGeBU7J5ia8gnOOmdYDbYwT+HZpX5pCLfEEn17Qdf7P
W3YypmPekWtqxTmoJnUG5Cxff4wTcGxQG8cJmxvMBYnPYO+Qaf1xz3YZ+UhVnoaZDiudzWm/7NJU
0iGz6YhtpzYojELMTSje+8/JcDUmrZNcefQFr1poDqquwx3+evFgis1nySZnpLWARDMS6b/zLwKY
nLs9BFEn2uFNtXlfVV/vz2ZxQQj0r2p5WWtgtpklQDu4gY8vl5CmBxtN4QaEVjwtH+4ipejqPoa3
kT9BIEkvN+eX1u+AzdNLDilA0eVWKo5kajaV0C0bBP4HOhrYSyOqtnAiscY+8LE+jGxCwbFa99t/
mvHoQ1j064XPU32hHS4wct6un1WwZf4+RY+Dv3UveU3dnE0oWZuOKPp9r5VZB1TsYMqoJ3LoqCi9
OCXGh1H2niIZzPyJVL6NNXZONuXN5uWNIBgvmIIe6F17VK8QxbnBbay9HHlDKPUeT5D/5pUwJWzW
+GP//0pA/w3BW3JFvuKdKaKZ9PQab69arSdqfRBkLVKBv43Z9cPHTDltD3ZIEx3bQ/DOXnpaGb+L
6FS7zhFdCuUNugZ83Eiygfx8+YOxPFLwpetqi7+0HMHDeyOr76V1kGqBeT9AjeF8GIAXLEYSQV61
u+aVFSl1mZkxRjwDtE19ZoaSvktxrj4So1uJpFFSNyYp9qrPEizSq3FILzlX534EcZI31PRjnkMG
zUPTtyTzUk4izDf6LDeLqSvHh1P4+hdzKSBbUU3ZLoijr5hkK6MkLku//JKnxp15ZID+0/a/JuD2
jsOyuWaDoN3tjXnQLC1i58m/Y8T6BGmvhUX/rsLznEr2eWuJkQbYru2H6RstBntQPMRUnRj+ToWp
jxK1UjMlDGLr1/AyGxw526vwOUULu2nUzXnf/0SHzFMZMfwUtTFgSRi8Jgu+nICPgNpyAoSl+mb/
4d+VPZ2vIN16zWj3zRAbsX8ooX2oSo0VGwb3M4IRD0oj2HHJQzl42ryzou814/c2X9mYBaO6JHGC
cX1N21eRsHxqPWdo/TzikiW2AtBlKtCcmkkghOqJngfZvdpmrYk5wrJm5HH/A86jN0n2++YkyApg
zJIEH+2wAJ+WYtJyfW7aXy+mnZyBl1VGlr8YzuxTya+kMZUhHtENbbm9Wfo51Rp1GGd8A+MlDKgB
vWzRCQYYA0ZPJ0V/VKVPKiJO1Q0aH5P12wUIfGT+evVldbCBpYboe6VCmlVK4Kc2tAOhAZO4cofl
7YMPTDxbxowRc/CMpxBfM9r8+ASwHqRdZvaKhkHgSBDMuhTwaM4h36+7PjggB1NsgISXaZkjR6CH
FBRndY3sLA3aggt9RTFQ2N1bsKW+v6kVP3zQ3dgWQlVoRY5RVxYckzstkHIEjuaPpgArIROXIV7v
Fo8qDIVGaM6nx5ssA0KH+6shfbZdZV+Pfk3RxrD8cIoeTqVRNAjj60dFnC+iQO6RmljyGqX7rmZ6
Jyo3H+v3NIgbNjh0DVagTzWmki5QVw1lqiL5BsGKpJ6WhnAY1PsBMXdSJ8xMLLvovOyMj7f+otJr
nRoeGXzwE+jFDwjjydCi3ZbmP2m8IWESP3EfVNiCxmXwU+pjp3W9LOxpAC/A7UDOIRQ+TPxTgMoj
jAozBvncv7ATsuzIuv+vCyZjewG8ovwddcvhOxoj+FC3KYeA5F4TlLwFn02aYW4bXaU+o1RbLYue
8vAk5Rk1g2ClB+jDUfxhDk7208nvyVex2wJXspA715hEMnbtUudjQ1ywd4miXTP0bV+n7piX2kd2
x/jNhgUQS1fxT0V4a2+Hp0D7xcCGfnVbVTDKz6Zapwysj+lIm5ZkOotBn83B0jfX9n99MCvx6/RO
kzx8/L/AbTimdsRigRT82xWNnd2pdpfX5o/KEn5LqJfKxQ8GyzP8HQtBb6fVqsOKZKqYXT8OMI5f
FhcLrAi18RYKHsZTLKMLx5B6rZrvfAbwZGfICyp6BGK1bNj/SXg+VyaGJ59mBuke077xzP7P/XUd
8Zf3XsIo3WyrfYrgYmPpYKdsZhsikv1Z7MAsYJob86Kggdq4pP9NgoD5htvuCg9VaXmFWCTvzbtA
8HIQkuLb2nRt+9RiLt4OAMr1fmoEt1yvHGP98OH1ndzBD7Q1CVPFvRsm2W0iZfcffjQo/3j3EKEW
YOrq48Z29kG4UzsDh/e28604dY80Gzu0IDCFB+HXutN+s/0YIsYUjZZC5RVZA576TYoReUEuIK23
ZhcLUJnJQzjRdwo5f/I2hgJ95iBR27tPfEGg4GV4e1OWprGdLOy+ZX1ykBKQFW714jyCup1tRjIz
dnh5O2C1xIdVDDrRtYDxBmn5Cglu2OthvWxxYmnJtbc9gOumnuqQuCGRzxStiI3aZDMGnB4ceKwp
IYiiDi8J0wC3godOb4EzcmW4vAaYHr0imGxGCx38krzI7a4XtgMplwATDL/6f+Dy2FRsmmr43vJU
J3oPldUnzIh6AOMe255GYmVBpj3Ir+XaWuUg2ZStuTWESzVIrSx/6bWCaQLGRayCG7Qxr9wFLFOE
0UPuoNYwzrrPlQ5DMKS5F7RduxSWYmbva93ikyi/X2NbjmWkC5NYYHdsAjUI7y0xXgY2xULNQZ6+
UJXoQ4MG3PIzl0LHqzVQKM8SgOU8rzyOJ9rmx73/GJrIY2IjzwTk937ABjiezIf34fK5/9SqKmfQ
4X4iz5ZxvQSAZPL4cC/+uX6Z0q6byBV4xyn7E2q6pnUMc7qlUE1HR36ZhIrDLCNxFdUVWD4xaw44
vytlC4g6IYITkDhStLagrdgmBqkJ7tRVaEbgJCRs+uh77VSH0APgG/1aLufwAs6T9fjAcVc+bYrz
COTSdJs6Fih8u9M1zQgC996eokIEIK/21ltQqJGziT2Jd4k3HpC++rZF9+2g3LY/cdMTyAbdoVwh
L87niWLwx7K7exLgDHYphaDLWAm5/1c1A9NOaRy8lD5UEUAZMVz6PaPdVAj/sDtDCreD3X045IXt
2nNZZoy3DOBjt/6heWN6bnh+3jq7Cq1YXdas64nsXMLgXh8lx3ZsFsbwnna/vVg7KpKUAM3wdl/Q
OHyurFZQR/EITHVWGgS56++8VgSYXn2IkrNsxdDBPeJuUvuE4UKByALEtxtcqWCPvYrOL9LP4cjB
Y+2DN20lyR0ooQ4VbuTmHTIPADUCiGd8zwkrK1dmsguXukSp8zKqlahHg5jf9w6P88Hzf7+xxo/F
SpYWjUmJy7aF3OFGd0zECYLzOXirWFRSncqLw8D+yexLYDKeZKWp445F5WiPenEap/1/KSMKo619
5eVTgyGY5A3Q+ONTjjCFwR3Ojgiocz0RIjZZtPdMVg9B8GJPD9JI+cM+4tFFjREDgKI/4iqee2Cj
pE72VJXcFbDMx5hPDXombdj2QYP6L+czuvbgeCmDV6opQfjx5UoKKIsJbQqZTkk51RgxkDISzwuy
+/Oqo8A7tCItGQhWpMi/uH3WiADYgu+LlLT8Ap5WaAOmxueM942MV7eO3goXjy9/iDK/lZWlyfZg
G7joKZU6ya05TZcfoDHcf4Jxd9y5qmqYwqx5AtfCGLy8A1wgCRBbWVqdjbPbw0KS9YY3Vkybi6Xe
5vHLcLduTTv2MpLYh5bM0dWZqU208/rN/3smK5MUMP/4onIGQmsqFiq2I9MN3+i55xF7YXz/UZ1a
bhsMGiNoXlQaLmj6JA6Inafide6dlo2d9nPZqtl0gMDCFzhPs0vQQxEk1gOf+srxY7WXMKBJ2+9Y
eVmHkuktOSSXICQxr9+B1vCaCscaaR53xrYn0Kk1h+AmeMvf/f7TGbj9AU/2I78+b09o/5cW0ROu
UfBTEmxDOHYBNHvM0PVDN7StmBPvoSXF72lExE5kbnqcSAPv5FwHZsrtzmGXSbe0eEvfavZsfmIq
YBdA9BzsiFhPhuj0LDm+X48iipYw+QsTOXL6wFRsjf2Wp7Ulk0y1ZmREJn1t9MWxe/9uDQf6TRg2
WkeM2ogFyzcZ1a1sIaXSwV6aeyMKFOzszdLwYy86WnVd7xliJaNUpTzYMEkq6qHP6TTdpYWY4tUi
2Hri4/F4iw+pLj1br6ahAxHfeCdKPB2moKIwyskhLhTAiL3Ca5VhFGWOsl+uaGIIFNQAu1mf9u0m
xuOkETSvk+gcbT4vOv/1YrkTrT87leDNpm3qDrn3JIQm1RlAn2YBgXRsHJxu4IL5TUPxnC6tmtn9
tK+NGm0bsAAISA/dJweRmPNG5HyRnA5OgCW4hpMKlXI0I3+PdrznvcBbjHebywCk57mSt/lxFLAL
iv6fBUIKTaGZTwKW6B9jLcE6mPrKXhxdqG3FvROQVxhd0xA61C+Kq6aGdS2/j30zaFwCHZTftrhm
XWitu9HXYrAyh5YgModLJHGah0W5mejBoBlgBcaxl5XMM/cbxPq8g67dOfgwJHct/yN5KvYTj5lE
4knFf8rw7E7RDXbzkyKH6dsrAUnOv9MjsswOleiTUpUZLdaWoV+IJVGLAvA19CBASRh7/QmmuRAK
EB3UYlWTcQymZoK1olL+NX/u8JqrhSXfjnPTlZ9KdG2CyDHk2i9/u5F3MPXwr5oqmBonoliZ2cYY
GafO8zUcylTLMT7B+rZR3OEg7yE4lGYIsVBjZPCyyL7S3gBZx8pjKxJr4wCHttuQpZ7NRyYVR/3m
HMTC82As7ExT0KCg4ns0JkVfpnIwXlDh58mWeWiYJiSs0UaM3d+7KivByGH3xCZc5ZiFIfJQ070u
FXY2KeeZ2xdqOZVRekuM95IUtdd6OBHFacomy3tEg1yJxyGk4J5DSR0W25LwRfsReedrQMyjvMow
6/wswk9sU4Y//yem8aMW8rhpcOTmsdLRgDzOwBnpqEGJuOWALnvj+twmDmFvkg6PBDI/yWPhCVI2
4OedLxyCcdc6ttBiwyiZcxuRzJ3c8p3LUeiRoqX8yMDSdcSxP09QN4zDUtpSC7VdPoyqqoKNeszR
BRX/BVlKaE6r2gz3xHLfdajEym+jQ9WPah9FH5BSUlAWGzhtzfmxcsjNDkIONiUbgOy5Sh2OCo8P
hfOQa6efzbReIOo8+AfvnWoJjgI/FjjfvhDBzQq2X5ztUkZDFt1SEMDix5INNz0Ekuz7fD+sn0kA
FrXkaDyXlgj5zoB3nujemro/RsgvkatFpvGP8rXQzpp73USDDLHlbdCrJa0fI+quqIn+wvSjnNex
1/6I4nRLHGWoT/axIVs3T/hSqLQgtRAcyn6AoeH2SPUD56vdqH3XNMGsy5eFL2kA8b4U328+T35c
qtm2XaqWsbVnXJD38f15EFm1UqpQSRV7IBz5IVLOekFVCssOc7rZgNiUtkXECV6e7eo0az3RwLht
nbGOcBEbk2knbJIgR20+T5wh363UYM8Ake9f7jKvNstKXvLFgj7DepCPCen5/tTN+l6z41OtbIyw
aWfaiz+r0hzPoeO8z8kbAHnx5/tvGRvtCJByzWEYxla9p63BDGSuqNbwXXm/LEz+piJzM54Z5cmW
ZGoMK/SOoVfQZ1OCmsoJMSty5Oy4jKZpyWOHFJjYxCOJ7HUS7VWHfqPWI/2dSnX0I1l85sEcndbJ
0EIqFWRZEFQ1GvA4A+IksdyzpQc8hBV4aogXo21aKr984L4ray/CpVEJ/6i3fX3B//iRHcxK3HrY
MhBs+pwvUXb7AwnKZeGIGMHnj9029R38a3I4N62CLoiHqdsBKI3cex17Xz0dDfsm5b5QdL6eRiUB
a3TXV8fju9Qt25DdjKS1Bs56Ds+Dpft6pFPhSBW1Cj7KubSX+Q9TzthhJBZo/DOWbbtE6sB4hB4r
oB6+hrxbC+iiyXVeA8F9Dq1DauU7zuR/YAThqViNMJ5VcV5iqK42doQ8rLEwL6T7A/yJMW41mLs3
8HLJAWvv1IjzqnCvvTFIt9MIzsMimR5F/Q6qg3mRGn3wO7VTvfy/f8av8BK2D7KVkub4kGMeqtwk
BQpF4xSW/AhOZFb9pp1NoeNqzG5GPH7RDkqPUVkA6NArB6VpK3IGELtSuIIpELY/8H1BuL2lYAbz
RdiHh3LPya14kKPlEiSsZbeSdnVwCDZ3rr5R9T49hVp8nhopZlmHRkr4LTo8md88vyOIiGtYdAbx
tWV07tCwFcERn7SqJ0g/UKmor7rbFv9NsQ6ofGzQvf0FrsXL7A98bUlrwfxK+/zjeAB93mnp4RNU
RnvygyaaIM2IOjldaLV1hGiLIeOwcsevSzRTmkWKnHp6LeR6h+F3zaeA2mHiYd5nfkH7veluoEG6
GYKsyLJtTDHzFWGzjpJkaX/oKw8SoZAYnZf36TJKfXEp0UFnzzK9tNUWI+hVMOVuZGmuDyr20EHz
YiD5VDLigVZqHIxDI6Qgaj7lzogdT4elv8MxP7me3YZbEXvF+Pcl/tEg6BuFoPnSTUKXP/4lbhTV
Rp0ylWeaKJi+pWTa70oMJnqKLpSTWhKZWQCGoCbbqE3xVwWobcTqreoE6Gc67d3mhwaE9Q6oznQP
qfi1x0pTKtzogMkMf/Igq9rEox1kNafbFhq/YG67ls1yT/selz2YA8uUGIaKFL/uUqIUDd1t++7q
VgvJzcanI+wxifyRPe1QT3P5h3uyx9hPa6mLVUeRPqZk2RPV8g/jWMc8f7iO4+rJSqB7x6Bxe7NQ
NntFCvY6dmRNpgo7JuzuJz4UTmPDAuzG702rM+WpqNo7nfNKLgsuIHXY+TUcvsy1uP0kTEOzWdnQ
dniqVnHEA2ObnfMzjxqetn+9UjFyREr4VSJvk7XyequVFJSXBf2Mbs7eO2ybLpJF5vX0zONtMv0l
mzAvnE6McMTho9IS+iLkH7TnKsmv6pBIOW2RHi++9RXI6nXThRKiADCt9wtX9a0lrBLLLqB0Uv2B
ZdwW1LjMCabpon1U9DV06mOpN8Sl7GYfpv7nThlHaaj+De0vlNAET8EFL2iwH7XsvcTjsiMOTxBd
EH8KHIswjp+yAp7SjVnJq+/uII5mcnGvpyAAqLy5TUtWq5CwxCn/MaBzWBwesl0VCjx9LKromchQ
QTGbf225cftDkPxWMVzGMcR5w2RcycyIwEhG4zyPuSklQMcAJ8ZbdU+VwTqCgJuS4K5EJ0NPKfiB
NI3NXXyJG/+cyUeW2WxgbVJqYy+bSgvd21bdgc0l8hKgAuDfAB9UlXL6D5hkhoDyPFCD90O5p10l
8Uxw4EbFU039+hdPH0RPNoTWTuqSbElTcmReFg4n7OToZ+OOM60VAfCri5QDd4z13bAGrxFbdp+P
/nVbvCtQGJWu0MK20H6zIx2aryoyKrNJWFDB94zRbwbnyLOgHH3/patWUUcrU+JFyKkYWIYQsdJB
29EoND3bPjqt9Pe56nIiATUqR087LMOGojo8Y3Kj8XP/U+n2MuBwEmgR5c5VeTGOOPrqZc4Kjd+a
XWO3tF5T+zrPX3+0Fr/5O/uKKmucYiQDFO1aCc1X4zL5dFlYGSuC1WyovBDqWeJYVYC128P3wFEm
sBT8wFFV5Z55b6C9s2zkVp/Rja63qa/DHUPhOk5QypyzAis/AHkD1ZbNGWxbwlgMHrSq07lNjWrr
yJz/eNZ7HwMFjmS9a/pALp9d8Ob1jyEIV8tmoUei+fcjV+6NnTiepTW+UupduqVliDE69bk07teW
9ohKqU3iuaf0Ni8QLUl7TldHSR8VtNKQgr+Qa+eK3vub9glEKQRvc9FZyynoDbBZSc7imHwXuUI/
KX/DdPIrbMLWPjtXeC30Bb+pLofJGQ8UtK03rc6KzYuoK7EStWavxe7y1MRjCWQ6Dj6jOSYzMDv5
4bF7RKhfeJKPAXV6GjS59imU6m7moleHpLsrfu0/9oT0iPLUfEm4tme4zcllWVfzTI+hrL0IdC7z
36Rm3IW9D4a+CmCeI4kIfi3Ediu8nZD7hw1uh9GSm3qmw9mARw4qZgFbqBhK5qwMgsVBBDwILhy3
PTneIgdM/27jXI3dzdj9DKshAsownVj2Ivk6j7hKeny1p995WMoyoU4w+Jcpl7tWcdEi5Ha3ERgY
LWrv86wN9kJuSV0deOekHhduo1JLUh8vVVHadA7TP642yhaAhlEDLZenelWYs7ILPYlOKVSyWeXv
bOzScp1X7QzMYspQYBvIFpjxxLoBACHTTZbeuCGuxol8UXcVQgrlGHD6W/pt+paHuPqj9sc+VCjn
ocDveKHPWr4X5k4OZsQOZmJ5KL4QZZYKcF4BiDjkMhjpV+CuocZxPLDSmQYV3TDaL5+Vm7coRMwi
E9hI6POW9Dp3sgjT8Z8B6ht7L+VkmtLdGwZ6fxvrF2q3e4qj4cbb6IZN6sobzlbGsnDfsk8DYbJ9
9SWzq1ifzjeV7+0Y8fNq5ipF2mdQVl8ZWAkz9WkZKjK7v0NSbekyk5XCGnk/t48mLxhTScGXRZK1
zigqevxjNHEi7A31orzpbl0zHthuxAIf6duM0u1aLfBEIdiV+WOW2TzjBTllnfMUoegRM96mL/wU
U6Sk+G91BZm7pbXOBE2noW3x/PL06Jo1Tc9JvwCDHaci7pMeSnRBsD1Zn5QiR+/Qu1S9XnhTolgq
3u/w45RtwT18q6NndvmLRkzMppMJS0sD6QBTKUcLBEebbDcpu1cIgGRqOU8l9SBGEKuDpMllBa2k
dDuBfaAmGzWFTbRw0/EEaZAKsa0cAwdUHo2tn8ZQSeyFdmwOK6Ed+f0/KspBLKK+6DcvHgm8A1sd
hyWW6eByiOgmgs/Ey0cZgIUO5y4tr4hKuC0XsQk5YXGI+CLibOx6sM1Du953ICtU3H1bkYC0vcsF
x9Qu8ObJjEUYI2EodctnyS9Lj36zx34ea/2+pPRfcL+fRVvoyCDfj0SR82PStMnfARjClYz2laZI
bcjso5BTEkjjS3zXyOacTMmrFmH1yYKl596USCmDz2iXo6SFzZAR+1gvHEDaG3Tq6heIL72m0e1r
EW8AjXx84jHclntE+uoB9daxyO5NRht5U3+6u/OmqMGnvrI0WAUIvTQkB9TyIqUuVg2XgxBuj9Sf
MrBWxLBHbNQNieyuxmFeOY2U3rNJjIy0E99Vm9OrzeUeIUpmtEPfopPYU7Em43wYE3+Z5DTyOdT6
yhwx1JN9PBAY7bU+FyH6cVpq3ecNNHY032Fa1ZhZ+e7Pt+Tc9ZyRGn3QAMQWpjqa699ldxpfvpy2
NF1rWggk5NJasioIZHBqFDiYr92MAJiIiDy/iiVdZ6TYf6NFLsQHHPVwSz0Br+GYgbMINZoaagTr
3v3paXn1/Kq8SkxX3CAG3eXNp9lEQZByNWmMpBmTz1xxoqzTxmz6xlRJSzxYKQBpWyWGH8A337DJ
cUmWXUzURpT8ONyUoossveSHEFX7uulsXf6BMzZY9FsgCpuJBWED6srMa+DADwqyubZmqNjYMDm8
fZ1jlXvzOQP45QdOpkarHPqKuQH+0L6v4fkx6QaP4KKONWpL5lBZQbOv9XzREIiHz4y0EsP1Bb6I
vy14a8usUIIOu9cv9T1WvFrYntq3Oz8YxQsI2ZidKTHdGWr05laMfWvGlai5VkQBdvn7SySdtY3w
4Yj+Tj8tqPyI3eav4MdsxuTLsAXYo4a93DMGzKPRUfJaLLsWmpEW1539W9K0By4IN7nXxKCLYpVX
KPJSR87NzexNoTCbzP2eGviJ3DYL+cryzQFviKondquK1oovv9yc+GbCPntsFnG+AEA8ZjXMdZWz
+iUuyb1g68b8exrETF5k0FihBdI9mjoL2l30Ncoxpsb+0IADUggyPH1PYSaJ4phNpEsIKJObTtUY
ZYX2JdN61vgtWsBG7vlwfJZrHePsbgbFIsWSRMQrWvp9NDNZ9C0KMOMFc66TsI0D9zNZdwbvSGyf
L6kBxjTLsdEthGBFIBoVi2VTojwRKCVSa1Rws2ukMemgr9RxN6q9T77Tteoex9DbUWr3SiY6WNF6
Aj8NOht895vrBzXMOL0fxl9RT/V+UvvRBv1V5x574Ylpw8Zt9SjwuMjYnKd3iTTOqcytQQg7YRI7
DrHFVbejx0EfRUL18s+kMywbTOEy2cKVzIgCaL1+NkTadycp6ob+9lfFAxPwJ2IB3Pj9bpXtsUde
Umd6bxCzso2ESaAk3ukJXVFtHEGuxQQF8COVFvfaiMcQJeK/P+r44I89LBb6wKeznoCYBoAc26xG
RNVMQLp+eVzLqEtGfmNZmPHF/Icwu4fc6I36gbe0bG05XbP6bzsmfT3VrNWvbzhffdG73S/MSwFM
lOHpm8yoriAtecubuKuZYbDhEoBE3dvSOH3uHg7+tBNZVSlcdr52BRYWVaory3VDekFNFvDc+i5d
VRRDphKQyf0Scfbv+La4QJXOYOTfz9G3PjsTdtpKswP4NrKykWJjrtAg7SPqikzOmVFYPVvXTWXD
PHab+pSZsgz7wlvHyi0JUqDUPgdQjSIpV+tymc0MWezpjTXI1v4Nk1N/5oYs8zpBlWWSNtOHk30b
3cpRBUrUOaWvSKEyIHoW0BEjMYmF4oXWEppdzi6YHLYEdD1TkLgSFORqIV6xfLs3WJL10SdSEuYS
ox4W1PE0tvpoKnBJxTryoKg5AHwEWVRGVZ90e5+5qacj8+UkHv0kJ4VCnjYw0BWrJN7knbf+Umj0
FShs/2RkmVX7lols7Flllk88mVA/Xhl3bRB6tKa5YXVSMM+hBzTXuvcnzs/+gxxYRLakO4SgD8TZ
57W2TB0q19mVfZEP4glIb7EnYu18YV25chdwVTU6R/vp2wVapbo9jDo5nr+RiCnWQBvKZ5a9UNUR
XqyWz6DHzi9cSrUlGOnOuaEHmb98yAYEbs4Mv9oR3kXRO4dN/dD4RrNzpKIpi+Qq8ec66bnYTUBS
AD2YL89Umjg40wmOCDhCZdyPlZygQC8e7kBPb4/PW67CisYH5pjaORlHQBQciYrX8lWQf+2/dDPw
EgU9dOZM6BH07iYwXedfPIj32sM+NPZDYhRObtON3yZg0ULp45HJFQ8Yi4oyp7Ttix35WVgBIayV
yl/IU2IQpR7Q+s+pa+sWqTOBVgy1u9TuIW9iXQQt1Oy9wULAMXZhvfZbPpeH5kjAYR9qixLOxs5/
CxZ+qoRn5TZjqRu3+qISXb/SZMoRb0sJ86+3aj9oUmHXZqP1xld1JrCFheVu75Fx6WBVgTIj/DwG
F59FBw/XYCJ+8ca8+ky6umKhNw0qlB3bXqUw8LJwIrZDexkcNERsHEYIZUDIDxMN6ao/HnLkGO49
pZfgdFoq2lLeNKRi+IlU9yZHPamaP4+3AHpBS4sWXROirpZKaclE5I/xKCwlv5IBgahbpvTLShYH
WUFf/aHDVzZr3PibJem7b2Qn7rtT87gmeH6Lyhy0PAV5ztP+X+tCPxezQQSEdfmMRia2KUYyCwoa
Ua2y3Vac7aMVU5q7kSRilaIe0uORPHLIlPF1d3HiSTK0FkhqYP0S3IeZ99uanlBrEWvHx+r4WjSx
6zxhlq1St8zwvLMBld7SUzCb5J1sYJq7TtM6nLPMRCYfbKFw+ActaeQBqL1htYmrqeHKpKB83mGx
/mIQhVUVDA133F6Ih1zTsG5RCpZuO9Qk9tWLDShRuXh3rm953W0eTY4LsiRQuvzw90mN+RosNudx
Y1/4jNXezIyvr4JPGexR/P4XY17u9VwsrHCMpD7h/clCeXlZgBpk5fBE7wikuNicoel7E6BVstzg
JcV7A4EpbrnloELEnPCzndL6Uq13rvHiVSY8gfpIHporqtgPCb/s16aRtADuequo+tdHJeQqTYHD
Y/c/s9aRFRykSPeysOFffrd2qtvOZK87YHjisZT8+QxC/lUT57vpdL7+FdB6IyVBVxo5jhOr2Uu0
PP6qkjQAQ2ttZEj4O/pN0jw4aOPohiRFhJ05cruIPp5d6qulInzH+NbUDmlVWWhp0qgNNJGpSva5
4Ybz7EjMJ+x/E1X4gPLqa28+G6ZZilqoveY00BekHsBduGq/xljPVvtOxcsz29w1+3OWcsG0pW3e
rVqr5WpQinqDEqPeX3i+dQA0mkGCbyVPuOxG8z+zVSYOQnqxAKjIZacglM1qfMEFnF4oDr/hzx4p
x+FqtAEAPWb54XA+/VhYYB1kJD6HBAtCdWmFv+0ca4F3B8XvIm03r95ENkaoCsDdxutXPYJpLyZw
6wxZdb82HMAFQtb3eZHJvzAcDooCskd8V5xjieF9vJJD2JrFPwxtkcb1NJ+i9WanIemCwOcqAWnP
7DOrvKVULsqHRvmjbBwWiKwS5m1Esbr5qjI52osTfDSbSdQwYSVo1ZesxN/hAXwxGjOxNku5fYK9
ZwKskOjphJJlb5Rxg9/yoLELFjnN+LjCvinOqsTZP7KEjNghd/S8UqkhvxbvWiZYZz81/lDsM2K+
Dchtl0fSw9rz//Adbc9r6QgAL0QhFO3KmFa0kYzcqB1sQ6wr9UkzGriZxDfNYn49XCFC4+xpapkd
wHSqhP0wfdvNYUV9tIwFps2hH5H5hcgNbFGzIws82IMjkoTXIBG8ZIYDlB2MkyKGT+OKjBm/xFKV
I4S+SBNxGZcWh/Ne6lIEDOCwmpVyyERqjfutP0mPSsoyEvwxNCCZNbvUzMQBBKs6dSGn5g9GyPXG
/1zd0alzVTVscQeSidvt5L4T7sjEhx9bujGNrgKHHDCdiis6tLrd/UIFy5p3IARv2hUUyOYOLvH7
jR0GrUzIz5ub8GNPELo26IWg8RW1XUuWPhZ7P/t59BwV3eBt0LNEHsq8mTIZ98uYG8+PQ2lW0NqC
HTeFDUWFpbqvmNFqNvFivcJJ96x+VM9jT3N0ZJ/oawbC/XYwOglyX1wW3BB8qV6gqUiSTiWT50A+
rUtC9Bc6jsBjAP/x/MoVsQI15e/Z6utdBZJwfP+nC0Mb30onkZHQNGlMoOVVgwMLJ1lWhav/erx1
60BEHkjDTtCDLTiNRD2NIOtEuqqVMk5PIxtrG/yMqGVsdeS5HF1gX2f2Bf1QAoOqyQ4fwChSJBO9
hBp5uINbqmMmQOQQF1mnVN9U8sSStGhXNSUq8JPONndK655sGf2jXMdOMaZAlSHKNDf4bQFsfeIH
nJaHSGjt9xgM5tEK/MNYdSRHge71oEXAOV8kX3nV0qeFu5Ax4/XfMwGbvFtHXQJyzRWQKYt4xwS9
oSAvO6FNj+4lWOku2wj6z7ZolbRiR8UCnQ6xepIODFcMsjP88BFZoBXSRo1DjY1WYjI5Eg/iBTFH
zTCjk1nWlnpLr74nKtVF6iss04b2HbwOX6m0OOlS1PRzDs7AHcrzy3P4m2e/XiOwm24rMVefoD1J
DXKKrsDLsIoh5k+vqFoM3jW4Xj5ufbCFnT/653nY8/QP6ElQL1oOir0J37y+wmmxov1dx0Ht5Stw
NJqxEUx809MDoj7yzx0SWBtZ7CIMIijN3mrkWjq6ZBTE6ERHXe0YrcK6yD9Wnt9t9DeCOj6ExsYP
RDdRzMJyUBCQeTRFSmPN6P92+qhHpFoZxlhjbkE2AxdGv2p462b6VYyrrZ7vRtoP/PYI1730f2er
rmMd+5nnCulDjDQFQk7MB9kvMjjfMbAqy14o2C5E0BXRR+QFF9ofU8+bzzdc5Ox3wm9erMUcY7ap
EmE29btmiU+b6G/Vf2SOkHM3X2cUuzS37d1VP7xa5VoXQcUaTsT8Vr7DJZ7vffqm3DYoC/HZlceH
m/bGzZXI1kPs+eegopSsE+P5mbTyt364/Xdh4ku/u1CLCyNH8tbgal26JJihqPZHNfrBG/WQQTwO
JNiBaH9+dawqf79UqUqQeESjg3aieEFhSt9DKh7WaW+Vb7uoCfBI3oVHcB9YacRzXxtsuo0vpov1
qiicnkKMbu1mbI2l4f38YAuxrHq+bU7ZKh772ETmPu7t3zSpdnVgT88ZRYg5nDLruqtoKmrWau3x
yzYxDvVKaT/nrkcH+PZmmz+wEDLc6x8EkaTXb9DEsnVIr0rjHBn7jt4OiIAlJjyVydKrgbwhRyUo
pGEGkIWFWYDUf1S/dHynh/OLf+Vi9mc4I7BHRsZBor+BbeRwpboY2Xz2SyI2ezO8uqIcBTwR8uxc
SxCurErMZ99QaunbWL36RabVnlLIoO94AMXYiXqY/JMi03iTOw8OlMdMahygBQTRlKhGt+wS+3WI
DrzBRhKm8UCZH3UI3A/WmmYL+7khlfadDiuQHL+PBEaAiUm4/4r1+7zkX394EjekP4wo2VtE39ge
ePtw1LUMD773vovE510cYIKZU10mZD/sW9wxOKMBqotg9dx34Y0njZI5FsE1VyAZyzitVfhZsJqF
HlrXVbkNiBgLlLQo61ye5S5WMmYNmDFjTpr/+cnaE3xcgXpRZKmU1A/axoFc36WZzfjSFiGxHg0j
xKHEZlVBIwmQPbk4iJ/uU3aEr/sbta8DAFkQ2Nn+PwGeMKTmrQqeQyt4OzE8hCCRLLQOp3J3nl0t
iAIhZE6kZPjIf6YN8Xn+l//f2fv5byyJ+m0MB0ZXSHILjPhX/Q74nD4wBvs4Ks+WjT2JWXpo4jLv
9Z2pjM8HyyEJfxK0MSDijbQeDqznv/3j/Jm5pCQc2FpNAUjPw4QXulFWIfLyRwhS/pYpzeHRb75X
grUkmZqFhUnmA89hZCnABGW0e3R2n00RH7EDygTQvIDdf+rGBV2Dc2khQ1jJCrIc7vjMmJ2HZSh3
Du3nDWhTwYEyf4Jyy8J+EbDEr8ZHfPpsty7hbdMhVZ84ep9843pWAO8Q8WkwCtn6Uwqmc2N9Srwu
5C4Qfq/HhtUFPUZS7DA3IG/SXyFmjQPPy9pCyZSExUmfskYxrpGJqRrZESQ4UTmHKtNzoNEgrDFl
YDy1Hv1TCxOj6KcB0Q/CejthjWc85+FS2YDCW1bumt83m8XyIpNROJpr+GtPLSX3jxAw/bIqyNuc
dFObD+xJgp7rTs0bPGDGe8VJVsomLPitD76F7krC5zR+xqWqmu7NFazMmkvRqvoBujheW5F7wmJ7
x4Ueo1YwJ4b15vqt3lNIgCikwWPn/LtKdcToZTWUZVMqNZm++s5RIMVPmsCrlkKxtHp0LJtQKHKV
RguquBiN2xRyVJfxYkwuSiBAqD1c2BayKN5o5nSgl6xd5bvwau3FVyZb68HR45VYe/H+lHdF1izT
jCgJQ6D38Alz3NxqqbcvYYY/V/4pIkIIqQdN4mLIgmyxNS2v8ShcbE2OCX9G5RcfBudHLIRjZ28K
7xIq3li4N5fpcND/G4in+K4GlfTfHztMz5siBhxpDFcwvdeg3K0sphAG7xLLLglfA5YJRPjD1q2j
1Sm/RPUgaskmtDxdcTzwDp+Qs+gs7ddK7dCEroeNs6mlpp9oOKH+10zWEnMwis2hewLvUPx11y6I
7GjjCnPKmCjLH/hUPNWC2p7fCzI6E9lPIwv/QbHkKc8371K5bvRQvA8pu2UfAmaUSXjkZ4R8zEJk
oXCEItsGoFhcRIKukwnyqQ+p56ik3WrZfVwtYlrceFpjtj4VSB7TdnU5wId1HRp32NN3ddluabHh
qRfHow82AK8PFcOtduuhfgdHadMJXiOCaVjhTuiXlRV5/RtCC6HoVBLzA/sG0v+EkwcbkPDX7NWR
RuJQ8HjIB9LAtS7iMrK+UnPRy5HEaS67q9+9i19qER1ZOVulF2zVH8+9NFPwVptGY6cLSC/izZSs
/2H8OQvhZFZQx5llb/Cjj734QoyfMJ3H/8cIot/D1InTCBNA+UC4AtMa1Bh0g8CeZJgCbw1GyZXm
L0wPnUmlOGKWKZrx+tu95Tf2kBsrxnr9yMu/ZlxJV/PX1F7Z6bF0901w0A8IceItVBXcqB822+vD
NbABXFSbmUjGeNtIqNYBnNfZRMwjTMrQYd5XmkA9uQXV4ZEnPba5eF5ot7GZbLqFYZSD+paeGJuS
p/1aEOLgHqJ/aE33WpmNWQqXEKZWuAhdn8CDeJSawU7itqAeQwwgcOR/Bf7ra0EddGZybwLCGK79
Va6GaSrj8VUPfNXFi5GWijFzdAlsygvbBpORNsTs6Am1Qn8nMh1RJdI98rv/VImxWpGxRJz2K48I
NrnnTpBe8lIDSTpAU6oj3VVKG3WbtfEHqLxT8mJzVlr6oXIM4TL6Jiw9nLy4FM8EVk3ZEAnq0aEC
0grFOGS5N4Gdy6XT7VQCSFJwJUy5MuEDPzzfdOqlUJNJzFo7iInYnn0AjhMQarZQ76DIrpA7N+0Q
Qc5L+MN0VkzptIiYni9VvAp+97i0Ct4uDQ4vPPttstRXxRwsP2rEmtSYp/hWp7bsDhNqFKSYqPHA
+JgywuVIS0Kn1mjGUC2c7rNc+0q/DremcvAhZnLPaa3EDOkjVS3z2buqtyEWgio5/QNvC7K2XZla
Dbm64TKj9lQYmXjdDb+UUtPiYiyoM2m6f3GCOkVuUdVT0UZIOTjwX8q5OPkVuAicm+CUVFoz8F53
yecSeVx8zPaLjvFeYkxv2+poXC7yOFvkM9/zpgT2/IyaPSYKNuq6aWJTYxjVgQTD8Fjn+PuCS3IF
19czhWcThNvErVM2y8lM4Aor6Jjxz7GFnAZHfARiGYHj5vMjx7prOAdnvlDRWfPJVfaOvxFkls8A
F9fTIslrA0e2xaaEb1I+h4VaZ1rDsxqWepYg1BqW3IFyd4aBBaeQIiSAt2fMbG4FIxxqmMKzw/Qq
Wp0i9PTK32kJie7XSpxtMySpN38Oy1qc9G7JXtQ8Jyzy8ArrSP//AnalJzXMKEgWju87YgB5S5gW
oFkAwgTDBhFpRdcbKBzvMdjppLPMq/Gsd6K1fZREGNhORuogpJd1NlpNRQUHJ7fEatX5Q+whqugq
bD6TG2xVzbEpXzjuEnWUC11ECaGtFXvjqBxKA4YTQK5pRoU7rBhIYvEOA0u6MZvyUzwcMYf1npxG
4UGO5bVrEURsDzEYhSuXSJnVIhrlU6Juwqf9zuB88z1PA3Ywzr3fAUBXBkXCxNJcr+UJcU02GUd5
ZUAJBSS8Me1FL2TEVklIcdpybyLqfQ+s1fWGt+N/rFfADRUdk+J8gJBP5JJHFffvf51F9UM4X+BF
i/5Kv95gOnv0jVKWctEQvsvXZ3Pau4gCI9X3KulJCV0eNO4TCoNZOaHEoqMCN1uskiSgiRX3x8md
jttEMFnwefvJNnBEg0fAm7SsgVMEfjKVnAZM/1MZLTSGdAol0WomKzJB5imsFXkKKso8PVS14q10
8DKE9wSYnua7tzryshCRcIgXZ0yviROT5O8AtFS48S9cIOVot2/CGJyRFdHZphH4r6N0myMoHWdS
Cirxn1CJ16Q3D38bIiyWtgsBqHF8F01sYbNpg/Rqrx/TP6TjepxC3cjgIPbrPQ/uSh6L7Ha4wIiI
5v0vhJyhwVvbSbQoOKnM8P5xbep4wWjb3xZLzDoNawjtmXra62sxJWLp1+Q9GI9P/aye4C6wwAQ7
mc8l4yGkns2Kl/TWnaBvDc4Lyn200yUM2G21eDGS8OYRsu1f/TaacZvwltsRyJ0lqMJLRoFalHtX
/Ku5ph6p16MNXXu7isKber9Y5RN59biRXqYwVv3kdQzH3ArtvSIQYLzB8Il5k+FIiw1FNzlZJ/TL
59YGb1ZZCjeyAbnvuWUIxQ9/UudQiuyS7sNIwULQAcQV1qCxaQi0b+Xh3c8l7At+W5IheA0+bOSL
s0FkZf0FiRUug22mhZ1v5849vJoM3Uciwjk7wpaQiuXYGeUKE+Mu/F68OOvDV9ATkT26HNwdtHMw
/zeL5nhWeS2/SZtB488fgwpDN4IPmVMib8HWK4wuNVIlYW0hBqXgejbFxLlFr7puKXmQFUBik1I1
RDHoxvK1LvKWbcjkdhb0ifkygYH5nyClmY+j/ym5o/+CrnAOOWPR9zcVfb9dhjwCmR8YU2vgzdbo
XXL8gxVScBZJrbqZVvNfgrT4eFtO+8SpiJ+bCBselsKyvuowhjOsMTgNdut1XA5jdxnKglENxuUb
40lCOlL8B2SQVaL18VS9dWhDs9ZCMavte/sepb8QtheWbgHiXDJ1awbMSltOjWGssvfbrg4W869M
c1tU/NobfBLdsT4/1a2kKpQ7Wobc3Gc8MJiGEkIK8Tl1/qKYyfZF19v1wNldXMjB4LFb43NG81Id
ZufmSi41kjhJWpTcT+75vBbp8b+1xcYBPe8NyzoxUBWrZFh68uytSkvncIUw1N1/SJb96Kdo7Uvv
q2gHOTL/vD1+5Z3s4Z1+DTQmqHOCBhcq+fZ1D0BtDZbklxgT1UEBUADB4wTYIyL5LLIW4sw5EecO
Ed2TIoeowBt/bhwjZ204iTtU0Nd5X1KJOKaK0UvibDy70Cb/X0lD6MOhAc4qJZF9MANGk9H0O5yc
ZzgkP8qb9gq1hkwNdVV2MGvxDfwQPm/ZG1Sth8X2hD9M1zdwaTWl93/+JsoVXQuvZQlMD/x2EWBD
XNG7ZJscw5Pti62hV/b318fIUUxn7Jth15mMVtRKo1MoxBQnFlfXNFImAGv+cpntwkExmfEEJKf7
cra/eSIvenjCEUIwydT/S3oYbuxSzFgotGR+1gvFEujbYXFDo5l9a0O13+IhziVY5IwXo4wPiGnR
iF2GjHPY8r7hMGiS65XfCCxQDqH/u7xeT76z9uOy3GCEHa5rthxOth99a8KiVA+LWn6322L0Whn+
PDTb9dI75rX9TTfRjivI+rmrDJncZaGkfcVTpd8f6RMVasBfhenj/Re5wvb21k/ZCwyC+GoB9EOE
WjNW0qhJ3E2QZTa12lZ9hBWCMfkeyslP2Cbw2Q0gpuc0j+hebsI0aXudpgOnKSeO0pFfRslkZwqB
U550nFRBaodPyq310Bp1rfudiUSBGpYEtU2c6mU7eKrnffd2rQLXo6O1ZAGHtp6pPCDPvf2Q6bLl
wEhLIz1uPvHddE0Km5y4qbKfzO1iutCxoiMuuty6a1or2CbU1wNXZ+cmzli8SCZFufKZSTuU1tJp
sHlXoANuKYO2uNuGbwQNW4heglnH7kGs4hU0Bi+fDotW3ein1dYelZKWEroOzxMhFjOywLb8maQs
KD+3DsjwTXwoWp66ouUq0rEkXeeFoki5TI5BELtI5Ni9qR5ge9eozzWfMuiNgWReltqmvoim7OHb
TjdnXybi2F7ypLl3kTyn46MGIB3LuJ9PF/qAGG1Wmb4GOnTwaUv1BnOn6Tofn126/KeVuxNy/N/s
TcLKkGSCifTvX6a9zwmEcjzP+eXp4mQPWrESmNYml2cosZei9LsE7R+F/dmeQR6SbyE6zNu0zx/3
Ijk5QE0q2cPXEP2nxud9Tj70cryp+TJ2jL9EXlFxBdEe8wgHzdDQfczmAUJ86ob0A0XG+j9pN4I7
UTp48ASrLCCt9dFgahvTISNjaGxt0lL0jGQV0bSjnA8=
`protect end_protected
