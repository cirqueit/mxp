`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
KGYiY9wWdmTl7p26QNpaFfPTWCr+3ZsoJTeB0CBFulR+uUHjyxWl7SUGn/Cps8bUMCCeLXpn4wFj
IruXSRdFpmyDI9xioO3duf82Kpp5BAk7JM9gH2IBJ9spAQnHyxUu2lMJ1dszFA1AY0aaK67mONYf
ave+Eme7CerGnmuypI3biN1iAr+SWFyXeuIQqjbIkckRhthqiBfZZV0N1cxXyWJojUNjv/3LyJM6
f/gdPo6mLL6Ki0bCEGr4g6Fm3/ERhUmdYcB8jY3kWU5lbf/nJ/0xoc7GoZ//BNNYp8EjhvkpYcuf
zKhiPi/atw/ihJWgqQ5wRgWUHCMJSeNo2SHOwTbpJjv4Rt150Yiexl/m+MPVRWYfsJAqzW+bcI0U
epRrdfbU5rXFJNeJxTQNoQnKUKG/fjXL/pPMJ7xmiODBcQQ/tckQG+oFAJ6PA+1NyUr+sis0HX+R
QsxILbLuc5EyvKmSy7hidrMLQtDGIu2BZCOPiu4LdukPpVG1vOS9rSvmIcAnTiN1VU3MHenGE/eu
8oh33HA6zcpqGpraBclsn5tDpLyT+wf6pY/8lNu7CNF23oK95wWphecc0QP+nZ4ihyiwMaBsojD+
4dynGCu5neMLcrk0vSsEWiFkV1KavjO3XiUN1TueL1JEjkt/wfSUC5b6nJg5ps5PPKGJHK67ptTn
Ed0LFfCBoSGOV4b1iM7iE/eXuUmQhPWA04UURWOXRnHNq2YcXY3j0f+NBPhivqOLB4L5BENbiKjB
BLF85MwwZC1gNRi9kKALsJX4x4DKTKHxfUq7wePdnKeJQJgkZKF6xIjQMRgzme1D5Wj61+zARaIg
23eqa+SYmSGdj60x7nawkTEnzK/QgV4L1SSyljyWhst/CIju+t4JykcuZvgmwtkJieCvD12A0s6v
fYG1DEuWuf4OVIcwQ4XppNZLyo8LMTxxpmzgRrmN2g6jvqqo650HY8expuZTmK81mmHSTPkVxovf
/bPD2f493orlO0WoMKewGfs+2vIWgunmcyITSEYDPLmWVZnSUXqjRWRZJiFR9g7x4IWLYioCt4NS
xv2EgUOt4XGU606ltAKS5o+mfSCO9e/r3sU9FBjQXucIHXB5vLzBmtwCYb8kbRqEsalidfnnkSEv
ye6hfSJSzdhCIpqynmS6DlSm8/hCsE6vRZEIJAq4KFtjw9LzruzOScd4eCu4VM5G1aUmBlJBen07
1MKfttJKLsMtCOL/p40Xn1mmdBf7N69l4IazWgC+caqK016cr8xHdh/5C0899ing3f7nVRGPTfyM
WlOfT7HhjUbjhai2vMKf46sNeUv3RzXsoIn0Hcd3/NRWGwCYuXtEEYK2uq6avwap5Yy0UeD5jrg4
mlQM2VQUJI4qSygfC/R6O6+XXAMkqCtGbJJiQ/OWCERJw3hKrbKjSkKe7I18xkDBSHsK3HfrqVJ3
mjm97P3cUEB+l2Tktf0+PyLJu85GDRKmcXrQj3JLVHVvOw3Q77ufqkDrBukfJ1Rqicki9BWk70lr
0rCGjHNvnUckqyHhRBIUBbyk+VZtEvzXV8kYAmX/CU1eDTxvrFakFphOYOcZprFNFz+9uqqB9SuE
SN+UEf0jPSQhD865I/+C3wyhL4yKvfLIyMw1fPD0q83TWdS90EISVDhvdRNcuNBENYzPU8MdpI+E
AZsUCindOnlfBJjecN/31nLwdaCs58uoyzxCWnTkKpUDFEaB2CqO5wRq0sWBHtgTmdihHKP4FfGx
UbBP6yRVsHbUKJrC18CCwP/ivFTO51Lthk7Uvn9zjDyQdVmVpIglvOWNufSUrmdKQOIMDBDq198T
fbH+SMRynuI3hZtaSdK9jHSWi2YNcCNajR/YDTmW/78cUo0dxvBdPDCyABZyesT7E3j+XyPyw2ks
ujMF24VpdS2HqY9xO1ERciLj6beqHw8tCx+jh0EyM3tiUCCBdQ/43d5Abf54cgl0LxAIbUHDbgRb
arwd/ixlVLBRJmQu87/eIVI7zqnNO3Yrqa5vfip4CkRBYgbB0tOJUWbo6PIdvzewaDPYEKNTweEA
5QT1L8qCBeaiW7J38QL9zdltyQ9eZsH4fGrKO4v3Bk4cKySVq8KizjCxSURylpKD9awpp4Jl+CYX
n2bNNGZChQOdQSCx78jXPMdg0XoE/S+g1z+0BG/sj5HBFEfsgUVyPmd1IhJibpTqBvPibOX+97O0
Q3KSefh41dYBSMw36p0p5aSo68uWBmgD7QGYsK4aKrjIv4Qn0JgduwqXhbaqpG+k5FjxsEITT0SQ
zV3f43RPeuXjGng8GsuDeljxQlky7dBY50p90MEddFcYp8XfuGuUFiSlvC+GYU8wpIt3pkUfNgVG
OAHi3L3mIw+7B2VT+2WrvAjTH5OIQ+zkD+E0pYNyo0MGMOjBAsB4T2b/MdyL7r4yfijY148vDHsd
UCK6veTUoNtBV4b3PElAOGcrzARRGFghyqvb6yNNkHjIuc5xyu+2R8CPUqkToA48mK1PkAFDSL5H
mq4AjYqay1xeDhuBZf4vJr5b/QTJnA89y0pkHfFSvBFfL9gk6DUm3YK03UhoaAafr7MMf77Vc0T2
junTesVrWjXK4sDxR9LUb+YKtvL1dKGqWiNpRS7n7mxLOkT/tUakhAffnRe18UM/D/kqjK/kShEc
Ca9MZ9nblLNrgKh20ReP9gStL2abL4MlvVwP/LYIatu2qmCvVolFizUQ5u4WCqnFkzeRPwnM7tf8
3Wgotc/g8DL13HLshco7qijf+OJkVJDlxQZgNXDUOPrVyoZPwKlOHcYj0v60Do/e01YU7hr/oDW5
7HfSE45bPr80lm7xIdvrjL0Y76I7BKuJo9tzIwDXRKaNMp5xfTwEhNZz9pW0Kzsmczc15q2dXhrG
g+7nQ+xxuMO+VrUbNoCwgX6gjih2qmW2FV+cSrVxLo83rFm349mmuo06TQ0nyUUtxIBtkvzsiW1C
pRohx0wGAK2G1hmRJ4vjNROget1T6LLelUhiPSnpMlSeHtGODM5oWVm7IELv48nScsdniBobcryS
Tztjf1Bk0KMTab8nld7ApFocHvpR7F3Iazz5Q3262vYT7N9UCEms8rSmKyM9NctwYs/i19MbJec5
THfh8iBxAMaevMyS33ungGMwPDI78UBheBcq/VQhGvsv/sUjdO1P7e/kG5nB99NtZcqKZOxPrQak
/WstW1GSt8cqyXBf4nGPf03hLcGFSlC9UyyYyOp1+fLgQ9dDj+VSXbXIF09Ub0VOCMBz0sqpiH9S
oaeTFWOk9rqRPUB8TMK3M9WtZaoHlXk8bKrsYp7G78i63KP7OkX+8JLZO/OSPjMrNjIQlZ8p6yhp
izmvbHPjxYbwA+lqAfpL0nhpgPFOCI650YzRRvnrPEz4b+PniBIDY+l62hgEax5uZ5V14/cHxNaZ
sFAatsnKnfkTSRNsh2dmyyS6GQ3ReB8r/PTYFq2kCQPj8LufvZbQWs8PGhUPpYvr0agEb/rBzCn4
hRmc8xl45HutrSpvSXI++eVaBpUwUESBN/G99Nq8k5gtO4h+LhyINXNNhpOm1UD+yevM+qVwZ0Ok
RMTIpNivKd9zZ/AvtRIouhmimmWjUVyowlj0sXg6H2UYYDe/um3Qk50FGKXpLwkPTS46CPUkBW6U
djJjeG0NqIjQvlmDfVwwOQjpzBhKLylG1umqpbrt1RhcZ7iR/EnlYy/4FoK/5wZmjv5216trXzKg
t8Az7I5OOctwDrxoTgCOorFI7ZtZDUiEy3/isfem0DtF0wfikWVEH3oz9ZuHgTs371R+lEGPJsaF
mTJtddTL7b0sQEMg7pv4Jb0Qaf4dAHY3JYtV1e4Cxx7DoQ7g2qyiuAvxFpz9i8yLGl39nUMreAXF
32Kw+6eikVk31cYX7agtlCISShTA56r8yAgH+k1QLLJKVfuNI+4oqsXI6l+pme7mYiOJytsP2lq4
pK1lZ0wOJXIUQoLjauZ89lVE6yk337bK+DAZRRlO4V6PqYSlzJoEMeH0zYe/mtpRnU0cm9uIpX88
6M2aVOdp2afDK54O1xv+FgTA0JK1P5rdQjim3DgOV/BDiFKuFVUEPAXUBuUK/dSf2xmI1BATjTZv
Rprx/RY+Hxl9nPYNzCKJCs3+n/9Z0Zy+9P8sYPk3yP1y0RWLmPy3XzU/o4twJ2RFjZlREetYf0OF
NctFb0qdylnFQSK+F03ONIAjzbTo2neX0b+REHIA+EQettfhVW+C/vS033x1dBzUAY3z3ByITGb3
gFw6cZs1PPIo6P/2JWsudyRwyq0HWQcA+3l3lHxzyIXaL9oKENt26R9fA1c7Aw4Ih1YnYPPcpEaC
sz+iiIe/YTNVt+GVzszCpQnFBOjW8P19omdiNRh6tqWVaMTCnWL+ZRvsBdcoP/oRv3LtRqxEUIPj
p1Kf9DLNE3J4QBHQNQe6k4jUoacvas+6io7T9AVpMumIQk0dzyoyPkvz0D/Ft167Wnezjw/pwVwZ
LgT9UzzZzCvsSvzgyGo4U+ZqsCbLQFc7J9xZVLTmqByk4fqibnREQN+DAqP1YVxR8oIr5iYaCnBn
fk6g2B7DR1/6NUxwVgUREobH50T/CY/CQYHVRWbLLtFV8b5+nM5fDixpYgajIseU6FUJgGnrNCRQ
xybEaAAiQalEUZ33tDupuTbqpMdmLAJGJg2u
`protect end_protected
