XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6MD��6W��m��;�.�-�(ڡ<��q��D����>C^9p�U�<���d�}
�_j�����?�ݜ¯���L@��S�ھ"
���3�<�R��?:ꧬ����\2�����$���xJ�+:����qu\C���Q{�ڍ6��^���*ҳA1���|�'r��/����BT�C�����/^���0 ɷ�pRk���n=g4s�{�[Č��4UvI@h���e��������P�.ǬӕHk�3t��l�9h~g�_����ϙu�]Uq���t��!4a�����|-HElCɞp�5ܙM����Z:o����ucIO'x���:>�F�l:i.[T�TG�Ŧ�kޟ]��l7J$y���u��L6<��Ї�ǣ[O��1mM���=���((D����$!��k���ʵ⫝̸[�^��G�7zO��¢�L�.Ź�]���L���G=T��R��Wx2M��}���Z�1\w�b���S�Z��W�p�?CĢ��B�γ����Ap�e (���)"�2K�ʍB2�EY�6�6�q���鮐/C����M���>�p��^)/����:�>M^��?��Y�g�a���f-��2B|�]���nܮ)e��ˢJ �x���Z)CX:eF����@�1�c+���g�T'J�=����"�_�:44ˀQ>:���O��к�_	b�BRMM1��Ds�1x`��wF���Q=���v�C͇X�'�f6{����w
��ϑ�w�KXlxVHYEB     400     190���Ӄ h���2�ԗ���mC�X��-pj�RF?U��=� �r�70b�>DG.XȆ��>�Mn
G�����-��2�<�ϐ��6<v��RvF;�*஋��9�;�.Ö��K���P����$�1`��U�W,0F�:04�9�Y��5�t#��D�0��x�T(�J���c�����ؖg��8��)����\Þ�݃�Bu%���D������R�����.�1h�7�'�7������%�R��5���Y
�J ����䂯Zh� �z����"mm�iE2���H(*�5�v�)�
�;�>�r���"�L�]�(��́�OC���.��T��f_>�#�ʀ��QY2�����/��/��J-?�*]�;�|��1���6W��M��c2���6 p+���H�XlxVHYEB     400     1f03������\ڴ�{x��}o�I���zc����ŬZ�~m��-�����+��<��62W�X&������M���6�P����!Ph�^L>>�� ;�g8�D�/#��b�8 Z����S&z����t�G�5�6C�7�����|Tuh$"�(Gj�pV�%7��gX��!�.���������1�S�X���C�9uqA�y՛��ͦm�E��nm��`��/$]%q����>��IlO�j@L<Yō��r�y��[�k�s[���:�m���1UX*���^ i�}"`ifv��J��5D�]�\>h�_�-���A0N��W�.N�/��I)�M�{f�<S���+ԋ柠aX�^�N;��K��4��W���x2���p�&�������?;���_��T�P4�,�(�E��1��d}�����|/)��S5Jx��,��Kй�n8��ȴ�̄��F��@��W�H��.�g3$��̕<��2�W�t͇���XlxVHYEB     400     200?I��g����σ�%�]��?�M�U����˝NG�z�Z�����ɑ"��E�a,��%�fB��Q����ݡM�O�I���l��6�84�x�	[��(>���� ƣ9��bA�(A�P�Y*zI���l|?8���b9�:���]�7��>Dx�Ҟ�qUU(��>�@�F'��2^����GI�Ƭ���=U-�֍Lf�(�~�$�n�h���Q�g���ۏb�{W��*���!ѐ�������2rďY�)��$岵"O:�ݢ;��J hW@�מ����t��#�vs���H�b)�l�17T7��2�f��L�Qj^eumК>����;���*�G�l	AJ>kq���u�����ˊvΩ��*���b�D�`��q�0�a�P\5?3p��� mD*�$i`vO^�4�m���}�.����$����V��جs3G��z-r�ܱ��V� <,-G�Mܵw�6�E: u�a����I���L|ǀ�~�I�����۾Nm����XlxVHYEB     197      f0
ۨ���x,����>Q��-f�tJK�=�E�+!E{��E�<,��J
}=�&;����Ma��J��l�H�N��I���K��ܴ��aB��D��`��]R�H�7��hH{@�wg� ������M�0%��ؓ�kBP���SX��L�_�.{��ί:[(j�|^G�eO�/�j'���AC;�1d�|J�c�dBD!��VOiP^�Ƃn���Se��QD��%2�M�;���