XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��N�p[���/��遳�Ui��:�G~v�`m���XUC��s���Q�K!c�N��`�M��/	�3� C/X���h������Xm|��g�XW��6pݑs?�	�݄k�V�}��������O���,{D�^�#�n�!~���zg ��<�������7�}�<U����c��V�,4��{��>m��$p(�qm��lO]�Oe��7pX�ߢ����?���e�>s���E�����@soq��6a��/O�)�to�x3���&*�2��bh�6�<�W<, +=̏�uZ��lFH_���6#�8tMyZk:X�.�@�� ���]�ę�A6�9�D��V�q��ئ�O��%K�-.����;��)���SO��f��e�Q}+k�p�ԛ`���TU $+I�쓬��?l_����0t�?:�R��Z�v��,�Z�K��9[[לے��V
�'�H4=��p1!R�S�7�t
��q`�ͫ���ZZ�C��7��=��l.q4��*�����v���2	�j��J�>�M��3)�e����{�ѢQ��.� )���ˋT^*��G��C�!��?���1SG3!��x1�i�XqC⫆�%�^��-׮䫐���ޛf�~kU~�o��aʦ̯^�~�ⓔf��z�ֽ�I�S�=>ŝ��ԛ�r#2y(�qAĥ���uK�Ĳ:����0�Ũ>�޷��<���"����vbҝ\�S�J�p23u^�4�1p�EcX�� ~�죮3��3?��m��XlxVHYEB     400     1d0y���ϵ�E؄Ŀ��t�y^u�Cڙ��~,u�^"� 2v#�]P���e+ڜ�]��m�1°��N9ޡ)`<����6��H�#uǅ�ig�It�>L){��%���a�si�B�<T#+e����l�9�v��A.o���Tl�v�o@_s�Ԅ���d�M� �ho险d��i�3��yA��H�m>j�9�~�Qjo���~l�΀�?�{���� �H�y�0�	9X�8_֪�����S�m�>���i��WZr�|��~���&C���� ?׮�-֦O�D����s;�Hʭ�i�ai�b��0�|a�o�[����;`�q(O1��9)���ry�h�������<�@D��yI�[�̤�U_�dxϵOx�����*)Ԑ�F3�u�?�\������a���4��a�TԢ"-�����8ڗ���j�!��#�Vy��b+RQ���rTw4�L�XlxVHYEB     400     170d�U��Ԫ�D��l��讔�yGj`X��
r<�!��S���Y��4�Y�R�D�@J�U�/u@�<�I�?'-��"󂬒IB!L�sUd3��
w�yq$�]�����QB��歹�c��f�ӡ�@bf�*�����B��8cK�KIH2�i����r-ǲcC���'�=�Z*fxGƅ�D9����D��y��F�ˬ,�l�~6�Ё�/��T2��i�����V�*1�o,_�/ۃ���������WX>�wD��A���󋹆��l��A���?��E�n��!��m0���ܲY*�W���F���Y@M\Euo��6����>��}�:D���h�N����������mc�~�������uVs�ۥ�XlxVHYEB     400     120FD��'�f�xn�E��}�f< �%m�F��]�y��y�-��LQ��j3����k��[V����e2�&�U����0��	�}i�\TKݵ^u�j�%�Q�P��@�/�����e��J�����s�Q(��g�^m����d�!Y�=��?#��ksh�F܈���:�T��c
�X#�Ebk*��e%�<�¢M�SoN��ǽ�Ayn�Dx��F��e�j�Ğ�[b7yh�V*g�[�Ø\��K*�eeﲬn^`������4�n9���@�l�ܽ�=�~�l���HB/��3H�XlxVHYEB     400     170X3�ƧO�Q�Vt�'>xz, @c#?M7P�7��}|�\�:����>¶��F4����b�5{�Ѱ1�*�~���M&0�W(�m^��5Ӽ�5:5�#����8�G=�W{�w`��BBh੹����G6v܇����!}�əh��d�Q��a�D4>驹��� ��/J]�,ry<6�a�𴲩0?=o�v��<��?Vǝ�a@Y���8N^N�g����W�7(���l�9�B;�����N2%�29g)��l��հ�I��1�2��u���W:���|X��Ko�^����^fR�@��[�?�ɽ����m�B�Y�L9��]�i2=CKq���e�-{��;-���2N�|�X��]�ܦXlxVHYEB     400     170�\^��˪��?��bU�#���O)*z��P�{X�9͊�O����8<wl��(=�6�%REl�N�ſ
�pv)�a>q�����#�n��F��)�J�I)�0Qev �J���H�}������vfu~5o\���(F��{2��0� E��y�[?�4;ٙ�]0>$���~���x󾖱�_^��/���]�d�1�~QI��H��p�z�� f���r
%�r�|����u�.2��NW���qKGe�y�r0�Si�����J@l�8SN{./�ͱ��"�2�NG�A)F��@kC#b��o�P�X$dQ��:�ݖ�G��5;�v���g|(�5+�D�18#�=�t{{�bhS�_�ىXlxVHYEB     400     140Aч��Ћ�E4ҐJm B��ꦑ��O��"��|��k�=��j�#��T����ف�f:�1�y���P��%�J���Qx>���Qn�.teG/F݆����:�^�AO*nE{�m�t˰�s�ǌ
�0)4A����y̦��I��Y�Fe8�5f�+�k��Cv��D'h�oV2Q_�,�����"�-���Wލ�W�F����'��y���HF�0�ɬ�N�����Yх��VZ�7��GF�1Q��=9U���;,�9U��N�7iA1�\Oqͺ��Q�u�z(`_Q�ʍ�x���={+�fgyXlxVHYEB     400     100�m;W�PC��Ė ��Q����)���N�#R�\�S}Q��u� F�^FPS����B��IpXVځ����K#]Cx�P@�KV>:\���{1c�j�%��tԳ���=���95N_�3�K#��r&ƧY��S�_V��&����.wi�'� �R���M2��.f���>tP\&h$-��OuTz���/���`�aX�J���KL��W��x��*j������]�h�i+�G��� ��q�����%bH�1f����XlxVHYEB     400     170��*���k3~�S�������^K����~�T5B�h�؍�"�eLT��+�Dy��wLtz�ݛ�?�j�&a��Ux�=�m��P�圗p�|�4�p��FAv*�ڧE9$�j f��"��&���9�y;*-��?���)2;{�=9#7M�Q���B��. �������5OQx�9��#�"e�U&����
�]�����'��Է��<�ؼ8��q�Q�e3��P��"�IT�Y�6U����m����)���_ɶ<zu��>t2WX���.�a�����Z�I)a��(x/��4"F>�X�,�{m����� �Ov+3@��ٯV)��g�jο��sD��`��Y\�Vl�XlxVHYEB     400     1b0�pd����-N�Ųk��"� >\���J��^WQ��*��k|�m4���:���Xs���k�p�=�4V�u��2�ĺӥ�AƢ[�xK�ˮE��m��rS}�����ݤ<C v���
�eG�{g6$	'm�j�hy�cQ=��x�O�A w�̷y`s�P���I�W{�O��ӥ����1�\�g���6q����~;�a0Kw���Լ��ڝL.�؁�/E���ʨ��0���v���!25c�4Cy`�r�����1� b��ː��y�,����wNu�ܾ�J�`��^�5e�%Xy�G��k'"���'�>M�z�P��?T�l��1(A�P�P��'1��m�JȲ��{�1���<'-aq�uժ����4��y3���.B
�x��1U��l�:}V�Tly�65��K1f���g���o2�Z8i~'XlxVHYEB     400     160c�{����DڲEd��?�|2#Ke2��� ��+�J��2!����׾�(v����ݚ?�2���iE98)�����c�[;����?{<V1��%=��	%_*M�����&��*q��F�rـ�n2���s���
/$8h	'���f� ��G�:��̥	*[�֡�A�>]^!&Wx���X��NI.X}-l/2�%K|g����y;��w���n͊y��������A��~��AK�*��e��EV�I�¾���Q���������C�Lz*�*r�hyT�K�f�a�ADSE��W��'䢃����K#���Qv������t"�k���IXlxVHYEB     400     1d0ρ���'
�<C/.�y��E��Q;�� r�l1�<z&�ZKJמ�%ր�]��M&=�� � �&����0�L�ذ!S͒��zPL��z>𹂶!F��[JFѪ�@�ir�M�2"!P�a:yd�:ߏ�T-�W�F�Daʢ���͍����&����P�4���^�Z�l��$���8��������bu��1�:7�x�u�U$ϻ�r:!�$;�i�Z?�{=k'���v�F��P�rA��{̈́\ru9e����"����K(bʝk����1�<,ȿ���0Lgd�ym�R_B�,��9��z�T�.;�a܁/����W_�V����t�=Ƙe��W�:�]��b�EZ�6��P�%��V���[�%��O5�p��ە��b�Vכ$��_�n�E�7	����� &;ǖ2T��u#�W��q�	-z�2�Z�֝9��x�����iD|v}��#XlxVHYEB     400     170��9h��ݑ�w�f_�2��W�U���a�DC4D8�7ہC?1�R	�UH�h<�ݺ�>!�����w����i����䪀�������o
��)a	%�����-�H[a�Tǽ3B%��S��=E��x�n~�
g�
�oȣp��/�u��=[#^1�r>[<�/���ՕD����y�J����N��K���	��)3��� ܍�aR�~�cM�^�x4K�����Z��P�ݘ��@b�q�]��nj�"�т�C������� ڋK�'��̴���G-��-�gyK��L��̤>Le����?�./.A�(M��|�{/�F��0x9�+N�W׵�V፵2�
ƛ�kS%XlxVHYEB     400     160�]Q!��Ŗ�ӿG�}|�I�,�V��c�Ib�[{�� r>�Wl-Yҿ�#ǉ���	��8Y�)���7�8
�~J{u5�S5�4�6�<-�n7Z��?�c$�)�\F�Y�V��;P˥=��âT0=_=H��YŊ��^�<�;g���	i��뱽3>��׃{Uٙo��=�!�`i�{�VU2"�z����49�=ĹV�{������{A \'ذ
Ȅ��� �dVr���L���������j.�Dk�n�]B{8SYl	Q#�-�L�ԋ�*���m�"�����X�s�=[�jU�K5����1�u1�f0�Z�=�w����b�戀O�w��|ۏ���~��!��5�/HXlxVHYEB     400     180���]��;��ͧ�8��u�b�S�_��GU�)P`��Q�o�3R���]��n����)�"�,[�(�C�c��U*t���3�����Kz��u��e)h\������ǋ��'�vY��F�ޯM��z2C�w�3�c�E@�ؕM�&���f�@�x3t�@�*��y�G��&����&ãdGGnV�s�e���"����<��YN�:�l7<?�'�_C�'!�����A|Nf���o1L�K�����4� ��ɉ���l�Z!�:�)����@%��t���V��Y��<`i�|6�|��Vo����Xnf���ɥɩX�;_f����o�/���PՆ�yv���|����Z;����P��1r��
�XlxVHYEB     400     130���e�UຨOL�J��qw���y��߁�j�r�ۣX��|���tq�$�U!��V)��[Xw@[��$�g~�	���(�v7$�;���lX�e���\�,+G�F������4щ��1x>4_K��2K����E���Cz)���OU�||�X�v-��TO��1��5��-.+�X{��O5$"%�+�[�t�!�)�\�x��p����P�ύ#ھ!	,���g����@���]�tq����Tf�/kٱ��`�.��*��bMy{%e|C�?O����xm�9�XlxVHYEB     400     160�Z��a��` `ǒ�0㜹��Ym-��,���ΦYMb�o�(��5���HU���G=��`�!�2Cw��#X�F�[�ݕV�=�y[)Y">ߖ�*u�=�b;-�s��+����Swz�������$�ʁ��of=Y���ޛ�=��;�S۠�zyb�Y����W$��(I�߻)90�Dp!5�1��� �9�=���B�j)�=݊gP�0v
�v�V�O죓f��Z��(��YM���eQ��ó�k'\��?�1# �81��C��plΐ1�u�*����>���l�-Jp_����"da��zk#/�d��OA���&l􈿀�*�)��A䨻P����ItH
�XlxVHYEB     287     130��b��*�w�Ǥޥbob�#=��JB/E�`�|�?��W�0k�j� x���a?|�0�CM�{��\{ ��a�D��`��*di�E�Y�����m�ڞ��[�s'Y�߂q`�&I��FU�j�f���1��X#�n��Ʉ^�^'Jd;G��CQ�d
��7����`\'���n��,�����t3A:;h�l�0+��˻���Ҷң`������h=V)Z�H��2�����4X�kYb��pdx�����"��A)|�`��<�f���Nq�ħ�
3vp��[��`��I�+R� ���`������ppϐ