`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17472)
`protect data_block
7DnNI8JJYqmOkL+yUkQRoeznDJdGUZhGe+T8/VUkfpbcY17oC+GdwzmrO55m+3bUx2+F4LcNeSjI
Ho0sNlaiWJCoo0X5oqYvQ2zFshxetRTmPMJoMYxldzP55ZKWCj1zaiEJK0YVsDPU3XEaiocQ7gCo
QvFzMdtdDNiTVQ2yzoirph8klpWi1HoJRZCEVg9QID9dAlXBYf/cqUKxAVtJBhq2fDJD4ugOWV5h
uV1Hzp+jB8IIWvqJb6pF8+LRWVnneCTorFt5FomTHfoagAc5rxPf1eLpGPBa4O6WpdnD4eMMpC1C
ugdYoLxCalXbyvclvsGQRowtiDYGZs5ockoVz7BXfL+7W+/MRq1zUa2aBTGCqRP10ay06tFsTGQS
1u2DTTSyOv9JgDm/A13H84M42ozZcq6vE3nz/fhUj1TJm81gfNpkWc2lzq8rRe5MZ2V+1kIlKm7T
9XykMx6KmRduwTLr///+jwJNsuorkPkwKtXEhIHLFSbJm89MStnX2rVwGA9zY1iB4JJ+di48d7e7
3xVR6raHvYqY6D0Ds28TFCnQhKjMzdeVfs9W9BiicI5tMYTu30ZlPhJtA9PlJf3h11XOw4C6pRWC
Pn+yHgAAfcsA+HTsoa9fwad75ipTZPaCuvwruBoCMKXu8Jz9fEeBmAc58DKaS8YzFGjIXSR/rpnT
n4FP55ukPEKVMLvCLBuJ8hVQY82tmpz+DRFtJmvnZ8G2Nxq25xsxMgQtsTDwcbg1Y6f8Vq+mHBlr
3QdeDct1BgX2otOkbFewJzBWycrBDxJUm8Tq/ayzkxlt2nbDpJrHk42wBYULsLUHW6aRmYGBuH0O
HUQeqpsWuHnrDifGYbRNajdMmxfdDle0rfpDoyf/EORCr5mPQ2IaZHDf4OIgBzHe/5ygpvuPW+XC
vPN91SCtg1JVh8yoeqBY+QHeEatbLfhWB27wxuzFpiTVLICTw1/tSSoTdxBLLvq/Bncy8GvbC4kx
YQKNT5sGfKpH7MbHNXmBXmbnDzrKDkg+rVXe8/VgVQkSkOUlTK4ghh4ZwYwCBDJ/LKN4+j8Xdfuu
XL64YFDiuwkAwW4WaG12PvVZ5g0GhgFkrzkhLglD3EMgwy9ddL1CIi8vc1puv3BfVx00shXy7HkH
9zfng/sxA9o8yq7wXbh5Zs+0cyP+EQB+XaMjUeNjULfgTPxR6T5FWSegtEa2919T06XhprUNuvZD
LPiFlPnUuS3D7Sx0xYb0Gd7D9AWdT/8bc3JsyqFvUuERq4vW8hcs4cZdlnNOhycBuYZBeffPIYhN
gF5RJZwJmw013esACVriN4uJtGI78hoCVpPYmtATS/bu+9g5Re7Cwizv45+26K86BWbp0F/Vv3q1
fdlB4pCoN5ByjniiTzb+GmBTi9Z/sASmUS1Hat/0W3U+vwansFSdfht25UMorPsUKQ4GotWWqyx3
irESHeQgRWyI+nWam8gwhsuaNUUvp6/J2gABkCfUMMqYmZovyI0/NnrOA9/G+WsH/8mzSHEQxELW
Z/2NLbTpHd+E1sBXKp5RnIoGMh5/M8vT9/8XdoKJygnEZQY6tLcGe7OGbFleOONJOr4MhpvtQJGT
iGwAtfBjgVHq7G5+SAYjE8HUxhaFTsl+lcg/mAnLxXpD4tW2yqUftJJjIOvyDF1ks/72/buOIfn1
vFmFjTwSDMi8oNitgfIwDPbuUk1Irmmdhl2bnh56zD360So5VZXdQs7p4vLor/37SRsEizClONVu
IzfO4DiD6G4VTYeofaHYFUlFxc3vY5fF/ABnMUqJA7BP+I/fjJ5YDRbSoSircSK48u82x0Mn7Y5D
TiYx9czbMrTT/5DV7n0hjIHr3ume6umemBe9L4OY5EJ3qQBg1w9Phfu3QXdeWKETI03sYbvmcjEN
PcS3KCCX3oTNxeZom8w213BDXgHWuV6LElmxOZyJ2x/sGS/wY6CHPS9jq9noKzg1bikAq4qZm2kf
9rnD2KU0kG8vPw3uZMVul8QDMG272J525CVriSu5RMiep86P7dZI/JGmOdpFboYusyWie2J0sxVi
LGZwCCYgXJVpM+BYSSwHvbOuSYSq0e90qcDAka/A7UlseAeJiywCeKLyYSXuCASz9/9a9/oicWco
4ajvWkPpG4w8hf0Q6/hddFkiWmhKQVyva5tHfQGJxYY2trX+LBkx4yhBooUtzhCCjgOJqa8yMoZW
UhZJkSiRde4+UBDpt5/SJxq/eSUPBCxTsRIlBrfsFPbUD4w3B5XEVuw980e3YaWkAdnGNGtR2klp
C4pv35oODgQEssfofeexnG7bTxacWYT0wlNS58xRlrnoz+JLtyvxUHCZyVpoVW428YmDxII3bG7U
CoiBpqIUHw1DO4pkZ8YT3eUSzoi/W4KqVR1vI/WqJV6WBpKkFOutdre4KwLBmkj9/OtuwEYAxgbU
y+KfNEA3K/e9Ug0Co6/VL9cokXwNjVOxnYn0C53P8PJoLgf9k7B8mzCg/z9khuvswYU4MlfjR6pI
TBDxy7/oiwYp2j9sbKav7ctlte+ex6t1RBemAXYa2hcjcoB77pNnBBglS4xXBvoIdzfgI4CX6y5Q
P/dt04X/DDxjNoHAI1Aoflx1EJDh+BEl5J6YWm+eL6gafk3omHiGWZB6CLCX0SQ3TUDrZ4+LeUzZ
CAFtaFkFsU6Ao5Ga71pqg3nJVmyUeGTJlseRwT+mprSod0E2rw1L8qAwi5ggrikbIIjJwPLVVt2h
8JcuQMfrm7td56SBlIopNcctk/h4HfUQ0N0C062ewRhJpspY3lqwNIIBrkjukwBEA6+F17XJ6w1G
Ziu2M03JJGr2sE+Sy0B46XPUjvQ6sA5n8btdgNTtz7CVk0QvrQA8RtafzzMlyURzfSpgnI5k/E1E
bbG82cibuZThAcQmBkp3WM0+Hj9XkhOvQQLCoIysFGUp4AjlyCJoqGVTfq5MhZjAVYUuti0iyVMB
OzDR+51gE5BQUzQKyco3lQrMfDITNBn59DdxZN46ks2wHU2UN2OA0qUjZWbAfYkwLMkwRJIqrG2y
qXWnbJPvNpB8hTlt8N4xo6XTy2k2a4SZjs4LcuXLge2rrvI5RIPvaMyuc/NDIeV9bsDAlELjC/pX
EsKQ4VyMU2yk7S71SBMrJ914uBlsr8qvXy1+m477HbUYs1bDMWZUWGNtmJF9CwVUISFfYuplEALS
u2EXiAKhGWUbDPUl/ajx+8gJ3ctX06mJcH7PRS9f6sxu9PhU1ojlGvy93SX4fVMGEJ+GHO04B/Qh
b05rkfoX6J370owkW5BWpRqpZH13RBx7/XNA4LSF56k1PXsjr0+FtxNyzXaJpwcy0hSyBt5/9VZl
PBkez9dA+90Pce4yiDWyWqAJmIkgDNAzkPmvPhbKkASoFT/uLLBiyKUYdC1ccC9J/tItQefSur3g
xfFr4UP2nogONn3V/tMr1r8hbp+TdHDyv5Qq9pnFWcqUeFQF0hLG5o6WiAda6vorWPT0AsebP8FK
fdpc0uoj7+YDTbR9v6oVneEFZj6yqhbW/hvh9BFG/P+W5N1gyHHVOYODoHmD+ZDcBQ/qaSpyYwzc
vLRCQRxm9BQRgGmoakbJaSNfDc9u2+IzAroEq9iHxJiyWgjE3siBiEnztJM963tm+AjNPorONZGN
FAJEV5JzQ9xkKqr/a8JrQ7ci8GfwWmOOnEW1pi24AeCIutVv+QomYiL1fwmRdqJdWEy6C5KgSNbi
i6//N6A+rpr1hqE1lRlBq7wXfic/0OKllo4OS6g5vdCwGdPHH1eC+j7syI3dNmR/MRzQlzC/8B6X
7bf9esiHPiszxSJcKdaPnXN6zk8WJ410eCtJyrWQcVyABg51u2GwncLmVTnzIBP0ADts30yY2tFF
jIBieNf8y4deZqiKrI4g7loiMZqrVe8aTQy3MY9tm7LImZ391MUrQUaZ/4Qa7tiGtImmXHFrjWYQ
vYLo0L12Fqf16MdzvhH9Oyoz8Bb2SeBmAOIkvSgKP63ugv21h2lXTiban3PnlTSol/q7CuVcUOgF
PKIy24n0hhEltRbwABLaOhAZca8yrmk3G38rJOVaRV08vQVUycSxfwOWgChBj5GBfVEsp/RBy6F8
quwj+OTLBwaXbKhJ/g4CXhKSa+TP7l0NvXe5LmU4cPv/mK9UU0ev/5j49sjtrWZjO4D+Kroa4Ze6
c7z+s28Ow3T4XCVgEkuKpO+sI+bJ/JrFsiZGS+SL9Gy11zb9pwrZGq+W07O9joVJQ/tt7ExbsVDL
XqDOXh6Tk7mKDQLO39AGQoYaY3URJAbKYrp+Aq6k3rRfCUpyvLE4DJTgEYCUKiJP/LTXvcXRaFco
tmBALKF1QuuSiV1p7HXqFKLDpZopOzK3uV+bkjYdaBCDFbQojoaP29uFB647R71ia6EJh4saq3uv
0MmCU5EocLLeVUAvnM1tDuaoMf4wIwoJ1Au19ovcV939kI0WeZhtS5EOQgh1jkotgE/ZGVLa3IRu
WIBwzGuiRiUO/Nh6eDKY5NnC9zf8tR9GI6jWfdUA2McznRjHBnTjKHRR3gIR1eSfavoR0N/0+L+m
na8LRnn7FQF3p/eHxLhBRbm8SijYPtT9Um2JmonCOAaSdB6lpQCKLfiMSG8n/seZiK1DoA716FIF
smaZpIGFjfmFq7IDgA51fgVld5DpM6MqsM1wwWeglOzBJjLpT15gPesh2fGRhHU4GkxoLZo1OJCs
JzDVAfZ0B160/5uyrYHv2vXx2MdsqSesK57XCuyeJh46aQnpYBHK1IYXgU4W+02hZQFRvvFhGAau
DHb7nr0LlFGzA9ddhT1zc9akTL2Czlb/deQlEVe28Yj7OP4VGKkg7Ooto3tGxDNRAiW6S4o48Xu/
L2S9wnZ33lgJoPYAQkP39dqb3JX686Hns1RMp1VDFHsB78OcG9iqfraGhTlu9BEPV9bkwG9OwFbl
a+HXSNJRWqzA9v9GIe1oWA2YyMGPiNPHC9gAPcgrWehBDf/DJbvW602bkTk0YDqHgefVXKrWDh7F
bNtnwdnXCzbE9fR0x7RJ/NY+08Q+dhHsLaeemfwQXCh2Mnkfv/MjQqM4a2HaLzrsHn+Q4lZ70h5e
nya6QTlbLPgidOJuHrX8CO/3/eqSaMUZadkbXOXpmyO6LDFLaFArdpaz0YpdXfHscidT6fxWRcOa
XDxeIeAHHP5wqfiwybYgqag7JLswRjNF/uU1VNwt4vIh2XRRZxnVssOHJRKnoRM9idigLZjhxUcf
k1HHAaMq2kFG3+b6iBTb6o4xn+3qjtDTYV/bFyXeUEQ11MzMESeed9BC6FZNmojkTGkyiLh5LS/C
mYRjuzu29bLs3FfGCUdfs4S88nTz84xKy5GGCZJ2+gIXWLSpRoLZu43oDHdVCReAA5QT+C7E8KPh
Ug0Hc3bk7hrSgwVnMocB7I8iBm/rtxHipUJFVxKsHPxncP25+0UnVa3FcHiGblfK5qe33P+PP7GZ
F0kA/0XHt1TaL+NimM9y8k689oXk29Tt/YcN5HxD78fKP8nlgRddBcnza6SxShqZHfGIsUvLxDwc
i0oeF6/3zrnXe6DnY763WIfHtlu5xWrFLV2ztR+l+ofZHaB1bnLMbI41xz+p51d0QKzR5mTH4ScU
xpggK53oOxD+i+/UM5STUSxxBE3M+aFc7MJ1KjzdUbxAMFt6Q9hVnHvjsNjzBmdqcNe/YEMlNuQO
JUjRH1a+eXer9sjeyCDDD5T6s2/xZD9jrD0W7wHUD6HSjdO74fSD9AtzkU29Zvhp+Wkho6z/WNkY
xHeu1Q4NlyDnG2bXmKz2BrAzTlAbRrIoKGohbvLP2KrgjmpeiTsyefbHPC0X52qF+Cv9mDClXnH4
RvYgt/vBWU7jX6zglmQb/mQP0JA2t5t0AqPjVIbnYrVoj7evXRzpmiGIXGD3IVxc07Dr1wE0Kc/t
pINhjFDmYVgnhpuZlPKw1WLMNID9zgvH8tjXXdGTvNGlnUhZYyl1OOiDi2z2cuo84AF6uH5A/LdR
xmpU0Lq4v+sSle+HH+7EH9Fey3nO70hl8jeO4TdKagVGVJ0Mfe28oO8/llGl5gFlVbz98c3eYMw3
9uGf8PE0xaMexbunDLLtQmkoMCPPlp01bQUWvu9cO5NZTzyJk6dWBb4/eElX11Psa2kUydvXSWzJ
6zWLbvkl411kuiP/kH3P7hAjuHKpb9Ehw19gr6y1xCU0F719cBLzSFmyMPlepQZlupOzBBg3KJxz
cJbfIoGM4vg49psX3OsqR+Htpf3sATW71UGHewv+pW/cbDrtCiLNr2/2fgg8sob5ajYjHR9ITN6/
2/AUWR+TTA3bG/uOwDeo+9AML5y4fdh5h+LESYCXCw5UkZW4L606B1ClW8yCSc2DHZbkRxfzs55W
TVP14IrMwo03ugaeuNU6S2vY6o20sjmNiVv8fYjL0uwXglQujfv+8LzmLf2aQms+zx2+m3QDUGCt
QluKlNpdoc/X0HCLHfUY3I/kbN/HTglvVNhcIvmPgpc/Wd5HYd/JIVU9mJhqo8aTsyhkFAp08x9g
wzlFk8wtO4XlLm0iO39AO9K01V4ep3Vd47gj/UrgmoOU5AYxC6+EX4EX+636pBY8tiCps8VqWe/m
RcWkkm7hptgtvxHJqGCzoDHaZf8KYrpsp4f0XtkVuhT5yyERMsPAk+UDaSXUlCrJEUM/lEXCTdF/
0Rr2YNIZGYKCoyVpP28kEhqHHT9ONyFAi7jr+LEbgV69bHvOOo7Hxz5086R04Ro3FIQuesKEqscz
YifVkG9a15x34kcVqnzDKxkUs+Ow3bRyhlYM9km2RNsPevwMlsX9H/8CyPw3/dnysjRAQNxH11HO
6OBht/w0z9pXwZ6jGz5bsKIo1eOBlVI+8q9zKM+d6hmUdSO6Md8zqkShLlDQth2pI2OJctQ0pKp2
5MFsCg6P5fAA3WJcnROb23J11UR7dMYVMq4w2+IGauUYBEfdV3Z0YjA6fOpNXvFb8Rr/5kvRjU3n
4Hg5K8Oltc/39+9ocEgrTMs2hMy8nHkuafNYbbwctJaLRQnHR+l5cVg4m6Xv0acyGdS1+YbTNZwb
7QzWuHTzPx19bf7kIpQTxVzvoSdXABHDJQA96wr2n1hEMYC8SAgfOxlM3LHfFv35RnShsy/0x/Be
u6y0OMFr8XoO5rJmoqvTDEZykkfo+IEBF8shKjyI6kJAeIAJzFNYbQi+/Oe7x2/hzHQwDb8kyFA2
s7ElP1O+eKKckDfiHXUCld0Gmfgv3IbzvLH1ddhQ9093HmCZOJZXrf5oF5HFV4KgAHf+0InmFPSv
Flm2kZQ2+FeW9J/KFd5e4ffKE4LBc50Rwn15c2WzbylJh27uVe+HyFooK0hag34XvLxK/+X67kiz
NoEn5CGgolL3oFaOXljmFf8JGMNKEkzbZl4VZjpF1R7g7PvIaSxBdtrk2RG9p0efmhyIDhpCNPPY
ICHL0D/8j9bnn0agfQih7ytJe6jEFBswKQyC1yKID3ZOHUHsFoqWw1vWurfG6DyEp7KxyUeeI3Zu
awxT4k04PbLKho783yXpQlE8Zh7vkg0h/SlsJ08tuT+XOkNnqyAw2ALVOj3Boa18ineES7xN8COe
ufD7s9+TP8weMyWYyz8cRtS9rn5U6aaf/uUywIBf4gBBOpF4bcPp2oMp5361HWFvOoiw8vtFtVQk
MAsgR+ipzBr93CM/INhnd3vAnYDFaQIIquCCgNrTvxjb0jPat5mBdQ02b/OQqVNJRL+hpVCz3p3l
0NQ8IH9jtd64+2MzZMLOmCdR2ZkmL8gSFuf4yKnzYkSiU9WrS6uCHmY/mb2S5sYNk3xV9mn/s5bQ
TNpCluVxvv1cYBHaqGfU7ny6n2gcBas6LIjn5fSQqeF1kDilk1j4H8isZgTFQVUV2zCtlD+kspk9
7vGY6Kkto4ChFauDtHZ2x7FngF8+QGb11zT6gsHm6RQnOF8iSfS8U15XGdrdYNaTn1Ius9P46tIQ
4MeIUljfTf+OG95xBPlc+e7LkSseKAYq/Gj2YGq9+UiAZgMdT+dGkXxQuEmjBMQNw1H78vAgovmc
zPaWovVKurOG1s5ovZNi7pAUycFPxCeqV22LMt+xtqGauTPG63S7U5ffADso1v1Q81/YXpZ8FTR+
MytmzEIz5hrCUl+wooLvelV5xqnngCvNkKY9dTit3rnJTV+Jni0oPcC06IqwLNAjBCJLYe2EIC33
uulb1S68WXzO5dzjFM4uMeSp+eFQ83oSNBWEmhTGqJzXMQoHMVGmns9h8GJn6Tevf+NXAkdLT7Je
O7pw/tVO9xjy9COGbtWab+8dSfA16l9DVk4617zv5R7yDJyiBVB4ug7Ky2lzkQs/6OY+SnZ5UZn2
/Dja/OePXxJx8fAzZB2jVanWaJPWWoJ6+kjQhZUJiSRWycOffqLOblLBz/PlNlX4UhP0jO8ZV5oF
uTCa+vjKUZjKybVuSQrGY5it37yb2mUxZaYeXSaj6CF3S/V8i58heEDoC8crfcMOup29Sao9Om5k
8qa4GYVLaIPe4x8uXuCTW7OKsfw6jap8jleDLPtop5s16h0W43b+nL8Id0jrq/hZ/4+hA39KYgnG
2d/16C9HltOpstn9wOZVCbYFq0pzCC+P4RwlYs0t5Rt7qVuF4TQ7Cti7Eqfhg8lzAGyp+JPqvd8K
DEHpUqmyyLFxi8pkb2xFcNLnxR+eTm+2LRT4+B2+ZnEncQnCqltaextFJD5NzUcMSAAJpc72c4BF
tgcJ2BK4sqZC8X1vPl6rt6R+urOhD8XVHbTfnE+Mg93VZIN/hbLpG6r7c1RXZh3OCeuLBwyQhykH
SMOqZq9ATgZ+xe1xEw4IQcwbNHb9DeZ8AgkrNZQNwP9Tefkb+ymIiy6uX01fVjI+WpeTiUMJxrH7
aAc5C/sdAN54SL6KRsWH2FPOcV4lSsnI/DML+f8HUwnepAAyWoe6qHy6vepC5al5uUkMxgSkPAKC
kCWC7M6TAdDaw3kRIAukoiJRQIxi7lPNQtGwR/XqVCj1Ioq9C6RfDpkzVxbmmr1X0E4bpLKMdSHI
Hmvj12M5myZ8bj7NP3iq8wb1lKAimKT1qxyVm7wdWeLu3nunUT+PTelR1ObMDr13o1SOBR6UwE/D
IiF+XWMpGSCkSRVELEOQSKjpy3Wc75Rn+q0YQegWXkvJuaa9aNsjlxE/t3lRS8xJMP2afn9QW16+
ZrRgMZBgrdluwF91d3cIAM6RsJRUGi/gLrj14zaEzA2InvZGjvkvPd7go4cUdoQQNU237BbQzRta
b42llmtRgcjcnP1BAKFZNRA+RkON5Q+ae7pXUYMXHofeFuTCXLIcXVNlWEIfw40HOG0B1I8WRUdd
jYUXD9V/dnpsMXi/78CGWAL+bJx/NuEOZdV8ULhe9EjklSW9W2y+Wa211yaStiKDNMVzunouplZv
o681v2VnSUHxNIqYvK3SVWO9KzD0ikCvAUVaqtGDSeQ73lwgdAD1JYBzdHXdjn6Gk83+TDdGZIxL
pQeylGEyJFWyeX7EJzPHjmPCPH8Th5+c/7KTkjYOvXeoKhuBWxbvk09mL7UJiDxin5+8NHEuwhAd
Dk8Y4gIFaDtejvyQcPlb37hTCxpk8MzaxytIPIQJr+9jZfl5C9wxanCoqxpnMCTYZtEJ69bswvcm
sjNBTr1+uXTIrRokOxR8pH/NmTAwXTlE2xJVgvzvNCVgAltgev+TlIi8WCS7w8u8n2BoE4PLG5Wu
lud3nTq+38yyqnC/8de2AladDzuYkhXc5Aq+IojcQu2FFbcLIAd5WP1JgBiLVeQFJLEW7wM3ex+w
S0g2aW50z/GGJiDL28MhhJdgX32Q3qsJ0Z4ru7mxUZhrniwEasF74Xmy0op48xwpatZnYvP6Fsy7
Ioy0DNLYJ8GmLRw+049+eH6M+Jaq8w4j04jJ+mz+V6BOsiGt9TRREEs1mewwQ08h3i+UICYjTaAZ
/YuQa/HsZHyKEuhUYTjn8giLGMcYMH9YqcIfl7sEzUu7uOjSIwYU4H2ecCfKTrwvKMr+AZYDQCe/
zJLmqZuJAgSm00OoV/dxOPVu/k+c9fnjUlHj0BRdW1k11nXAhOaFdnamRyjhk+NfKTT31ATkvkY9
fYBSTreoqLYucFLphSOkBIZlnf8mGcBQmDdY1nrMMA9fbwbJn4AKZIpJuw63NOO4Rsv10ZRrwtJ6
7Op5ulTHI2Of3gLF3/5ZXSrVVRMuqcbgfaESK9d25BOP/zeX2c7eG49ExGFUcj5Z+u75MXCKv6jy
6CKCGIvvp1x3us61lijFt5BxoTQyf3j6IVv9zcOpkK05HgfLQ04Z65MAPoMqKLFXZ0Yl8mimTvko
3/NZhLshfNuMwIlYV7zjMvpHm9LYmfT0SU8QhTd0W+qqqf9urm6o7mxAJniCZLGTcYhxLKlSbdNP
ibegVDuv0f4Go+NZjNDmeZVzwl0q6rZj+8U3fqBGLUvv5xK+E+KkjlHVnfhDvH4JY4K+wyD5uTO6
QIVLHbC6p2o2EDSwrHz+qv/qtHfGH8fVNGZyMs4ZcqYH1I+JzwFrqEhtKH6d2+f+yf4Uz7OtMunu
KDQi6pfUHyWN2oQlZxQggl6MG2AfQtiHY9peRrhJ/Pk4Pq1jPV8F2pYeL1yKAwvj9BVnH3ysZcbI
IhgUQVK9ZCrp1Ui7aaLQBssLMTj4/Owkltu2wh7V2/ZW5EUaTQ8vnQocmxbel9hI9NvG2K70msCC
9OnffN/59YGUi/xhFebr4oted6rS37P7WEXFKBbYxBaZGHEZe3pvWudNaPlYQnqRtseYovtlYMhJ
kDS1qK9y7UBCEIhiZDtUEnRv0rltNfq1NPSLwvzUX2025qOrefPqa8yfXdhl9jaVFyrAzzelNHkN
YAWET+9GqXKtip2CI3JItiwql4YF9Z0y3EGswcRIZf3RGGIcoOxpm1GPHsnLywYq44YsVGLQo69t
TnAEkqu6d3TXJs05K232W3S3U8AnyXebAhLUOLD9+cabmUtiuJnA2o91z4tvQCmR5RfXdBBSQ01a
ddsGdN5i/uTn0l/JOEhY5kjFFbPlmAROPB876iudZKOVpZCoOUUWhlSzg+Z+gYMjOB9iXwREKimB
Qu63zgCaJMMSXvoAKnFMUnnXjeijql5TaPxyz3UCAfgTA0dnIzq+cle757TNieTGvHdtkfvcbGNf
oL++wTf0SCgFfXFeNlIeoGzPiQ9KtxUwiXN4jFdCDcA5Eu2m6ePzFautSLtf5Wnl+LsKO+o7dL5A
fu771wDdAScEZw4jur88JxBDOf7Q8Khm0Q+38cQYZ0NFegcOOFHjPC59JUs1bP3A9zDyyIMlDtvu
hWuRq6NftmD3mufIkquEKtFmPtXtb1wmCAvBiokErYMvLOhpsUfKLyq6i/NMu1R29VU3jZuY2ceK
LYpMeS6WFbM4cM4bCfSuDjDsKPZUB7TeWwnePiDqkc+QhgO3X6m7M33o7CuZ+8Z0AtAN4MpyOXDq
SlS1ttLwwr671iO479h7BnZ17Hd0U82Xwmi9TKUMIBv5B3aZ92hoUR/1oGf0P3yeLyuGb2wwDfIg
1fD0vAdINYzPn0ob1xcbwfaVIEFXiT6VtasoKb3Z5/F6t5l9qXf3ED1HmDuVbZg82lztQt1ig16j
h7OlnUcE00w/wsUJofw1uuwEzNlDXduSr3JBf21UmZqfI6HcE+sDBsaFPgXK5a9r4JSqATQ2TrOS
0w2z/ku5is+AoDd/1szL6Sjh4tFBTbNXLWmK4k/dA3QYj+ShleLg0L2ImSj2yaxf8QIypc5RhJfQ
0Q2vddekQj3O41g16eOeGedjs/GWwCqYXpYkSToWShWu7W+TnHKcR5xVc+7/tljoHASTkVKzqAw+
Vl51ZlurwgAbwTkR5UPE8yLRiqrBX21lBX8pTVdZCD7vyPAaSWZCGbBOnkANDhdzVcRdtxJFJJXU
74lolXi+SXUiE0qfIdHlDxm9XFdQSHASRDzlkYO1rf+HeZaze7nFFDFgeBswOdHOBWSXdazpjK3T
D2g8Et6skzVpknIBRM3/K8Fv4Ul1Jp0nlHA9PPmBGEf0Z4pWvTX34LgBho1WeirtOtvP5jyFEU9d
FSdHmbmZihN2KEQS0wY/TMyQKsS5vb8AqekfgVCnucukuE7cboRd6ELWgCGfTL8zxg2an4F8U34v
8mYHMJan5CvceBE1EMFOpMdD22JvmbmJSlYpuN9TJelM0pMFEx2NOnI3BXIzk2nPcu4R9DybxqKJ
lhKyAkgmaymDyeaauHIchULr3QURaBzl73+2CNUDaYtz0Vyf/7rr0jMMFKUFy3wtaRulB6GSBQa2
gFGXlT1I/TpDDL9CD+wcCVe0BYdi/yV4nSAlkGX5oRwIu2FqAz7+SoCVSWhP9eJoFSLOmzxxhywv
eDwD+ldGpL+e50xb4vRNGV3rKTA0N4EwMqwuj/E4lKYBGkhhNaoLrSRHaFZqrBWfc01V9nlP3CPa
ilYRbkVDIQ5CFrdcsKu4loM9ar21zww9qdKgHT/4ry2YAvaUxSzkeGkkWUMYJkJu8Pj7tUPhaGu3
Kv9FmxqU2KFLVVFIJhuAfFx2YgMWV/9gR4lSPS9dw19FSrbXG3ICHZhAJNWjunCvVjV0eWJGWBZJ
8DDAQIlcrX8HLufZdt9tgCa5wXOG4Sy6XpPKRTp1P19W9lJYEDZnVIUuap5pxrZK6h3K7xDE7D7b
lVtl5MbK2cwgwyX5tySC09SCXUkZO4Mn9Qc4myny2d4J/F+c3LdXDZD6Ly6Y7LBdpNLO6342yVdA
MpRUD+CGhKDFJd4F0dwwRtbAl/O7eDJSJ/mGaQozszHrNhZz0GEq7EdzCzc8jW05ijp/YWr4l/oJ
K54N8xQl1vXqmsqIe+UdYHz7JJmPy3UoefTE2Ibdcqx6Fl/sywTdEAmTo1dQ1juETnj0tJ3oSPp0
0w82Dze5ZpmxsfjDGyJ2BlWIEyjyVulwrc13sQgvhy7Tix/FGeREE0Ug/D0AJzp4k4JbHxOkSjgo
5C8SVF8cgSY6tgoefAJdzMdLPopf2p1My2XIE3MLSfE69ZsBPpYqmLzvmdHVN8P9a6qlm9TiJUgQ
9Ad6jl5fcUqfdJSI1+QgjI5LWYoARVRyiKMpy+oiRTYcZEWRdqkc4F6MuuQd9tKAZbUHii8Tydt2
8iIPQa6dGUTxzwwdH1XI8Ejb72D7MlOIvRd3NxnLhihBfwPXyEmPtp3TXGVaVAbXxn8R5SstliMQ
iJ2xEcWjblcxCXJlR8U5z5zsgkyrxLTafTBnB+EpBlgfY8slqSUlmYvI8VBZhexZDPVIODGmdTQl
XGJ/peUJG9653HdT82brzUvbGvvFHibUq7sPwzUXluQk2W6CdeEFQCP9LlK08UfD+DnyV8VE+/LD
WyAxR/edg441QVxHOCgmMHbGVaV9VlFoeM8PQU+QqBn7f93bBMpenVHSKCSCT0Y1IFKXYQsig58v
eH8kw8Y8F5e54ahg7Ofc8pn7tLsjIWuSXLzalRrRxU5XYq+019uvy80ZYTM5nKT9GIB9jUh0BOk7
rJWQrkS1XOHgCmgePRYJ+zXl2uMKvm0Dyg4bGIJ+x0WeJMky1NLEhGP3qjKo0F0N7INttk/NwNfm
QsSDj45YFZI++xfGW7FllSaD64SBD+GYZnYlTLvWAk2p9UBo8/lbd2XKQkzeBRSAuQ7F0t9/OkUq
pyLpbo5nd1Z4AQcJoJmHpwAqsGAUxwdWRFvS8KqjRzculVoqPZbW2tjeIDm1m3hK7eG8OdPaAmMY
8v01GLZPPk0L+zLavGLVPjfLyzV06P55ZttYwRhXx+IHV7oZWlla1pzobLN3KNzFx12vQYqQhG/n
K2wUFqm+HhLg2D9BJr7bMJC0o/G5Tm0OIAxLQVL4SbFC7y8gWE+W+MenfGN1qHnjF8KLJwIlVdzs
CLtG+bB3a7GNCLZ6Dk/jPoRFZmdWL/BkOM/0TOOLJLds0wggngj3/TkiisdqlfBbN2DcBVEO96er
x1BklUT3PRcfkui0+4Xz/i52sXZpqeQr/t4wcGqJeH5ri4EYv621XzAEaUO21VA+k/ivzVbHO28d
mMQ+0zqtSopvr6Ihdst4ZYIXsqdQdc3yftTXgYfmZmkBdC/2uFwVr02NDCtsrS0O7PTr9WkvIvRE
AU+/+U4wWhrx9OMLthMN4RgJCZGfhSUYOqZuImd1/5L3gjQ/mowHz4Ih/IWV7c4LKSAcpg2dLO3w
c5cXu+iTa/D008Z7vuGJSEEp3BgZ5jppUslpvqy38ewGQQmzode1SWZVWMSL7YuR9BNwXqujgThf
QR98Esx7hUCSCYEMN2rCUdtF0Dyg/ZBBQb9xhjaMad27UzuEmbowTUxqblYO7lDGpmnb5FE5DK/D
3ruZT7794TZQXIgRJB6Q1Fs/OwbpgVN/llzeq0ysHoQ3c1vsW2NjbxViKteQNtiY9Iw1eR7XC5Ry
aTPHtFpKdVHIhcwi3P4pGQ9rF9p9OHkOL62nHd4JtvUKdoNbugpiaaAqVxR9UGFMadRpL0p4o6FZ
VRAyRk+memC53ORuYf9usY1Gzu7jxGuFOBOvilMxdLlSW8UMO3VzZAKpulJ9Mm2phxEA3S+tcjLZ
Te64Fk8BlchPBk2vQYpGdwYqE6vBnadsb7vDECEWvcXZ611NBWmpx0X/c9Me3LYX5iCgUfK6N7HD
nDUn+qNv1L3SQGjtTjRgJtOM4UwpzvCQe0GVl2CjY43+WMw/TBx9n2KTxz98iSRuYxt/HcmVuKBW
GwG5Zh8F6bdDFqM7ad0X4DAIkrXyKphkJFtB5xCrrGDdm1YY76PYmOPaYEqDEiiGhZqhiXw29y2q
yKl71doCxyXa6+CXSC3c5Hxjr+SoqMOPeZnBhCnEu1rK0o1VyMwQIBSFEKqXhxqtyZEP/+0A+SnQ
uWCcWu/51QagVy7DyY32qAxuJULEdmi4KfX/dWco1Wib8wf2qnbvCX/5EAGT5mLOn7/Zlym7WmEt
vAhgj371+VXuaH2/tnm47vqv891ZCCSJ1oPOZY/jcix6PJehZF6ZhHYUnWtcGVmSYR+xlmQKyX2j
gnF8wJZdbJpiuvpws8s1Edfg6NKR404tbnkauJsgLYQWDiOztcCO2mfGMVgzieldrpkGlrCb43af
0W+dZY1SpX5jD4T4jQxJo0G+rhzoc3pM2BgjKqpGLlAZ0OpSQFx6MrTtJG4YCGye5u4UawKqKT5r
AlGzx1wZ0B1z2fKHqJegGMr06TiFfwjpxuCV3lLOmY37QFThxOBC4arMWp/Vmnd0lWe2J9mFPEmZ
hufKnzvb3wtW+noo1QHw0LHuKboYG29AZqwiyken3jrANtP2/TOYpoY+2VAkRRVlAFx3NWYV3X7T
aEnm8Tcgx/caL9zRw9bkXscinpW0bUsYgNuvEkXikuZW8QE9ag6sxnBHDDOnyuDGbQNYAPKv4SKK
BAa6MMtcjvYJ1kTfcPgAUyg/2mTpehkG9ixUUZMvYhEjNhkCARNAN2QBVz7cf7T92ynZ3FM1VSwP
jURnfOfcuLYUgmJH++fGG7yFo8k0W000HpfEnDJIRWGn7HRazLr48CJ5U2VCTuvcYyrbn+2oFtb0
JQsNDG4DqlHLIacV8u+i++Gu064Dbb+aN2+uH2owpRhXevX7qXWOJ6O6+haO81OgdDmKSiFrh7cF
mmAweNuL35nGxv/4hd8kOY7pIrP9pD5hUR17/hKlhWiySus4MS2zV6+zEmi/p8WJlEiv4BZ7DLiL
uovvwnZ/HrRxm6qyNB83O9Ad9nMCue/j5RGi0Z65RxC1SivRzRKWr3phebpUrSOGwnBZfFL5K7nw
Uj461K8+xJAasK1oNdHljdylDhYNfZy3uk8s8rUddje1KHMVXWHtdj+RFKw2QGH9MLuLNinBMwds
TGKXLu/qT349o7+Giog8uHvYRxIeYsCw0JROShe23f4Ud2LINBH9pDl1HQIcChOvpif1pwugukxz
VrgpmsSLVXIm8Slhbs4Dyf+oDBG2uGqrGQ93EnIFje3QOU4iu0zdOUwcLJTHQaOx9fm1OW9zeGN3
tdzC9XDuUGQpy+JYOfAETpz/WjQPlkt5tnBEQKpuzjouAnrI5RoNop+jU67IOnNWb9AvBj6KkpY8
Jna4IjWKVUIo8OW27i0uvgK4r0Tu+J18XS8w6yKuuN7YLFRt4kj/+uyNVxKaWZBDlPcTe1eQmQdJ
I/AvRj0uEuQFYkc+T5h7MNVcEWdjN7DCuXFdPsj0O50DFsxGqhxrt76gPXumRr9wJ3zLYBDTIY7I
Onwl7lY6QZl+LzBBrFq7rKR5HtpDRTsCKe1DF4+kejuv1uS43ZySiDPcOF5eR8oIYAJgauCKMjIK
fJmZTOXX1kL9hkVMejo+OEYGdtD9EG+lOWquiTlNDFFx9ETG7XUIXlUN6b3BFJw9e9Af2GvaXTnj
3dU0AzUTOwp0YIuxwf2wwFIZ2+IBaZkz5gk27pMKWBtxLxkOOPjHa8wQMgBy9DvOq9K+JnYNlyQy
IE/Z6CNDSDhXTEbTrfEEu4rDV1ioeI4dB/c6MXtYEEwiABI+KqD0qfhlh0fKfWdjM/E5IweJrvpz
1TE9JliF39Or2kKk81tbWTF1qZBATOoOU4EmlLsyNCK0Zzi9Dp9QW6oMtnBJ0cRStHkydryFZXku
+bMb1n/DpO/JfjwHJredsIcS1QRu/d3uYMo1FIovKMJPEIqnDXHcjppeTuZIhXD0G+kpeKirM655
xKHIyRHS1guqxVNSyRmKgviFtvskx1sMPwhFZ5KTYxYapAz+Q4K/KZwCXMIXtRcBeCP3qA73RE7X
l+gzr+xoztB3YtCd4PKv34NLve8j3ArPDHv5KMuubXrzLENxg7wslPxVIWDj0dQP+29/slFna74s
4DD1JetaDZLliTQsV25aM1RL3lRw9ALUXU5+wJSP8BJc+3jKE5uDbZdGcbhEJBVegvQ2jo8eRdjF
ebhRJFrYAVpKKKuHbqa52pj+RQBCwXEVVYyOSU1R2dLxboC+mDv6asfokA9TGF1GLBC+bgJx93HA
srDNCjg8/bGmJturcOX2VbDNeFMMsS1T+KSEAINLFeXqnDhIuX0F/ywPORH8HbaVCq+toAaF97r7
hbvbaBze6ezT1Ph4ITZrH4GJtg5Sq/zLE888y/X69cbuAtDlXDmw3OM4bxAU3AxDlGptTzuACuj6
aaux4gyRvev+eDYKmhBzDjjJZp6b7rEcqWxP87dgpXl3QMLPSpQyIySYlkqT1HvTmfPEncss+KdM
G1ZmpwrXHSiKnVLlAW8IY2kWMv+HO9CCsFjcKEP6tp5X7C0SpTzTZpmnOOWhYfMXwOFyz+4vIUi1
gnBEFjfQkFDkVYcOgpJDQq1S76oLBz9czh3qt27F+76oFGXkZd7gJjFBbttemJvLeRKIj4JR79o6
ZE+WXhP6kpG1de4OTTwIs9104oyvr6uFfl7nBbbPk2Jyeg/H9Pw8qPnPd1MOi+hUQ31DOlljrcfX
6LP0wB+UWh9DongECKWkX0+5tBEMSngrivYVTIcnMwPYHqz7l0BvC1Lj/ogxGY167CQ/2/aX/TrA
zhnTLfp7G6BhTjV4dB6hzqOz1J9cUQGxW+X2M4AV2SabzNho7xoyO4azr9WS+pP0RESZh3rNRon+
L9+zV4HgtKA0tjDgLuFNVI31lMfHtliBkswAc2uoF20U+adYvisljms90CDpd277FKxCy7OctzEo
vldK1lqNv6NU8bUQ3XnlwHU5sn6gtHx8oCnHyZi5DRwU0TRLxD2ZzFV4fnM05l986uKzDIPsU/mm
zx0JtPGly1liw+DUqV7honVfbJ1+VEJ5mIR2jWonb1/7vS73ANIa5Bp2yuYNec2xcujrO+YvEi+O
cZTU5esnMbKDJKVs75uTcf3k4Ckwt4rBPfU18IhvRUDJgTKbUSwnTxAD3XIi5gj2Nb9I+s/zC0J/
18m1E+9dC2+l4yS4NQRX6zn70iBCKoNA3d68pZV+wjReuopk8kBYo52gXn8Kj9XHsq1ggjv0XaCl
I9ws6PrhHqKrGfwHawooSeAph3yXkue6xCRF1u120qjRycdlcToQMGN62WBg18Uxp1QaM6RUUSzR
Wsy3PH7T81rVWFULT1fk5TH923b/dZyyqKKP7EF1RKl58bV0j2yW5Dq1VCUAdI2CidDEvzh1sUKb
L052YisOjbXfSicNz4gYokpL2sW9bN9dca4NIY9OWAPC72wZyXreiJfhnSiGUaszA/LAhSRYUKhs
qi5Bf1IyUb8HR0HStw9DxxeU04OgpKqqc7BkxTyQC6g1CNVzWH8S0J/vjoSLhBftylmv42spImlF
8HKc7Os+zfxuL7x6zbUTq9M9L2O1xqaPO0Zx0bs4X/TKvpBm3ObMp0yTG/N2clFXKiU9FHz21V9x
3PpyLXsQ36KAspArr1IKhA7N5N7hkU5Ka//WZhtZX6xvYVxRMgEXum5hpbmzpsrPCO3mxtLZv0Hb
9EGWtfZ5uRnn/CUMoIFnNnHwkYGH/u3KkOS6USlqfAtMw7F7/LWSmb9rbA/tcToKrGn1irN53Jy+
+LhnhU4MyPiw0a04KsRZH0Qk2e/z9fSSaTYo4oG6LiCC5sXI3Ql6N374tT25q5AzPAstVHqJ5r4w
+SvmzgA6nYseYYVN1+jXXzn1/I7ehR/BsgFu1o1y5welqq+LEeQnPM9H0pL42Bx1IszebRKZkkun
gq58o6VVXO6Ur39XNzSvm1L/ZSenwNofLYxEs3+XDfaGXOlRDlcWrHqnDzkxrloKQ9oyDw1BalVY
PEPresOgMX+QpVYpetK9A8I2X+YwtUpDH6geSfCHqiMe4ikmy16WsJRRHbGSU+U+gmAtPhVWDjjf
WzLxmwvCVR2xnEnXWmqq2Ax5BQ/6JfUOFVYW79SeaPXpc8tVXpk/V9UgMAbbg5ZitGMCbbb+uP9b
DtmG2NJ4OkOplPTNqD/WRyZ7VAa5B81g/iO1GQamtekTNVQ93gb2KonhzXvWgtvgYF5QbiGLco8m
woZh9IjFLDNqhlBAZebiBaLxTlypymatxyLyPCIVRhJZw3Ubor/WLJOrR8BLI4uTT5JYfysY3uqu
RF2/XXOx3tneXmDMVsoi4h+p6M56clM5lZkRBaec87BulxZ6/5MmM2vO6IMd+L1UUchyq7McYg3x
OOvdh87uvso05TxO3MHphOnOtF36lgExHXnL0jBG0bizZwBaDizGYAcv7jxq8mEul16D5S7XhwRP
eHr7qx0tmjpjnG/oRzNby/sVF9Mk8trziwZqkIF8PS6xKb5GbMpa1CSICHidhljc94rQVInZc3Hv
jt6SY9tZKs4/Co0EEu7pisU+Ipd7DYmNB/JuKlEc4a3gh1WJ3T6ty4iGTuVqOQ7iI9MIRd/UpePK
NUxFFlFoSH0d/+1JSAP//y9612+N2/x3qtpQ1jPr0dC/x566SKLeXBM6+KVhH2MzqSlQ5+8dv3dj
IAZFeIwNTrKz9s+7eIlj8iiIHM+G3HgnLiECB8Dz4q7SkvD6NZGeHmOahGWqpn6xbN89YXvwtqxN
ddAcGht7hWTarPc40a096v/xQ863s9ID64rGb3uxgA5pWjfrx/FLvA0uPqC2luVViiCVVtr+VI6P
Z1lvPPLICaUQP2raxsBLKJG37kgTd3GT6LW7euga4D2PoAkQpbbt8d29Fbnw5D3HSRMWdV1sKmVA
Qx/VUhdlx9iXb8cy9sZbh87XKhqCCv9p5FlI8OzwcA+bIG4Mc8OBXCicv7D+Lzf6JJlTGVPEEEJw
pEjMwHo18TKRET4DwEmy04vf6/HaYsADV0yZgFs53vprMFtmy9ue+S964aMXtVeJuvVZ+lKRYiSZ
srpx9ES1oyw/ZA300iM37FURfR1bG83QEQX0Qa66Da7RNUYUqGbA2X0HxpsgKK/Il2x4G7E+yoC5
thUElq4POOGjbOeSiRf7UgmnYicFcrsirSC721mQSJPioirUoswvVs6HFOFJcCwQ9biwSbc6twol
pa5DaTu49XlB5xE/RX3xK8ItqRUgE4io4h1ukuK42pNCx4YNlhndtnL/LgdnszhJAzmHGYe/wrPK
tRB+aYD+v9wQ43xZD0llahUfSZHpYPXDmtt9X6cKn+6Zghke3yu+bcy2Uz8QyZb8fGPnRw7k4HpV
BNxbBzRaeFjMtFpqsvCt1BMHg8jIF3quW2GN2EUy/cIdyY/hnJUipH5M+EznIdYV7Hse6fUL5jI1
xQnFzXYrcxXL4qBD7buRLnf4bazbiKsXtagr1zSmUzpE9VYGJEbOtfu1FLwA3XQs6/iPh0PMCSyc
XOSDaFS7WnDWsCP1HrxlEYM6dHWimMVddlkNI44MuaMG9DNnLvWuDm3UkXzBztGFPMAiVGE3EAnV
3WS4TSf3BunUYbb4DvPM9jn6hWwk9MFyU6q4/x/C8Db8AnNmxMKOXpPQRzOXdug5tKvuafu6/KdH
nDkTMGLlGuBEGAEod35W8ZIH6hUmOl8hnsZLLKgwNRREb3h74Vsl8GoPfx1nbApf9ckbX8srbxeb
qiD0O2Utxf6NUk1u3ChB+QCSZ1AbafRNMLDTfaX48oO4eMGHFEZlJkStfNxv3BzWjhgr4572rTS3
0xlOBBwfDQ9dCP+gEdaOG6ilGX8R8rwRCiR8wfq8coUw+3DmUF37XUmbB7rsEq9AP07Bw71yY+ef
Q/R+mLCJ2d+OyVwbaH9S4fUciiyxTXOQARVG0YXZpvrv1cjW333LTNeLrnWv8+yS439htC3nDm7l
Qpd81tgwxezA0X55eq10wPejxat974/mCNbUflr6ZJNeVEApIcwd+EuZFVt5ssD5q5U9fluXfYho
thStUTpO8BbGgzv90HbpTmjSo3Yt5lTmOBBg+URPCGjnIOmkrAFrfhU+2ApLRgQ82VOZEJ40z7Cs
y1h386MIUDz8q20tN+Si2SSu043qAJyOpztoI5GBdeU7dkcF5Ot1birxvacy+kNDJhZ91qsPgzG9
7kVt5K5c9vXAo7m59HG9Dx8QlmcvuBnBy22tM6X/JPn+Bn3Cd8U0MV15dR9THsdxCa+HQcs/sE2O
6y6Sw8QdN6M8idd7cu27dR6YAPYnyv/6h0CJbmhfcWM102CCMA9TstXW8HImlfBvomCJhSUsD4aW
ub2D1vCKowkSoFUUoTPvLzrhGD5AyS+e1Qvj40MFGYnNc4xcZwyG7xvUtC5HMpY88sINOSLWRtLN
twXGbJmC65AYHWL8pm3SHK5V0jx+iy6QfkU52ilprsSyyXGFfUdbIQhwksd9KrLTq5dD8mZj5Nvj
4oE7yBlvWg4Cymm+1syG0nZoOYGjEUrtjSMSRzQ+v8yRVL0+XuN+uIJUvh2Whxzk10DrjlrYKTWY
Y7TZ5PRCRg4MRMeyQT+JGE+SpSRxA2WJ7OfXmHUyAhu8zzl75zBhYWo33Bbbh7OVghWPkwCSmebu
zaCzgYwJI56t1U4Xpj+ddU/cnfZIXhYcxWqKT0RvCwB/VYOhJ8C7fnxi5b7J2ijzkiM2ttMUEoKD
khQhlIqvHW+jGYTjsm4RKhDEgxme5T+lZ5HF/Q97IlXqePGwGeCHs4hKmDjCGegaS/ftczMdN4ug
Ypo0FD79GvuzB98J/5we6D613m0W3pnx0y2Vl9qqO2wiVJMVXunWwJQ5GSi9vgVcwiP2qWm16ZMn
SqQPPFdsIUBqikbXG1h5BzFvi608s6Qytyc7Saq5OZYd2OFw11TJw/XQa7WmZhjrFGtWKhOAiIbJ
/3VagKcHeKSCQ83zUQJlk5KmPEngFrF5irLt75Ox0yRMJ7DHDF0GfP2XnKnOcda8vRzoOTQUSxpQ
XJf0GAgWD4OyF9llObmb2ufuuVmihZVpfSAcF+ckDA+M+Hewcmk71IvtuxMkqHup6+i5KURsUHn6
aQeV3RVfxp0Y9lyM4nRK9zSFepeULy++oVDco8OPgw1xakEgqNhH57pztaFA8Isy/wOi6HI3y3tR
bZ3Civ3wqeKzKsb8qSJhbtxNNliJgs4nKzBpK8b2sG+R45lgHiAYfXoQKGsUurhtnEtsBOWA/fH4
nMhOWUCcMKJLugXfWTLcPdEIK1kBzTJh7u3HoxIP3KG2hzYc3ftpYLyDBKlMWZZ3w00AFgxXYXgj
tnhPhXQr/rZ/Twh/LfcUF0ZxVbxv1lpOG6f1iQ2/i3x1SPtmhBTV+F4Ug9P1faFMGkwpZQRkRKtm
0sMBC7jiZ5wQpFK1c80FZQHBWfVcS0l7LBr2CoUz227SYaOybmO8/z5yzu+fhM4pcwL1N17isolt
PHDso9x1q9qc91K4y7GSe3BUF7UM2Ueib3lb10cr0RzWXlSWK0YpdA/42iKNDmD3rOdt4aqn5gNk
YeHnOlv3YUOsXZRiJRBBJWAimamHjgFfg3E7KaZlQvAauKvvYs2p5ISm3hsY3GL6Hpq8ITdnJtEx
/PSi+hWJpZuHcyhySYXV/4/Eq7yA8WOCKAC7kW/QIFRSHmr8TKEFBVzw+jiElCq8i5IeIJ527Vtf
jqxV5XnlRyQy9hGvwyIkYya8TXR0o3iwlUNXPBT82SWBv2peODKMXJtFami4yloo/TYQLkiCfnC2
in/nhu8oU1fBlz3f7uxGRZqR4fzhpiBZ3IOPaFrw/+3yXxrfhHgSOySBgrvSF9UpX+h2E6zCUHHK
aItmxUxT8vvUIzEb8wuSaI875EyKsiruLWgq8qeT95ffD5nDcz1hOffu2yZpzCM1bOOAgVey3r9e
f5Z0foVO9E3bUH3GBu6XYhu3WwxCb8pKrzglYUTLpjLUZq3M3AyYMzME74Omiw8xgODdFVFP7FEY
hdr7+KISmdWgUB+G3+CMxOhWOiFhFiywDCf3DnVq5K8C27KJusLdKL+c4YErlvyPYWAx8eoJOcqN
Nmrl0n5CSM5tOKBN3mJXB3cRhAbkMniTex1EKExY+1/DPf2DaYJFNGM6YF6Sqz19ATO07S1mBTDg
b4oUIJ+OHvGiG/Ct2832xaSB4jmQZTarIxPPughRV46LksuViYkyiTbeoUjCrhLwZZslpeIlSwwR
xYiagi0YaGL7ytKTkwmGnbKunJmgrQOyUbHR0Eulu2toiHzj9vdqY3JU/oHnmVDLCgGZy1wWTvzn
QIk/IXzj3/sHAPzK3BpeAjQKUFp//2jBG6aM+Y/iMNNBrRB86B6B23ywt+NJf0ZY402PbO6Z5pca
CNcrFfoSSIxiNhSDEZyBN5o1M8hu5sQ/yHXFA8b8S5+FsCg/TRIRVgTFqosDLkx3stXYkh4Rlpqy
RHbNny8h+dWRv17OefGeOp0VqEsfX1stuuoH/jIQ
`protect end_protected
