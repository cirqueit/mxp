XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���_����������?f��N�jv��>���:Ս?���y��!�S^
(M���B�z�0�$>u�?If�\��y�Xv�6s��	5��68��A���{ޝ���7"O�T
Ѷڶ�Ѓ�f��|����A��ݮ�ň3Ӥ����b%��NzI|f�D�BeX�'�?�̏$Lo��]94"��<z`SJ�E���Zܧ�?�3�^{�Qx�7��> ��}}��O�)���W��K�tꉶBEa�����M,IZ��+V�h������nh���� �h7ի�3��G���t��X����%�`xm+� H� /D� Z0vq45�%1���o Λ������ɉ�����W��M��f0�"}co6{�Y>+��Y9�ݸN���|br9оC����V��M�l��^�3���W������^��H��1u�M�@�#��\$��۫��Q����{�=uNG���O������7~jM���W�Q���юS6z?	�U4t7��#e+��ye?�f�y���75^%�@ �Ĳ�	j���O�pY� �5�o7G� e�v�ۧ��md�ä�X.�̩٠!l)�B����]@�6��O���"�	��dm=ѝ�Գl��h����[�	��|(#ؿ�;DR�J��+�{�q��t�3��z��FB�%����d>j��*�#t�5A��u>�.O!ct)`;�9o\Q���C��d#�M�fT�eR�up]�ך|@XlxVHYEB     400     1b0��1�^k�-6��%�L�cE�]�}�*�>��� 4�D+~z�g�pb���rUW����䐩�f���<u��{J���D���t��b���
��euF���� �z�Fy�Y[]�Evf-��XC;,���<�m�M���z�N��sK�$�k��]\���b�H�o�X��@�o��'K�q��|���uC�Z���|�
�3`�b�&|Mf4�N��R�d�������)9^+n�_�gV��Q߹m�U�Vp�DsZ�?��B����>9n��k	��QD�I��M�G�=�$<whWRV /#[�VN݀� ��zpC�~L�S�H�m�[}�&X,��)��۴*;����S��NsL�co�~2��4��x('�M��m�h�������ۋB��`�P	���ޱq�l�P�����Zj*�XlxVHYEB     400     130$�8�7�&�jWUvO�u���=lGI��x�SLW<�L��_�]����U�^��,���S����,�؏�%g�뎠��1���;�U��(�O2,�d��Yu�B��˓W�f�<|�C�/}��ܺ�B��vc��%���z�9��h[��J@:ʣ�#�Z$nhN��� ��� �k �~.�X��k�?������a`(�K2vG����a�LC��1K����|���J;�����
��b*�A�Q�+/_�:~N��2���ŉ��T�&�cV�js�C{hR9�-��}W�A A�G5lb��M�XlxVHYEB     400     120($��O�_a�$���O솮��6�ї���W��RwJ��Wẞ  �Uy��fI6���&2���Q�)�����������G4A�+,�Ñۿ��'~i��k�Uf3�Sg���6�唸%ƫd��
���H�lC�]�d1~DDR�[�6O�p����݀�|���S�E�H�R��g����&�nw#��A5��+�Ҫ����#�$�h�T���h(ւ�5��HUC�6S,\�����'4ȱȱ���Ƌ"�.ja�r�?����c� Wj�,���D��,�\&v`��3KKXlxVHYEB     400     170�f�������L��7�a�K��jd�v0ſS.3�|�L'� ��)��?͇'��/��N�x�p������"��1��1�"��ӗdw�LE=����HBy]k '��c�?%1 ����w��'LO[o��<��_p~����)�tpy���wܮ�AX�.���W�!tq���Pr�!�J2���������,����T�vʑ�«�\
����u|o�?w8Gq��0g,;�ӽu���S�*]��*��#���Pu(�`�[n���M�-.�T��'BT�����x.� �U�.�#4�vG>3¯�|&-Ƣha}������}:��7$�K5-g% _�m
��P�\��&��XlxVHYEB     400     1c0"���4Ծ{G@*�v
w�@f��::�i��s��Y��'����:��1���xpn��k�z�0z"��͎�+ѪĠ��!���6�2�B&qٿ��!�<I�G ��EV�
%w�;���Y���v�{��U4�g8��9�c�\�����E�X�q�@27I�a�
$����]�8��B%28����-���d�U�iڃ�e���B���ほ���q�:ʋe��u�P+��R���^[r�0��v;�/���{R_3[����_U�.02U��Ihrr��5j�����z*�콆ج0x]�W�R>��ۙ�4�d�a�9�O���Yf���mZ��1����6��c�`;�S
��F+�=S���|p����c� �O����hy��;3EM��S]��&2uE9\H���ź�~ZNw<��)��v6�����侗hFXlxVHYEB     400     170)K�S#���m��*o�&�J5>�r|z��Eʀ;Pr���/��
`7r�g���	q~he���h�ܓ*�i�eJP�MݜB{Js�ry����Qd��(����L���w�mSu���2��-;�f�CoNV��Q�蒀��k�Е�heS{��Q'��5R�������y�u��<��(����j�r};+�誅��23��胂��w,wVq�yn�e2A����!Q���n6ټo^�烫 �����>q��Z��R��F�w���9�
��H���S�/n�	�U�Rs��&�kZ���Tĭh��Gƽ��еɮ�#��a�@t}!�S�4��cUf���3:�1~�V�w�����w���e�_XlxVHYEB      5a      50��h�9�ꅂ�ޚ�����ّ��H2'��|K��l�H��<�TL��%�5�!�M���>���� �r�DF��N_�m�