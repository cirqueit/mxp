��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����ͫ���c�T�#I5Jâ ���q����r�ǋD�
�g��;͚Z�r���m�R��ͅڅ���p��'����
uD�a�בyPևT�o���w���,�:��y�C�~��d��s<@U:�q��IUR�%�:�����Rs��q5ؽ��4�eaٵ��>�QؽA\�����V!�W��B��6p���<��� ��V��n�WC�����\�Fg'�IA�A]�-M�s{	A�R��J7�_�D���~��	CL�Fh˳���Z6cX����a"\t��ŝV�ӭ��\�2�?�`�<����G��ƣ!�5GI�EV�bt�W��u��ep�!{Lx�y!PL�
L��z����]��G>f�3��"˂�W%��C4���0���]�Wpҩ��%S��=F�ATb�Gu"O�:%|# �Y�sʦPF�~_ڑ�����!����~I+�J��-A$J��j5�����\;xYj?��r�}�``3�i;�	���*�:���`�=Ν�EY��Q?�~����eE��5�t��b�>Ϙ����n .�
Ͼ�����ˆ�y�l��+w���Rn�0�9gE���~Z"�C��T46��w;>��g���v�=��_�g�`|�Z�`ɷ���6D�1,G�zp��+������}���1�(8W�*�}QwmC�to�8`޴2z�sփ%�3�8F0$Xqb� �(�`���(n'�{!T�$�����m�UV&�*�0{�2T~��M�TK�6�(����ץ>�b^~��}�M��UA������!����it#���p���]�p!Zn��l�XfDlN�6�w>��c�'T[c����i��� �ظ� K�'ٟ�yq��ђD3�����z����>�u�o|���n�;��-z�
L�^ux��]�qs��QD�� ��� r��<dr]�Ej�D�V���AM�'0��g0,F/ j��t�ޥ!5��t]C!.03������d��;�s�a���������S��v���bȲ[,ѩT(�Z��o��J��iC��c�/�4��bz*�n d��ih퉝�j�r����X"�>�Д̲�BW�˅������#���tV���a��8�
��K�Foi��ەB9x����r��c�sb��+���ׅ_3�d} ���� V�G�û���n�|Isz�B!��$ܡ�"�N�bd�^U6E����5��ǭ�Ծ�h��p���L
��i��Q$���nc�&n�"�z�^r3/��.�*���D �!� �O���VPd��֪"nѐ��f��'C��3�~D��@���\ ��9r M�X��#������{|���D*����5=���^�0�9M���U��'�'^D>�(�(�x���>a�Ȗ�G���w.���S�X�n�P��	Z(t���}?ܡ�����1���}0�,$�F���8�i��>�J5���\$u�ywwY�%f?)�v�k �f.WQ2/�j�[-�|�h�U�Q���M����6�a�2�V,\�	b�hɈ]�Q�H�K�8Lz���_� [I����W����-�h��A�;��(QTEc�$�o�^ZHaT �z��K�Sݍ������؜9��\���W
f�m!���^zR��zȨ���`�6��3R�*d@)|f�9��ߥ�V+��>��;4�8�:̝<�����Z&P�8K�W�;��i�(	�2#��1C�D�*<F�Ţ����6Y�\��7U�+p�1�MU������ޡv�rĺ����������ױ�[�I�ܿ�:f�m�Yڮ�����{켆�Ǩ\'q.�CT�J���{�/iQ�_��ouǾ���{	����-�f�������y�뺦]��M	�+���:�fC�X@�Nژ����X%^!���+���0�w� 4\�Ϊ��!�4��.�Z�1���5Y���u�nl��W�D�q/�(��O�S�����g2$űg��L�;��O��:��e�"Q_D؜��o�r�JAt�1'�,���k��k��w�tsZj����WWbj�^���#��[�V�/h�<���������F	�����!�cT�5�������Gh&�p7[�٤�E�mZ:=(-�@/T=��f8-��<b��2�Jf�m����WT�ݣ��a\ӑ�q@���F����6�O	�*�?��6�&��	�5���q-S`�j����S�Du�k�b鷤�6F�Q����n���>O��n��5\H�U��:Xњd�=Fe�1^@9}a�`��d���4�
[̨��,���d�>�tv�|�i��t�:>T��cp��T���0���8H'~�QL	P����|Z�EZL<�i���_�z�Nn�p��,g[�����:#}=m���vbth���w3iui3�����y���u_ͮ{	4)�JNOWq�os� C������G����`����$y�)�9)�h)FX�4$B3��.���S�3�T��֔:�i�A|_���h�x�j9�rG��:�*��	1j��sl��ҫ*�Z��Oͦ(b�5�)c%��H�
&���jz��1��A��[=���Q�̦@�"����&��[�t�#?&v�c��d���a�{���*��xܹ��Q@��$Wo�N���d21�l��ӭ%8�Tp��0L2nKr	�?�E`UjMc{p;6B��V>7vg���Z���n=B�mh��*��Y�CAC�K"Xղ��h�&m�J'O���{RF��u�IA��|f�//@�=��{�v.���V�'�X8E ���_�h�J�Ǡ��w�^ɋ˭�Z��9xR���N^w���FΕ�D��؃�F�{U��5G���we��J�$..>C'�K6�v�ç�Zu�mBX'��J����f~��%���L�)�E����7u;�k(V(m����?}ㇼסLzǰs� V#=���������j��hV����ՓtƉѱ�Sʳ�7����m���-~��~���k�4�\���4_�
�U2����.N��;�!��Xx�Z�,�0����^����8�V9�^�e��9��{Io+���+���π@���ќq�F �ʥ�D�m$
���}�h�׫	o��:\ Bɑ\P���cV�F)���?�'�X�Y���J��-��6�ɧ}UEY�XКc\@�D�[�E��k�z]���⠏쪗P6p.�D�g�b��MF���_�>�t�t��P�����"0���7MaJ�LT��+Bq��t�Q�2��J?��2Fȇ���J�<:2�������I A����L�b���2�u��鄗C�}��@���G%���ؼ��t�P2=Bl+���.��>Kn�H�\<m����y=8�c�W���(J\��Qt��}r�E�s-�17�|��������O���Q���������i'��E�LC!t�G��:�LwIS���j�]ɉNXo?�8��;<��M�q�	�;���7о�s�B�w�<g����V�Nz�r����.w�Na��Mb��;��U�p�%B���;��K̗T��s��H$wQ|J��ϳR�c�e��c-Ф��F��o�wO�$:AB�M?������D��dZ�=.�n(?��5����W�/���q2�� �m���]O�}}k�j��oFԜ���"qz5�G<v�$�'��DuL�@��b�'T�'�32|��J�72>�Q-�I�nO\{Y,r�����#ߒ����2��EU�a���::Vx��b#B�p^�v.�$��8о���K�=C�
ʀRGz�3�׸<5=`���?p7�c|]E�[&�0RL����x*�#���
:�R|=�FT�6V]�ᤋ��������\X��<T��d�=�z��o��f��j 
���K���c��o	�")���w���#�D�������qvQΘ5�����r�X=�<�!3��7Sw��f�0!�J��@�F�*��U�x����>L������IA�dc Pq^���§�w���3��z�*@����d3����P�:�0D�%RĦ�FHb R�ѭ:q���r��p9T�6�ߧ�����aT�J��9�������# �8�/�Z����$QT��<���AВ��6�4��K��[�t��nңD��7 6��~\�98���*J�d����\��H��J�ٻ�%E��T��ۇq:���v�(0[흜b��-���yp�� q���c:mX\�`�!����Z�hds�H_E����8�%���'��U����+uU,����#"xT`r��!����T��i-/EȽ�3z��!:S����0�p�֟�6��YH^	����5V>p���Ə���]�e�#H���o�I>�G#i����F��G�>�_�T+�����/��ng�s.	��#�rcx�7[�Lz��6��[[�w(BI�����.\e8�޵�����f�8��xuq�+RSM1㺭�u�����X�T��{�Ot�I�ʿWz�k�'� �BJw>�������0O��T�|�~�����(�sø�8.��XE	�a�ϻ2�~� z��g�Y�ܢGr���_��L��ᤠ=�,j6{���m�|-ƪj vl�<0��Ӵ�U���W��ظ�+=��0�ᨘn������Y��8If�te��1�[�����~b���Õ��㷻�Ռ���x�&��`�L�T����V�X��h�{��|`-�������oLޖ@S��8efz��W�Z�nF�����1*������cWZ�c+�p��Q ��`���W+����XNf�~u����x�h@��'{����9~+V����KdsV�f��0af4Wmy��~j�@BF~���❳��Nv�h���!m��<�7"p�(�y��MƉ�ЄaOF�� k� �� ���e)�B�@��\iT�(��`��S2��?n��-#��*����`y�|�tI��.�.�rx�20�0b��Ch\��{ �w�����x9UC���K��v�=����-�'��0�|�-�Z3�K��(�Z?*j_�=ktn<�m4���H�WX�Rk�4�e�6N1{.��-Z��5yT8������p��zL�Β�ڈ82�&FE�S��q��	�\����B�ͻ��Q�� �S9g���S	L�j><���>����::��T\�8���_q�1K�RF&�)7��'�/٧$=b���������X�g:�MA��K;u�/K-y�����5K_�m���E���;0k�ͤ�F��j'����8L�#�Ņce<��F�ݹ�q�E�S糯J����C���U��>	��3��R��+�F�z��+���f��k\r�)L
rS"�ŁI�Ƹ�fɢM�(��2p��6�~$�אl0%c�{3��mv�凎�����'�&K j�8x���rϡ_�j����A�e��i��(x��.-��\��E��jv�ǡN�8��я���A-�0�=^������v_�Ӣ�Ѐ��_@��23&��t��l�&	��jU�����u��+S<s�5�g�
en��b׾�h�[��%E��B��{D������|q�l[�Ƅ��,z��8�P�Z��p��T��g�$��r�}r0�QE,^�P'L����%��3�W!]ht�;T�45�b��]xu�5�dl���%��4�U�9ȃ���m�������!�
��_�+W-�2�CZ])��kq�㎿��Ҏ\G:PT3�3N��u֗���L��A�f2��.��.������׮M�컁�2�N��4��b��	P�BB���˜��2�OH�^�� ��_K����D(�y��t�� p�h\����n�̇յi���Rzf*��+��0�@�㲫��V!�"�&��1�q���e<��ڝǨ�Z[��e�֯�̇U�8붺��	sU�/�˝�d>�`0�Mi?�~n��|{D¿��q1���CU�IZȾ�BN�9�H�ٙ�N�_;m�7|y�:�V�N{�~���\#��܁G�X�&�B�e�K���"��E��$��L��`�w3n\��m,�c;J����J�.���;H�?v<�v1ԏ�'MҐ�_l^g�I���ݖ�� �c_7W������.J}p�����:��C�&/���9��� �iQ�,p߅9-?.R{�g�����8�"�Y1��@�m�bn�yp:��ȇ>`:�G�0S	���!��i�
�_��G�e� ��E�sՔ��y�"��ؚݒJ!���p��@���f7�uf��@{q��	? ���A�DIq���i�{N`آx�bk��YX?h�16�uA6�G�a�4�=[T�:x�t|$>]tj����1��s�P��+�b��%ڿ���oΨRf�Y	����?�B@�r��t��
X�O=uj�g0Y@�c049��x����� {a oM���J��zn\���9쾀���Mti�-;i�f�͔(NLp.�A�z�KX�(P'W��h�"�y,�==�o�,�M֗�A[�
H�X|m��A�i,�F�YQ)�I�� �=e͐������.d�7t�~/��p�In���o"*�c|$R�,��;kZ��9�WH^��H-�~JUL�6�׈�V"�p�ppI	_j�n�˜�U��6?pFQja\�9Rӿk y�5�u������o	q����������>T?�]*�K%'��|���X�ZԖYO�D�M���}�k=��t��2�L��!�TP�Y���:!�'�_~u"����􆸜�-HO6��-W0؂���`�?�O���Ȗ/�K�I/�۶�u�<�s��a?�~�)'���=�%]'��ٟ|�v�.΃p�N�[0��ƞH'Oݖ6�m_�ٍ����,!�Ɋ �:u�tk��ri�j�M��y-!B`X������
�+6��N��)i=uV��Z	z�K��w<��ܫ��(�|,Q��&�\��>u$��O��|����r�t�G��iH�H��tP\9&1"�V�7��Z^X�����n5��rc����A���	{��4z�e�y}���n�y*�g}�;V
LeF*���x���J�ޒ�v�{/�nm�8=��*�6m�EW��\�'B��9�o��;�	���B�7�������@�1��"�+�f�
�աk������'8�r/���L���$T��2�g��i�w>��
�Q`��'n�6J�&=�P>�颩*�.hNj��ZY9��N�~�
��[}Э�\%��#9N
��C��_{.4ĚX�cmv 2	bZ�`h0���,8|�U'J|͍��Cқ���/FQghA��4ɴH�&���U��f檡�
�`N�>�I���J+����UuGh���'����jc9x8o�