`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`protect data_block
LAUX/Sui9+QS3F3FSQaAzCVewINs2bIw1Tr6ADH6YRgCzecbIqccA1gM1B3JYZylUfEHDijzagl8
BAziTNiMAnSoXzWvwT5ijdy7nHkPk4L5Hue0sE8I2Q6RVS6Rs8IirVeifyVkoR5KZewqKetEjoSQ
vw6Bxtfv8KULZd/v7+Xb4a2QpNd5j6HBoi7U6QXUCEf0KLoK9l1+1FqJ4o91FVP/ohAwZc7G1u/s
LBZoV2ekwjhdhZ2SAG5830hsJkuttLrd5bNDxtjsa86JBXGz8kHVVCLSvVT04AUQmHVYebkCVB2B
v9S9OyZihnNncdETBheysskJIB9KbAhjaj1EVLF6yzB0MuyQp+f37W9Yv/MLX+293chFzcZMRb/L
gZYFvmQGQQmdOUb4r9ECt1P5S1bysfwhatjTZJfhQ47jAc/PDuupjw2u+6d4sv6uagL+UcOwuha1
HWTezf0PitrlqSFZUfA+F1fpD8oVGRMB4BHJXVRynj7ti4kOuV0g9/fZEh/yRdKiAXRdlkOePxCL
bbpoGGkpHCU0+P0Y/dggeC+lRyNxfAkVePNsHEqcsGUlg6iVbFzG6A9kcpUQeVcqvFnSD/yeapIY
acTZdu9bjA68wLKB2lGUjF2WZSRdB50BRJRbmXFuuw0nb1BpmA/u3zFDq7XyyQ56UyfSrwTcXIF/
SsET7D8ELHWHDTTNHuoNqGhWL8QQerSnRvCQOsMUaUOZc4YO2dsew+kZPWCpbLjsODc7ItFq46AO
3MpVAUJiJZSR1EXvcHSPQsAisc6hY8r6hYrYtP+TacZ7yZXTE4XKJijKBGI7h2fVuee7g59djzSJ
ZBMTOvghbpsXZCTr53a7YYJlMLQVt3DsHYmG9afPkeJr6J+VBN3BVocWEpc1j1+1izPbhiPsQX2w
jKco2smQf81GjGczS8vtL/TsRC0OG2SmwlHKuZOY7I+P1PCrTv82tX7Qri9knU7j07ofdYRD0hbe
ScbVL6d4BeW2ZQCOqhaJzUru2o8gFIohBxcu3EYquvdB0xXC+FwrI2k0KRC54lKVrWxbkWMyUQS4
xSBsVwoSHV7h5Bi6nWFoCCEFDJeVtiKtyBqyR3lj9HZWgYA3X0n1Fc8qQspGbq52Drhkhan41dQ+
N6zsSec37wJc8LzmQYl/6LTN/XHlonvhYG0u1zomXW8GVDnZdgc7LgpzKYg+aEJz+iSzckJ3I+hi
NA6qXoeK6Bk2zsIASTSeD7Gj/NXvFq8GxM2zxzqVTHec48SdwsnyXsKalTipqt2PQXEyjWMpYpxQ
jzaxaBrJDi69nNxmYHXM2MWmneXexkXW4D+H4TfdpiPMz/Z0sZI0k44C+WNPYunxmFeL5EVYzRZv
YCo9fJBAt9Ta7Q+siM8TAulX1LWspndy9fMbo+As1xtz8imtTBLoaKMuczK2x7t4SQ2mSN9XH0To
PQTEODWCLyC8PYkKoIl4Q0wb+myUwVxKvCemWOhTHu/uUh2DazzRKySx6uKQB5TBT1GLxneRkrBy
L/XbEh8slUVct10MIlL/C+EmeuUnpVcnfcZwtfkMe1z5LsyCP5y7ph0JdeJRR2xJgZzW2RCmW81Q
+QrhrniWVQMRJfwiIuuh+0/72oukes0CuaCaBjFHLrHWSKJ0nRlhKzIFrADouIIzsESr/AWPFGic
99zjNXJcVnDHq+VZ5GUHW5VcpG8XeiSxV8zltjS6Ttas6Ni/gequ+CROoESlRSPfSZLQw9Nxcqa0
DnJBNAUcVMkgGw/xmyzTAJLDJtFdygl01nfpaaPrwu/ghetD39pwjCDZ5sUF9qhaZjFaBBjJUN7M
p7qO3l8VgdO8j45v7k5B72CialX11AVKiQ4l2gMpOv8Uj2KEM1+rf46+FKlHi7ge/Y2T+oR8W8FV
ltwqEh92O+7iJgjsVER7HvhWS6vXbcsts8fFMeBgNDQT+rrI2s22PBnVZdH5xwrEAIQMXigeFNZp
yvxH0seql1j9F1agFBeVp56p0693nFOAO9xm2+U+snOwaAqYXw4MM35sEPynwVVcSmrmDuyaS0Yt
aBnS6iszlfU7sCCahYVdayaSYI+rT3XlzaxP2qRqqZAhicBSG97mVQeUeln9TAJED8sn3mf3C/sT
9kChqFKNfPs1zSEcMA+JkrK/DjcIOsd8bm/o6klO30MFDp42SyZdp0djI/BjVu/h30s9LgUFU6Q1
G306YI1Q3UH8xpHKwLcsz4z2utuEoTH9gW1Zq1cWoCeEri4hmaYH7PPOQmAAUwVNcVeYtqN7IPkg
VoUsm/2udXLm7Z2x9S467iqqEp/YYYlvzzzJKjHzrbK0VXw39r6x8piYbpW7D/ilJsrhNgMbfQJG
P4iRkfvfmtwpWbe0dWmC6uy0hK/jFkJGm7vGOJaBGtBqENA4kvE4uDmU4DErsbX8nuhMnwVFPNIt
Y82zH3rlUgIw1L2MyVTdcRHdBJx6qvegTJCJGBYshHIKEnh8JdnW2SoAoorFGdR7SbfKOuV8d2ED
1QZcx49AVLvguOcyI3j5sGyB05H/966QCuEXx5iI1I/VwNaFVqsMczGzgw40CL6vWP+FyBmtbHpq
0DWoB2x5TvkDcdGsHO6B2Rn8/aKGheWQYLFl34b44DbXA0ArbxAXadlHOcid3ZkV8Bakkq9KubAr
RgJbmUeOeHKz4j9s1Ogu5k9YmJf/6XVMAXGSI5AKoKpSS3Bi3swj7m0cYmWvmzVP8r+uTuP2jZd0
GOADDfNoEDl5wTaJfsAUeIXAPbmiMdQaWj9yvkGfxAJRm0UVJoqrdmPoNcvEdxDKHZHzB039zY2u
+HMTqNXMZnSj1xNRVMQssvGVFxoCBltNgeXYyu4Jc0Kl2qY1QiGYrSMCdGAXHc4qxaR4
`protect end_protected
