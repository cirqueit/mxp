XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8bφ��k�L��peRb<$�Q�.[�&=�L��sAl&�^8�"�u4��:��J�2�s���n��W�Z�5/�w��M!$/�ˁ�b&	W���J�,�V��*QO��b�R-��uįE�*8MhHˣ��P�r��ιu]���b�O������>�P?�����2e��Dp&(9�K?�ʧ���SrK7cw�<M^�?Շ��ָ∍���;R[��S�����y���L}۝�VV���6��Jb""}t�;q;���H����[|��������A<��r[������������?a-"�)Z�)��َ�@w,]91�����������`�xVy�c~�a�{'HY�za����e𬳔�}�?�<k����PV���Q��5zhw�=[� ̭��5(�2�O6u���⫏]�;�W�U�*���X����j�TY�j4U\�\NTRo���q����<���-�gg7(�%iSs+���Xh��]�7�=�.m�8q�QL�޽|q������*v��g���;{juh��Pϝ�Gw[����,�%�|���|�i�,6�TB+8��F'��-��n6as��˭V|�:F�.YƛU�(�!���>N���m�}��}7rtQa�#�VL��&�:]�#�b�2��[��1�~v}'D]��(���id��Oƪ�,w*�0�jA}S��U��Ѡٗ
��A���Ę�_0l�K�$9�\Bc���4
(���[l/�����溡�"�j������4!��g�xr�+XlxVHYEB     400     150�p5�r6ݚ��M��n��ہj�"o��~,�=�_j��fة��k���ܭ#��D�!�,������0��e��^p�,��"qsd|+�i��1���dK(�Ë�N�=T=@�myn^�o�׌��ΐ�q`Tm�3 U=j��)X��4a'0aj��>L��SU@�y��rJ�
��N::�"�nӳ�3�a](gb�ɢ��$���%�H��g��ײ�]k��.!U��>��3 ��M�Jz�:����DP�P�O?Ö�<D�����V��^%2m���n���9�r�ܔ�}��a��H�'c\�>���,���H���YҐ6�XlxVHYEB     400     170b3Έ��`���Z�e"����Rk�FlM=s�xM5�j?�5Z�C�� ;?�C�B�S���2���j��x��p=r�>��r��Y�1����nT��4tC����Ü��g���ز)`���Vٖ���ئu 2Z�2p�'3G�Ql!��1��jMk,1�Qm�N�q���N��M�h�?�\�ɒ��7�*5xT|.޻hU��\c��)���S��e�?&�#� �kz�vI�,�����S;���kdy}]V����xS7&ɯv5[���b��b��Ŀ�_�;����rM����E� ��G���*�a�ө��U)����D��v]�퓺ZL
<�yy8��@6jY�6�>��äS�XlxVHYEB     400     130ZG�a�T��*��>N��A�/�� Ă��+���� �jx�6N���69Yu�KB�����}�G���|lT7V+, �>��K���#KL\IB"'�ov��{�uHf.d�r�E� <Н��"��hJ�o��Ͱ6I5zSޘ>���<�ߵ�/�qrWd�P�,�KOWi��?Y�����Q�ˀn%�&��*�6ڒ�z�d�Ń���A��<*�-dD�#���#�bu�M��&e����]��s&Y[�"�~�t�_�=t# aݭ",��e~��з}Z��󐊮%)��-��b��@�+���N7*nXlxVHYEB     400     100?�V/�g؝�ų�Ѝ�<��0��*��A��,V��>��x�����g��Ḹ��r�[r���se��e�d� �N�r��@+�I����9���C���G�!'�@����6a�% �M�������<М���}�UA�%y��L)Xj~EQ��B�W�v�*Cf�V�(G�@<�.��HWl��.;L_���K�6�iHM&�e��B� �(��.�G������O���f �J�H�K��3�7Y�k �zXlxVHYEB     400      e0�}��ـ�Gݜv��skC���0�������5�>�KW����W�^��Y!e��1/u�4,e	�:
�)����:*2�4Ila�oR|ߠ��Dۧ�.��p��hb֙���)Ű�}���8GL�)��,W��rA�-���ylar0Am-"x#!�O�C/1z*'�Z��A7�߄� 亅A��,n&�N���>�g������Z��l����Gc=�xU}��E'XlxVHYEB     400      d0L#,x�����A k��2'PyQv/pz_��%[cB�}S
�8`��(��zGT��$Ѧ%X,�؜�5��Gz�>wu��zv��n�Y�6�uh �l��T�(��ǍwnP����h$z����`��Q�K-����UU��ve��_9���v�b5�N�/�,=��Z��R4S.�����(F	f��j�+k�?����Ñ�IŤ+��-�]�i l��XlxVHYEB     400     120��=�р�t��t�ݓV�gaܤ�v�(;�KQ'Uvz�����Ϝ=p�De�zZ/S圛������s�J�v�R�Qń� �	�98I�b" ��Lַ:�]����"q�}�B���U���w5N�a��²ƿޅ&�r����Y���ѝ*�!��k� SsVQ��~�)��&F
�z���ީ�)-�,K�g�n@�h����}�Q���,�oi�
d���R�����>k�2rʵaˀ���d|���waM�|��t�鐐�RK�\�g0w���;��	�����|��9XlxVHYEB     400     180&(���;O�Ǌ��ÐkU�I�^!R�&J{*eYI��O���p6�����,w ��
�&��x��l�]�t�w;K�%�d�'�,jo��H鍅�֛�K(����em�vI�|?��`(+�ɮd)����?d�q��>�>�_�no��*��jw%�a�l��SBj-k {R��9>�c��$�&{5f��w���r;H�,$�Q%�~�Nx���8�
���Y	p4'FO�Ig&l:��B�}q;m�o��⸘ϐ�?X��B�u2�Ϭ���JD�4(���9�����]�'1x�������o��,KS��E��]�}m�5}��t.�Đ͠DU���"�j]!z5�
ˆu�қ��H�eFA.b��/��o�pT}��o��XlxVHYEB     400     140@���Ur�R2P���$�Q�V{��)bP�"xs� "�Eܙ8��A�D6r ޘ�kӵY�l���N�����Fls/��x��p8�°P[~��Da�We����c�s_�;^��}�2��'�"8L�70v\k���
^��둳��s2X�A�
�L���2�����D4y')��&�QN��~��h��k���Uk<x[��A3o� AU��k�l��Z$���y���,i��D/Qn2˯�GK�1������|�v��08�*a�yu0����P���#Ť<�W';M�st��ܩ\n/ßpv��7n.��(�ڵ1��~(����c��XlxVHYEB     400     170WYH($B���P��,�5u�);2to�Y��/:���LKx���4q��%m�4=F��mi��N���� �.��岩:2%�笊2�w�S7�g�Y-��6}7�U�0}A4����\���`c)U��J0<���$���Vd�M��w=�A*h	��Z($޻��F)K���x������T�h���d_�Y
X�M�&:d������o��<��Ȓ4����=��9`�4}YJ���P�G�����f�D�g�����~�1<�+�C�)8ގ㯄ެ�ժ����ɑ,�����s�}��y�(v���z���8tG̹�oʶV:���R���|p�R	����(_��ꋀ�j�����KXlxVHYEB     170      d0}���#ݻ�l�����H5� qW*�{m�}�n�����q����F��8�kև'��T5��w�c2
>Ӆkjc�F����� ��;u��-�}����M���Tq8�:D�ѣ�]y_�C;HyVH$I������A�,& ��2�j���������*|	{u�S!aZ��.z�B�y��B��6|������+�S�4�m�u