XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��M.xl������bF��Ϲ"~���y/��Y?m�UA5�Zu~�F�6�R[�Ea�2���`�W1td �(��<T��#>1�Z��2T�?���!b�ѫ�	�|��J*�x�c�0q�������l�B�<0o�#5��~*�zYS,�i���kǻ�T���s��WP]�)��ݤ�d�����^Y-<�4���Ҫe�3U� L��be]�������aHȮ:�I�mo��C�8��X3$�]X�2(޸�_�]�Dw�0��������!�3�KնD���g˄���f��H��X�s(�%�����@�K��o�	��Q�Xoй�ܨ��i��P��:�.�>+m�I���lε�� U��/�*��X��lSP夀��'1�#d�Q��8����	^���m�2�N4�t�I�i�c2El,���KD��&	�IH�v �)��;k]q����9b�@��˻���&��&+ԅ�yu����9�TM�zc��%4R�`����Sz�������v�����m,�� -.Sm>�0}�(��_��W�sw��[�����{?��ew��5D7=aXm{�uSU����E�� �|{Wي�k��gGw�]ƙK���Q������[ذ��&��lGq/F�C	A�1�N�I�2r70_1u���-���h�8u��1S����<b3�t�
fD�<>-���/lW^?�s
��:*��&E��U�;iiȦO"��>���%~ǳJ�N���h��d`�N�hUr�g��@O��Ak~�:�XlxVHYEB     400     220A/~��- <�yѦ0V��w>
n���7������a�d����Δ<(7���뵰J?@��J�$��~j7����ǯlޣ.U�y�9�J�4g�+�{�Q��?�)X4�ш�}�d��Rڵv�쭦O��;8E}��~V�inm���+'��DI'�^�5m�H]$sF{���1��ܱ;f>l҅؉a�el�N���H�dl'���6L��V[1f���F
a�eGv����s.�
.���c�6������!&<,��|�E'�֙�Y ��P,�Q,�` ������jG`�W< �P��o41����5�9�6������i.��;��F���@�X�#��$����e�fqbM���t�3��C�'�Y�DG�����KB�j#����CIƱo���?���E\���d]
3���Z�~o��Pk�YY����z��S| �7��A�$�_=��n����s����X�P[uMN-�����f�S|zp��DLi��W9�^:� ^��*�R�%����:��t2y���q�}:XlxVHYEB     400     220�[N;-���Sb"3�M3 �%mnҚ�l����e�W��sr0��E2F"G�gy�g��Do�T��6�@��y���z��O�*h�v<P��K�p(@�{rS^B����({��7���K|��[�
��3�8p����o�Q\#O����H2"�� �{\��b�P��S��`b�:�;�� �S��S�1�"�ת-?@���5V��jKf�f�@c� Q|-R7���r�W����Alˡ���R�x$x)��(��j�v"�j����A/#
Q�u���Y�S�oOU�z�O��ռ-���xh�p�H9�,_Z�b���9��S�c��4��Ϧa��=��f�;?i��p�:$Ӈ�lov�[b�l��ϰ���4�}�	��i��|#�l ��d'�,�B�,��ݱ��tK_fA�N'U(��t��9�԰��=C��ʐ��U�����6�I/[r�6?T��T�?A lAQ��w�@����&�߲��k�~A�s�{b����͇rހ�Q?&�q2n�}�-wJȫ%���G����j'XlxVHYEB     400     1a0��O�}�=�c?SHEu���4�(E2�D��?F��2�=gp����b���j��h�x C�*r]�b��Y�3t(�j9d%��g��K� �u�Ԑ��	�v�kw�*+V�T�ó!_�А�y�ˮr(&���v�������9�yy.�:�c��!%&�WV{lhO��xiS���s�X�JS>N��� T�p8.p���cN�#@;wI'��� ���r�Tg!�M�B��Z���I$H�ޢ"�w?���z�S#�8͝���.���f�Xfy�2�{�]���	�YLF�0K�7g��y�Ms��4�1�%7�[��a�߽*s,YB���'(#��&�"�X/8�>laK~ڂtN3ܤ'����IS��ע��fy��"[(ˆR�׺�7~����1�ԭ�٤�D�Jw��XlxVHYEB     400     130�2���t�6>�t��3��k�~x��	I�L���\}ķ���o�b��>��
8��k�*�`�k�w�+R��&=��S̍�[]Qe3�����o@NA;ջ=q����X��_�� ������>���ڇ���{��\ߵe������[䊛s6n&�*I�)p�R� �y[ޢM�q��
�fr/ ��ӄ���W�q`��C��K��K�����O�"^bLe�>+^��\��o���ӎ�4�i�����H�)�ݬ��H��ЩR�G'8�r�\��%Huy�V���w�-��h�Y��x|�d�±�XlxVHYEB     400     140�?�_\�&������@�3�6�4Q�����=�kr�P��m�����I��7S�_��U_��V};1%�3^�/r��AǢ6���I��R�����
��|Î�)��ޕ�;Zg���g��ۆ�����R(H"����E)`c=��
9���}�ee@��L�o�2���{����B�
e�D��x����h?*����aYI�G������ؿD�c{�n�����u�kx�n�3pb�=E��a��E�����V�r���w/R��O��h�o�Eq"��~f�
%o�j���C��|"g��3�?K�_h�`(�zU^��+�XlxVHYEB     400     1c0K��30�#�еO��ɡ-��W��a�-s�b��bb�T1U.�ڰ��jkO3R�zd�R������P�(��L\$�=F�X$�Z
��=h���Nk������I�DG�!l�P[ e �􋳬���G�I�(y��z���ߊ�p�kgx[��U�+��~H*��.�&�x��I��s硢�k��V�W���Q�_LTWH�Z�*]R�J�?�}�dme6{������%��P�C���|+����3!���9:��x�2�^�p��;���<��ƶ�7�_�S�-�YZ���9'�g����L L�bi� ���<�B}Ga)o$;ä��>D_���o���X���R�=�s�|�"��?fd�(X�\��0�k1����':���}L��TSj�8'����B�����Z������
�'�{l#h�pQ�D�>�kxP�9�<�XlxVHYEB     400     200�e0^4c��ԚM��9"�mrT��� A�W�Dl ;?�! I4
@e��j�����(_��a��N��Cm^�rCK��Hp�>�%r*���X���A���^���}���*���$�J��&)�O�|�4f��Ђ�(�O�+���ʒ
IQ�xPl��q�gq��+�;|t,�
uv1��?N	��]��3 ��1���3怜ˉ�bM-j6ޓ�`��`n��OѫSg���ύ��0c-����&�������(y�;�:vNT�X�X�}+�9R���s�����*��5O�M�a����ڨ�b���Y��:����,��z:�>e�r�YvU��E����m ����N˚��Hd��?7!h\hdb�y�<��s������[Z�k (������Xx�Kd��xk�	;�U���͸.S*�gB\
�Z�ҥ1\���,S��rT��ߧ�?�RN����A�(�pb�/�6^,Y��y�/��^&�pw?qsH�r�P7Q���R�8��/�XlxVHYEB     400     1f0��u���I10%5�&��[6z�����������V�O�	k2��f���`#�Rt�n"�Q:c��i��ӆK��m6�I�w]QV<�/*{�%M��P_���$r_cd�~�T=�b?�}�Ȫ�V�E�%��y�ئ��a��#�s�W�
W�h���R׉���l�F?O�}�[��-��#�_�]lLKU�Phn���/�g��, ?�΍���_@��������.�*:N�ū�T;�g�ئ��]d��_hsZ���H.�Q�pw�E@��?�����j���$t[<��?�mA��`�؎c��x�@x{1FϬ�m5��Å6�.?_P���ObY8�$y/0b�fBu�yR�s�Xv��1�Ǡr�Q��'���U޼A�H����b�g�O�}��y���^��Ӓ��ZwEbp�����F�	Dr�	��H \��}�"�8�~���5��<������"K~��!ϐ� u�y`!�'<=�������+XlxVHYEB     400     1e0�����/��FQC�J|�ˊ�@���I,￺�s�{ƌU�0	Q#Y�� �����u��2R{��v����)W��w����GmN���g7h�8�Va���b�=SE&q��5.��!�g��F���9]��l�C����d�FVv�ߋ�\�ѝ-����.%��W�o!��ݵ�,��P'e>O�4K��h�{�o-�=��dm:�R�C��C->��Lm�0���y�W�f������?q%BjS4�jUG�_�B�Zg��읗�͉L�bK��]��Q�?]5�}�M��
N󚧾h�doNFk�X�wO�V=CӰ�����u���TV���H֗IJ0�{ŝp7�a���c ��	��B��IL�-�Z�I��H��ԃ�L���'Zp!��#I��)��{�oV�`�����p�3wn����ӋԊ����P1�=c�.no�Wu|<���DsQH2�%4�	P��5�O�1�|ц��p�XlxVHYEB     400     1c0�;�*�8�����+Ɍ�ܬ�Xʿ�8:��S)T�gW��������g6Į)�6��K�B�$��x(-ƭ��_�(�=���u�Ͽ:Xa;��S)�VI���=ݗ�k�C8|m`D�;$>,U \?�#�ǒ�\�^����ƺ��?j�	���nW(nASa$���t(kP��(5BT�c��?��V
g@H����T~|d��w����4S��%��b��mV���3o��<U�Q@\�K «�Q4����s�ԑ[�2��,�ЦwzZ8<dy��O�/3�B;'e���u�Z@�����^�)P ����&��41��!��g��#^##tJ-��.��\���X*�E��a��N?�v���h��>Zb:o��=O���+�����)��c,��o,��Z�u��$�r�ɾ�<i�y鰔ߢ�Ey8�`��jN�2��e"�.[\"��/�.XlxVHYEB     400     130H�˽�9�{���*�U�I�e�z���Y�"M��5��Α�7����,2nm��g�սn@�&�ct��j�WR����t��J��>�n+jF�2�p3���Ǩ���b����f���p����.��>&�I�2�H�Υ�\1��a�/�Da�(3C�
����k���L��A#���O� �T��[�pN[m�YE}��R+m&a���8S��5S�#�HU]<(�S�����jB%`k~$V�?���hk�\��+(o�1��ZѨ�Բ��x��!�ݮaS �e�{�����1e�e��<]S��6�W�ę.2�XlxVHYEB     400     170Y��?����}�B�Jh���uO.tj�Q�E���aݠe-����W�$��������I�w+M�|�W-����39J���QQ�&,��b���<���Lc���D(6�����e�UY��3&���{�j�!L^��*�	�0�����g��HHgY7��d=�ˮhn^D����N
���������I��s��䒟�l�M�p`T�.Z&
攧>�QJ�#�`hZ�+�E�TCHjfXr�2<�s�ZRŘS�+6���K�E�O�*	 ��Q�oRe�3|��I�C={�gĦ�PHhΤ�<믑2t��Rg:��Nw{���EuW�B�W#-K&�g�o�SN[ol�=�)��j�J�h!'/t����XlxVHYEB     400     1105�6j���ՒA_	�L�0< &p
�=X�^��f��v".�Uo�=����Z��r���i]����ᦑ鋣"�2Fw\m
�N�����
����?}��W���.�O�*�_�Aˍ��@Ol�Ta-�_���-�
ȶW<z=J�t�W�1%�욊IC�,�E�`�D�)'�ʧ9JO<>7���E�'�Xw�c��U�����砡���!F!��%xG�V5W����bȦ��K�~�~oY��D�PX#g�Ͻr	Vp�PK1XlxVHYEB     400     140s��S&Ѿ6V�\��R�S���J�ތ�>+�3�]f�p+u�氯_Q̝���L������x%Mp��n��-7vo��i���v홲��r��FR��%�hIvG!�`�0��7�*�~)oV�$^��+Ё^��tl�1'K�y|c�&�����OҢķ=��ӈ�V��>xts?�%
�B[@�|������a���qy���[�=���C�4�CQ�֦�y#1=�u����<������H�L��-i0�Їr�#x��r-ƷR���s�
�է�Y�#�&�� jց	W��I��܇i���������3�"��Ȓ�3�XlxVHYEB     400     130R���a���u�T�3,a1��ψ�MϪرYzC?�&�x�Oq�%���4�<�n��=�K��v*o��Έ֥��̗�9{�cV���ˬ��-M��H���\���9�и��b>$Nq~�Ъ����S���'}6{}���ʌ��֕�tl�TjL^\�?���g��i8�)Y���O�
�F���%E���ʀ����
�<���³��W_Ц����'i���]�L���hci�]��x���c��e���|`���e]T�Y�x�ˉ$��s��C+�� Ҟ(�	ս�c�K�蹬+G��'N�_�XlxVHYEB     400     130�&5��^�吲�NL�y9��.�H]빵e�jv�ކw��ς�h5�@��8�CA�h�Aa�ç~p�����au} ���E�0-S|3���Pd��px��@L�G�+]�:I�|�z�6#
h���aT��ޡT��߿�!�Ҁ�qv��:�T3 �S� V�޵��ո�'KY�Q���V��N�d6�/n�o��G4��c&�U�*�Mɸ�����}��}];nԡd��-���?Q�Ӝ�|�&웞�T}��b٪�{����>XIn�dH���~?d��{xt�2���xO!�O�,s��P��B����XlxVHYEB     400     150���7�i8*B�<����p�F�a��b���=��8��d�Чk�P���(�V���+nF�_WD��c@�f�ue�a�:x'j)�g�w=���2r��*�nҕU�$=b<��P�
��:��=ҫ��ls�6���K�h��[2���7�i:��d��KZ�9myկz��ǬI}�. *X� [��Q�0"����/~���y�����p��6��J�V�H� �0�������Zg
`�0%�U��C�\�	h�^~���9>�����֟��[�>������.T-}�ՌIlS�}����\͏���Ρ�NB�MasؼE���GXlxVHYEB     400     180����(�H�CR���MM�H:�]i�Y*�f�u��Ç�S�N�������X��t�>�3EQ�g��䏘�#�/qG�7��-��Z�D���z V���l�#�d) ��%ѣ��75�8�_(���
Jx����4��ׂR3U��7�~�^L�O!/��[��1��
�}�Z8�-�mt�W�T�w̳Sg=�9.�#G)]�_�lE���'���
������:��	�#�/�+�oV�0B���R	��i�ih3����&g�1e��<�8"9������(���x�� KF��˙3���c��b(�pa���]�X��K�kW��S|u��F\����@� �:�e��[�x���R�k������n��D�T��XlxVHYEB     400     1d0'�e���Q�e�k#�2��Y#[Q�K�=��Gȿ�"�m��I�v3AxC�����5t;@#Rl�D����R���
S��EA4���;ȋ}9��0!��/<7ш�1�s`��I�"� vM=��E�M-�� ���s�pg|Q{�?o�Q؈�a����V����-�D</t�W���hǲ��o%ă��YR]m]�E�D�U��&z����y#��\����cn��5Om�;mt+|'��$���{jʷ=�/�	���M��Ju��w���޳�� G]���8��:�&��V ��~�{ʷ�i���|lUJm����&�[ ߶���h��!�h		c2�?��M����J#xf�Ȇ/R�D�iR����Dn܄	�I]�t0�~Nvn��ןKXС/���/�kմI���p�;�����%��*'�yH�d8�Ed��)h�O�u�ⴓ�K�+��������XlxVHYEB     400     180Un�NȆ_\��2��'j:b�IȜ�P�wj�
�5�XG���x�Q�f?d��x2��N��D�$Rc�0��,���٠�`�ɀ~�ά?o�j�&����=wx������sD�r܄�nq�G~�@B<@�G��ˋ ܰ�A9�_�F���e��2:Cj}�j�E���w0�7|��*O�K�e=����Ĕ�A�������]����1�*M0듌0�}O쎗D��=#�;��X��8d`JL7�|o1���U/��s��"2/N�[�T��.=�/�$of92X��{XԘœ3���6B�|��w|�='�����6sj�~q�Nc5}��|���G��tz7��Z������f9���0/K" 9��y$ӹ?��D��� ,�SB�XlxVHYEB     400     150�ǰ)-�)y����U~�^�4a�<�('c|�?�D�H©��\����j�<KO�y�=��֒-@��޲w!����N�|rF�_�޵��I
PH%�KbJ��R�@��u����R�a����/1��	�:ͣ�n�3O+�j �v���W��$�#��S�a�
�܁õ�G��v�j�j�">9g٤��}�uEk�
������'�V��F=���`>����R�Y��W#�	('�� ���2#�O�'�Cp/v��5�0�0
�C�F�(�^�2$-N͋�<m�w�/N�E�!_~�Ԟ���o��7g�&Á��O�?TJuQ�wyh�t��3�XlxVHYEB     400     1f02�&���$��5s��no�i�����jZ���vd*����w�A��#JEk�&�R�k�(.���f�I����1�i���7�s�s�������/���1r�N�G.;���}�����S�|�szh�p��9�~QX3,�Z�(^)�?s������~�O�R��>PtkmF��v��N�w���#8�J��.���������t�O6��ˎ�㺬b��N.�FmP��^V�bC�K��Z@AL�,�����G�N$3h��9��ɟ��,'N5����-��G.���{wĀ2��c���*:��9���5&BیҒ��b��aWNN}/���@з|���u�3s^��g�����|�����Z|�(U�`����k���R���ڶ7t��ei}�������)Y������͓��(��=�<.#��A�B���rq\�E�Bzӝ/e�v.��ol/�}�2�o�J����k�~�s�S[�`�'�����)р�#1��XlxVHYEB     400     190�W�v|�}�,�#�\B���*��>�7���p�=oj�T���u}8C�/z��E;�B�'�%��P�N�d�CW�|E��`�p�
.����**���R�]�.�����d����=��-0���抮�A}��T{\#|/���8\�k4�m��Z�����z&V�RDIn��(�ο󴣬��j���~�a���?�XBl���7�n�m���1�,S�CFK�`4<9����v\��A�t�}�换�p#O8���AL�v��E�Hm��J���L㽄�T�Ȥ#��o��,ќ�ޫ=�zZ��YH0Kd�i�l%#Fį=7p�wd��'Fmԕ���IJ�%Q�Z��p���� ��n��*_!�/�h�.�l���:�W3��8�9�Mj1m��/l�@���w�XlxVHYEB     400     170o�ȼ�~vL���#�q����h�'�d!w��q����V�����:�^���J��f���<�mni�~��fU�T+�^T��y��`�xP��l���yYD<����g5U��zH���������?���"��x;�ϕ�qᭅg��$��G�*ۮ@p��d�f��<�J2K��sn���2�t��c��C���kd�CؑM�i�mVp/�?q��| k���f��^sb4�_� ��מG뷙�t��<1��B��W]���zل�d�5c��GW�- ��iU2<�Ֆ�����>-fvp�>��lMT(<�)�4��B}��O��F����>�5��5���ݖ�(��ғ���5w���6��y�/��XlxVHYEB     400     170Z$��KU.���2tWq���Bm���[o�|�Č*#Ę���Xd?+@l���6��"�[G#�=M��RV�ЌE��I���@F'�@m��������.6��I�aEO�*ٕk�ͭ�	u��D�ߤ��$x>+��v�@�VqĬ�G
���~[��W[�&Ʊ�a�3�/���Kg�S˾�r�+����q�
��ksu�7b�#[�m�Bc;�T!;Sn0(��Vք~��EeӴ�xz@zB�=��r����P4i'����w�]5Ѩ��J����	!��es�c[O���L{������x`e�ٔ���)nT����6�@TV�;���T�E��+<%/1�iQ�a�|K,�&B�`/XlxVHYEB     400     110h,������������{�ׂ>i1�-	��p�p�O%��f���½;�\ar�|�Xl�$�aZjG�O?h)�6S��#��)p����9�-��o#7��bY��s�z�<�:�ğa!Ӑ
d5�,��Co�[%�~��B���^�S�{�,%ur;h����k���ŉ\��7@	w�O1n�ra1v
m��ss�&��|
7��C�G�ȱ�
�������y��0��	� ���="���A[�e ���;.4�id�w�v�q�3����XlxVHYEB     400     120 �ASXY����w��N:�L˃5���%B
;�������N0��)��?��v��u�U3��烕u'�Wq7��00>��oV��w%�[$��
�w��9��I�TfM�g�<��c,g��CU�qb������r3 RҜ=�ѫx?A�����,�㉊�����@Wt��ag?H+��s9JT/S��g�%����e�G�t�Í4������?�R��%A�x��0��KԱ�@�[Ÿ�O������<-ִ�r$$�c�h?[�J��BG��dI�ϙ��+�XlxVHYEB     400      d0��j�+���/����բOb���>�
��Df|�w��� x-D�B�n�����gje;�i�Pif�_���#��!LB���ߊ�_|P_�	�Q�Α�:(�;��#4���I�/�=���Eb�s�N��?(�J�!�1��qe����AȚЪ�q8j����#�_Xȿyt����O�fݸ�e�O�ڇ��0"��άǃu+�XlxVHYEB     400     1400ӡ��0D����R���6��e�k�������� ���!¼�Ğ��QA�&�8�Y�&����n���1�ӪX������a�0y���ho�K׬U��}�pTX>׺��&k�<���M`�ܯɮ�+ݲ���ש����Xs������bԽI�y$bf���w��7�֟T��_T=Ƞ3�E��x)aaZsj���x���{�aՍ>d �O~|�NH|xG<d �� p6ҷ�A��;��"Td��_�� ����'���?�g�!uX�(m��
���Ŕ�����3�1��S��S^�O1���g�I��a�PJF�0��~cXlxVHYEB     400     140�����جh �`�؎-��K@��bL�|��]��u������N..<W�/>���ݴ*=z���)�5:h�����d/���
� ˏ�tV��� ���)�wyg�{'L%j�S>nU�X�PE�PYB�ʚ�i= ��H9A�?�@?G[pOp\�9%���.<Dx?b���gҝ}��*���H$
Jl�.�QdӘ�pĔ��=1,�	��V�a���%h��,���Q��'�kw��ۉVl�F���h��(NA���k�x# EGkp�v�]����{(���5T�[���f��8{���d�1�$�J�XlxVHYEB     400     120���νc����r4P����B|9���Ad�I� �9�o��F�����-
t7�H}dk���ux4�qo<#�`y9z�2��q�*Ӓ3^�dH�������
�=2��n4:s%�N �u����}����l�Q�׶���N#e��QL�q�.��Xr:��S�1����P�+���T��E��䲹�|$�0P����*XP�Fy>1�ʵ�$��8z��Y�Uay�M�O�	����UD�<CD9�	���-rdB�Ti�5�e�����?	�v��-nXlxVHYEB     400     1a0~�%�����"�������{��pe��E�|�:/x��?��˕���W>���8#+�MA=��a��w��v����jW�ͤ��e�}����H���~�O�hyU��sTA�����N��$r��ޫ��Εr]*w=����`�8�ߘ�
n)����H���'���lp��e�3�q\����
ߟE	i%�����b����`����<���Bڔ't*k]�<9�L@�����e�I���������xl>Y�أ�p�.-�o?����b�����FQB�-*w[Q]�X����r-'�/��akz��`���:q��֓��t� KC�/D|J�`+Y��.�U��<"��s�裏��-Au�r���V5��ޟ�����Y<������U^Ӷ�P��1)ń�!f��u8���GQ2�<`XlxVHYEB     400     120�~��M�Ź��,����2]�R��%T�R��X�cnvcrI���c�5yZf!Pİ��@�G+m*+s��IoAa�����8������vz���o���<�i��T��=L���r��l�ؒ�V��l<������Z�9��a[��1���o��;����'��`�rR�|r!%�e��AΫU�1�r��������q����<wm�\�2�+-�7u�^Y�3q�Z���i8���֪C��D��s�FR�t�HN1 ��_��b�s}]-��ر�w��fE1Pŝ/��9�H�XlxVHYEB     400     180�tҔ�F���w�7����o�ƹ�@����Ĥ�'�F#�'����d{i���/�dl%�\�Aq�9�hoݣ�*���:�?{�L8�2�S��#~�O��Xw�d������7.�{�<�;���M[�.~�D��!�<���?r����x{N�p�>:�`@zA�c�a����D�N�^��thK�����O����x1��8.�����;��#�_#k����b���7�M2"&�%�d�`'K5��*��jU�)�� ^I��eb��^K�G�ю!j�R�{�K��s��ߋ
Yq]R��ʝ�q�-M����,�4(�a3E�} �.r�f=<9hf�'"ޤ��ֹ|��;�U�g�v�m'�j`��"����"N�����&I+�f�|��XlxVHYEB     400     170z���p���Q�ꫡ9�0�"�i�0T��!�!I���6��X�{^�W��B�_�|,^8{��]/�i�^�����)���ʳ`@�3��{�%�si�15����G�Z�[��|�0�����\�wuL8��Fy g�6�D�,��+U~"���R꼢�3�%��&1�uJ�;%e9��@���m���A6�m�{�8����/WmN�h��;�6v~�|��a�g��-�A��K$�i����[f��p��	��[�.^N��53bc�l_f��Cy���\���"���֔UN��3��3q^���{vSn���.6s0c��"�MH��Dt	�J�j���W�k�=L�����.�k^sl�#2����XlxVHYEB     400     1c0�:y
��q_�d8D���G|�)^���̪���������|�[���}e�#���o�늌�؇��;��&�~.��q�����0ic_w%�����t���+�FW5�ܸ��@�c�d|0=�MV�vq�c��ţ��ѹ�@��ѻl$I��� 8}�7�)Ԁ>�c�M4< ڽ�;S��>~�̼�s��~��̽{��]֥A�%�QU�'�Bx�D���Kg��1�����_N���OQpg�Ϊv�pF&�����ξ3�^n�Z��h��sTVh��CŨɾiXZW�_�2H:�L���-� �eѩu[h�n�����R�c�_MeY4���C��PJ����p�)ϰ)���u�H��O���~� ��<D��4�_#���A8�B���I�D���a؋ gRV,e4j�0Ća����/����a#��l�8*#�eXlxVHYEB     400     1109c����>*|�"��7�T�a�?$�'o?C"�z�_D�:H�U?���oY&[��{����W���G)�t?|����GX̛c����F�~-��"���46d�&3�붚n?�v{i��%3�8U�Ā=vv�IgSֲ;���$�e~4T_��#�>��_|E�$��e�(��E]� �[�)5&��&��xr���؟ʇ��Z�4�W���Ȓ��3�r�qDY)�-���.RR�7JѯF�9Հbt�6�/�����L����� L�RXlxVHYEB     400     170HW�����W�W&%ٸ8��Md��d���a�+������Ô�{W�f��^��8���D�8��u�U��P�YFO�e< ��)��#�ʌ���[0�2`��y�#��%hLk�"��Bh�E��4�f�H�%��^��/��hMcq���VaD�7`��Ô\c����G������(e�0��2��I���
�t>��Rѭą�t�ʻVY�����~?Ɵ�z�lki^���O|��X��*���TҊcٵ����H�|��-�Ȇ_ܲn(�7�r��^��!�X�f{�[7�d��V���A~�;z������CM=�uI�dt�O3�x�*������!Y�W�̾���\��;WR^Bop�C���XlxVHYEB     400     170��n��1���y����Ȼ��)z�yʌZ5)�~[���Je\��Sg���$$�%`�f��������C�Zdø�s�
)�.%x�d��� EO�y|c0�'�p���C�?����xlW�
U:�S�"�_obń�9?�^{����?�Tu3�<,�e�B����R@���=^�H�7O��A��p��>�#;�Ëq�n�$I�+
�%}}��b����r�x]��$_���$�";N'���P�]D7��Co�����uy�NV������hg���h�|��1��9G}��f7#a:p�BL���!�����I���
����_�"�SZ�V^ �����9e�+���H׵�=sj���C/;�˳f�R��XlxVHYEB     400     190�O���+�mC���"�B��תH�JAʗL(�
Q�X��//iG�_���Jj���=��1"��?l@�냤�������7:Yx�:��M���uz��+�X��g4�c�M��HAɅe�%�
���<��y�cG|�AM�AA�LN#V��=�ľ\�.���&K`���'m]Q'й�&�[����6.�����{ o��R��1��Y܎0�[��u2K�eF20#ӭJ#3�����~=g�$uU��q��M8�Ы��V� ^��e�Xa�J7:��%�:o�u>�0\�r�z���-J���"�W��L��y�W�'�v7�y���V^K�W��G�ڠQ�	O�b"�U��&��Q����,j�����jΣ�y44aj�ql�����Ō[�<��XlxVHYEB     400     1b0S���8w��q�E}>�����^������Dipږ����ֱ��37%Ԙ�kɉ��f�'��.��B�a����'�m8��TXY�L�ƅO�����X� ��j��E,
�$��^��胻�k�;\���ak�\����e7'�>-�E���P2�@�Z�
4WH��-p����K����.LC�)�z�g��$�1j�d�.;�|_A0avN|�8�M*	}l�]�<Ô�%��Z@3�_Tq��mcj޿C�@�K��tJ���8�(F@M~��m�%_��r,{���#�������P������Y�f���O��)+�'�����Y�;-dx��Hg�f��R"c�����w�+$�k�D��;��b�#ܳ$���}nX�@�r�}��m�L��n;qߡp����E����=�CC�BCZ\X���\t�XlxVHYEB     400     1b0�:�d���
T��xr8s#3c	
4Q+�)>gv� �BhE-��%��p���>���O�	����|�!Kfv+5�sR���\��D%�$9����L��W�)a,�d�>_B�-��N2��tor-���B��Dv����w�}W�d�����l���e����b�Q��}�-�=58�F�fW5T�F�l6,:l%&ՇIj�*��d;�_L��{+�W�50q�R�$�/��l]7o�]Q}Ogh�?�T����xM[.��_
���hi�����/����ڦ��QԲ��a�cÆ����ۗVu7B�����zDȁ����giΥ-�bvtObd���h��P�N��Y��	� �G7���8�x+"F�8�yS�����c �VL8��r�:�6M����$�}['^;����wJ�y�bΞ���`YXlxVHYEB     400     1c0������e�'C9�;���m�E���\v�&u�9A��ymbSCO?f�H��H�����w�$I�to��x
��`J��T����q�8����<�Ӗ�KrW@�����f�n�*�:���pY�tBj��U��>� �u�����2�ޥ�ۇ��(�J6՚��F�B���^nHMx���^�y����i�V�d�a�'�4��K̬��u�!� �Bt����8�z$NM�[�l����n�A^ƐG+`�r� g��Mx�@M�Nw�\r�S��J׸����mi�<\��h��9�T�׎��	��gT}6;"����-Ո�=��E��UJ7��E���G�e`�'�@��F�N�ln-;K� ꫭ+�iiL����=�����=1]�B�����Ec9���+�iؘ��F���ư7����:�C������f#j�N��Y�ADE۫<GXlxVHYEB     400     140��jz~hH�A� N}+�#�H���,b>q�A.��h�B��Ӳ�?�l��M\ �=ƃkm-ž4�-r�7��_��a�a�' �D�����뎂� ZW~G�2���"T/0�� �^�:"
����g�K/��o ��$��-�U��A8A�u�.��L�2#`ܓ�2�����ӛaIH�k�Ә��b��}��4>��)����7`�8�X��~Jj����d�����:�O����t��v�n���c�u4�k�G���Ԃ���ʊ�9"�S��C�g��q�=��=1)N�*xb�o|`;VI�j{DPi��Dq���XlxVHYEB     400     190��`Dj���uQ���l[�r��ͭ�I'1`������*p��r? �D7X�i�x����@0��10��߇���M
�|f��	��J>ԈێFp�g0�gLhˉd!�Tm�_xrΖ
PTh]�'}���0>F�H�jǆkO�`�&d�y ��h=������:����*�_��-�Ez��e���uT0�5����S��G}��� Hz�208��RZ0jFK��t&�rվ�27S�qQu�^O�"�ݒԀ���ow�s�j�)#<��FK�ls�A����(����VR�>o��.Ȯ؍�/-o1�5]�����+L;_��Y��������s(���u/*E?�`�P��Ⱥb�>ø���\�#â������WL-����$yd<>ʉLaXlxVHYEB     400     130ȱxhS2��6o�ߘ���&��u|d�
#Y�w��ӓH��^�Lc� D��ӌf�M�~��� ^Z��u�g��^�#e�ئc~��{��앰4���|ʛ����Ǔ���DOӉ�3�V~����4by�ј�6�"eUd�V�M��&�l��{y�`dhU�t�`�A]ԩ��/�����9&\]��A�KU�#���u_�(	�����^�d��W{E�lsY*f��:����P<���O�ۯfG�*������!``��ᕙX���Þ���\���8_Fv�9z�h��D��XlxVHYEB     400     150�������n�)�ѥ�V\��Ka܊Y����=7&N[N_PB;�J�����(�4�Џz΅���	��2J?�]6QoS���7�C�!�R��~�,I� *:H� �����\��
�A��1׹7��?/�͵��w'S)י}��v��W2\��:�������W�A�W7 �J��D�,f3"u!�i�eQm������}�2�lpb�]��6�&�E�G�7�UU��j\�v���{~AU償�4�LG�.XNÊ�`�33c�R0�=��Ԁ�����yo�d�jZ�A����`�֞b�^@�cN�L�*%:��OհS��XlxVHYEB     400     190c���襭\���/̠�=c���/���&WS#I�xa:���3�i�ߙ��t�B]����%�?�Fo)g��L�
ۇ��j-i����h������ma�Tu���vn��*�������j��ļb.�tw���bC��r�{Z�a�7<�lƴ��UT{o�ȟ⍖\ǂ��J H��ICV��!���QBj���Ds��󆜱i`��~0��e��%�#�*���1�Eu���@�l��D�M�C�/�3�h��K�z���Ț߲O����G�M h�ߵ�)>{�2� �c� ?����N�h+�\~�V'�W�*��������sK˦6Q�ޘV	���x�5$:惗-�H��s۾Z�xL{�R4P!�A����e�i�y��A�|$.��_�ܑ�XlxVHYEB     400     1303�V�Sٌ�>�i�35��N��;,���58�`��;"f�/h�GE�E�@��$s�Ar�:\���_d���Rӓ�9+N��l���B�����.v�F�[��Dp�
 ?r˖:�r�ߙ��H̗��$k
Uy�IoKU�GZ��./BkcӍ�2��F�9m�ZW�� [+`���8�_�y�1�mŀ���r��dp����/�4̎��)�n˔�i�$|ꪜ_LE�si����8��R\3�+���ow����c���/@ ��)�HhH?�+%p~��ڒV���cbi���RUr$��pEXlxVHYEB     400     150�˒}���guq�M�A�)� �ӱ<�bҳ�
@��J�	�S��u��t�WA�q�<'����Tͷ��Y����~���hy��"�BSCN�oĳJ��Uq�ò$.�w2R
��6���x$�V�������d����P
��*���w��7����؏ ]��g�����N�M�>Z7!N]��9�-.[�o'�k�d)}�y��{����劒��:FՇ�2��������
�ynv��^�ceϏ�%��v��z=�E�,�:��Z&��f�P]��Q돖���&����4l�LQ�\��R�r��mi�(PlE'�!�P���Q}��HO�2��XlxVHYEB     400     1b0��h&�/�2�`�L��xs���{L��$��y2!]p�'��xǃ�爌r�ht�g���B=�ۘ̏�5 i�+I�"'uq�#��ءC	N0�L��Pf��V��M��0��oR�w��b�F|�ۆq��;Q��D]ݽ8K��w�7�����K�
�b����7��2�s�CTe��\\3�{���p���7e��������R�ə���١m+&��h��Q5���m��]��3y���gL_���x�[ē���T]}UE(��BH/`�i�`��]}�A��s���nw�xY�@��?;-�lt��C�/�'\�:UOfa�v$uM�@�P�6iȔ+����Y
%������6
&���B?�%���]�p�Ȫ�иü�}���8F����_S�S<�#��<l��K�!ti� �����4�a���4};���XlxVHYEB     400     1b0��S�=$�/��N���T��������橠>�����,Ƃ���w0��;����2RiHm��Eۂ܈¦���+F�'2���p���ڛʿ$Wb<3�\N()��o�0�m��n�+�+�ec��(�w�Fȫ:�D�������>���Z�t鶊�?K>m�~WM�~(
ױ�ш��>5����'����Wk3��FHq���#uG�\h�ll��6<�C�ن�t���S���;7i�$���CP�^�il��^�^�J�4K�3�H��gW;���� D���V�[���{*�"O0�HDecfIϗ �;�KR̇��N��	eQ5Ī2T�m�%�\>MeO�Շ�xQ�H�HҖ0Ƅ��g�YG����56F-Q���;g��+�X�%�
C�#�Y��
���ˌL�'�XlxVHYEB     400     170�oY�DҐ�&�W��E�Dߘ2��ں�>����1h��c]���\��gGˠ���,q�����6P�\�Mav�m_ʉjs��;%���Y��ë����22o��i���Q�!�n5���CE�ݦpU�#@x�>+2���@W�xՖF>
���bW�M�B� ��L�%\�������͗p�1J�B��3Ndb0;�f��\,�:����`��Y,샔�ɪb+]U\jf	)@�]�v��Ƚ��� �/K���V��;�b����Ϡ,^���W�c{Tl����[h�Nr
�M4�BO�vR��͙U$�a�H�&��>��(>��.��k��+d��H,�Q��@�������6c��p��%лY<��J��XlxVHYEB     400     1f0� �<��5������,��8A7�������E�����ŞeϚ��P
�E���WP��Q/�>w�U�{��8��|���_�r�P��}�����	����$@ca�o�8�s�w?��O�jh���l
�����NI�K�}s�O-�ߴ��̀�p��Mm��䡬>��K,��&�y�˻�����ev5�[�D�JM@ڶĳM�fܝ{/b���To�V�>�Nh�����x��̤��u��+�/G=������	���ͯ26��%�V�kG����4�q���o{�N���&��m���c=���2��V-e�:�.�S��~҉V�!�|��ci�������N8m�a
%RP�Q�8=�.ŝ�V+Z �r0]s��`f�ZsM0~����O���V �!����ȸc��x��\�>ٷ�>6v�gQRr�G�2K73��	l�?��Ԃ�8M-Z3���d!5"'��so}#�w�8�ˡqRj|TXlxVHYEB     400     130�S��K�ڮ�c��a���X��!_���K���w�a�v�V~�~�%���&�w�E����$-s
�G�_k������Ro7����̰qo=�}-�'G*�6z�֠����dv�)9�Ykpa�Ǹ5���yiV�CU ������g���r*�йܼ�E�Đ��'y�X�,yz�d8Å֞[.�W�1\��`�K�/���#4 �
��9��'[{�1EAv~dsq�1ly���תW#����<GWK78�eL��-
���-�
�_fO�S�<��8Y����A�.��Ɓ�
�ϳ��y��ߊ�XlxVHYEB     400     190f�๾h�����!��@�K��J=ꇃ�3n5.�T�R�p��ީ�;/Ϊ��NZ,���F$�I���i%�/�cYZ��Wh�#���ӥ�W'��T�Ѣ�������p� S%�4��2�����v3�2Ǻ���}8�r��L������{.�i�uϙ�������"�W�u�˺]w�1;�~��y���_�a��#�¼" A��e�@�^dK�� �g��C`:)9�z�]�V͟��7��?�#�:e-z�ym"�x/%�nV[{�FU��Q<��E��Q!�$r��	��C��?�qaؚ��w�1 ���T���E̋R�!]�{S�L��D�:�?ҷ�$�;���u�2�'�O���v4��k^LB0
ꥎ��UԠ�9�$���9���j�XlxVHYEB     400     190�JUT��I�H3�/i�V����̵��Lh%T�����YwN7e�t��Į�8Y&_ہ���hv�.H�\���ũ�^Y��K��@��|��c�
�Vi�D��a.W�)���{��v����J���%�U�7Vwʫ���iN.�d�S�*g<��۝N�\�)5�\ն�H�偖�%�`�o*m]cTo�wq��'���8��k�Z��#dUMi0�ڄ�#�G�r�q*�Z�b#� K�دD2������փ�u���O��o�Cà��_�޿��@J�\�����+�vIj�����lAgL�z�ï�@E��t��]3��9(0eF��$����~����N��`?q2@��Αg5���(?L����^�
���O��/w��t$� mF��HXlxVHYEB     400     120�j����ף����=�{-�/�(�w��{ ����U��D���_�P���' ̋ɟ-���bN4��:��V����3@	�����A)��I�8n����+��h�%���p��5��6��O!��zW�_�at9c)Q��?A���`ܤ���_�����E��a�Vj$P�L5�"c"�4%�7�9)�n�Bc�O�\ʨ���M�At�4u�;�����0����n�Ԣ-"��B^�/M��3��Y���U�x��G5[�?�@i4
%[��WJDX�{	�,՟�\u����ΝXlxVHYEB     400     170��]|�ׂLp\:.
�7Xٍ>н���_����#p�kY����T��u��}0̻���$�C����r���������W�H*:[~kߌ�u��Z
�������8���4���Uv��a���C*Ha�,�.��?.�)� 6�8ڶ�,Q%y��i������Ƥ�@��w���c(���,��v�������
�.�%ư�xN=�!E�V-�08U�,�:r��2����cPJ�Yc�_	8�����\�5��5�
}&�li�;����k�1�d<��b4c�b�4�zO�Xv�/�$���������&��Q�@�W� �9R���H�L�@�Z�/`��\��d�{�W-^@2��XlxVHYEB     400     170��e��c��
�B ��ʋ�F�Oh�r^1k�VX��o�L�S��r�Ns�ᏹ��_B������|�V�Ŗ�((��c��Sa�xa�k_�i� ��{�+ZQ�q�~ Ips��E]ܤ)"	SPb��	l��b_5��8J��|�>��tsj�pF��΅�OB�[��n	�İ�#Y�5�f��KP���V����_x'&Tsg�s[�(���Q�d ���8���@�-De�
s�)bಘ���hL:�����
Y��X�P���rqv~0��Gq� �e��h;��.��Ś$��i'4�rB����Q�W:f�&٠)W��i����7���$T��GR2��"��?hh(�\���@�XlxVHYEB     400     1809��dad�F�i|�|O �|3 d��� ���Q?�#L(�"V~:�eC�]�+�J8�l[����5��]�y����\?$�}�捸��XC�������Q�w�T^L�d̐E}�FI�w���@m,h����$���Pg�(���gf�f6�o��."��O��lk3�� ���RWv~Y�ط�J1<�';������N#�88>�:��u	.�Uy�z�K�U���A�S`�`odwe��!��{9�%��/T�+<���o��k�#/�`�BBs$�A{��XͮÀe9�xU/B���:�80��h��6���y>0��u�k-Ө�|�/*���+P�9��,AȄl�N\x%*'*��}ӹ��E�e�XlxVHYEB     400     100l')�iX�t��k��rHkI������[I��Ǟ�P��	���W��#�]:3�KS��Du��~���. U
����Nj3�.�7�_w��h��Kō� �o��v$+ W�+&̝��.E~�>���F�b� ���.�퀶��O6m���L�&�\�}ˠ��-�^�e�PvbIh@�D�Ms.ۜ���C�(O)!�z.4N5��8���C �n{o9X�A$�T�3���:��(���w1]�NXlxVHYEB     400     150��bϣ��:�>���O2�����t�Z��a���R�q�^5hܖ��p��Xo�{�O'71��3���e��0hi�	D؋.����[_R�ZnF��[R'��ȕg����	��D�iT�Ǝ."��{��tmY���3�o��Юp2�KEЈ�a��7Ӆ�k|���"�Q#p��A`���&d�N�dc66��C���nHw��Ě���[䃙ۃE��P$8��eL}Xa�Þ�c���sě��Т�3, y����O3(Jy{��@��T(�x�S�y�<��c�J^``���Z���=?Qw��S4��� 3�j�,#�@[`?XlxVHYEB     400     150ԡ�@E�Ѝ۰c�|(5��}c�g$9^�2�hl��xuW3&�B+�(��V��鵣��f�a�(��ޗ}��I%0��s<�:G�T�e�:u�K��$����ڈ�^��՘)Lt7���AA]���Q���fq�歯�T�1/�-rC����CrL�퐱5y~�iGs�o;A���4��盭S=RB6�Q"�֏B_�M:
|Y�$]�U��}�i.mf�O`|�6��r��0�B��fU}�:AVR���"&��y��h[��v8�tp�
�k�Q[�1)EW@�0%%�xt��&>tՇ�4�N5��_Ŏa��Y5�����C�<c ]K�g�ޫ��XlxVHYEB     400     150:-�T}��¾�h�I���5L�\W���cԠb8��*�X�����y���� ��4V��T�ÁF�nU��io9Z�J��6D*Y��q*��Ej� �Os y3N�ۛ%Ap�M�_��6�f-������>r����Ƽ�j��IV����I�C�$ E�]+"���7��=!�_,�����΍rh	m˭»���!��c6�F����7����&�H���M�pF?C�0�i1�;�gH���+�U�kC�	���S<��O�������B� �7yuy ��M�-�T0øi������Xq�\�Sj��=hg|���
&0W��6��l��Y�XlxVHYEB     400     180��Ʀ1J����tNG-Ǭ�y[����<����&��4z籂ؙ�(�B���K�[D���c�"�o�\]0 #��SK�R2�V�g���1��H��\�(/�)g�u���y����xM8�vڋ��L��I�=�|�Ay�c4ܬ�y�F��f��f����41����T�m։+1k���ƞ�7�����T�S�!٬���\;s�xz��"B)(� i`"j^Fb�U� K���Ot�>�(�HZ�E�]��!��@Ū����X��s��8�i��ĵx���n$��i[vJ��Y��ΛQܣd���kp��c̳�6ё0豋��z�$���?���s5 �Ac�]�q�s�p$&�ohn������	zXlxVHYEB     400     160Q�h����K��B~�8���R��7"xY�����v��~��J�EA�ϳ�4<��t�n� �=�s�ꂲ��3�@�D ��iBA|�sw*\z%�L�
Kپs9�:����Oݳ`���1?9t]"�=�Y�+�6gˈ#N٭xN~�(�@l9?�ιKjeS�-z���8W��'ߦ�Hv��~�0����{���z�$�Y���=m0��I�1��Q
2 ���q2�2�����*������in�jq��jˑ9���%P�`1��:���p�]����dPg�y�-C��.c�{d��馨	��Ys%(�XP�������q���J�zSܥ�)�C���ìU�I��w-�C\XlxVHYEB     400     1a0L�q�'*мڠ�ۍ��ӓ�!4	��3�b �^��c䤿#B�9ol}���a�܋ٹ~2<>-b��k��)�$�˸hW%�j,�r�����?`���'u��p`� 9H��_���<~���I��Pp�Kc���~�\j]$�/��,�?���|�^8i�2�XG�.�=v�eHA2����@:���S}D���I�R�m��{�<K ~��j0-�R$��H�<�����l!"ٕ8��m���9�:��ZQ�HfLrRQXM�)��j��L�#j\q
��h�-s�1�̨�?k`���ʬ�B��|�n�9`Ĳ}`CbbX������N�[ ��9�D��`Α3bq88������̠�k�W�'j��!��,rƱ���>��'�_қ��<$ݶ��J�0�?{�����5<'�gO���XlxVHYEB     400     1f03�Z���߻�e8����sp�<d�wNXm�e�6@u�mu� �5^��_P�����b���g���k�d�g@mǳ�uiz?�a@���Q=c3������OO�(�b��j �pe#2��6b��V���si,{��#;AW�����VaU(�~Vr�\���b!m�5��Z��6��s2�\Ȉ�\UL�r< �g�7�1�ՊHW����tn�&L��a�H#<��ڹ|�.!:G�@o\�7h���b���I
�V��FJ{_���w�س��R,��׆�x﫦��?�x*.�/���9.`$�h�>��t���aI�ѯ,�����_8�~PwW�ϕ�!��R@~Ȕ�xWQѨ"�7��*��׶��"� ��k��*���[`�u�̣��O�(9d]�᳡�{A���T�54���^1Q���ABj4�ދ��~�Wl�GU�L�W�ɨ=��1�Y���:UCͻ�j4:fe�t/g�ɠl�c)r'~����XlxVHYEB     400     140�ӊ��m����o��x�j�QG�n����5.+M�G�p������Y�P�L&`]�,[B�~�<%&33�r�H&�o~��;@4�����g(Χ
7]��`��� ��.r*.�	/X=*�㗰�� yB�%C~[8x�����qw�;����)�+b��+ōҠ,'YW��ep��׿�[a<�<�(��g*��<�v���X�UE��ێCz�������Π� �GY�[{<@��fe����ѢIX�ي\M!��N�<dW�
�W(\���N4����&�(�����x�mq*:a����t�WhL0_e�{B{Ln(�VXlxVHYEB     400     140V���L�����n=��}�Y}E��D�u_��@)R*�7�
T�.n��*�p��ǻX��# k�P� vZ��[�rY��H��=�����9?��}uL�$:��"t2�m�y��r�� b�E�@���B�U�Oۼ�eWm��z1Sk�6U��m�$N�֯'J�C���S_�]p0C#gu�dN7�^j��dH��hI/�� ���Q�Fx!)?lC�ʸ3�*K�h��;���x��J:�����V"4vДgQI���kk���&���zH��R�qA��p&C�^(���?�z�xH��'Uhp ��
^�(XlxVHYEB     400     1e0A8�� ����b3Q���na�FK�,$��o\dFP� �VY�w0B�"�m����  ��#��ɇՒ�����b�f*ŕr�]��w�Sd�F�e|�����(�CH�uhW�=�
ն� �0o�+^,6{����=���?�٨8��&��=�E�0�B�\���|�/g)u	��εj���8�?�������]�x+�X~7�	����K�]jU*i�Y�..�lc:��}�޹�MZHw`��hM� ����/2@�ØP��,�ɭ�	�����ĸj�������3��H�z��Ol5=Zf�B���~���x��"��6���M�x&iw��fs�P�+"g�f���kΊ���H����|Hj۽��I�+x��z�SkΘEK�:w�B��R�g�ޘ���-KWj�I���&�'�ɻ�<Pc����G�˟�3�nm@�/�q�}�3�S��v"���ѳXlxVHYEB      90      90"��	�1�.`u��'�lI�
����(�A~�%m
jAt���Ǟ�+��r�O���Չ�j�����-���.�$M-�%m��L�S���� F0h�}�֚u�����}�E�X����^:��7}
�#�<�e��;B��y�Bχ�͸M)'�N