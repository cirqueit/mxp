XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����nJx�d;e����5�:l�;fw�I��J��&R]�!�YN^���sn2�J�iP�i�m���(��.�M��ٞ�r�ۈ�s4��ʔ_�	tT�G�������$�eG{a��MY ɰ����ON67����m�����`��W��qL�HEWn=�}�Xd�Au�,[d�O�\�7�;'%�,����Ǚ3Of3����sjz�1I�\Q*ZM�X�^�����Nua֑-}��z�ZW��Gp#˽��\�+&��=)f�H(�b��C�T����fׂ��1be��X�uB����%s+�d���h2����$�fwcQ�	˶��;b��$'=9����2�6애�ߜІ]��IoĘ��{����ć,��D��Eo�-���>BbK��Xy��ؖ)�����������>ҋ����!�Rn��/ � ��+�bL�M4��&������.����3���۶h�@��χ��von����z`��}�sG�^�P=s!�����1U/�\{��ۈG�ѬC��cn���rB�7f��Y�8Ī@׬�Κ�;��;7�8N��Vh�8֙ܨ��}�����vZ�b-���X��p��E@����c$>�$&h��k�� 3Q�L��N��N(�C��]��]�f	��ez�x�ԴX�6eǫa�T[?�1�Ƚ.�"E�&"�0l���̉:��w�h��ӣ��¥��%��D�@�����x�CtG��d|�zȳ�zFa�)B�5edV����G�l�XlxVHYEB     400     220P6�l��#���r0��a�r3圆;�C_T\Is�h�,��X).����c����6��j�}g���d�e�Z���ѥ���<�J��Ɵ�S�#L���_1��?Ak�Q�������?��\ʀA��<����խ�DJzX%Ó��*�yIf�F�w�l��U* f�U�U���%�
�L�vsn#��|#$�����䦥Ɨ��Ĩޥ�iG%�2Y�%9�#o#���4�G�zϳ�I�x��6W#��}l�j��B(0x����$�au�Ҹ̈́�����[�f8�{�ա5�ت�֟T�t�Z5z������,o��N�D����%�W�?�t����_" �+!r�nT�3�jEBo��r$�xL���<�GP]��?C���?٤�0tQ6CD���R!�� 埔��=z��7y��AXA� H���!�Iש�\�qc�h�m[P#pnI&�����=�d�(���먁�K�GU�S���$7�V�Y]:�{�B�JQet���VP�5��S/̬�He��'��6�}��W��W��yN'�۠~�9�R1"*�Yt�XlxVHYEB     400      d0w-g���Dy�p�7@�65�h9�!�ed���IQ�rjݸ�����2�$ \�<���f��%��[�4ݧO��=�el9TDB���92�}�i��GD/��E�E���~\b�6xxסKU� �����t~����Sh�)1ym,R{,.)&H��l`��P(�u��]^c�~L��I�XB��?{>������!�>�c�AtXlxVHYEB     400      c0��@��bi(��4E���%�Y�k�lE 2����0�)��B��mEu�]֔&��O�/��x�r�&���=���l/�S7#��2���Ozg8�ad���O��e�%9����I�*�h����)N$/t,�J�#:��c-���1�t�~d��]j��m�e��~��g�%`N�҃�+����w��XlxVHYEB     400      c0�J��\DdC��q����{�+F4 ���Cv)�}�b��i�Wʵȸ�*���.�:�V�_l�0����������Qg�-t��4k�3��ciA����7M���S��ڊBb' �!�]�pH�ܒ��c������?3�<�,5ػ%�2qn^1q_�A�Ÿ��gn1����#m�ѱ�C����ЏS]ѮXlxVHYEB     400      d0�~l�z�i�y��>��]�	4�� ��ֻ5�M����D��Y�TI�R@��<�Pq$��b��^���>[�<��L��P�
u�n����J��Y�n��%�R�������Ŋ�3�%�[�we"���E��':W鞀���f�nٴY���-�{^矎W��� ~L�+P��f�k� $Cn����(Ϟ��F�ز�'f�#wXlxVHYEB     400      d0맼Z��d�y�� %ߩ���]+E��6U	|�S�K���pt��GZ�!�螇��UG+�v�:����#t��r�`��qx�8�/}=7�(���<z�����m/x����R2bQrj��O������%���Z?bz7i!w�v�w|�0ҹ�en ���GDM[Bu�~g��zf^���swi�yƂ�-Xw0���/QҺ���}[��_ XlxVHYEB     400      d0���ׁ�����hڌ�q��*��X��&�z��ڴ<���Z�?,���.��W3�����I^��ڄK'�a9%�~Gwy�ڹ��䪓�E���_��^g��KC0�
�#�T�"$����ȾJ-�$ո,���JV+R7�af-P�%Ɖ-��<����1����1O��ٮ,W}�����a��dz@I.`Ӎt^�TI��ħ:|�4ċ�~'�|XlxVHYEB     400     170&�ZX-���X$�(�|e����>�LG����/�@��TP�T���A�E�4!r��3]㽀G�����PI��>���6d���x7�~��~JI<��o��#�]����P��Z�h~�2�ƫ���y�����1U_��t*��)˺�@T���5��Q��g܃���wx�Ω�k�ݦ�¹pK��%�Y��R|��P4eX�f�&0���V��p������N�j+��)*?֡V�H���,ެw��w���߳�c�@��}\tf}n�1!��^s%�V�CS�<P�,�,�:�W�J���62�6I�.�E�g��5ȞJ�i���3�V"��q�Oe��:��m�qZF K�J�� 1�vjTE3����#r񗒫XlxVHYEB     400     140d�����녞��~U�t�G�UD���=B^<R��u�O�A��:�|2 ³"�On0�0��W6(�"Bāa%��c$7Ӵ����`Du>��e��j�|�o�j��sj�!�&#�2���Mi'��$">��4�H�DK��a�<mv��oc�`�D[����%q���5�b{�ܦ }����L�[�hf�����QΫ}lmy�if�6��~�u.�z%=��:��R���08��<�Ԣ,)�M ���{���Q����}/�Y���z �y������hV�{�W����X̵֝w�=��Aa�:7)�T�U^����ŜXlxVHYEB     400      f0��!�Я����`�~Tz�b���T�+��9q�n���NX��YǯE�Ix�G�}��CB�
G�Zgu�A�890a�k)������b���?%*6����.r�GR��S��2i���c���d+[�V��5��C����FT���l�<e�jg"��1Bɭ��j¦�vW�3�g�)YV0��g͏��Ad�ȇE���C�P�6���E�m���p4Ύ��:若"~�� f)�@�eXlxVHYEB     400     100�}��,�Q���Z���-���Q����k�.`%��_wl��}�� �;�%�"#*לFu������:�Zc0�\-�(�haX�{q���� ;�b������(�[����s�9�r<~,ߩ9L�1a�X�Z˚�������'����ꯔWSCp���Lw,	�M19<��(Y������<Y.?	(��i�ѷ9������ R*u�ٯ�+�=�)�537�mT�=�	�ߊ;��ҭ�fyC	��𰦒yy(�]�[XlxVHYEB     400     110?jIN�ἂ>�A�0����&���T��E�&�<�pwJ<�,�,,%e Zޠ�kЫ�=���
�g��ƾcVj铘�͡O���~&���_�bS�����s2Z�o�������s�u�E?���|�E������N.���`xXׯ�Z�>c��f+/��xb*9�#���t��bh�S*�q�����  q����>=&�U)m,{uQ3�����pm�P_�Xq6;�@���+V$=�f]�����͑�V�vE��1�D�fl*���q\qcXlxVHYEB     400     110c�CΚ�'�1��b���'����lh2�ӠD�8OǶ���"������[}.��.����}x�(.�/�w���|B�b�y@�̷�s��-7���(���&�=�ж���K����IR��#���0F�!ΉK�m��<��Hc�!�����Ɲp����O�_��<�/\� ����[���;La�yA��7*�wA}�HS����Q�v�B��� p/���ɠ_޼���%�D��^�9�5�FeL�3U��H�,���y��Z^] XlxVHYEB     400     130u�\�ɯFH�G�T�##z�q#EH��5��d�O_e��_�ÖM�6L�ϸ�oI/��R)����Qcx^�9��(ٿ�U��H@Wj�c	�ϼ=!��f6�i����>�H�0���Q��f�3H`?&kr�zo��K<&/N��=�*��<i"@��;D�m�.X=�������g��X���V�r��Bm�k��A�����,�������G��fs�}�����-R5��<}���,�����rR⚊�W�z?��D%f=)�jx�0�x���؞��J$<u��E�Vȃ����XlxVHYEB     400     100wT/��v���g.o.�����'K*�-]9⤨IS�[x�e0G�������0��k�Yh���=��xh�p���6b.�l�U�y}�g�ki�x�y���h%�3��tlϏ(Oɼ]�����|�B^p�gc��sE-�e��F�����&�H	�� f8�@����g��FLf�t9������������wa��!�>4����Ae�������L����+�Έ�.���M����Qt�
 �[Z�
��0?UXlxVHYEB     400     100�	�;�+w�-e������r��u(CĝX����{����KLl���qj0�̖���D��hD��Vd!��-'�c2�6�١5B���c�U�qW�F��&��+`J@�y���'��^����������͌�I��B�C�6 4�+gt�ӟ�.�"��I�H��f�Q�u��g��N�a|-�W����dT4  ��?�ܦ����s��Jc.C��u�B	�nE�%���Z�[K�B��ЇS~2������	�d� ���XlxVHYEB     400     100r����B��Y�]m=��r9C}�i�y1O���]H�9KOK×gdyԅ�� J���/�lN������/ܼ���J3k��"�lk4M0�k�!Wh���%Q����^����^�*�C%Вv�1���v��x�.D'd!��q�N
S�$c?
�����������I��$q��M$n:�e���G�<B����������4 ��]�e[;o��(�[,Pm�P�Nȴ)�=�8����FX����B�ֶ�%�!?��XlxVHYEB     400     100�Ӑ�����X��ݯ�nO��uWL�J%(�c�H,,V�Ujb�Q6�o-��H����=��#�s���U����� �qz�qp3�;B�քf.�kI��^�1xbsy�VH�O��m0���)RL�#�*FZG���)��$�U�o(�Z��������j����A|%�7/�*&_����.U7gΪL�}���m���p�1~����O<QΎA���}�uJ����"�Q�? �Ϧj����9a�f�H�p�l]b��µ)XlxVHYEB     400     100:�=}x�r"]�
�i�>���L�'?�3̌��/6���|j:���Io�˕/}z�W>Ɖh���8:]�B8�1RCjQ�c��]u\�r������ r���*�#������5$~y^����-ŝ�p[O?b�t���q��M�ϳ�͗{�`�X�I	q1�uc�O��Ŵ�T[� ���֥��o��F���yzD��(�Sj�����j~���*{�����[���e2���������,�͑�¹T�٭;�0���"苦�XlxVHYEB     400     100#�ˉ�T����9d�J�t�/�e�r�VmR���`�w��<��/��=Ь���A3:4x>A�����2A��Š�`;���gL�a��"tZ�{j�\LQ!�9C"/�)�nc���$���j�#z��鍏Y���$:'��ݠ\�^#49S��Rs�|fngn�7���F�"҂o��jf�5t��m�V�$�W�<�YA�Rv] *T`C�BE<ѯ�mB�[Fr��	�wo��>����30�|��s���ҪXlxVHYEB     400     100,������X�g����]g^5��D���r,�|�;��`7���%�W��X�6w���u��x���U �>��4Y�}3m'4q&��߳xY�mN<�ˠ	>N�ᓷK��Z�n1��}��B�NNJ�u.3�k������'9Ce�`�����?Ħ*=ШY�ǅDGX�i����:KrY�M��B��z��[�L��m	�L����ce�c=wN_�L������:����6�6b�"��m���ɋXlxVHYEB     400     100z�x�Y�6V	��*��O�<�{�}�<���$-�Ȥmט݁���o@�6����Ƿ*B���#&����y8ǧ�}�S��m�%������	%sR�ƺ ���f9l��M���I����
�uc8bzօ�r¿
���!�5��aE�uAX���Y�o��<��TH�}D7������Zc�u�qt��y{�zt�Z� ]�g�_wڢ��W�9@n\؞˃`�9�����;�qN�m3�,�~�R��5�k3���-��
XlxVHYEB     400     100l����<�d�H(���x���/��δ�k)/H�U�Ი??��R gOD�w�������(4��w���Ē:���C[�y��i��<�ۑeQ��V��w��4��'I�r�S�^U���?s8��B�u��6�7��5���9�t������)0LYiς��X�]d���ugm孙�wTB��	t�(PQ�0�\�Q?�ºw�x_?gk
A{��C�1C�y���br�04+_�����d���� �^ξp��/XlxVHYEB     400     100�S�S����\ y]��cs傠X6d��/(}=�t�ha]�Bl��o-�.�T���5{�6�ceZ�e��-՛�t��+|���f�Xrq"�/���2����/�WX����Q�GG\�$��g�unk{��F�j,m(�(���M�ײ���pK~�i�'C���Gh�K�"W���wʇpu��ȑn�� ʥo����k^�����a��� Ɩ�؈���=Rw�!'l�3�gfի-8�� Y�;��6XlxVHYEB     400     100�P�@p=����s�^�S���W����5x�&��N�-s�s
6t���/!���8	O��h*�םBE���H�	3�@��!��!,��]�(�=\�
���Z�k��Ŗ���5�D6���@Ty��'��~�ŭ������i}���2[{-��^���}(���o2#�>�ze�����x {���3�uK��D�n�Ҹ�b��ex��yq7x�����p6�D���Ύ�\�<�9��o"���!����XlxVHYEB     400     100<R {����@�Ф�8���-:��Զ�|�槺s~��L�Ʒ��/�,:PT\�7�6��E��il0L`�4�
%�����=��r@D�m��v��8��H��V�G5�(��^�Y������3�R�}6����vti�"������i�4p���#�Dm/ǵ x�]�1𑘬-�L������L�L���L�J�f�t�Lzk�(�dy� 2Qxf���iU�R�`\��M������<M#C	�y��٥^�(�P̠���XlxVHYEB     400     100�F?�*��Q�^ ]�7tt�!�
�SI������f�Y[�*Tw��~6򹟜Z�w
��X�<�L��@S���}ζ2��ȗ�mh9�##l�ak����wGo�+E�_��y���E���>RA��d�����M����PS^�]2ҿu�:V���)F��k-�F�!{�Z��rws���9b���߻t�i��l�c��=����)��edyf0����j;�ھN�R��nf34�}~�vBNm#FX;UXlxVHYEB     400     100��G4����`x�\��� �&�ד���j��W��9X�Srbk�B����h�|F�W�
N	m�>v�a�nnl���*L6$��C�>�#���(�����[)9g�Ǎ��7�,����Z���a7h5K�"V�I��X5���1��kt��N�SzpI�6:�\\pb�Z~d�/Z��v>XD�]/<6a�1���(|Ǳ'6������f �8���QdUY�A�.}�p�2�f5"�ၱ?��8�a�>+��i�R�XlxVHYEB     400     1008�&#�"��k��ߗ�-��9�����=�¿�] ĳ �I�b�����@dȜ���l����ڑ2(�L��[���زN`z=XW{���$�n�/x�<��ݑƣ�J��d[*kn�
���<��tB ��+ܸ�H�z4�v�n"R��c���8�1@/�˥nI%��}�e:�~�??p��'⬔%knfg�-c����s��՘/K쌙��Z�Q�Z� ��9H������z������L��jXlxVHYEB     400     170���GeZ{%7�����8��Zt���H :V�e,hݽ��IwI
�	U�[���=�%�p��G�z��!Z��rY���w󕔍���X��`@8m	�d,k^>lVQ'H&*���|l�
�e�8�^���vZ���F�g�7�q��v�r�7kp����឵'��E�#�n�U��ީ>����Խ�K����B�{�c�=]�iB��&���ih�b�����޶D�a�L���7�Y(����a!� ׁ�;� ���)f���˔T��O�R+N愬��@��򾪩v��`7��-ʜ�~��*�Ij� ݱˣ�?s�*0A.���&T��Q�� i6�W�@`���4\iv��v�+XlxVHYEB     400     100�w��&�	���G�����Я�j��5�����O������A������r�?1L�?q~Ź#2��GKԒ?�R�-3�
�Ǎ�+K��,%��H�#�1|�{ӢW�t>��<�x�]`PܱF��9�jNS�^����ewP6F��uR�ށ*�_�Q_�#��^���?ϟG�V�(ZfJzT� 9b�{�j����Kð�=\�E�o�xW��Jvb��ԭ��zSr���D�/�4唍����˅is XlxVHYEB     400      c0{R��J�z��Hf�F�t8����(d��N��(4��o�]�������p�V�XJy{����kR�m�8@a��&Z�_��,�r���~G0�Ud]$G��:� .��$���̕)�lUEM�rحZz��BLi�F�XQ|cy�n9�f�UP��pTjb*�5J��@^�g�3؜k �G�F�3�Sl�0s,ոG�l�XlxVHYEB     400      b0������g�p�݅�S:�݁(p_�����ޤߚ-M�u�Z������\�8�SH�ݺ�X\��ƪ�D��&���
ҲEG�Y�-���F):�'���$V���]]�h�:j�`�&�p��.7�F�׊�D>��(WG�M_���L���4����$Ru�r;طeXqM^�XlxVHYEB     400      90��׭E�D6F��X�ϲ��)�����J$7��;��9W�1��s�a�
�k~��<���Aaא+n��
N����x�]o�����D�<�\+X�4�;�pNk���/g8|�9�&���!�ߛ��ʮt�?o�N1����5�XlxVHYEB     400      90������^I±<d-ٮ#�K�`�܎ܓ�	;���\��i�@������� ��M�y%8����������Ɵ����A�'�D�&է�Ɇ"�ރ��C���93����)(�����lKf�ٜ�������Ur���3p�����XlxVHYEB     400      90����Z4Z��}�R,�v���'�Z��֟ZF��KG�/�R��M6��y�e���Ъ(��^7,�}�k�8�]L��h*⊝��0$��o�u�?�Zd�Ҕ,=BP��9��� [��Ք6�V��/xY�L�O����]'K� �����XlxVHYEB     400      90��Un\��ZA�������X��΋��8��Q�{���N���&o ���v�(-|��4�g�T��1�\  �k7�Xݻ� g!g���P�4q�i`4`��Y�����M��7ۺ�%y���~^t�G��5V�+XlxVHYEB     400      90�11^_k��u�\c`ͳ���xu[Z�(?6E���gg�v�8��Oo�h�tI9�B�"v�"�kH?7˔����.���N�^Z���uI�����{�3�R>��+M��+��H�z*��L[��ē�}���j)`�:7�3�XlxVHYEB     400      d0͋0��z����g�1��O-����,�ܣ��)�uL{ɆF����K����r��֛ѕ6�>�K$M�?q~�y�� �����[�9��`���e�^6�Y�ﻠ�-aΫ�zj�ž���X�@{yi���
��ǫO������H���Q�j�KR���R�W�~�_`q}l
���p���� 	���Mx�ۗ0W�iE�4=(��[-�XlxVHYEB     400      e0j�/��w�/�>!�ّ4A)D���ј�#CڮC�26�DX�jEz+KmG��oC��3�&_$�PQ�@�"�A��$��*X4����S��
��Α�������X*r/��%̡�a^�h?���)M�PFk��2U|��h�r�Q�;��#����#�]l1�Ş#�no=�K��^�e����?�= }����N�5�-������I6-�\��C�E�੟E�~��.2[�}XlxVHYEB     400     100�d�������Ѽ��<*{�rƉ�
N��� ��rkGuB�z�o�W�i.�7��S	:��kAejҥ�ݕK�q:�-|!2P9��s4�h�s���Cp��;fƮV���E��絽��45�vP��j.�Z@�H�������G�g���ׂ�p������f�Y�4Q�p�Lw�8OA�"���8)�su�z �Nͳ]�͖R�Zȳ�\=3������#���M�����*a�DL�ȸBUO-*M�'.�bd���M|XlxVHYEB     400     160B��,�M�6g�!L#��\�ښil�e�����2���t�X��y��4抠}r�F���dC�X�n���lb{��'N�^hn[wZ���'s!%}zR�`���+Z�Q�f;Q^_��m2��A�#�d������q+3`�&�$�����~�6C�ۨ��M�|xr_�_���M���n��g �B��t�
P�?�k���M�5fR���Sa�4��f	bn�Rn���7�,*]m�2ܖA[��4��;�&�^[��l�F)kMGeUH���k�HT9W�X�����A"�E)����1%j��U��&�Y�Uu1lUUj�A���r�_~t��M^'�:T�'�%;������ҝ��{�XlxVHYEB     400     160�w�t��G��E��2�ί�J+Q8����Ⱥ��-KS��c@�J��0ܗ�xv��{~�!�6A���nrI�p�h��V�e�������h�j1����8׮���l�d�ڨT݆/A�>I'�:��[��2]�6�}�L����k]i�o4W�c����i�J�Q�qAJI�Ń��Я�1�1CN/�A�ۘ 2�nKd����a�5����i�Q�gcH�S�[6�b.�r�ю^����6�e��M$�_�K���զ�\t�ZF{�P�CWlv-��.L��q�IQ�qm�#d��l��ȕ.d'�� �:��i1gy޵f��b(~{�$t�
~�����XlxVHYEB     400     140�w����~��%���9=%՝'��r��6
� 8z���R=��-my2 �{��~�"/)��v�y�r�#[T2��	���]�����79?E�BT%u��W���/�?e�������}ζ>_��DTT�m����X�BCxv���e�t�il��Q}iT���L���;����E��
3
|jT�����W�6Ұ�/X���-�����V�V0��|�]T�E�&�=ןH��V����Fi�P���O�+��!�20t�S�$���j@#�8���ÿ�����~���>��b}���עWD��p�l�(�XlxVHYEB     400     170��[׭p�?�tZ�]�1xx݁|����@�2��ف�@�Aٱk���v'�ʣ$I��E�րxUCXS�2ĺ���i���.�\���x/5�vt4qqp\�꾴 ��h��a펏S��Y�,fa9{ޓE��� \���~���V��*f�Y�O��U��w��^k|7�B����]�K����6�	�5�@��"�d��G�B��1�� ��!o����lٙ�,�-j�V�5b@�^K�8������ߐ���r�J<�v����>�85_mM;�A('8{Z��[�]�0��v5w6m͕G�9��������^�1�������A���xt�dQ���B�w�
LţZ̈<CY���-c"������g�XlxVHYEB     400     150�8�ߤ���a1,li*���'���[U��rK�^�ʃ��j
���Y
Ef��яB$P�x�c$đ�׳R����F�3�s���
v���5�Z��k�.��ͤ��;�F�S�"�:X���Y�%�(�����; S�����Y;���ve�#�����Ǒ�=y���N"��	V�c�B��y��������h�7K�.	�`���܂�&�G6�R���+��?�w"=��\�S�~��jݖ���#Bþ1���,��vb΅g�B�ݛ�����࿗�#�2\�r"�4/l�lp�����=Aq��܂�L��.̳�aY���ۏP���qXlxVHYEB     400     190>�pc��!�����X`LB4�[�"�mr���!؜2���]�p֟;HB4$�xZ�&
(q9�GLc(���܃���nS�>�S��i�^�  M����o-_�.A�s�f�q׻P ��z��.)�<8��Cl�2����&��O:7�Jun��]]��?�@V���i�ҠW>/4 �[ �KW�y����b�N|�mE˫,J�f�!e[�� f�r:`�*�(Թ��в�C�9�@[�`���d|F�$O}�"]��ݵ�����5(��4oY%��DZ$��3.�fΕ��ťfcՍ^�Y�q�j�D������~O'͌#�Q��0Z�{|���@����X"sI�K�l��a��_��+
<�>$���/��]i���c�Â�)�}��XlxVHYEB     400     150_[笢n�$�x��C^��V0R����T(����*��	�&�1��G{�!�թe�~�5bD�ur��~x��6���4/�M&O��Jн���ȝ�������l�a0u�/��!JmY}TvCQy�&�f��`hIi���Ҵ����]��Ԫ)�~�N|����GhA%��I{?�!����Z�I�'!<x�R�r>�(0{��\�MY'Py_��>��p$j��:g֞,����QJEaE������GL�T�x6>�%� �z�qg2߯&����;�Y�Y��"�C ET4�+�Ǒ>���gQ�9qm���~�{`o1 OB3�����1Ę	u��Rnԯz^�)�x��XlxVHYEB     400     100��bH��2�*��a�M�S\M�-�][�*��[�`���߬�������}�����E�ua:��u,��&��w�>C���s�s1cS�ai`�DQ��U�v�x��>�r�{�
Xa���a�<n�[r��!͚e����J�D�I��?���Y���U�� �:"�
��΀�o�9\2�l���T��??���Zj�;���.�L���}n~O^�h�����8���)Ii���aO�X�*G���Ԓk��KT�7K?�dXlxVHYEB     400     190�����8�~������n�rӥ/��ّ�kV2��e~' Ղ5tX�����
�m��{ַ�E�ˋ�q�T9}�G�����-�L%�nC�J���+�����1Z��
<Jp��v[[~�.�pJ���9O �uOL�OJtnA$0�����e.���]ɀzZ�3d�ą��X�c��T���Z|��l}"@K4�L]N�L7�'ا��J�G	���b�P`��<�����}d��8�]���=�nC�e,�b�Ħ8؆�-�U���@q@	�-@��J��
(\n�[΂��foV�w�s����NL����n������HX�1�ʆ
T���iW3�IT
H4=|�oN/�>���������"��m\���9,�|�������gz9�nqo�XlxVHYEB     400     140�]Jd�ޣ۫J��N	������m?X���������y��#ا���q���8�8e0��3k'h�h����=_*u�j�� ؊�h��'TE;
%I��a8�^�(ڲD�zM8�z2�������a���P|_�`(��:�5`���o&�=G҃����yG-����K��C^�Ɇ�r�`���A+�ҥ!6}DQ�v8¼�ZPyOYo�w�oY*�K��J0�9���j����"����$��sS&b���]�	�y&���<��ʯ���3E����孙�D3N�Q�
���?���f���+7~h��������PK�v��XlxVHYEB     400     150��&�J��#��/�5��[K*/��wjqf�ሆ;	wT�o��d��fm�҅1�����GCsX��>�9S?+
Q�F��ѫ��WR�>���E�T����>�z��K��|�W��M��X����iַ��Mк��7�a��۫���=�Ls^�A;xi+IQi���o���or+ E��=�a��p�O*h�3$�h��*��.��m�%��T�f;���$$Bp�����I��e�T�p�vA��DXɤI�Te�s���[-��w�����\�����"�����`ѝq8o}�
yT4��{!C�3v7A�	PE+XlxVHYEB     400     110@+�@Y����h��[n�SBO���9d������ld�i�v�˛�.�c�T�~]l	��)��$_�x���*�({v�5��(��Q�T�(z�A��/��W�\
���j�;�U������:m��Φ���m�ka��jO���)]�~P0�XsZ���H�^���K�S%O�|�W�	�0	�y��2P�ga0��'L��G��a�&���hJ��?2v��q)}�!�62y���4�Q�c� �ʶ�C���R�a�b�鲂�R3/D`NT��'XlxVHYEB     400     160S0r�IAa%n�W���NOVɶ��n%��*-��JR�_����A��"V��ϚQ:�����|�I\'���扰>�!>N��]���q#�/|�<�d���;����Z�R�c��T����w��6S"��%��nI��A�� e��_6��9�no:�A0��� �8o8���z��L��(|�M�y"
FKD�GՋ鎹ks��d5)�
�Po�]��f�;ˌ�#X��5����Pᘜ��*ъm�Ѡ�x!�h��h���YIv5�Q���{hj�T,�'R�S�5����,r& �"CI�ϒN�?���?x�Ie�+Ln_P@�ջ��Cr�����H�d&�dH��U8���)%XlxVHYEB     400     160���b�������ʚfY��s�v~a`#d�t4t�����6&Q��T����f�v�ח�︘� �u�[�Q�gJ�@�$(�ـ� ��A�]A�����K{��`���|���u].Y.wձ��Ev ��L8���i�*�����'(����ڮ�~�G�O�"�?�9��b�&�5��
To=�q�~=�gK�¿C�{ě�Ls��,��v�翎���īB��J���� ߉���l��m���q�G1�-��]֔|^�V��I�/�p�.pO�m�u4u2(�JS4���K���1�Z�*%|�̠ǵ�]y��Zq�e1�&�9���<7�&SA�(���E<W��m] ���s��sߨ]�XlxVHYEB     400     150����*`=��+%Y�pa���Sى'po:�0�e�y�C�F��cq��/E{��������eh�෹,�3rH7q�F��Z7���x��Ȑ�Ю+̑��H܄��k,-L�I�ʱ)����{��ǡsX��T�!�Dz�> ��O�'�a➋����m3 �¹4ǏN����,c �4����A>N�M��}D Q����{ԎB���
{4���҈0�ߋMąL*0QN���2�׹3�Ƒ#�U@�_�S ��W�#���a���A����q Y�Z�_
�x�&l���G�ԓ�@�_�����M�;'��#Q;6XlxVHYEB     400     150�JT��4fxkE%��L�8
�����Ǣ�����;�A�ع�4�NϹ;�+�N#2f���9?ʽ!BR���d��o�e��.^�6æ`ZӴR�����L4�����W�]����hX�=y�CxF}���R[�.p�t���UF�U�G�rj]�`,=��uw��+��D�AvKd̋xr껊4�\�^!�p�&��7�.�iZ���6�k�ӝ̪ZP���P1��1��R%q%��=s���E2`vp|;ʲލ��'�r�U������:���N>���@K�����ؾ�91~A�Bԫ���e"^<��b��FXlxVHYEB     400      d0�I1�ӌ�jph��i,yfn���*�HT �z��X�")��^6��)���ĉUe����.�܊C��6��$���bnZ�X+�KBSQ�ic6~�C=�'�D;�I�6עy�^~���@��(�s��v�i�>9%5��0�a�r�S�<|{���d����T�&~QZ<b�T���%:!V!���9�\�Y�-Όx-��U��
��P7�XlxVHYEB     400      c0�Ǯ�.ɚ��%�Kx�I�
=��Ռ�F� �QV� +P�m���s��6x�d³��"]>�(��lOЍ��o�7��@p`���kM{&ʻ�Y_8~.L_��������K)TM�/\'�P�+�����2���秸*md�ᳮ`ߨ����6����Y�����ɥ�.�-@ח�Y��>/�E�XlxVHYEB     400      c0p��,�\D�@?��+3� ��Z�����_�S���z�����p�f�%��9����������T�J��2��^�圠���(ܕ
�D�&�3���Ws��ʊ��ZSO�R���+"�Ω�G�\f;��eV��Ơ{Y��U&.��l��'��e�P�C=><�?d{�SA�%bTY��"H˅�(�s���XlxVHYEB     400      c0C�`Aa[V6�fu
�B.禃��&�n�N	-�$ݡ�r��d�8���j}�b\~�;P���C�4�C|�~5���iY:���%�Z$�8<g� wy��"!�S��/���јc�Y\��H���D�. �����i�5�b07S�������q�%����<M����R�n������e�<��k�l2`��Ϡ�XlxVHYEB     400     100kRJR�~8��{'�i4B?=8)>x���OƨXW��e�F�]`7ڢ��^�����3�=@g���+�r��\��gK=^�fS�Q�(zJ�M����tz�'��{5�bh���su����3f�^X�M��mW��	��FJu� ƼaE��#��L�Dtc�ʺ�^e�q���8��G��r��
�:p�ˌ'2��(X�D�&��Qa��zˏ�C������e'�-g����>R��S�������P�;�](��L?�UXlxVHYEB     400      f0� "����]u�f��5kK�͛]t�ʲլ�?���ʭCjQ�����@N�X
|[�Wѧo���ݖ��^J8���so�˺�N�64�@�����1��sak����֛�Ǡ��+I�$�7ݯ�zh�AU�L/9i}�A�y�Խy��T���K�8c�������U�����7�.�ojGOJIi��aw�����h�j��o���7�-X�;6����bw���F��}36����XlxVHYEB     400      f0��;9�Y�F�~�
�`[h�.���˙�uՓ��?�43	�y�Z��N~ÙjW���Glغ���Ë:p�-���?���7�ܷ≆x,���g��ӦP�ŉ��+���~.��u��uX�Vkm��$�_���m�β(|��3(�nL�b1%i?;�u�IF;�L�{��˵�!xQ�N�f�,���G�9w�c�à��t'�cP�tq�똯�_X�p���4�I���[#k���r���ZCN��XlxVHYEB     400      f0����X�ʎ�����.������5�c[���nBJ�좈�	�K�G��K[_��� ���d�n�dW�Ҥ�e�V��S�f�\,rMa��a_��`̹���|oGn��fz��N��2���kB�G� z�z�����D-+袧�.r�[|P���xC�(�=���/�L�y�"*� T�|�<��'x�
A���\��e�4}d���2��g��pt���'�����B�I11|Y�KXlxVHYEB     400      f0ٚ�{���V���t 2�5��Uƙ��-P��e�%�������3��i�g��~��n�G����!��SkbuuE�އ�e&���aEԘ��LȆ����Id(�^a������8U|G0;逿UӉU�Zu����)r�R�R9P;�EƦ�]�\������X��p�{���<!�+Tܸ����O,s��\,���m� �����f?%-BnZ?����4�`���F�>�����XlxVHYEB     400      f0� ��>d��I��������L$��K���_��pw��U`j�A6˙辱*���j���e�Ga`:E�V���SL���`��_��ˈ����8��pM�A0�n�D�i�6bS~)f���<&^��{���_��i�M(4>�ӭ��ap|�����]��3�� 0��$�/�Gb����8�4��ȕ�  c*;~�!Q�)�Ι�z���h�Jz̷�[~~�8
`���h'2�F��o(�M5�C5XlxVHYEB     400      e0��;��~Ũ���x�P"��|�>u��c|�n!�;G���5TF��4A�u著1�-��[�(�x���7��T�L$���fV44Bo$�ɁjdX������������8rl%�l2�w�i���g������jZ�Z����y��%>�TL�S�k��E_��S[W.��h�5FI�K��1�t�@��y�A_ͽ�����EA��׺�׿XXlxVHYEB     400      f0����ְyRNے�[BF���NA����-�9
^�r��V����^�&8�`=nQs�]l8�W�!����,��t��ڽ��E�N�$�h�$��v��j�5��d�ܰL�u�+]	so�m��������j�	�<��Oݠ�^�G�_f5��t�Eq r2X��%G�|X>^+�R�~���N���z�1��D�̊,\'(��ъ[�������UI�'�4v��x�r�cF�s��YXlxVHYEB     400     150�@�f��đ��L[� -�%�Ե��e�������~��fW�P�FӪ�*�%�-lEb'.!�L�^��	�0��O}~ze��C�)�E�!/����G\�)WB��1�b��J�+)�R�7A|c��a�8�=�|��
�{3��mu�:��e;��F*�{�L_, ,���g��Z��x��*mR���0ZOGj�S��5�S*9�䏻�q��W��s�M�F������j�ze�� e9n������u�끪�! �E�C�9�&�<SH��Q�M��b��!;(|��!�G�;��3h	+��X���.k��)� #��B��ets9��SN~��C�:�GRL�XlxVHYEB     400     1a0 >5ƫ��j�-�~}lM���m}6�n������dћ�]�	a�	�Β�h����
�t6T?���|	2��)^�`�+��GH�>Tb
��J�0�y8~X���Y�_�Ȳ�o>UC�RnW{�ʐ<3���"�ܒ:V�|y��K��B戥_���|��?	ꠟ�-G� �#ںMs2�P�E�~RET(K6�.��������3��K��Z�������{��\��N���V�5�7����V�YA>9�����>y���)/0�F�sP�)��~	�[���
��fOx�U���z^a�\c��c]�������o��<�&�Ln
���ǳ����(�����4��h��}9$bN	��>�H���{��P���9�p�8�RuҲ����Ydl{��;�#i߀�rSD�qj�M���u��XlxVHYEB     400     150cJ�YC�������^6zS�4M�dDO�Ů3 n�q��s��ׯ���ӝ�tE�­�W��JL�����L������0�;y�pD8�����+�������,t
h4];f�����Uv��M@�[����t�1�Es�[1y�'���翚^�+uGl�;p�b&I^S��J���|�d��Ѕ �-�%��;�Y-��J�]h���0YT�kyb��0	���a�6���i��~(��O��ք$]�2W4?(2W�_/��s��H�J�����җ8;G�A�1��VR�'��~�&I�?�d�\��4�L���"���XG������ך$!�XlxVHYEB     227      f0�3k�AKh`9E�Cׇ�ݿ�ե�×���'��	�x"_��ղ��" sg:�1��!���ת�~��jh�+x>��&P�]� ��\<��,�X|�O/�wh���D
��y��o�Hw��q��J.�sJ���1!��ywq��n�Rr�����4<i���=��V��n��C���=�u�\S`�Y��~�4�͛:f�4$���^@��U����B�7l� iU��5�*8Td