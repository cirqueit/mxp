��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����¦`����\X��+�[�t+v-]/49��V�, ���0,��w�tp�R�ѹ�v>b�_�������m�H{
�����OW��S�AKC�4ɇ��Ӽ�&��|>AP��f����A��ų�Q+	Q)��]�᧘�·4�V�)`�a�P%�ו�\_�̳vւ��P���c�F�[T��rq�4X[nnPG����T�mP�(SF��{㴝q�W�I�Si�_jz7<9�����jӵF��[TY_�Y�Q�A�s�_5��]]4ŷWX�\��y�cjK�In�iWH#�ķ��<�k��봞eu�FqȤ�0%���L�u׀4�m�c�(�'\3�E�]�s?_�k������ڥ��;�Y��i�~��Yz�4;�O��TW���-�R¨+�����,��;�[1�ҕ����W��7�`��=��m����[
I�:�Yx>
m��������kfb�GF��S�
��v��S��T��,�ze�9��3xvTUĽ���tPeKߝk3n�g�@_Z$WL�̍�zO��T0"�U;a�4���h�.Au�JS�A�uf{����e��V��˒�D��.�E� ;�t�k��IއR�q�����wj4��3�Q�[X�XI���N���ߍ�4yZ�.b1;D���ݑ:��56�֟5��lꆨ�M1p-�Rb�ǓAP��|����O�V5�z��*�VBr��(�H;7/f���/1�V�S�u9#��5*\����]�o����T�:ճ�� x��R񟾋p���=���"�����-�6��m&e����>^�A��)N���p/���jR�{�Ѷ�LIK�Ɨ֚�R\ ���Ei(pFӤh߷b>G���t������SHl�*-$Ŀ�����&=,x=IE�:���e�k�΀w|��4�R�E�	t�pY5^��"3���E̥I_�
轥K�KI+u+ |��_�Q��a~M�>�������)��B�~�Q޹]��`������H�%�����) >Oc��c��z���}�����L
 �O��������m��5�< 0g}B�.W땐�Yh�Xd2���6@?#3���xW�#��Ѱs���O��۠������ki0e��6p�Ƹ��c	���=���)���4�ۆJ��:cxqZ�>�7�t�p�-g8[�?+[S޺��q�"��S�V#_���D�f���,����uMBm ������4H����Uc%/��W�OF�[�bBec�p�tM���(�~��/w�/5�3%̝����c1}�"� φٔSEgS��v�RB�/�rU����ȁ�$*�����=�P��g��3��f|�w)�?�/��	�tZ��j��kJ��y�����o�a-�*�_)�X�r��8q^r�E��/:�U�TZ)��䢚+
&�4ɬ$m\ �_��������0�+�h�ImT��շa���2��7ɽ!Z�篑�ó��Z	���0�F�����C<�7���/����[}�]��o�2FsG@a�}7�bC�%g�V�5��N#��1Z2�߈����7K��	�:�O��FQ&k���x�{��P5)Z�_-������Z�8�5#���F�RF��B3bO K�ȈI	{�:'{>����m�'�Y��Ap����Ub�q�J���3�b�K�x���i�#�{�G����M�����d|��p���Cd�������B�"�U������(�[|����t��M�ZrM�ٱSD��u����u�p";�x$-�ѶċK���X2G�l˧�aT�IOv�< ���m9�[_�/���jA�� woHg�<�40�dgSf�g�^m%��~J滫�<���8�P7,
`��dv<�a�CFY�P�q�(�R	�=������2�{?���OL�9��b8���"�3'x�=Nt|���� j[��������E {\�����e$w��Tn���O��?�5r�g �<7����]x����x��Z#�J�x��E���2�:b9`V��GY�.*��ՙ�N��𾼵��:�Y\$^�P�B�����b4�wdF��g��r�V��q��6��ڡ�@�L����.~����v{1-ʹ�&���h*U���-�a����|k���;�&��j�q����y����T��8+F���5�c����\�z4���&vL6i�S<d�1�:�9�����u�b&���KX�������z�r����;�ݪZp���@S��Z�^�wI�����z�e�<����(�Jz��y��� '�Y2;�s;��i5��c�S�F.��K��2�3@�f{$�X�^��s�����X���WsR��c�S��ezul���utSNb��jd ͧ�:��X՞E�?>6��e��[��Wf+�(�X�O��!���\'��-ˠ����ѭP��A����~��Eau$�=��5$���Mq��n��,2�?g�QI���=	���[Z����t�#�~(�X	��4Q)�C�`�ϣ���Vm4 .'��B��p�L���b�Ix����7�y[^f����� �ÐD��\�3�T\�|F��#6T��L�{�ZPo�7�Z�%��zT�+\�^�d��S����Oo�r��sJ�?�L|��Ay&�S��,�$yƑS)��S�Ͳ�����:P����t=�KB�.E���_\�Z���5Q�Ԏ��װD%��e�����ٯ ހf�?����@���+�^H��HDY�rE5�fW�K(=ܿDǝ�p*�jh�s[�ko'�h�=�B[䰽N G�{�|`�ي/�'�3ߢ�z��ǉ�ھ^�5}����4Z��ܜvɽ��;�̜��P�����^b�*�y�j:��
��;��@UA+R�'�O�&JnL�c$�B�x�)'�i�^Vޤ�&��\��Qt�C����ֻ�	�/Q�����3����?D�:�A+�<�T�q��10�&7`�ő��qt�ܽ���g����Y�W2o)T⻏	��>�C1k���VJ� �|����