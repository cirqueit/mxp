XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���n v�ڶ7U~�g̍k��f�V���j5�p���	�Uh���?�ȏD�� �r{�l��21A#��`�[8�|��͞r�1���c��k�{����lz���>"s=~��d)�ڴy�e��۳�z��S��]�[��+:��+���dF5�%�9�W>P��f�%]�r�'f��e�.��mR@�N��j�:�B �ej>ă��o��j#��[q��%�ܥ@� ����B�F@���"1�lv�i�hU�X�=*�3ߧ`�LK�c�'V�g	�CG�Q��HK�=qT��sa� (�kj+,����1
mae����b����>�E�a��ꪦ�S�&X�l�):�p�������ݛ\0ux������	�'-�L>�QWn��r�fp��ܭhe�x"���d�d�*N�9W�_Cl!�%޽�Z��NZ�\�Δȸ6u��w`4�X���C�|4a����4� �����}�?rm�"r:ʉ�Xq�m���FB&������B	F�5����L(�~'��y�x>� �#�
�᪵r�NIt�M��~��t��ꪊ�����;39<T�o.���$n���1~s��M2�߯S��]u�C����{�W~T�/S F9n�����D��7��S>"&I�C@E��sOG��ѐ��6G�j'���J�i1��j���lh��wvģ��g�2��C���m�9�qA|] �ݾ�#������%a����[I�랋�IWx�B�̍��XlxVHYEB     400     180����m��5L���o:�� �!D���DVɺ/v�uH:K��0D�-��MX�e�7��&h_)�յ�t�X:{4���4��o PO�B�,}�3r?"�s�]���1��3�f�&!q`�81�d�;-��!!�%O�%^\����Q�Z��m8$�ѓqQL�´N���t_�{BMp?�Q�Xx� �N�$��	#CtҎ���*m2������pHPb���F��\=�J�Ш��
4\�Nh��0+7!�*�f�wԢ��$!B/�cBGa��#��W��s�p�<� �& -A�O�M(��S�ŐUy���zbq#�V�h;>z�@�Nz�����s�-��c��_�M>\#���<�sϪ#|xS��OL8�z%�.�k������[��XlxVHYEB     400     160�Y� �.�e4�~��<v���w���(2��C���;��:�+=ڿc@��ʭ���HOC�?A�+Ӗ�;�XOV�(�I$��d¯�B��߲�K%Ed������zn�l�)��%ewb\�u�5i8�>*1�`
 ���fr0����K��Ur�M,"ze�0�Ta�ң�����~�!���k�:2E���D&��]B��{��+�o'�2b�#���r��}��m
���\��j\����nB�jF�Z�	�1b�N��������3�fMUW`�z���5�/}C���W�i��>��Ԁ�Þ��|�����H4	�S�����E
M�Y��|�Ֆ�p��BpXlxVHYEB     400      a0vW�}�[L��ۦ�7E���ء�dM<?�Z8��)7��G�b_���f*>��b v����zOė��M��L?a~
�3��z��*���a/iR?>]^5�y2/)�`x�u{�����t�f�(v$bm�צOfu���&����s�N
��`g��XlxVHYEB     400     120uk�!;Yd�+��dB�[��}J���[�#�����e�AN��OS�;M���S�j@�Ӱ2(�\&'g�,C{��w?%σ(��?˂��쓼t8���2E�#�0�2�6""�|�6ǜS)��q�qa�.��|n�W��mv�<,^��������c��=�'�<����7/b�7�]�Y�ƒ����j�IQ��q�?XH�ڳ��`U6t�D�Ѳ�"�����:�M����;1$���t��B�	6�P���V�8�P� T룧9p6E�wma�ߖ�Q̕ �XlxVHYEB     400     110@�ҙ�L�i�8�F�_bW&�q�X�ƀ%��$e^$�-绳�_lvXƟ�H�	��7�o�a���v������~U�i�a&M��S~U��X�@�����Kg��|d����L�V�%L�<�s�h%��sߊqԸ�`��F3nJ7�eu��\̐-�I�3����27�=�)��������<��%?e�"�ߎ,����s���V�"��Me�{"x�2Q����`)qѼ�B��VVmĄ ո�u��<��U��V�ٺOb	"e���-:�XlxVHYEB     400     130@7��M-*�,�)ẻ��[���e�Z-D.n,� �����5��rQn�@�[O�����hYB��P�W�E���>�B�KJg����A��}踝����Y����I�:�_�Fad+I�7;�Z�{��V��S˶�a}�T3������׍�[S�tkBf�yZB4�=WSm�	`1���S�[�z�=����@�ເA���o -,=��-����#6���Y���1�X�	�i�rկ���M>v'�g�8=��EV.��1��$��>g��lK�\��+~�)<u�\�d>64�ض$��XlxVHYEB     400     130<��l�9��LO��C\"F�NaЂ)U�d�!O�^p�k�J�u{f?CCk/��^����`��&��,�J���y�N�(l%��u�.�3��*xG;�h� ����D�@ISO�]܅i�u�t�o6�\�f���z������p���I�Z��wh�l9�ը	��\qqV/�@ڼ��Al� ��	�� �E�fKABQ6n?<�v[X07|ފn�E#�5f%Z<a��q�y��]��Γ&߫�d��/�?a�<q)K;*��NqN�q�C��h�D���[V��j��96M�y��@�XlxVHYEB     400     120�����	BF�i�O��˞�ޠv_*��i�r�C�)��X.�X̘����,'UKv{�3��vKs�a��#�Kl�&���b�����o�>�w�²;��
� Y~�|�՟�f�N����D�*�����Cۄ�>���M��W:�'+?�]�y�nW���\��.ΎhD�|�9f����v�~?��9���Q�87�+��~�'��^��:�n5�ޱ��k��.��!�s/�d|g���[mALO�8��e���_+�'��C裩֖���<n����v�B�XlxVHYEB     3a6     180���<�QS	�p-<���F^�`&x	�U�a�(��u5j���3��;S/�����>�u�7���Q�ji�Z��1����7e�9dE���>.����uƼo��Q ��Y`"%^�3�����[��خ6�g������Ex��Z��)'��C���wI�#(�|��%u�z��u���݊��k�+���H���z�>�X<1��2и��`���e�d�oa�٭�*	)c�k����X�Ρ^�����t:�zI�����bb�?�8�P�G缴�Ф&g�����ϭ[Sa0�j9�QOS^$�mG&��:�\� ?Pk��y�x��M�!�KEB�k�>�uU�9�07V
|1���)�e��n�jK9�+�kZ��!�k�