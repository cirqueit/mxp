XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<��wѩu���[�^9��žu��zәAkZ������2����,�����" "�dQQ_�
���ݷ�yC�����������@���&�ѓI�k/ʱ /j�Y��U,�q�@1I4=��AQ��4f��i�5>	�^�|;M����ѱX��M��Ig�F�L.���u��U�ٷ�w:��Mfjs�Tl�dG����^���{��,��y�v����dR����~�Pk_��02I�L�;_f�+��1_��W����� ���O�De�^�H,��$��x���|��6�$s�D��@�Pp��8/O�Kb���-�z<�z��/�G�œ���ON�ל-�"�� �;A��BR���w��0�M�1ϡ�9�iyFWd��a��Qc"[9C
\_	��黐>�l~/~&(���#��-m!����]I(��cQ��*�dX&-����qAX��[�qr市�������oLf��,�*�>D'����R�	����D��3pà���x6߮��$`&�0���s�+}2B��Gg�����2$W��)�)w��C�i�x��Is�����^�ZP��5&&5�� i��K��*���fx[#�y0��w6���)�
�+(u4�	ѻnT��4@,l���?��E1g�z,��F���~�c��BemzV��a���q}��DD����3N�pifR�N+��st���R<v`_��ߟ���Si��/�w����<u���p���P�XlxVHYEB     400     190�>Y~�;WOu�4Jc ���Nȏ��X*�%Q.��]yj��ݬ���[y��j�#kI� ��KЈ@@m>�R	���tO4��[pQ�@/7�^�W�/���A
�������8F(�N��6��0�l��͑$-iL�YM�%�A�ɤ�1����J8��	��K4��DL��)W�E�Fu5+� �JF�lg��nP�]��w�cK�a����>��,h������
�W��'}4Y9to�ǔ���}� ��±�����Ŋm����?�\z��۴?v'�kT��A�?��yO ��8Pȁ����I ^��)1�FKp獺u�ս��٣rt�[�Q�a� �1�-� K0bHF�ǼV��3�g�u��?�˰���P�F�p��Y%&|3���XlxVHYEB     400      b0�=4*E�-�_����O'~+�'`�L�f���Ǻa��#��8�+��GCg�6S���`,�V���sS�k�����Q�w;��SD�Y�Ew���CC3R]����_Z�%�eSݢ?E/܌{ڽ����S�`�˝� f����N�}x񛪺���Y�ƹ�Փ �n��ԏOXlxVHYEB     400      f0�z��AR�ۄ����6�L�%%`��;2|��^#��A��UqF;Rł��Ě���_2ڱ��$;U\m�u��lCf�� e�ֳ�@}���
z���]�1)��a�믶	v7��,��r8ҩ�ْc���:���[��6�ȳ<�~��'�SC�2u�wGvJ��OWU& ���e�e.�P��G-����z�X��)��Hm�-��6���C�O���R��D��g����q1C����S�XlxVHYEB     400     150�)O7�,۟����&�:wT�ś&���6;�����=L~����XS:�}�uߪ�)�-�r߼��]�^H��Q��N9��p�$d2v��)T
��?搧��`�=;��P�H6<!����V��h�Ry�<����֋���G��{�l(�c+X%�ܒh�i����\���Ғ�|��r�7rO�#�4	m�'j����%�xK���V��/��_��@2�PT�/Ӿ�>�j�K�(��QYqz�!E�+͇���P��vЩB:TI�L����M�٘.d3F��9�V�9�!:~�vɖ¼#x�M�P��>��:7_f�s��:�{����̏!27�����XlxVHYEB     400     160 �x7�l�S<	���;\ŕ>������mIL����������Al�J�7���fD|���ʂ����s�y�g�GO�x�m��R�0I�GsH�<(~Z6x0����Pe�����<�@l�6�8�nT�|�^n���rr��cn�m�<�e���/��y��P�v�c����=v,�%J^��۶��D��T�G���� ]-Fޣ�,$[���4P`�,�HV�����k�a|�F|O�-��r@Vf�K�v�!���-�o��S�|$T��AI%�`�)d�
�Xփ=o^�ߌ�b�OY�f�D8xx���`,2��I�>���+5z�"3s���N�yXlxVHYEB     400     120��!9�ե�����xw�ϔ���5�;�*�@nn|66hG��]N� �{j[`��f�Y.B�10�p�,�<P �9-�O�����a�b�a#[�1�)��1+���p
H鳐�KE�\��{M���=^���L�Y1����G�6Ě뉃x��3zƎa�]'��Y�!R�&m@�쉓N������!�t`ݬ˻�R�`�W;�Y"C�������"�j��4��,��um�8�iT�M ��22�M��D�}�zkix���\���!xo\���V6���3jCpXlxVHYEB     400     110�'7�¤�<��]�q�جS2N5�\�'�:E�F?L7;�I���bvqU�V�b4��Sd��ӏ�p�J/
e�,-#�e�����gF���:���c%&	�Q�z�0i�G�XQ�#૸����̸1	�������uج��;X+��|�n��璸T�[�8|	��)
K����`�x�3�2e����[�#�{�˨]A��]���|�Z۟býK�_��dmk�g�:�k��8��IU��)m��@��U��*�����|#��D�ɴ{�2S����XlxVHYEB     400     110��qz�~�7,���<���gg�A���g?���s��Vv�&P	lR�}�:�2_�"
4\5�I������A�R��\A8�ؙ&���,�_.�c����؊�$y�"i+�!D����%��/���\�{m��S���g�JO�F7���T��/ȩ����H��HHY��X���G�u�L��v{�ryY]��_2�����R���Rl����[r�8��b�Wu�*���KA��3�~� K��j �,� �����ߎ�&��8XlxVHYEB     400     130��-��>A���$��*����EQy�*��o'�b@Soe�F2��V�Ø��@�����u�����g�m��r��I.Tȹ���䩸[�>��Y�)�o$$����K��F�m�2�L���K�y��l3`i����X��Z��`�Xz�R�^�D���Cʪ7���S~��!�6/K�b��S���Eb��cմ�Q9(�(c���:�. ��蛣�u����eM�0F�|��J\{�{���3���+�*\_���N��X���k�@i�Z�����m����	���]�XlxVHYEB     400     140g�t���8_ي>�!�)�[�eʕ
��1k[�g d��YteB{=�A߭��i ꠯��L����wܑ&el��I���'Rl?���G Ru��m���zÑ����N�Kɑ���:���,Ӭ1��7
�C���YݯJDL~߁�Nk���}��Кu����G���}%�W����փ�ra���1������	9�ά<G��!l���w�ʾ����f�=sf?nqc|s8�;���σt������U:j�<��d��5�y2�P'-�qZ��#���厧,y[��/-7j�����C ��K��fvڅ�f��:��&A�9���*XlxVHYEB     400     100rXO���h�����S�P��̢� T�Q?���oi�V[ƠH�7��(	�joe�(���Xv;[ ˆ#r��j�C�r�4������z>�M!�X�2���Um#(�{�&g�<�ځ���d���ՙ �a���i��~S~+=T�WwO���x�@��v�WID��X�r@��t���DW�[�^��>�t�'|Pd�����F._��ij+���zܡ���ESC�d~S+v� K����0�@�AXlxVHYEB     37b     140��d��a���c�ʨ#���8��y�����XM����Ch��n
#��d�>���;��uU�Ͽι��t��IY�Nd��IF|��v��%QP�m}��9J�*m�٢8V� ��K�P���&��#$��Wj}�����l2�x��a�0B<�'��!9�����-�U�=�;��B�5�������vie���ZP�%Y��t��%�P1�T�SYU7�c�R�8e:�	���P��^N	���A���֖�q�����ZU��A��ʢI���	��,�o����x�O[�6�_�R��&7(�3�)�G��m�