`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2448)
`protect data_block
OuJ3PgCf48Jojb79rWrD335a4qwoQHbNqaZ3XDkhqn0jzZkzIqJOwIMhKnYB/pN6YA9/PdLTtkif
dwvoV4plJupGq7UGpnJhz/ULFc/5SF3+ajeE1QHJmL0ujGNjtkm6TXvSC9DzBCyQB0QqneJpN7Wk
qFiyUPJ3EXrJqSAQQUj1/OZL+o0CJ2lqEJmeSofwZYl5lCaTIRytJzFYlpGEcVF7gem7X3RffEf3
EKg0V1YORBq6CnBlG8m3NGup3I3sdrdyhZd5N7GnqLoyY8tzN2CiPkn25WsHsqNeCZzN2w27fmTn
xcnPcBAxcTFCj8QWWYH9iCu+By6gE43JKNCh3Fd9rTmqYotwy57xn+2xj1+7HvE/x7Au7sbnu9sJ
CadDUlHRufso8kqfb4tcaAoXSZrSgN8AxLUcwO3XrPQKXeORMoyKN9ka8zdtQNZSgGECgsG2U28o
dXAae9F0SwQ5sTu3nlWLHycFfgEWCNhKKBSPUJ6STgl4YKnEmxuQL4zcDU1ifYmaB9/g1CEKck8Y
UzNXTf3kDDjPAaibwUeOBNu2TCS26oF0IVQJS44/gZjFf5ybZEeVrYd+DAQY85znDrvOsvkqAYeo
RVnZ4Q3cxX06YI4UvBwQeilctdJe5Df03oxZPYmAoLhIlHUbaEVzgP4AO87D8qx0Dh7p57u6ypsX
dcdoFvWAYVBMnljE1I6zOKQHq99DMdwGjMMK2lrPDSjy9FzS8lLqoK9HjHqitJD7yGg513ZntoQk
Flw6ZbcLTu8+uYQkGeqnizicLH9Fbuw7tZjf3IFn4L1W9SlcgtPpjpfObrk17N9+alarO6JU3+T5
JWQZyJKTS4D7ag5B9z5OjRsSISV9HInA1WdzPuXkuIT/lzxYjkFrd8KJqSJ/3eQ61iSO/rBoSY6D
aPUAzxkKm6gRKDnqy1fGUjZvo0Gsuaf7gS52nyLd2Yhv2p1s7blC9f5jTVLXeDd0NRbkLTgXMznd
k3ykS4iX3dg6aIuNUZdSk36wehuprxB28AwFFRzftPCkFxosciHcxdFeHM7sgzD5Do/yQuTnkRxv
ayzNvUfRyn1SzbHDMq9lE/8K5oOPo0grw6SAvWVQdv2UtaPZRg4nEPL7hsIZRrVUh4jaw+mg522L
smomviSUqdHgx1SR8Tzr6zG02yP+tvWAk1XchephLWabjwQgaPAK5K5Prc0Qq4H8EYs4I7MOWDB5
MD3ijANzegrzgpzYtTQqin0mRD6H0aMSqdElYxGIYcr97o0iG/S1GZMEmMTmGAE/fcxRcxictLQ9
JgoqH/fzbKmdpypMYUC+ZSkHJUB3AgbLZSLsKEfY1KRAjdcbVW1DJIO7TfYHgtkKjGLJK/1puR6w
86TW8soM/Hj2YizLUHQP42VqJ1nhm8Y5lYB1fkddNSzRPvxrZYsAl09PJWOPECAlhF8Yx80bLQf5
UwXVPW8i9vZbPrhuDZK1d/9TbHg7uweyOM7UXtcGX8oysXsAmUgNhkVGzdkfN0rqOSugU6ev/vY9
6LuWJ7HQGd9lDOVeMSHQsALZxsRApZ9gldHThmr47jcoTELxnyDTkB7x3nbWaKL+0aHp6ckCxoAH
WDPPjH9GoPq4le1cGt97dR58+s0bg3f/zCMCITeahfejtCGkyWp8nHM9/FpilEbCbRa+XAnF9bBH
braMOy6FbbsAqpUhswOpM1DfhvFgG6mwONzfOQ5Opt9qT+lFCuXVIyJNJ2Fn/E3MIsUqEIy3PYtv
nwzUkDRufT7JMb1b/6oTuBb1zsRKZxeDw/H3ZwRKab59H+PPsz7FJcif8sFB7fw0mOD38kEDVcWH
eMy1qUeXLQJKWnCjFpY10dLcIXxf7M0HnlXjPKDGcqrJD5cEvIHRDqHMrPcxkOkeqXcNXiXPf4Uy
2i/LZGvz8Bj60V7dzRZDbpvtAJx2o8hXumBGQ+GN9CpLNEs0CbWXqxgcY33kK2e2jsP4Y5+T3pnD
EpfDtk+vz2flkvPg0uWL30cKdLR8K7PnKvT3sa9kx9sC+XenkkLe72oh3e1gNI0rD/9eSR4tZhRq
0d3j5xM/pm4123u6IH8XurRbdLFkNHNxtr5USTVj8K4qvQ6YphzSFvLmynWNT6c2CjDufmS/J48d
+vHCdP9uRKsvwnVQKmAQSdNdPU2N95VMqg8G3Bsp4u0+80ktJkuKqbgY4jQAXRuZr+RDLBuXfap9
vu5gp4q/UT+0TL8aS9Sq29lStzlHOzKWoKe1PeXE2SxtgVEkLi/c7EVJZNpK+HMQ7kYTezavad6g
Y+SHDRZe/qDvGx2Hz5EqRetQ3l0DtRO8bUWNbmEUpnreqt2oEQ0JJRRRDuC9VE+UYUQmPYIoRzfQ
fD6c4XsaK+/931KPwCBGjA9gTbkygXLgdhckPawtkCZGvAZCb4o37WEcozDdlvGmWQdSXyS/MZ7a
JFtFk+hqpVsaIoiELLvUDyCAmhyo8cVsaRW6Venc2x0mH2kNi5qdn2tNMHu+J2CTmQqthdgGjH7c
RIMFSGdVCFIpwUhwNiz1tOmXmqQdiOnIUOxKWJiW9E8jlSagzfkqOSG0yo8BbHN42Wzv+yHYPiZd
NMEeqA/9OgT/TMs2fkPnaVV+xoJxXVU5Ep+60q1JdrRu3Aa1ACXBmljerZmerA/sNoUcOSYp7NVF
A2CFjHLyFa1tZ0wiOh5jlKVtkA7gasv1emPStMGOb/aOq4MjPNEWnSiu1guy7Y6ybrBjnDIgxRc+
HwxEfGs0dN+095QrVLaATKE+rXA/d09A2KRZ1HWtCikrVNPmBmFwIlKUcOIa/rksQfqor/yJDlqU
LPOfCslPQ9HpL25ZbU6MaG26Km0Vsj6dHNpvK1exKdhl7Jjb6txLw0D1zJZqZtuaFahBqFBDpHfR
/4BtX42pqRaBuhSKbD12fVytxxicQQ0yRQxyo93knbANpL4HpQw6ybpXyX2p45hquTOrSVvD9UKu
on5nhW9jesRtZLJdEIHS+r1m4XQ6Kt5jWo9RoRZA0If98Sy857ZTGiPK7RrAT4SV3/iMW3vaLAjc
12KbSfdGO51DIghe+fK3p+HSITkDzLWQNsjItRDYcFMgLN3AXTSOVCrEjp2uLhPpFgPg5cFXmwva
PmikrJ2fM4gHNy0W+brHCYVsq328d3nP6Cfq1RJRU8FkpTNcUynbitLTk+Sowm+1DxixKeleVBgF
rPCzz0n1+vxLDnavsDdCHOlB5egnPdhiNVk5xA0UrgQV1+FxfzeZNOI+ggd0k3eH0yrUDcN4
`protect end_protected
