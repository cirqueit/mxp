`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
fzppoi9uTuJYXyrqjF9uW10plzLzx3oyhKctrsK8BFUxe3zH0bdf8z9UWvzrQf9Smpj8nAwzGZQ5
1t+5d3oal7zvQRnuuIGV1OqpCQweSrU5gTkt1yj4Xe9zHGlRfviMdJcO+2MMr2g/egS5LZdcf65R
91eFAmmNOy8rarUpB3TNADHEBknp0H7npMLBsAOJQcm9eYChXWIjlLywupOrWPIE60UYWEMVt+KO
8JmGDmrlikziYMgn7kxkn9ej+pQ7iHtinNTuGjgXFA6suNwjr6sO+sgU/Kmhuim1521VzsdhG+Xw
pfSOkmzNYTUy8ea8LNYMCwlY+HuY9n8Ot6CdRGa2IRcovIRT5R6oh0x2yar1cjH2QrfkKxINCHV0
KiXPBFUcD/Qr23gp/WUPe38tJEZ7pwfthLyeWj7M0TzlpQ6c1sHCMkfYoZTIJ/p4nLw7SMnZTY72
aL8IFA8YRnvxq9xfpmvbupI8KZo5mD/UbB2DcjS8hIN2+9gpa5wsz8JrFJegMWGkfDlxRq03edjq
dN0Tmo/mT9fZhof7vc7k6358GtxxW82uq+Pr7504LPttPqnejLPe2LAtrB6iqJLnZsXN/7yv03TZ
AXdwn0+MhsG2cmL3RbAGx8EAIz+xzVtdI6u/2LxOH31P3DzNSMh/WnSbxWq9QEGGDmjWJGeR7vrK
zUhQUVVKXNU1ja+fdMYVbe/2GSPO3X4vgFoX7mCwZaAkobqB8fdrhCAuFKYSmkbNR0tK+I2tl8h6
nfnLpy0QnaPKLlehC+1KC1J8cqI4cTvadrWh5ladtkdE506LMyCIYZzsMDh3w5KvLZ31JNhGCNoL
JEjHvOVTgIQVPsJC+PIchMoR8IdaJ4hkuXu0GPvArmWpVAD29q5nlM7tnlQykxhMmUP/mDELRtVj
qodvoJI9wl1j3ByWZhkg0vOAqxWEuYuuJO+rez+UtfO7B71gF7QxL9e444iZp47a/iKyQAWOuK1U
o8i+duzoq067GNrlvn47qfhhsBeMXyX1tQLpri+g4wtWG4ZNAitPtwUBoe5GSUYDlR8T1ICBvnPh
jXqraS0Tc+novH/tlsQO9ZFFvY41OcQZAcYpBogVJ1n75lv4wHR/aMYVk0obZst8xHC1PDuXfpcg
bEXfR8YDGVqW25aGNRGL6CmF2RhpzvFnhisPnvqrZdlzyuYdDl2kR9OQTDHHe0ZLv+NnqrEnMfVH
CBPSp0hLo10LeEhiTIvVvizR7sT5/ZmlgFT5dKbcucAdt3aat3osTFpZR5TNGvQX0lICAOztTeut
pLTZ9UMu46Ma6KLWTBhc0fDaT57jmIS6N7RxD7uVqRgzlwbEowGWqGtCnYWHn5AP5xzFWp57nd9Q
dOuddiSnC/jRE4pxc0M4q2WdkC/eCClnEZzX1dRXeD13InvsKdwdRmOZdPatVJ0Cup0DKoIq2pdZ
FZ8NVzOzg8wTE+RBdbN9aTB8Q7yBV7G48azToLBluMLl7dk+qyawokWyfU0BiUcWOAunp7fv/pTi
ANzyECSikoID0qvGArWdq1zHSx8CUtvhOdQS7zIR6lReyelyXNCg82qY150lF8hLjglpwtVm04+A
GCwdaeOkyp7JM8ADcdws12e7NdpCuNewb+omq2wK/AHaY+jnJoQ2lw2ToMK2dfKmx57cv8QX3VBq
erbdVir3CqoxsMfYDz9xZ0x1mgVZ32+VpcFI4R3iTzyT6rt5rNCRqDmvHwU0Ke4KTxshcMbwUJWp
MIRPEdxzH7kc3N5jiooSzdk1UZyTWBg9IjSecygRM0qnDhv6g5F653hb2hPGk8N8hpEFNodrjOjz
RxHzMcbvPTpOijLufArdgZCL5NJN9+VO+0aXpXrlpUKybwlAK2s1spHJwVv8Oabna+Wen3An2nq/
RwRWWeyNbYybH47qhKhR0y+VTKFDDHQl+MsijtVB2Zi9otdFe+9LQ6MwqR4Zc3MM7wF4u/YHP282
X81lE3/moxRY8zBwY4jS7GWV7+3Y2h3gjytlRO2GV6QlKNwlKaE1eitqy5jllhe75lxfksbZRYpZ
A30xPmgGkKsIexG4ZL2eq28uEYassrOsX7JiIYAQHHvoI0uyp/GY5yS3u5+tZkPH3w4ddys306ia
HA4O7egzSq56El2l0C/RUbl4XGQXa7+x996JKBYNTs33D4oEfie7f/kd2yilOELX2EARg1T4Eu7i
ebkgwubosTnBcvOJ3fLKXbx8UOz1dArNzphT6W7fL+2Ku3us9VH5YNzVExVUelsRZWl7AhcZj/ue
HtkKCn8yFLjwmN28y7FCe5AcF3XKKuQeEftV29/pjdDPJh+YKP+EKQa6YISZtK12vErCbYe7YUkr
YigTkWsb6457PfYktHzVC3lNLGlL0TOpeXMxxwbUfayk4hnRrG8hiS8BCXTYyqFfBDuttFjw3Ncp
k6SRBUPex/WYX/h9NmLdP6qaIjuT5PQ3uupYrrbWCD6CkbcqQKtOtJb5FcmJ+Ee0Ta+0ic1YZeke
+bMfNC+U36oTz5h01T6npRKJ3vf5/X++XzMnForcgrvUfF0QXwJnjSvrcT5UUFdceBz6pqHs9Y8h
jcJRgWB2SN+In3fW9fHg+Lkgju5gVvwggLhUzEDktLn/gry53kpgPmqRKboAGV84R0N6KiO6l4HG
TVlW0WMpEre7o0rx5NwamhMoHHZDyV3rf4fkrI6FhmlC1qVerWNBQ7WjIgmYjQXlmDI1pQb7aq1/
woqDGUjgKwISgwHFNUIKL3F1C+93j/f3mfb3QoI7G8WKx4a112GI6xv5aV5HPt1S5Tr8o4RX9AsB
JNA6yE2XoL7x3ExEwzXqDFfAWtXLDDdvkq99GjuiL1IUtxINZPU2PBe17nGA0F7JU4gUo+h6BUhi
bwENtpf4C7hE2Ls3hXU/1w3JBIxUlaZ7mMJVf+rdQHSRheyYe2rAYgpry24tqdPmkPkj2dwEuweW
TV/M+NjMQp5tK8BXDcZNqX60k7EtkgVpvm+cl10/9wm6GgbsqatrP8ooZvxE5xNvUkG9q8l3U9tx
XBpONkc7snDK0j7kaDJLnUmjSqL0jf77MWxuyJFPP77kgDgh10yIH5zFVnryVtTMEL8MzboW4E+s
esOzRNmPsyhiVV7yrdO6MCvN8suHUvvlVGdsfMPNmTBXST0bSQUrOKx8dCSq3HnH94vZYQ7z1Fn9
C81wVsWPXdGrvy+ajonWmQ6e7jXVGsz4XeFRMa9wYdJ9ief7Zm2BisnenBB6q/sOX7Ez3CqqDUar
sVRXMTjSMXuDTYZE2xJC41UZNPxTbmvXPeEtGpbNjhuJ716cjJIDN3JJOorsWG3rb+GCTOcG6xu0
Zzc7Txgs3ylw1nlpbCxaKsmIZUSjPcB8ZBSMuIHOa7wi3SUSKJaW1YfJ/zI3q+bQrYE5OHl6Jmku
WDiKqSH+NO4Z158kwkvCUqPRKDCIiWg3S251wfKpZ1Qid+Id8yUSgSsrN/5uvsNV4wdsLloBgXZc
Aeb9+1Yn4UiaZH47cX/dq/kAvE+CTuGMivHcRP8vgu8r30MldA8D57PI97BJWCftDdB9/A8wzotu
LBxRbvmb3azv/bgw/2ntG0Jp349hBsaAjPEhdjbmtqHMbNEgHVfpAf8anw4toJ7ouy59jeBOidL8
ijrN5f1+AeHN0GZPiwR2QrK4Ywsw+pftP/OVHk+RYUSgaD4np0LyHOYMNv6v+Ld5lANn3H3dazDl
QQmfzm6t2VLEp5S9m86wZ6Ivq1fw8PwnnRWJ87EdviwgIUVoBRSaL32DlNTVlb6Tiz25+GwGM6Cj
vjZMx07uUcmNx28V9W9tMT+pH6JlDaTIrGYSyWxIlxqNH/TQQF36m3eYRVoJrdOf1JFp5DuBi3G/
QiA6qz8B2sxJtF0na+oSnRuCCUDpqcSv6qcu/FsK/vXV3lUGZbyMu8Tu63WEZAg7haKa/aKoXS7C
saUUBkZIhB4NVe1FMXwGiS1vt/xj57pGf9PZCjrs3ceHAXHM9C7WJyPWz+F7qAjUNdy7OLlUrNRR
N98+uhn/Zpubf6DKUHwVoj4gF87AGVToDEvwl5wbHAf7P4KbsvIxw+Hf+ZrR84gxFAXtqYX7Hngf
wqmOWsXcKQ2mlDCUjPTNt/SlaBCb56P2mScImSW8tOPTE9a//wnaGnx1Jxi9FA4j3tfoZGGQF+Vd
cGn5US1MM8j8Em7ciDRFRG3HedpIMhJJ6jVkDXL4/nozRFjsX9UExkHD+/pDTEd6kutLuxAwyJwM
5d0hG+r+WOqhgbiMdCvoxnZBAf5SeB0dkMc9y8O24JxBBvtzKw5X52fxMidmduhTrJmUbVEPSc23
4fjiPSlSGDOHtQb9wdPgjPWIjor42Yv7eu0HX21YYLCUQyxe+dTM3xElnS/lAB0xf5kcLmicBdBB
GQ8Ja/bc7HXcbi1sbCj/fhfPB/PutpR60jeQzZWorZD+UlVhegC57v91fc87Ca94dmQwIWu4j80U
Q6/5l0DeKJRLcF48Cb4RDiFWS2CWd4sgci8t/uOpmVabUKERsMidbrh5JZEn35isO4cf7I4qzNWd
qnZDozILpQeBy022j18DIzfYNt68uYaLxsvB6bmE9Ur0Z+cIuoJ+hD9u2PVJgcvl2bPHTSUtRHb/
ze3Akj/cFqFRkFNg6Brk2ik9fKLGI96ARiOI2c+Utzlz+78YOPLNSOpXsuuMJDXYIo19uW+8r+U2
BvFt8guQSMPJWIkxRQE6OLfgBW6FPXw2U0YfLvoHKOqEXBCIauHE41z93H96vgUEeZ/i6OckcTwK
n6IbEbjIpWmBT/NhgLhLcxXPfdHiysuoIFyf3ripPF6c6Jli8zY4mTdXkPXOq0oiv/aogz/sBqAF
owZfmWyvid8NtISowh6gbojhnQ5YCmpAI9x3A8w1RL/HiH8ZxmBAzYT75yptXuo/LmhsX2bWS2bX
FQtrOTC6Ajcr9J6+oljPTmUS2LclJom101orks5+rXrOv38tMvmdeDr7EDiDle+5CG18S26HQJt6
7lGwfSRoj8xbtggGkGnl39YfthFrXrnDBUn8LitAX8N2gdPfPX4VEzTjTjq/ZnP3U17AErfeFb78
hN6zinK66E7myN0GcO5SMiyJupRwXP7EG5wy/IAYUINoPmc2/00AKRDSXVGZcU2A1e40WC/+MRk/
iRzf8pBJZH+eqagyPwBoAqLo3gL6HIzXLhw0Ryf2SqVW3AtKHoR4OlpcaTBm9GAerrOZFNNj21ON
p0WSL4s3HsLUY2ItEUXIqTOetwYufGWotW2FbIdJVATcIqcUdPK1M6euUN2STRFBHn3t3qq+FDmw
xuqeJmOP7sf9Z4V9wso69d/jyimOWruKxuCrcBnG+gSOOm8O6iZpdj5oUoBPYAapUbSDbRWBqcVX
oXZP4oHF6l3wAalTx2bUPnCNjdgn8ZKieQun2Nt2aHEGPI37bbI15G1lUT4qBAJTUFhzSv7SVVwf
QWenpIMmoeG4DMrV5wzDTlr1ECLdiiCCg5Ugm76HdPj+/yOZzqfP5eAdV4ocOWxOvJdNcyTrX5ZO
+LO51Xw8cD1LLcgMOEin8VCerNPElYXmI7Kl8YhmzTJpjHV83EzlpUY48wUY366cfUuA8FBnNt/x
nzVBd90VaVpwOwDuloQTYPeSCeqxa7mm8i30KId0J/JqcaarPwillD4m1eUtNubY4USpGwDap/Tc
9oXYHnnCnPImWc1M3A6A+d3QtFAFOnijBn3Z+SJd6vYOpQwSxrFZ6kad7vJy5mIJllQ2fjf0yW2A
AwTqodamHG4lWV0cJ2yS7h5pkTme7S8R0dLNOtcK/YEGKV7AhwrCnPNHIyyAWM4fVNolCEx7+SF0
dGTtAMPoqBwMqeksTMzLNdMxwLyVJGga/NQ2rXYs5mzcSVY0JVqtBlcFh5xex6PdQ/C7h+u7JnL/
73mKo2JIr/jlYPbraQNiOGSObsipOdSIgQCEXS3tuSIffRw7Oeli55by77qUznFfZkRAl7kfAQ4b
SLF0G7Upygb3NdE8rImAkCgMrV4ohEP3HiNYG/NDL/XaAxInWfXnM2Ere/EgATNA2Ni1gNZfpjXQ
KN7JbUdEhKT3PLBoAAlWumcM2XbMZ24f9C11gkzSUofVRoqTAKpKMImtGIGAHeibP5PDfwnZrksy
rRkLnXFFfbxTN+SdLY/HJrl8UJaFbjqd9GZjusTfjc1jfwo0Kowp8LRc/UMlS6a80ivB7axgceAy
yu0jEqBVnzMrbrh3TsRIuN6MENbgj/h9cs2i5jLXkRn76I8X0gDYP4Vf05e5a5OX0gb0hZoSlI6h
BUZQkP15aw5yXL56fSx8M+rXVES0DXdqECPbRxe6ub1L9ddLOuTz1hxsVD0gzUgHXPXVOQjQ5pYH
6+a/vPuZcIZXR/brjfoOzXfqNxcw44YgVZ3T307mq7E+MIE2vBFqZW3eLAwmVXXEymhr9BnW/5R7
uq50X7dOutiZ16kfmaAVTWK32J/qmFW+6pb3nxwUNR+CblCwTCqCVYqFKGZNkvTqCE7oUvP6sPQr
6ePIMQxY3Vn+gOhP/+FkgQWfnC5nB14ttFZEkcQ/yxdflrQ0SpLkTT8iyS+JGMQ2jj89fixKJksD
WAl8UjgRuuR4loPVKiElAXuWzxW3KAWUm4iV2zr/i/7CbvS/1M46oG2gt/umYsng6KOSGGnHmnE4
tChSxWJJIAdoQRTiIsSVFHbOPX4n+Ef3IvAXnF9iigxo+jdKkfqY1yqLrC0Dy7CUvV+K37G03KLi
WaOXL5/ROhQZMzjCDsjqx50AukdZ1tWfGYqzNW1cZQih7ul9DlaiSUZdloxCwfMZVvOA4ohIXOwd
FzlbBvr9htVmvteLr+aQOt6M2NquBElXQHkZgybxv+DTOalINHe2PvoD+Hg4oukBcYl8vgXvqsx6
0cvRoNKSRtr4ZcV4NSvMXaALku3RqsrcD+GpNs/qvYhtfd7HWu/1n/5jVB+h0uhTACMdqx803Qo/
4c4QUEpwk5aB0qVs5usDDjwcRnt4jTBsgH9+Herf7gVW3ClbKa86Tdj/AhXMr5lQXObqQx0GGFLc
3l8QPqFJ6iRhaG82XXwD2yAK4o3aOGYcgn4kjEMBALVmplfIgmWaaSmmeUptVhL9hKXiGODII8vB
frRwwAs1OnPeMeAZmIRI2RF4TgNuwQ0uMYrsuIaHtPPw2iz4CoqoIml9N0he30F7j5jBZw2aO+45
B+gA3zUJuLpRvJ/k7D2YliF+9td52v4+KcloRkdBmq4+2DP3TGMeffwZfH02569oOQHTvz4874T4
sMCqo6JOqQnU7jRelXy2xky/vdNbxDckgy3R+8pKGrx5oWBj2w40YX2C5Qo2WyMbLT5cjGPPdm6n
Ih0OMr8tkG5YT7QJ9Z96WS6b5G13flJsGg/o9gW0t8iYaxuuzqAMO6orop3hOHxhbBU1H4T9Z40a
/UJoMRFPYFMI4AWzjAEZDakQfeNDfLQQ5clenDyA/TLM1ZJsXT19pCzhAO5f0YFmAkX8WRmDkE4S
7mXM8M8S2vY72NWTqYrv1DElpikMQP1+TLFhTI5iWw0JD9S47O5mD5sIvpFNZbCXo6x63KT5sbAz
PMU1fFVy4lkrC0uMn3qSrcupXJBcNIY6YUqgHhgpmjbJH14hNsO7SmWGOCYxMYCemTAhskEorMeE
1iQAzw68kEj9O6ObLl8td/SI/fzf49ZONi/Mzrc06Z1LZK6f5bMvBD2nKKJAPN2TdjrcG9CVdMo7
1zJt8pUbMFjWfX/8uK6akxmtmi4vaZUVcY1MoHwcHZ2w93De2wVtBD1p93HcL2pIgTZbn6O2FMdF
whThAFHZN7yOKUjUcRhN1ciDZB4ZqvxFmW2W0VonR2KBtDSsC6i1snNrKNZ5gVc8Pvmd8gziBV/U
1hoQKNWWEYoPoIcbZ9EwzVef66Z7dCafTEl2/vXzNQr/UWu/qNfs+fa6M06tGjRdGvjLPfUax/aH
31JREOCmEILp/Jlh7DhSWPpUES6aChKnco6PpDA/xYDwh9jiIoGXFYZ9ESUR8OW61fWTCOEDuYNQ
rk8xPns13WPRn3KKDLY83sz7A80TOlW8RwrAPHYJMt9YJJm5Lra8ujKe/y6aEMK8pT7/em1j1Yyt
BvDCwp74vjw7UVaWLsosbW6cGzzkQS8uwoI8DL9r2OzR5M4dVStJ77NqL3Su5Z0ym8XgY5w7Z/hf
/JOB6vLjt/KEF9T4T3ZOWtZnD+P7TzqQdG7Q3hbY65KfsPpwDOea6sggqyDcSTjUiuAfLNzwuC4u
FU58rkIx4s1Om0gPVyVwQXmmVbBBfhfsr8iZDeXBMttK3XcKggwxtLHnUiTr6J9EaHKjXccazBue
8YdwJXwqJuLGJkHSzIAEJcy4WDXayuOqkt3dxXQVFrm2zkDYuuU4/IQ1MjEOfaNYyX15O9jxoich
PQiO+k+M1qxBRjqAIsncm+VxWezJcIx/OHAtnF8QkayBjsiwtY3sVTeqFLoQrrmW1W7baT5vtEUG
ks9qATRPJJIiLjkgrgBvUyfZ5XI8Bs+/EIHCO47RhHjhdsr10wHZ+i3kUHzzCBcd7HKZrXYQl4pp
Yb1nw/PMaKmwR0ITwLKjBXWdFKHzcaT26Wz/eRMeM8CozqyK7vhpTPPD7etQqPoKUnRUvjDmZVMd
4RmB42cbP1r/73ohMs2GEjZCPnJ99IYeFViFbdQrAoeocFb7dePZKxfFfjLXQbQpdO9t7i8bXSeZ
Pif+2JeW6T0iftjmmm+Fy+WjsK2qjGFWBQ1nfF0qMxSL5fvgiDurs8lDw1SEFhKUyVGlM4Ms6Ox/
CUjJZKjwVL4F0I22KHB9FPOMD7ncn3gDQEFy7x8pM6Xd2oXHuP/NvjCsUHOu1wdSCxwzoL3cQe5C
vEFc1vt9NMvYVmMToyPZFzw84aDO/UhQU8KfwjRusYY6kgt598yvuJmuuxm1H6NxcloquB4LXx/A
+Qok7R5O6OCxNl2KqGCQxfOrYUvjLy92MrPGW2Lumv6lTksgxI1J+NisVdZO5hOSTpacCsdyzioq
YBroWC3hDSTehv/fWdTg5NSkaTh5+AXgfMUbkkX4Yn7jIDOe0os05lHbiPjl//hAkrPrv0/HUJcX
3JKKOCEF/oIo6lZlHjEH1wA7nL7RLXq0RPXTBgk4KdgB2h7+4YI15FY7+Ku9vTJGPcRR9zJEBlLi
m04zfPlj3TTnni0UtBJ+mG0HumUIexIq1kA5jqY409lwBvRaMSIhQANA//DYSgmMRdyJMIEXGVqe
YZSxSeVzoiRnzZ1zqiJRUCqr8UCYDHz0EMiiJk6IX0MGz/nmOEfG0pL8ZZ9QUHvnrXIpmVTzQCkq
+mcqo1MPiXwMoWh41FKlbJZCvOLssOvdFGIumau9JH/HC6EwQHkd6sHStdEiIYflES9SP6ksVjN6
dO1kws6IgardmaSJkD+arNeFeRIaOPIrmt/5Gt7KhTgHWXqCq8KRzj4VhYlPCCMAZvagfPhojf2s
2QdB6ZkNcbfNMM9g7lJyKuCP6FVDPkZYgcnK6ncysI/kwGq46moglJC68o+XKJrvBzXS5FMjEWPe
He9uyjEHgjLq5BnkkLMs7K6vjLdl4gW0IQXawC5bxQoOxKl1isPyjK+/XGYpccZEjlC5/TTOTxeb
aGaVmj05gTOr+itYe85QLX4pXMQXkgRi3hl9AHjLGoNUUcJ6GwDaujEzfBRNUn1v6uanoVcye3M5
w1pgSAwYhWxzuORvg04Fffjh+H4+jZyh6Esexl6b4Zy5M8Z8gIme0kQRv5KQD4brWQ5ceatcEhvl
cBzVtBtT7ms2t6MoTndbX1JoGL+RVPWd2E6MzAO0zZhJFWSLO7zWffT/lGi0hzCpiz2PsiEjP7oH
r74HEQBMubqQwUP8m0eCCZOIrWjbMaD7Dj3w+CRUX+5bFbxqjQe9OAXrXrxoDLvKBG4U+3K9subL
B0e+COe7LTudbdPRzyWpUvhuXYFnw71KWGgAWr+fAduC9qFT14nYbPpYguTw5XlgJCPqt1T7yMxN
DubOrG+kGzsmuC752jX+bQxjQysi/ZHC89IAB3B4aSxrgulxyiu32rI/9yM5L5WBRoRSZydx6FQC
ETjYM6dqyouZ0+18I0KXiKoKCTvD5YQF/6LvMueg50soVrG4Ms6yFu2HSlemDaMKNC/AHV7BEC2E
mxOKznYvAsFjc1xaBrEXLbVCMI3IS8WrO3efvF0DcLa1hvgD9hhaSAEI9FAXiOXf9z3t/+g7ygfI
cz8XSsvUETqtuXaPrvFb8YLBe1JBPEUvnuAT2XH8wZHBmJSgRRrASt9wNmwiZbG1TtdcEuuhxGgA
bts/H68LeqQjAcI39t6vZESGB6ElaWOvnoRRtv/3v7+AbWUtZj6sAOvjNVQE8HE89AgVZYmeeC9A
6tzRWBlau9LIeFGCV7yAh6Hh3yFxuOr5Tky+Wv3d2g6phL1CKcMpEcGRO6/HA8wskyqBjD/Kb2/p
VzTvff28LCqaIwcUlPT1ezuxUeHZHybz+125MYUum1KOWajbwbkcTfo6rWGyzr68ot2Cedm05ikX
pwDtn9UARAGj/dBgPmuv0pvkijmo9YDlD2fPo7q56DtMZhqYXVkbeZvmlYyU14lo+/el79uTl4b+
WxFz9lVa5f/DQ8qMiHn5g+J/s756+TYFDYWCdKAWiAg8KFH3iXL7i+OpR2vvPrONPv2k8FSg1aYV
A3SZsSHEnWndMPo5ZVPKeag+zAGGOk15YF4OZVwCSpGOlDoIt8Sgw17lH0UF7kK/iBSPeEgivHdZ
ytqSlExOasFZBJJ0m1qkGumJJYsAtthrkqgLggrZ9QeYdWHZVt1H4LmCoK7RI3HRwqQ4Kr400R51
Rw5RtNg4sWlJqVvaFBCFmCvVvmwKYzkTUsjj63NwrmWoOMogBo0D55cGrNnV1c3I1TcyQjZCjd2D
7EkwWA/1ztBL8qPGNQtVxHrMV72+l/CleUqHHF17ByfZ0H5bKevfIBA94Ut4oWRAU2BvYV8t3dg0
9wQ0ytTAtSX6d0u7XoGpVsGaqStAwfB4lP2iaapBzH5/PYK31eTOulUC2/d1kAhaYsVtGsjdh360
1IjXImeJr+nfKDN+cso/lRjgeD3bNNDknI0DvE6PrWVJqPheoa9PWjwRI+yhfiVP9fDfS7Lp7C98
fi68+OlZS8Mg6cInx2Ptj5o4JFOrPD8bAUZZBkFcGbneHIHTIpwp8dyieE+JbEsEdQN1HsUgdLjt
WSDKD+saPhw2Ciw9+aqEvcBXvb+VmNYsySceS/iYlmgitxjj0Zby9yD8u/XB3kX0g9Sbxe2oeF/6
Kf5QeXQNcVGHYsPkQLBHrVDFBQlYM+yiRuoIBufKuLva960+GQd9yoAS6850ppn+aojHoUE3dZFW
7l4EZH3kTznRtH9CslMauSv5EDLBrI0c8QSVVdX7vHuXmUcI0/9Cbr6Hm2w9UXpil/H6JCp/0onS
sw/HN58MYSAAqcHp1YDSwclDesag7rwBvOdUIlBVzT0hUT9v0wv4bxi65A18RC4bLWYXSvFQ5HDT
eP1IES9jZ+TzTzCkwnZhUf6aIbhIBhMjzSvQP7MoZ943LVWPjpAAioy2XIUZpFWZ5Zggb1f0xkZW
AklD1JAc7JGWadO3DpuBcsR7ZQvINOzvdkee35i4QR9K//I2Y3eExt18J0MXZ3arADv3Ik8L04Q6
khqrLiCqfw56LACXT32ZjVRoCG9J8HAkU4v1yj3yQpQJpaG0Gq1Nxng4KpKSwybBn5HMDjipV5Pu
HTnvbvIFfkJM8lXsxqEnQa2dezhHsGSIXS2C/SVMRaqxu6LKXJKOTbGpth1ksMH7NKzFrWZRQsvR
dzEe/e8uVWllLxeIZXjPcBaVKhLhSfB1RrrKW1GgpvNowd+qjsHYGrbVmmKvXd5IVA8RY8+/uSer
IO3PSo35gyM3Z1JHWolVmuxcRw7AAjddxcnit9RH9KqM6n8/+P9dVPhWosymr6lQUFB8ghnzVVAf
bb1en+cs2h/BYrNebEZkiZym2jFfQE9dlKmZ4ALInO/peTlZr7mERVN/FA2IsNfgWQQyCMU/HMRG
K+D0YH0sXm2KBe/020Cf6gMRIpNy1Iunxi4hkLBsKBJzXaa2uY2iWrldWXpAuc/OofSrplmzr6Ix
LTzCqV/1StrA5Fqguth5KFl7BHqK6htXzsvijUUjsfVZ/7EpztL62LDk4iq8HQrno4YdUIWW3acr
ZRdQfj8ztT0DhcScOE5IK4me8OCFjY6vTNDo+neN5qKyR9RLSpk2VhjTHGU1kdM6nGPT+GNNNt64
BOY5dvo1GDIKcBFPMUoE5GSW0CCKg8CMwwz19QSUUmVKE1h+a2hg+/K5p/c7m+r0lC322Gjv1O6o
ShMezqj63ENoOyxrnBguYudwpb/5ViOve36/BNv5W3EGCBTw/V0Y3PtKbikiRoOEuWasljJ/rnto
1pfaQAZCZXXBCATNzAKV6982nt1EPpQis7PsydiAxMStxNBThS+KqWZT6pts91Q7Sx3caHRvVpor
OhAfqcqptCkah1si7VbvY7Hn7PCVkg6PEzLka8MZn0ieqpzQcqLJkutuZGAm9lrNxpYfvn3a8MhR
atZ1AdTpNfF2DGt9OUBXRI+sJsFVTRN3oa0y2qdbjIEDSEfLaB/pmhNOokQAXkVJ4wLQa2enU+HE
pkpgf3M0JX1g0j2m8gfKUL+NKZGTbjEJGs1lZmoZxikWD+DtR2PkHGIpvLEw7P12F5soNQCvDMQu
FG5P2U/b2n/wNl/6bSk4gylg1waRTIA6gWgMPPVVTZzKd3/devxTptir+YpZrerT1lDVnORryBeb
R0Tbr3VMGrwPR0e/rOO5KL7Wy0RzGkUNKDkUHhTreEpPl/DCsqB3uoCwUKmEdHBHt91fb5g8kNw3
73lGKJW4GkwcPPdAlOYcQW2hlqdGX7yjfCgINhsrOjQ6QgtvJ353XZQDLm8ydND3fNA+qFgrKDYr
uMXxEF0RmvWH4zspPp0QUZIqi6jpTJgjKxKbuo+VnpnvhCRlYfRYpqnba2k2IEWCj/GnVakJH8yC
QyIA9URBLq9OrmBT9D4NxjjoOzlcWVS7X62PGkDpEs2+g0rir/9hSsubzJnAaaDnq6b4KzioLwN8
xez7osp6KWUuHTiqsLGtOPVdbrA1Geao75RkmXbNpYvV2X44QTem9F1OZiwRLuKcMzwPZqRH75a7
Iu7Ne+zpQ6BGAm6rSdnaTeFQyV5s298XEuNt7ldcDZzqVuTiolLDxIqVRywPFj+Gon6ECaN153ZF
SOdoeaPTmmpnrq1oiC+Qph2BcrOrqZ5veQ==
`protect end_protected
