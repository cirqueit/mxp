XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������M�f�6_�j#�?8g)���r^�♹n��7N����l��t�>,,�O�n���^;q�E���/�zʘ�}�EU���2�n�~� WB�!�'Ap&�P+�
6��{���)Z�]I&Q���Z�eDĎM�.(ݑ$�u��]�/]*�cA�Nʸ��83M |��ŵ�篨5CP�I����WL��ĥ�)���4�|t.,5R��=o��|�::���j�ܼ��PRD�O����M����F0z����P���i�iξ_�����kD��B��Ec�b�<�k=e����r�~e����8�����&_��>�L����$�����x-#���+��S��.FRjJ�u57o�D�H����d��*~�>������a|�a����v��A��	O�/����@��� ����5$?��ۼ�Oc����ܾ�2�LEɆ�5�j--�>?[|��"���Η�R?�V2V�_��&���!2E�D.�����?('Qr�V���S��G�i�%������F`�)�T�5�b�a��6���Ś7�	����{��'��Q�c�Ћ}��
�	=b�U��`������LU�i	rg�4��ΏpF�Jد)�f��h	���n�!5�AC�}��K^�����['��D�dZ�,��7�'`l���W�+J�#�M&W�z�T�7�tp������.�I~�?�C
'����Q�e�$�����V��	F��RR���~��R��+X��4֞��3i��� XlxVHYEB     400     1c0@8�C�۰�Ec^"1KnAʍ���s�,;B���[�*#����BlEN�$ܤ����Ж�+4�m>:T�~��S�H��b���2��T���>Aⴹ�Aї�pB��)�?���W�t�����_�����?��#2�������F��x�������3[p�1�u\���4Xb���le�D$�:���@���/�!���˃�$���ww��mb[��&�T�~�ͯA`�wq���eM�E3fo?Y�fL��e��Y��� �rM���x��y�͔�<����Cz �X�g���Y��X�Rd#Q�����?�T'�S��/I2�y�6���#��v؆4a^bJ��fo�@^S2� ��ciϱ��Fy�q<�):|��y�"�hUe�5�xodo$�'o�i��2d�6y���uf7����]�y��%�Ɍr�y�,�u_��Ċ8XlxVHYEB     212      d0����	5��x�d1��c`C�K�/������Ԝ��->E��R������_�l�`o73��3D:�?u����b]Cq޴��=G��D���21�g��`|����7 �)�5�8���/����aU��*yY�7t��/��I�;k�$�9�?C�U��� nŬU����Y�%����y{�[�Hjg��}�۟t�L/�;�+