XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��h�"-ջvx��E�Ԏ�O�������C� I�)����f�a͚刓�{>�%w�J��ѳ�g��ܴ��.\��
��2�w4ݓ#v=QV����f �F���0�p�W���HǮL�?���8��l�<�r� �Kl�{�N��5�p߶�����H�i5J;Q:X��B���F>��GM%Om����h�9�@��~�xVrbG.+񤌡�{2jB�g^�����{!��N��V�&FL��ɟ��XAF�3r�0v��|�N�2�i�:�H�Q��@t@"Pہe{�|�����w^�o�0��*�[ �I�P���㾩��&=���T'"z��'~�Ȼ_2xk�юT���F.��sx�+b������$�V6�U��3�'�S^���%�5p�%����C*�@����-�����"���8��R�R�|����l.�����`���|�i�`S�PD6ӕ�C�G1
�[.�y�%���'��%�oI�!������R�CbFeє�y��)��C�V:ɕm����ZA��[ґ4s+�r�Adt�ds'U�Ji-���� �@0ڞ�K�&�R%/d�U��y	��M�n��OH8�eI���W��#Wv3&�a�2hS������m�7�
xԻ-�>ڛ8��qw���J�F�=^@R%���;���N_fmld6f�g+_ؔ��]
��M��xI52����.�d����l� ux�	��T��r 0D%�]���-T"
������O�k�XlxVHYEB     400     1a0��>{l��|�]�+�������������ls�bon�NBqE�a�J�,'	ǁ�D>�c>�E�%�L�O��]o�Y��G�.��4�C���	^���;���ǂS��\���o�P45M��1�Q>�TX!�jk�������QT�~�q�=&�$"{~bf5��GUV���T87�cX<*w^�
T��wTn#�x;�rr��/�W>wih��{�II�!�6�Bf��jݽ^�*5��ͩƇ�X��ǳ�����3.c�ݥ9pS1��/�.}!2c#J=���Ǒ�g�NN<�o��Rv�6�$Dne���Z/�m��`�7��1j秒�2�w�����)�4&ʚ�����	�¤Wf�3$��SD8�GݒHɮ8�q�b)���Q��eJ�n':]���p�XB��5�x��uuXlxVHYEB     400      f08�m�����~¡0�¥���־��
�㳙|�$�mb.b�2�Ј�k�z$�~	°��A�_����8H����%�q_Ss/����L���{:\%��1{�ٶ���0�onu�J�S&�^zr�7���a�`HL`$<���
+�MUW�L�s1����E���O5�O7i��4��$n�2~q�������w�	�;����{�vN�#u6�+%NE;3�s���el^_is���XlxVHYEB     400     180Ӌ��>�ƈ�6�]/�'{��� �yi^�z@���;k��=�͌�z'~�\n�Xmf2��i�
�6��/��>��JO�{����P��7I��*&�hR�(.���g(���+(Ԁ�*w�I�[	��O�e�.^���P	"F���Љ�'���ij��C08�_��/�sI�Ȉ�Ɏ�X%9�<�"u�-kP����(�lR���3��yPkT���?l��)����+�7�C��P��d�{�S��UI1���=!γu|1���S�M��F�h����6~���c�,!r/���$�{���l�tr$�zh8��_gԨ�`^n��J���6V�P!X��o1C�^0"�E�F���s�t�|��̹��{�Z,��+�
��o\��oXlxVHYEB     400     230ϡ��72Щ��/��s;��5���~����ּ���]!{���z�Zw`��ݰDK����*X�޸6pr>m��&�y�F��\�܅�+'�Id�g�a��j�Q���_W�̊�- �l!�=u	ۚ*v+5�'��ir��EoIr�cG���^�5�)�a��<���}H��^�jg����Lb�V��p�Ї�+M�X���c$�����GMO�n6�P�?9d������W���Q�M����:\��;/o���lO������b5]��@�%�qU��8��w�y��8v��פ4W8��${C#�|��x�ֻқ��)C�/Q�ۂ� ��z{^z�;,C�G~�Ydisهb��4������jA����z1tC�ϩ�9!S&���[3�5�3{��$8l��-�u�;�4���?��rRV?2�!ˇ�b�p�� �����
��-6-7`+0�MH^s|���*�%������|��1��pw����(-^6��`�v�łbq+�a|��,jKf���&�j�h��|�ݾ���1o�,iA�#�L
P�.��J�XlxVHYEB     400     1c0�c����'}8ïa�)�\\�	t��(��o"����T��׬o���&8\È$��^>�P�E�Fx��f���T4�]�3Ga�R��v��0������K��X���A��-K�͞��OŵJ�L��	i�1�m����L�2Т��O� ��i:y����K{�'E��+�I�+t�1�	�� Ԇ ��m֚%��DvcMZ��TVF��Mы|m_o�����Ly�����q�v�'R�A��Xy�u�*r�+�P��NUv� �?/Y0I����3��2��>��� <�A��r���jGʈ�k���M(�<�e�j`�@�sM%-!���������Y._$�~ZT �hh��V�~ Ť2�R\�_q����#��ܺPݱ�G%=�%$�#9c�40��`�g� ;}m���ιgj�"��W���?H�CE�+q�W5�z]~�+XlxVHYEB     400     1a0m��ğ��XL��@�����t���N��_��PY�s��$���3�瞗9���ny�f��*���24@J޳���J[1�-���*O��*Ye xE*ύ{���n������!XԑE�I�$7�B��l]���	/|{�����A�+6��wт+7|?�� Kn�Mb�*��"M4��
�����jv7n��X����8��`�I�q�~(��:O�?�M埸ԍ�\t��`1���ǈ����	�c�'ͧ`6��}h�nSBQ ��a5��t���%��:�)U� 1�R�uG.[�A�M�I/����DVN��w$*�w0��j��D�Kf���y��˦E�j�G92�1ΧY$Kk�T�n��MÉ�8�Z@L��?uC�짊�z�ni/��1m�St�^|�+�XlxVHYEB     400     1a0S�Uю��-[�X@(��k΁z%o![��y�z�TR[Ce��-i�b����?K�Y�9�?ۤQ�r��p��`,�w�x	ˇ\)��0e��b�v���3�Ǆ#ɻP�T����׍SYA�1�&m���Q��m��rg�Sb~Paw^�(O0�F�G�Ϲ�B_$�)��f�)�A�:8So��$���|C�d��`�`�oh`%?�+u<�Vn9���ڙ��Kk��� �@=&-�����ub/f��{` �y?V�0�`�E����g�G����XBWW'������ʜ�r�Y�������&^���%�
�ST�:�i��+۶N�(�Y�k�~�t#���O?Ο0���T)lA�D�C�ag��*:�Z�N��v�L�Ι��z�{*3���D�9DQ���:H��XlxVHYEB     400     1b0&��r�ʂ�k 3V���R����y���H?b��X�$h��*~S$�s"c������{�bP� �ь%O��QAޅ*��}�
x_�H��UXd�� =��}h�.Jg\�d����hߔJ��:��)y�
vV���*_1c��cbr�y	�Bq[W��5��
�a���u��ZT:l/��O�Ԧ]��}�~g���F��J/9�6JT�_C��{5]�T�2Ak$��'B1�d��2��ŷ�iZ�]��n�`@B�z�����b�"�m6�/�lS�a=P�2�t�nu�ű�M�@�.>�g.	�!@d�ks1�oG�NoS��y�/��R�'����,Ѧp0��u7cF�*�CB{߫	�p�p��--R�;�[�j������Yj��qH$4θ$}� �M<2`t.C��S�)���t#�p�zXlxVHYEB     400     1e0	�!���cz�����q��>G{�Sq=�yr��BQ��f�,K;.�YNTR���%UaV�� ��;1
����B��� Ր����#N~���	���Y�=�}��C�pts���6�y��ȌX{���kٖ��N m��'yu���{�J�Rr�A� �Ǚ��.�'�2�s��_dl9^l�c����v�lִS�q��~mR��Ӳ�@~�H��شO܀�a�����?"c��|�	��lmsӥa.(�Cc2ϡ;��W �7�Z(!*j���r�`�י kFY'(����d�\��x`�j{/��-K��ė����	�����
�<���7^:��j�gW���Nl��\{0$�&����N|���=xi�eZ���O�/�eʁ2!�Ê�ܚ�d@Q��Ӟ���-W�`h�c��z'���Șg����"jB�i>���Q��b�-���r�XlxVHYEB     400     170$�~,]:zaayT��(-5E+#����^Z"��|d�q��n,��*&E2������ܼ5�:�5����Q�B\V�o��*m2�:�ñ�']xuA��*�a�xz�r�q���j`�F��1Zl��:C�9T�S���g��Q�/ǈr!��?
�K�����Y-R�fXr����r3�����8�֔Q������"�:ё��Hl���;��ȺF|þ�"lK�bd�����!>�	*�I�s�����]�ʖ�tr�!��G��5h��]����
e��9NXȺ����N?����4��[�g�wH��Յ)����2SP3�2�;�9�qÌ��b�:��K�]Ō5�T}�3����ϑ}XlxVHYEB     400     140���Z�ɟ�D.P���Xv�a>�P�P������9e�F*�9$Z�|o��a�D�"�?��b��g���fw��uS��ª���[4h}��O45e�xRK麵�h��v4|'�4��Y��2��������N��?X8[K���T��� آK.�l�ƍ8Ȼ�_�X9�������X��G�B=�m��NP7FFJ\.N�T�=�J�0�r��5Ts? 9F�_ϑ7r�s��U�8��2?��%��B�o�B��
B%c1i��Lgv}ù����4�A���̜�ޞ�hd��Rv��w.�~��h�ER�]�5*lXlxVHYEB     400     140r�6GaU��Õ����x�`<u�Lw��^�*D9Z򨈑��:�p1��2Ž�(blh�  J ��Z9Y�Ɯb�(�匆���LB�q��O6��ˁ`�L�#�W����&>�R;WU��ZK��ȳU��H���	��3�y�R��e��)�2JG��M�}���@K���Xg2z�2�{��c�b �������,��7�D�nT,I���X!҇(�F��!� ���M&|l�,h,-��f�U���1䰔w�P��/o��0�c�y��yC|d��Ʋ�j����_A���DT���s�7���7[(�B��	�A��XlxVHYEB     400     180�a�'���X����0�Bi�7��b$�Q���J�O�J,��u9ħY+�Z��If�����4�&+�-g0U�G�������Ĩt��K?i���\7�[R��؊��%M3֖n2��Wf<5(9 |N�>T\6��3�e�Y-hX]"�Fw;a��P�X�}*쁗����Ğc���`洊h�ikdd��nr}h�9�3#ۆ�p���ς��nY��w�����9Z�T��n�K�Rc
|v���(�B�A�(v��֗�(㎃_��#�Ί���Hݛ���0���(G��5�_� � �|�^/@Y��>1b���[V_���e,M,��F_��g�S,�9m�"!Dx*��5�q�t�*��JP��j���XlxVHYEB     400     180�:�?8z9�Y����28O�DI/��X���	�)�1� ��7�OK��'���~i��yKGnc�M|C������2�E:e?���$/�f�� ���Ft���%�2��	�4��ݢ�����%9d�S��EI��~��_͵&?��+�q5�?�X�jEҨegUP�G�Ao"�@#�}����b���R~A��U<swϹ�%d1�<�L�mF�pe
>=t)��#�L&u�·�3�\���V�o8������2�л��ă�]q���ܿ(�r������v�Չ�tŧAOh�'xy`-Xͅ?�Qc\��h�-�@�(�L_԰�x����2�[[m���q'i����ť� ��s�J�=�9W>?�u�!��AXlxVHYEB     400     180�֟�>Vδ)$>�%m�K�vDe�Fa9K�1����XԸ�)�\��b�F�V�I��\s��pѧ; 팆՜�	\�T{�˩��}O���s��<{@�sB�W�ܢF��uq�"ɂ\㠔c��hW�K�6�o$�`�u���1'��H5�s47�B�Z��|�h�UG���Mj�b��I���x�V�݋'��kш�W�($̣�fFn[�٬��h��Q�M@�W���^F;Ǒ�aڐ�v9��Pr.
[�rZ'��i���$R��UΥ@naw�_�'ι�� S�������O`*��p��>�\�G;Gd�*#<�O��$��N�����>m�28LD�+N�Z���N�@65��0�@���o5�%�;��XlxVHYEB     400     1a0��&�y��e�mE��O�E{�]W WQ���1�[�K���G��cQ 9�k����$�4��1#]-.�d_�#c������}��Ā4`�j\_TaȐ��7�����(�ϳ)lpG����!T��}��bl��
B�i㌭�q��*i�!�}�۠������%%L��	�^ͱ��M�2S4n,��lA��V��yݖ�d��P�R�9澓��9�L'bKQ��,J��՚�)7�0�{�M�&�e��v��Q!E��B_Ur��R����o����F��­�9`���Z�q�/���M�U	S�Z(O,C�>`\��������K�$v�T7p=;3^[Yg�[�)RvOGB��2f����E+�W�F��#��	,�1�	�D�̖Eͽ�_b.�۹�;2������}��6�?B��|'7�XlxVHYEB     400     1a0�O8���?� Xާ�ݣX��y]�Θ�/�i���1h�U���,��Z�*��pe�"�w��~�83�-�lD��1T�(�_�3����T1��R���$��3̟?�s1b�`��aM1��l�m�,��yKaE�b�>Q����Hh�P�ᢾё�_aBN�Uo�6�$��<�G��?���p4�t�y[�W�S����E�"jy��>,o<�k�#և�A>Si�^b"%�Afl��_&
��7|kN���4U�^^�J�0=��@L�0��r-������t��s��σ�]�ь�5=�%�r9�O���~�$O���j����QT7�M#o[�k�n6�m�[��w;3ý�L��ڞMd}4���rh,4(P���o�?>\���Y�\�1�s�V��Rs�VҺ��gv	
�'�(�]�XlxVHYEB     22d     110����b7��'eI�P���"������]�&�ҹ{��U(���|N��P�,���s͟�z7La��-��s������d$HQn����&t�(�b�����<�n,lukc�}"��Zկf���$q��a1�1�a�M���ؤ�}p7�{N9�~3��Cݤ��7ϙV\�cO��D�ٷ.�.�um�`C:½�u�J�9���7f�ߔ�E6����M�^s}&���0��ԫK�z�_�%r�\��J��[�þ�tTK�����T�