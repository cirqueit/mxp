XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y�D5�ϖ�����E�C;�%i�*��7TԜP�fس����.�V#t�_A>�G;m����mu�0-�R���l�Jz���QGQځ�B��Yv�k(������WjԚ|�q��Z�SXV�{xo�X�JkS�: ���7&)@k�мw�,K��x}4�#L�,U�^����5W`�,���u���g��+���p���%��#�A?r*��^ߝ�~��n8�#���(֌���	�����+Ģ��|����E�>=�T��C�k91V�/�g�Q��I�<�<����Q����/��Ğ��I�qu����PM[8��9f��D��=l!Z��;z�$^̜KBc+q�-s�M�Ap���8��6�����w���̕��e�E�$����J�������)
}ݖ;�81�}a��2�9�pZ�88N0}p�c�	QpP;M���ҕ�#�A99�J��g�8��
�A>g��3��ޢMm���}�A����k��O�`BK1K��MwBw��y'4t�a\P'e6�����LSS-�H�ɘSȒ�7>��I�0��s��5�+�1�>�i�*��\(wԎ�)v�#�@ӗc��v�:�lM$�ˮ���}�y��V碇���9��b<���RM;�2A���K%��~b����0�ځ�Fg���|} NkӪ�� ��T��a�7�<��	=���DR������j9^A�A�!� ,�Ǟ�W��)է����љL��1{���Y1��`��D���V.��a9뀌XlxVHYEB     400     240s�������ӷ���,�Х�"Ovԅ��y�q)
��� �e�q�k���3�D�����E�/.$j0�>�/� (<ri�"�WZ�NSP220�c��U���2����ȵ���2��4*��W�Ȓ&�D{����@��
��J&�8��	.Ѱ����!渄�����$�Q�B�e+�=���3#[��f^[�:"d.��m��3�B:���$�A�ڛ�x�&O�V~����	x,9��^Wݯc���C�:��و��@}����	�y�շF�ez�LR���\�ROi�5��y�Y�-������q,D�@��i8�v��w]�ϟ �9�3�$�t@ʊ;�_C�8ggf%��xa��i�TP�g
F�v{����E0S3Vqz}��V��䢤��S�E���p����~V��p#�ݙ&&
�1��c�lq�ŗl�ʾ��')=�H���/���i򗴏��>�S�S)
�1��E{��2�r��Gq^z0�|�#��Mw}�m�mu�۲-+V"53d���≥�|�}U1~מ)���T�`��vc�N#&�:�?n�X�Q���XlxVHYEB     400     210��`��u-[��Z�<���$�m�R�#ňF��[ܽ����l'zRE�a��'
෉�S��_K�&g�A�Zu�ƨM�I��^��$i<�q;�����Z����>Ӻ-?"�')���1��V�q���'���V�(EX�HyS���.�LsA�B�HP`�S�h3�ʣ�/��(��c�1�=��pcG=JK�|� Fi�{ݠ�"L��B 3��ߡڋײ�]2SF�"h�%��Vs� �1{�3s!��5XL}v@��c+�V��U㗇֤�|���`��`�1��|��
pqXL>`�p��!����{�~�F�(����;�*	B8���<�x�7m���Ū�t`���Dj��T[���PQ�ݻ?=����$�\�Uu��U��ݐ��_���#��)]���2�D�)�F��{�V�3�?�Q�V8I���;��������ؽq�}ՔTZa�,���yB\,%�Pҹǔ���@gAL��t�H����p� Y�Y�_�&���?j�)�"V�G}#a�K��nVcnq��/O]�A�XlxVHYEB     400     1f0V���ߵ�7׾`6��d���֦�D�����mՋ{p��J"�%P������[��՛�p�(þ̛6f4؈:��D�(q�J�r*��u�m��3p��۲|���W�u8�*��gܾ$*��-�BO0P��������Ĉ�X�k�$}v�kB.j[!5���V�-�����8�\+�f�َCe~�\�sp4~�
�F/L����KXT����ݶX�s�<�:�;/�1�����b(�i}����ּU��UV��%�V��^ӓ� �>���h��(�fQ��w.ْw��;�Vٕ�L��Z��xy8"�s�jd3�p9�9�ٽ�[���*^4c*�*�ou�d������~��
�ל���_�mZ�~�MY(J����np����5&����@�C}_���	�`qV��6����ě��m�����JiP̸x�n̮�(�qB�!��1��8�A}xw��lw��}4g/FT�ZZ�����-��O,Þ��s�	y�#I�̛����VXlxVHYEB     400     1c0mSzJ������a��G��R0�v�J)R����M����sG�%Fʃx�n~x-[�f���O 4��\��8�W�b�%b�]�[;?w��XT.4h�6.)�-�X�8���A�5����n�{&����_�5r�+��)�c��у������x߈��xL��s!]B\@�;O6= �&9C��c�	�FP�˴ 
��PÙO�5�&A��ﶻ-eغ����zf�bR·6 ��QP�<�����m(pOD�7��i�CHtS�&���f]J�؝�X�"�*����!k�݉IV�HR���	��_u�젇��#���{�ӳ:���-/{G#�tb1��0E:^�Æl�ⱁrs}}��T��pwn�������zS`v��j��1M#����Ā\XA�)�|�Mw2�IWTvWu,�������cC��xЙ fC�;,:@��@#z�g�	quXlxVHYEB     400     200����^�C~2����8,3��6���y��Jse*�7��s�[lC[W�ܶb
~I ��Kpy�5�������A��G3ĄIT�<n$�s��|r�;6��W�z�7�L~�����O.R[�F3���s���|Y_׆��������0����^"�P��
n��c�N���̘�6���<����E3��(�����	Xd�O�0�慨�-��W��۝#I���tE;{���~�1ΐ��l����أ��zQ'&�` �EO�H*Z�dc٢y��$�x"N��r���_伿�=�Y��3��� k��x޷��3tY��V1��'�1{^���_�*�kP�U
�hI�����pYu���\c��CD������u�w�|��r^����[O4�Y#2S��#0�;���F�>�^1�.�-G^�J�` �t��1�7'�	$��&�}�Ѩ�Y}�J�����0Xv}(��3}��ǏCsJ>*�uմxJW\� %���=a=�����ʉ`4���z>�Y͔fMXlxVHYEB     400     120!�i����&��
���mA_�Q�jxk�$O�^����8�'*,9�~�&�n�QΞ!���⪏��nA6������8A ޳��R���� ��-�^=U�yD�9pF�P��4�>k�@�je2�;���H9S����n�B4�*�K�5=b$�2ی;��xj���<�kt ���V��:#��l���3CRӳ9�N:������A^�;��",{ %��ڪ��R�i�+.��f�͕��pX2��>��g�թݤ�r���հ5K	��H虲��ך����XlxVHYEB     400     1a0?��`��;�3� ����b�P�l'��po��	�^=k$p��� � z<��������Y
�m"v�4X�om��9� �(���/X��j:���˲��^�Y�{λ��$�!{���<5b�8�u�G��O�pӞnZJ̴v@+bGH��9�����w��u��eg1�0e!�I9h����ݵ2��cVÅP�P��aP�sl��[|�X�$N����#)�a[PdPtKM�e�������mg���p���;�}��U���/@
�m������7�����!�OISjVڷb�����؎�)(*؀�z�;v�^	5O[�m�����U�BG�>�94�	���Ùܟ0�:�o�	�ߨew$wN�=77!4Ѥ$&���2l2y?𦪬u
O��-<iwkK=�����YeM��XlxVHYEB     400     110��^�tL^�A���J�@���7:J�5��Jy�@��L ��x1����G��ceU��R�(��y� ��R�}N��Q���,���������C(��·�ٵ�P7��z
��.1{�� �#��n Մ;�q@A�`RU��A�Q�隠�Qgޤ��Ѽ/�U�85b7ǣٌ�2�Py��v�i���x*������T���z
���MI;i;�(L��3̜�~n��,FZ�PmG�dZ���$H�1}~��;kXlxVHYEB     400      f0�R�.�^�ش?v�o�a��˯0�^
����dW�~�T|��������Ё�6�BT;�6�8�ta�J�7�Ѧ��M	��ۙ�{�Pc��w��=|��,�*�$kcX�Js��e�s�zDa����_+��!D 2�+&B�S�5N�Bʘ�m	�u�u1p����Ȉf*�/�St�XQ�=����)a��m4)�����e>Ĕ-�D�@���mL]�W���b���XlxVHYEB     400     130	.� �1���� �|�r�jIgt�H��B�:ܥL�������ֳ4Ze�����C�t3�/rk�J;K���B��΋��I��)װ3��C��۟"����4K���w��������D��[ ��-�j
J����"�.Ӑ�@��0^�?�l��������/� J� 6�aVE ����i���C�|uX&5�2���_���!�7+u�
גϝ��������o-<
���P�w�&s��üX���b<�g���v��Xr_6���O4]>��of����	7e��Sgg-+|�Gn�XlxVHYEB     400     130 ���ϑw��r&8~�벓���h>Q�E�4˱eK��S��T����79�1�D�c�TW���)��^��>�f�:ȥd�>����5��}I3Q62=�Fg�mE�J������6�{_���툺�uΏ�9ip�
�c݊+�v�j�U�f`���A^�o;Hu�����^\�\�� ��	�~�U�r)�����o'8�x�'�uh8�81ؿ�hF��ǻA�w"$%Y�����������\�!rj���f�.�FT������OU�('��ү[�h��(P���u��_K�V`H���9XlxVHYEB     400     130Rd�8Σ?��0���h|A��xG�L��|j,�em��C�=F��I�kL]�<*���U�;Bw	���{���dW�<��L>�<L#RH�3�Q�ͺ�VFWБ�Q��0|9�/%�!�j,Ay�:�Q��7�zsv�fzY���N�����r|�D8Z�CW�@��� �G,�{�l�Sğ��ꬥ���IWF�LOA�? �@E��?[��pWγ��j�qZ�Z��c���|�3��ԉߓu��ܟ�Sh:W8_�{X�ʧ�*^���}3۽��f�f��Pr4ΏEs��H���טb5{�(xMͨLKXlxVHYEB     400     190���I:�?�P��E<GQǥ0���H8������S�7=N%�x�1b��U�ֲ^��Xf�f��g���A!f�oϹ-v;�VW:�7
���0;����S�̠8Rwǯez�l�)S�(훋G��<E���zC������ɯn�	6������2��@[��]=`�_0�ߟ[*(�{#(���b��'ǜmP��.D����x6�D�X�����q�:�!��mˠ��=N��n^�:�q��1��F=��9G����w(qi��ή�����چtߎ�</5`��ʂ�9Ǜ_C�6O���Ỹ/,��Bw~cq3p���Z�nȨt�_��%����:��p?=6$������-�c���oT9�$(�l��w�;F���6�0���XlxVHYEB     400     110�q��⥿��z�(G����H�K3���{ᒝ��:M��2��8�<�^v�Q�Q�.��a������E�20�΃;X���\CCS�9̒_t�|WeW���%���^=z�S%����շˀ0���^��	��N7������cߒخ�Pe�)~aw���K}���j8l�5,�N�oY��=��o�"�(��Q�/fo�˱hW�DT��[�<D�WNnIF�ߝ�����J�(#8���	�U��|�sZT �!��-C�n��B�#��nCH�XlxVHYEB     400     1b0!Z�y��*�,<I�Fi���s��dU�+_�iA�H�MUD���g7��B�k���'�XNO�q��C������Pr5n��&+��Za��H�$����h$w8�7'0�ۙ��8n
(��%��M~C��sĴVײ���4�=�$T	`�a�pq�걔�a\Wxg)J��f�B���g��L��nK
�OO�uz�@�Ce@������Ѕ4"�r�H�DpOf�ѵ�<�Q�׽����!��<�%�f�}	M���s���ML���?v�t���l|jZ��Eiu���]��,���AaD��qϩR����XH��*�,;%�����(y�'+�$��QB���R=����N.���I�t\��s����C����Vu��I���8���QY��O��ү�˥�}��>P�/"����XlxVHYEB     400     190F�v����[%D�se��dd'X.7��L�0"c1I�b����1���Z{H� ��j�8��np�w]^n�ݟɨ��l������̻�-�KV�#Bz^c ,;`c|e���x3{�I}�4�G�5�:�R�X�r[��%�K�o6��ZC� K�u3��T��g�/�.%[;J�RSI�nKC��t�g�R�A%ɿ���h�?��tb*��"t^�IA�b�w�	��:7&����L�i�xaS���I��*x��b6&��Ȕo�E;���E�v��97؟�~E�}��Z#�f��^��!MF�����hE�G�S����K2�6�:l����T���>~�3�U"�Rt�o���P�Ԩ?+�����CfT�o@| ��Ԟx�d�j�OT_���M3~���XlxVHYEB     400     120Vi;�c7D>�,�)��j���$�'�jV�^8pKw�c&|[՞��i����j��+�}���p!���QI?�;&��S��4_B���d<}�L��n|�渲��%�&\n9�aS�g6�|��n�B��V��iS�h��@��/�w[O���Y�g��p�z#`��(�8{�/��^���:E��[��o�����ǅ��iK��R)��]q�g����1r�ui����v�G�},��MLҢ�񒯔C���f�g;�%��OՂ����!L,@��,��Y�JXlxVHYEB     400     120E�z���P�����i�Gg�Z��	̿��:6	Uk���$�' �3+!B���V��qa�6�f�4��EV
^��:�#'z�I<�RM��ӈ"�u� �Ѓ�Wv�y�Vэ;��� Ⱦ���`x )h޿�m��~���I��&���u�z�V��=N)���{t�AM翼��W���֐ɒ ���`�	�n�Mx�T	"�S�	:w�~��r�����-&/~��:�w�h(aٍA��$�𦉐Ke��QrCd\�{���	Z���BXX0�Q�tH��3�AXlxVHYEB     400     160%9N/�1P���r��_��_m~Md���<q��l��h4�H�qt3�^�����B������	J 迥���K�Ø:��S�3�$�@w��բH��!	e���a���w�ma��sU�Z�P]W �H�>��U0*F�3]��֎���	ArS����������:/�J-q��D��N��&%/����Wm�5C�=@�uƶ����a���b!+[xGݑ�B�7c�ݚ������3��n�Os)?�X^ �M��c�(�����X��G�V�伤�+&�/�*b����I5���v��}�?}̟�#&-J9���4�z���D�\S����ʭ����/$�H��&�̜��XlxVHYEB     400     150�{���U�Z׊�N����Xo/��5Ԍ���7����]��mN[�Ԑ-����|B��%rS�����Nz�mN^k��ֆٌ�P)̊M� �t�+�u�<�&�N�u@��E��}n�)9���Kԧ'=}��.�@"�/����v>�gk��}�-�x?��&"���ƹE�����(\XQ.��r��)���	���?b�K�[����.ϕ�L�c�D����-O���ڴd.ޮ̣��\ȸ��9�@��m�*PD��7ub�t�^IS]��l�Ы�ɷiM��=p�ƪ]��*W�V��䉩� �JV��_��`�sΎ��u�ij��RXlxVHYEB     400      e0ّ⿹�(��,��ƥػ�=�m� �=^��cC��F�J���i�l��/���${����{d����{�.E�W�k�˿�A|☚T́X�}lz�%lM#o�)��z��_3?.��)@�5��_�MR�-c�� ��m�����|�Q�|)�;��T��sQ<�z���K��b{�ٖ�B9�m}6g��PE�!]����η�V���J[�AXlxVHYEB     400     130OTW55�"\X`Kn�lo(�1��yIv�}*b����^ ��.�u��gK�8�DJ��Ðda�"��\k�HG��q�E����%�ix␭�6�ٝq�ۖ�()��T��~D5�Y�����	���vn�~�h�0�7��W�J~.�f-S'�m�!�3p�=`e�s�"�ZD�*�`�IĨ>�@>�f��<�(�Hc�fŏ<h�D,d��DG��#4�"�/B>Q��q���^��s�y��t;!���^����>]O<�<�re\��ޮLIk�H)�_#�7�Ή�}P���] h*o��XlxVHYEB     400     140?�@fBG����a��XZ}s����>XJ�_"��`�=�憑>����Չ���7d�o"Y*d;�@�!�f�1rћ �Txc�:�E�ܛ= �c]	I���	|�(Qt�$o����.��@���m��?��i���s���8;T�Y��F�G���Cy=�7����ghZ��#j!�׌�RK��U��>/�� N����C4����h��@�Q�%�֎ϟ	Ѱ�њ�Q2����0@v%D���
3�sX�W}wjeg�8\�<�7b��`Ue_w7��n~���ѹ����������p�o��^,��N"j��#ͷ����7�K36�ǹ/XlxVHYEB     400     150��$�HP~�X�Y�(�������Z�T$��!PW>��Ix� ��D�͸�n.<ܙ�ٛZ�gi����mE���r�hײ�"Xb���:�<�t�b��qK�++UܳZ���r�!k�e�N��,�$CH�?}Q�H�$�kI-xQs���Ķ����_A�����]o�:N�Ӵz T�pߦ����x����qS�2b;l���؏I�P}�Խ��1n��&
>P�+1ph����h�X�L{=hb��QaD!/�^���鰭�Y8����a:ㆥ�ɱ=o���ۀ��e�A�r�ɗ�F�wSII]�S+��*Ms��[�����?Ntk��(�}w�XlxVHYEB     400     150{|.�rgr�_��Tk�m��;����<a�]����}O%�R�1r�=�u�3�=����#���9t+a[��`/�\b+�c���i@[��Q���J�j��b�o��L(ע��X ���KS����2����?�T����->���ɾ}���ߔ�P�R��>+�G�p�XE� �J��7w�&5oG3�7���'/MPz�I�=�VF�����:;����裼�Nr��҈����mߧ��h\�ֵN����[�>����F+[�q��Z������t���`�C�P�I87�|!�h]��*��+	;�wc���[G�f�=�%`$h63uk����}XlxVHYEB     400     120�$ق0�
BV���Y6�+銝3���E�N�{�X��+�tQ����l�'M��%Tw�_Q.����9�p��o=�	�Q�!�6��:`?��X�%�/-�� X�(����v�"X�G��!��Xq�d�2�fڒ1
<Iʖ���S:��#xt褟7Q}oK	7<������(B��0e�;QV��KԊ�E�AcO�t��{�hm��FǮ0b��	ЙCRӜÈo�Q�����>������Pj��D'}Lg�k0Dq G����{�b��,Oһ8�&*mXlxVHYEB     400     130C�d�C��^����Đ���֛-��~:��\�P=�`�y�-�%Y{c�D���,�&� ����'��U����N�
9������܄5֝��f���4�e�O���ӝ�,0�䥯x��2��kO'��o�x��s�I�˗9KV~,m� U����Wȓ�+�5%���?�(�?Ʀ�b�����e�ϓf����n����4�5�e��-􅑳��J;��+��N��/C_L�>�'��� EI})��C�j�%��]M�	��B(�A��3F]O����or�b����J���@�Z�XlxVHYEB     400     140�������Kﶾ�bDǳ��hOFB?�����v���Ɓo�����S*���z1jћ�t���=*��J��I8��aUJg���zo�����V�ڋ���kdV�)���âV�3s9?�f�8C��vx��6��KO�����1Kw�S%a����HC*�=�"��y���-T�Z�w�l�n/8l�Ե!a#�h�%9�`�)^�� 6F!5�w����2|����x��g�
����*�=f���u�Y[Ϲ'�� ��
�����.鉀HJ�)Vr�fL�,��`kX��t{�KI�uK��'5.��?q�69��G��XlxVHYEB     400     120يՓ��k@~-�,��$����m��;)YG8�5���%�Ν�^��\G*I�O�	�f���6�Yn@����`/�_��x�e��;OZ��L�&JQ�H1Z���;�+��y,��<��M- ,`�8sa���	S�?U/�=�z���'�5
N<�͙��l�.(l伦v�5�؟[�i�AQۻ����.�2b�@b�[�m��	̠�S�x9��w���)��և�sZY�`qA��!+�az�v"���x�c��3X�'?�X��
ږ�3mS��A9�b���nU�G�ֿo��:p�XlxVHYEB     400     150�����m�%#>�����z�SN�?�]����8WPa2��8h^?�5%�� �wJ���%Jv�
�S9�7V�A�� �h�P���n]Υ��//�Jm^� �Ȟ����a�&L�A�
O��RVKg��C ��_�*�ʴ�?�|�Q��w�%�lq��$RGE�ju���a���efx!K/����=�n�=Q�^�`d�U/DzՄ��VF[�QWpOGw���v���~�������[�e`	�-aԖ�+63X�5_�^��+Ȑ�b�2�Z����|$,}��w1|	�gq��n&�;<��.�"~��X�;NI��%G�;ᧃ��*/*�\�XlxVHYEB     400     150q*J�$�˘�t�2A�J	c�����IoL��8�u�M��{u��.���A�kp��wrg��%�~B�7��5�0U�!M��Kd�w�%#f���O:�0#X�_�8y~�D���e0�`�i���EJ�[�
�7�w��H�S��:������!�c4�W.g�]��+E�D�o����ۿ�!\���Z��;��6�,M��:��
b��~˼�I����bJ>Bd";��j�߁ ����}�s��z��3x�[�z����$O.2�.�n"rD(��S���bwz����k�n�����@'I~��NB�&+�Ս�ka빜�ҚZ��#*?G�3��ԡt�XlxVHYEB     400      c0R7��8O!���}b�!���'�~j"����#R_k�P�٭U	�f���l;q�o�*��>
u�A��_aړx��8���BB��7V%����&s�7/<c��JV�Vq��k'���ZP�4�>��_��;�*|��A�07����`8���7�W�hHq���d�������yگ+�&��g���U�uJXlxVHYEB     400      c0Z���æ�8dB���mhrR6R�]02�=F`�(��'�l��۬����X�.���	񘿝��������geO�
��?�g2�.%z6��y]��<(n%i�@�J,�Ŵ�;�[�$O~�1��O	쟖[l�7�b��U��T�V'�0_��Tr��������Cl7[�n���ޔn����#�#��i$��XlxVHYEB     400     130�5���?��}�c\"�hL�ޱ%�A�hhn+��"5E��?������%:��¥]�B��3�ڤJ/yr���%.NB\V�-S�gu��6�EU�~�fn�$�i����<f�n�5�e��a��l㗿}�^��8�z� "y�_������fd&��G'�� AE���m�)��ʓ3Fa� �v��p}&F�C�,r����\$����BðeQ��޹A��T �v�dtϣcZ���T�L:T{�}/����	A�ߛCˠ�}:a���N`��E'���~�ߦ�t�]9=�0|S&^=7({�<�XlxVHYEB     400     120A��$�g5-D)O��O��[>�n�%AS��v��Z�c��ʨ>H�]�����ֵ�A�}����/��f̖)1sY�#�'Ǣa�E��=�u	y4��t@2��:7a1:{X1mwc��"��WǑy4 �=���e�a�aj�N�I�{ފj�Y\���9H����t\��Ej������i>�s��P��f'H����u���/�+d��gY���.[8([hw���uqWc�s������2�����jp#�
�ӫ('�B_��p�)�T����3���|�QE�t@3*;�TXlxVHYEB     400     100�׸m��g�5���<�a��o�e���/���#F���tdd���,5�$�~�Z�CA��Ktޅt�(�d�H��w��{���-
p� EB�U�I��??%��Z�*��Q������`d�^����C^�.�<f0R�u�ff��a��Id+z�����(�<b�³��&�SͪD���`�t���j.���؜�;}��x ���sݮ�O�Q��)ֵ��Ii���Gs�{��B�0a�ףc Nm_	�+a��z�a+XlxVHYEB     400     160
"���7J�1N��nV8��:�'&���G�ȸ<���b�)�b��೟�ϥJ�<��E��_/&S�qr.v�Kf�G;4��=��)w�ś�i����_��}�i� �:�>�*E���tΧd�9p�R�6GsE���
\\$�X��G��5�J\8��j�z��(\�ʑa|��`\<n���;h;�b]��
�U�Z,���%*�'s��R��˃V�=���J����{�:�1ؕ�<�G=�Ѐ���z1�/�X��`0��� ��+<�L��" 
i�0��Xo�P,�ďZ�,�
���G<�o��� 7���"�� c���[�ˌ�m��0�~:�FTVB-XlxVHYEB     400     1c0m�ObL��8x��x�S����RZ23e��_�o.MsO�-{���9�Llq\���%*�%=��R�/:m��Q@��Ʊv8
�n]���5���b��ۮEh�CV���U�\x�q%O���ן�Xr��lS20�Intv�%�`�>c�b�_�5�
�#�)�����A�l��1BE�Ku��9�M��BèkL�ֻd��q)��C����H��@c�_��m��ۤ���u���6C8q���P���l��>��ny<*�e�dih��DN��w&��)|�W�2x�H�q��R_��3���V�f�T�\=qkl�hu�IZ�,ݒv���.:�vEd�8m^3p�t�q�:]M}��h��?��ur���
ߎ.��2�e�$�:f��
�-g0���z ��" �~m3UqU��QĖ ���F8_��t���Y���C�T�?���p�Сb>h�&+�$�XlxVHYEB     400     1d0�(I-�n��F��H�j�N�e."=����\��&�o�B�*/���4y��k���3*��e�Z37��Q�_}6�B����.�Y��C���A��)6ː�ο��y2�F��LI����������Dq1��_T (�8�����o�l�U��z����AT�yl�O���I�5m��;?���yr�K�����n4�(��B���I� ��{�J����=�梩������i�}egX�ZJO����n�� �=���X������� .Ӭ��6�s�������9 0u�SHB.����AV�"���'�b$�/*Ivxh��Dq� B�vǓ��5�v�0�j�0���w|=��¤�B&�����%Z�mְJ�8�"�nsd���	f�����N�JR[˃�� CC6feHr�_�2z������������1���������S��v��8��kҥ�p�z~AXϽ�XlxVHYEB     400     1b0,"E�TB��SGդۃ�Z��''�"�]Ǖﲾx_f
�BY�ґ�I���e{9��Z��tK׮rό5'}�mJa�޷��w�v���pܮF�������`#H��Q�iZn��R�{�>���c?��sj���8�Rl|��#Wh&@�{��n�\�b��p��O�p�έ/�$�&�B�dTm�������ȏ��������u����.���Ca|�8ox_�Q��5)�U�4C��U�D�K��vI�d�h�B�u��#-���Q^�8X��q���	��l��ώ�Ԙo��43�b����2��2uܡE�����w�s��ӱ.F�s:��ʞ)9�z��q�ѿJ�6IWj� w��J��e8	RW9�������g����+�c����ce���X�<$XlxVHYEB     400     1a0�'�]��v{y�oM��G���e��N0��c���2�l͙wf���)�����.qN�p����(8j��� pn�Ӏe�Eq�ɩ�}�����`}����%��e�f5���w�(��ާ��KH=��j���/Q�����j${�V�������Uq���*PI\p�ͅ<�+8�bt~�w���;�I/l�,���3�p� �6?�ZH�I�fTs��!fjmJ���CO�O֍�Z?^r�u��iOv�fN��R��[�1;��v��JNk��CNZsS�[�U �X��̫l����v��9���S��Tty,����s�$��-|���{�>6^�0f�_e��]$��!iӎ
\�8(�{B�;�̒��@�*�P�T(�2��u��{21����ST.��P-���7��S=>����XlxVHYEB     400     160�1��tD�}m��D>.%Z8dr��<\�-r��Qa��?mӲ�,��^�޼|+�܏� ����XDP[��A�@���S�(���Y�/��߷��N�P-�Ҵ��x����d��+��h¬�7<����}0�ו��A3gZ�576������F֤����2�`ke,���y,����d�1�
�
�́�1�j��s�d��^�������?ZPYE�&�<���JF��tY9���?�3 �V�-C^r��'�p{��zQ������Q�oӛA3{�O������va	�'��9�c��9~t }�a��]V�ޠ3$E���.8��#�ռ���~(|���	�ra�ƊPJ�7��K�4T�XlxVHYEB     400     160� h8V_s��pˈ�,%������>�.��`��0rTT�M�m���V����(
�n�M.$ɱo���:����U�J<"��3��5A�J��D�¹��P�W«h,�O�xC���]E��6�z�ߙ*��������R�Ӫ���àw���oA�)�f�f����w\�o�i �Ā4S����_P+0�켟6�ϤH�br��5u�I�B� a8�b�)��,vKGu�=~q���&�T�����Kz0��^�7�F&�N�|����YO{ca�A��!x���I�PH!К��b��P�{�Q�?��s�h�瀧ɜ[=F��'e'��@�i�}洹�@�N�b�h������XlxVHYEB     400     180-{y$�����^?�l�oFg����X�`�t�Xg�Y�lm�k�L� ���,���-��S܎}ʹ�\�W��e)�������{\i��e�aC���Q'M�S٪���k�����q�&�ۍy����3T��:?
]����Ё~C��2���?��E�Ye9X�6�|o�p������HQ	y�q����\NG�cF��3�N���(N��*_�\O�>wsp�5�ԤCop�/�7c-��(�.�
�a��/ἊPA�_޶1��
��0�&�
fQ�:ƹ�=d �>4�CtM�2<�̠2�Y�B7���VC
�)�u12bn�.6�t��,f���s9��R�{���	|� �83�q�8_�D{8� �x��������XlxVHYEB     2ed     130�m�*!@��񲂥��vl�QB~%r�
7Ubb��<���!���t�9� Z#~7���=Ƭ}( m�^��J��{2*n:������1JA�5�\}G�Wߞ�*��<�~Q�QB���d�>3*T���~&��T4c�I� E]���y�@���[��f��d���|�`r�vR�/)��!+4��+p�{��ṭ�u�2���nӢ'��q��r����v�D<�1�qΉ�[~A�"��`?]E7&�^W;K}��} 辜��G	�(cL��ʧ���@������F�ۑ}(�/[�U