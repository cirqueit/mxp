`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
7Gu2Gymp++fXXUvM1kCvnvbB9fVix4cmovVrXbJA8uYdrmLh8xhez+SZPw5odJSHfHXcTxRrQD8n
KT2pNIz4v/UwBDZpOJMVDyTGDNnbaclp5l5uNJsDlPfvCKgry3fWvkGiZS/e0vOwgAjnDVIIJ2a5
jio/61HoYiAPZGprfBQKoh/E65rP7BCXmB+nEzgJ9FhQUD3870Opl7tXUS2gQxP9L3/Ks12BKsQ/
rlH18zMXsBueIATjSuv7c2/iBJytszEgRr2IqenWoVFC4TMS3G7+MsWR9qCjxyNiB38c7Fc6aXIo
bFQ1swW23P2ty4pRMVJ00Ihb2k0eSverzU7AL7DZPCSHFEw42JBDGHvCtH6wPpsubcFiPaSCBkCT
yIQzaNfRLW6PFoBXo0DwAI7DVW4G868z6Sk1pW67MogjMGokKRDh74OVZ/rdDiP4WHIcqbKeqL3h
+g3UKi+B2siOWK66ZKVHm3fx6sXljMq/a4XVO+Leg0QHIbzNS8FeQoSf0YH8g2X3svIGf4nHlcjP
44Ir5tmGEqkQfRNZAs46ooGN8gtvYGa8J1r5RWAnRF1mD8Sq6kvpl/HOlKLYVklTILGlUAwh5iH6
KcdMslgtRpESCjWJnk4uZD7Eq+OVtcXTYUblEK4/Q7Sc/+qBCEC4yOJ3GW0pRVY3YxkFhmfyDNbe
/VO6zJ0UmrxZTt+7E3syOJZSRLqhqplih0KIotxWzPX9FbjOXUY1Ic1sJepC8VdoA1yNd4vUVphP
gy5AwmJkb1kSjcmfMoPrITZ6cfx+sPG7rOJAUUWn12SDbOizI4KJGK7tD40d1raK2W6pfir4liA7
HQ+QHK5dWVSQtO4k0UrYXF53fM/p/KjGuPxeac1AJQCEWD+jwer/F/pOuJv4H9VmSbBsB9FaD+fa
kfJIHYSyOnyT4m56UNDxD3Se88GOgQn7YGvnyvCmYUxgbsOXfVZmW9uhFFnOlqgugPsq0AZajunT
82jlDfmuhpP1Puw/CgHNxPuh5VN2khmMptwS24GafUI6mFyqoSxfrHFK16YaHtQBc6Ytzkb8QFXL
1EpqDBQm7P5TBjkbtY48Dajcld795n7Z/0XU5b1vUD7RhIXKcFQ6JHbXBOTVMGVXRXYi/BBdzZGz
U8WAhGGY3Kc8UUdz1nFpHXliuVIM/nDZoVfg5qnIUEIVqT8u4tHE6TOBxvoHDQs2o+AkT55a2vMm
BPpmUUKW3WIarW264NEHGA4oLfS6EAFpctXkLxAaL7KVJq6qLC48yDdzCSkbM67A7vFcg4rfPT6O
nR+cxzSCOszt4mQ2dw4rgVnbPXeRKHKDsGSlJomA5jgcudrfSYRuzh912Q1qTQgkEtYo+Mumd9m+
ItdxCUBSxDeTSke1LwxZJn2k1mCUVzEMolPzgACr5pQFkNKyrEoKbq7/DIktPvZCqJF+2pF87ULI
qxocxvXvITtsDcNNhLb6eCWVzoEkZRQcMfWIjN6HAV3aUzBH6PCy0mSRmV38Fg5edXBQ7y/LdGIW
YkApc4j/T3OT5sL+UjAVV1Tv1BrTF6B8ZEm9tBZ6HCZ6hLYy2Splu/R4FtexPgESUUgXTdgeIZ60
zYXFxZBUjhlB+j9K/9HSWeX6U1I5Cq0T8ra7Sc/x34QRok+p4T3dkjtk5YxTZJ9YrdZ/rVrbSG63
0jurUEQw5rFQfCY9fKTn7/3wrLYwFAFB1HS+TCzVrkk9H9VwKDWk0Gs310aO9jz+ohZuR+VQyy11
hOrK+7qcCHS4M/qmNPzLhjlX2+zHdnp3ZtGtg5mU6ehRKsN2sDPCjJJLYlLKHc9JH0shWCf3aA6d
brtjbVuKSM04VFjSGt7ZoEmrOjNoIPiQRieJ86yb7IuWmDyH49ycz6UNguXpNs3qM+u5WxD0a8Ug
OROGA9G0TNRn7M1+g7KEhEmxHADN6nHmGjwZnsIRjI9vCZwp7bNzhxd6poGiSCE/H65KIZpYsGhC
bzU61yvNB8qCkB0BlRMKGPtWw+SjCXeBj8ETi4YlMa8aC4aecFANHDpROftC22NL8DwQxs/8WyyX
AioIQ8uGXxLa0D3lbKCE/1Q0K0SYUIRDiOj/EdbvBzJ5+ro/nnOcblOAICtmwTy0tpDYis2IlxpL
KMO75+t1AyrqvRbotWp+VH746ICw8OkX6/YpdUY5zoKeop1VAvhkE9+gplPxW08mjI9HG0ZhEWFX
gKM4j/ksFJdrb/xk74p7pz6lAFlr2W1ibg7FuZyDMW9gmmxREVplx4e5x1KfzfEyL4VjKhCrkXBV
pYlZvTdV1s8N1WHTz6oOSXI31LGUQNJRaaFPVdq6wO7KrT17MOeoeQy/kwsGMRpZLmTShf5e4BcO
sn6S4ZDchagKtE68DMZCSlJrgRSYMHsaVX85aW6pAFe6Qk5UPnO47ylODM7RSfSVqZbeKaEt5a01
XccbPMdTbO6erVz0469tFvwypfgQVAwobrQ1SM8pBycluQ8a+ySKvijbzG7nNxTjqdovcHP35K8a
G8Y5LHXiTbdTgbvhc95WN1V79OkdaXgvZTaiWN1FVcHg2/8uqgzXYsQTrrf4asAmuA+k8vt6yceA
TRoCTJqMMDWFo7HBrjkSISDj4DUZ2n5hYUfhEzeI8t1azwdsCe4Uf83KTHuGtKMk2KhM5KgIumMq
8HkiyKU++cwpL5F478t8KSg6k9h/wVwnN2RulsgNCwqqb0muiMQRZrcCLM9xAszUElXAfcseohuK
r7myVmVAyeKLM75BcEPEgNKx15A9gid1RfcJmLFHF5NUllBrA4rCKtLWz1pW0Dvo3W9Gsqfcsuio
TOfXaq9FGc49XKDrdzfNXdZZZ3HtA0H+OV0ZXI/sa8wW9AJ/rqTqaRQNieVUQHPOlGO8BZ/8oZVQ
5MfkgZC6dOwZr57lucyd+2XH8DxkWr2BihxkCLOCr6U1FUSWVf+5saSmfvnM4+OoXNJap6V/2kld
X4pJ5IrsiYSGxDwAwTfzQigVMYpGzH6WZWJ+xww9z59kq3u2ze+bZxf/1FTZoBc8dNc02p2JpJlu
AZLifuYIzJbWQ9RBLj4qb60wBCxu+RFTl+xDrdpOYb5L+LBKkptFQ40UI0JAPH9DJRFPXO0tvyFu
o5FsUSwUJtATkaulw5zR/YFW9QVuEtp2GNQRgbsBFCzfHzhvL6bKyDHUP/9zqT86gMgRpBDXWsXU
NOw7BN3YhVqHelhmHaNJdcIf6iTh+fU5b3LIci5gj8ObJUi82aXh3/jv3wVR2f5QbThBkQ6LXO/L
HNyjNTHmcy1f3mL6BDS2diQYW2RuYqAuudwzm3AqjzHgezqjV7HXk+bKQW8jC5EjZmK4hBsLppz7
jCSIokcNOB3t8aKGk9Q1aGVW2vtZFdvCny0IAKb096p52AN6WrRB/ud6GLrUHwP4MTgDpVP6FoVl
YmydazBwC6sAetY8CW1ZapwKY6bX3zSAtsGRtGQGrlRLp8ieMzOCdupg/uBM9swZCKniWzr8ce+r
ScADybd4ZWkbYrRpLkmBNZgp7aYjldAm9tfuRRhFDUYdZr/CEXMKm5AvVfZwze+gQ8LWbos8lCDi
xixwbLHocTl9NMFQvckeiPeErdccMYgxueShrfPiXLJdjcm2jbZDLdaUZVi+LPR4XznBRYwXMYbF
Q6/l4SoPSsA7Egc1rmh+16c9hVt5pcFm04WjijoT8GKm+BN2aOMgtV80tL3WKYvKmwOai0DxO/X7
9GvMQ0Orr6Wh/wEDuOOK4QeO1KiAwAAWe+k7sRRF0dyfgGz9uNGrj/oYSDGU2sSn8ikbJ39rtpMJ
QRSX7SpwOmdbTspU9cPn++bObDFZR5CTMh/rtfgIWvXOZ6GGMmF+0rcn3R5mYOJQ6sYEZO72RNhE
hg0Bs+QM9P4UzpN5kwENn08J+7cDlYGz75ivctaF1SF0X368BuMisbzmIJ0P7xPG9LJV9ZBmgEe2
vJ96xmDE1bK1ukXbkNywwz4lLsgxHepAATkS3xQNFKeKSYzfWM3x2ogDbNFOFJTDUMB0B8Rbbl62
53M4bqoJN9kNZ62/FvzgG1KxEBvjlnTqhQV07Fvn8p/t1KapAofiA+gTkA42YCkl/mK1MHBFTcil
awjh2qCKMNxcpmD7eHXA8mzlokhzxZip6CoSc64kummVvtStCHetCFWyV/ciKGsMcgELfhiL7Fp0
tjFUsX/07/WFNGTO2OTfUxjjvgslR56kM6rosi/2WVDJ90ljCWo3244shHIHTScHZ4XWwe4nH7av
YZiK0T9GOEvSTr7Imc7eqhxUJzOTnug4rfdSTW8fvpHSuuHukBEven4FaQ8pcC+ChqlFdS++tnRr
lKLn2yPS3UXcK+Tsa4ih1Kn9Dl1p418LXPCjRlLeZ/eDeMihyQ1UEjy9/MhUAUKXRqAllHFf8QZA
Du47pWZDWAHCH4QoQ7AN8r09SGnPjJ/TmMsjnMZSHIWRaBsbDk4T8nhSMyI1OMfgMgCALPz9VW1i
6eK/t5B2v3A1Q4QE7sAUAnvn160Xi+MFcYzamAZAhSjTxYgOPu9u8fLUPSTGOCjWNR4oY7xdtbJC
F5jn+aW5/TTlrmMmRLGqLxvcTGiJNGiFbzKTfLQNL3cNCmWNQGLuq9xbcbVPgtYW+k98IYNY0kHv
WzV6DattFJRQ4q8/iZZTeuPgGQZ+FbSsZAj5cXDmDQ8josGewZfTM9t9sc5ZIauztM8+XNsVIK0Q
rkPthT3AcS7Hy8GQju9VUlQRUU5sDB/jnplYqzjSFacPStCR9ewjfxl5N1aKX1Cfyyq72NXB4gV9
qscdFn4UnYYe8vewBzMMPXQRVi86Lq3OPIbxtLnJdUVp8KQ0eTRZq/B4Hq65udYDfIyPA1XMOau6
qrtuPEZM5GOAmlkgdDUeZuIsDVyQaX7f9wPA0W4OQAyGwoNoe0xAyhjTvwx/E0IRa0VMYIP6BdB7
e8CaZJClWoo3OYMPgDcUwl2Dr40M3M9yGu4D/UZ7o+aAnGVHYoWIvCtzr9zr+Su5rBnrOZCglZNG
fKGBuNy/IVey9zSMwvxQq9cwoVMWhRn+OQsU+MeyZRiuIpCS9s9c1nhfg9EY7TENoNPZnmaw7u1X
7RdPBaM3SZlFYK0aYZoEk/1atVJOFYitVAF+WiqO2FOP+rCXE1HwQKGJugxqpxbGyFg8el5XHJCS
789cq7eTJj3pZvddZ8xDirz9KbqjlJoRt9WxpitM8ey1zkspEwQHM5HctDLP7IG73c/kMy6nG9iX
7nJAzb8RSC9UoLXtyr/S8YiUtO4IVppo46RYu3pF27NpLtso4g3HtoCDtdre0PvddhBAvt/nMvq0
yTJCNPERZlzSTkGQTU7UKVqBAx42SR2g4t+we8dWo9wIahluWsLfMVfhIpf6uyifgbEl1M+NmRdJ
8CvUra/p/1V0z6TgubpDKtTfEimOvNIqdLuagm5fLv8M1t+E+hhJWdpLuCMn39O28f3VwwOwyRlL
c0bwq+J49oDirNFE7SAEZkbEy5Px/kJd68lt+huehe/TdjUocrRxwqTwWIluTl6lKvTZQsWfp0Ye
ekbWrWEMqI/GqyWuEOHNJIGfKduG5RidKc/clzL7Ya5zg69XN4XLJThGjqzMySkUZECAiMzXxbfV
0pBvjBIewLYo3+E3+WC307F4Xhuo041m2G40cLxo8NHsl+MtkdYEhopDFxr/jZlAUuFjjcuBXpME
sQEzUT6QjolqC5fJ+DQRG4zqubf66APDtAo1qanpxPLkI6erxfdMKTdC1BFCY+QJGbys+PtRLkq9
zX94uz+SAjlugzB4C6cr1jxI5+4qBkJ9sUjLzUeA6HIusRCjv5T3xBLaQy9rCQd5MOhmVM/qsw9s
qv0S+WB12DcTHr5GbwzCCiKL6FcU/NLvWumn7wp8C7eogBY+oA3obU/fJglPSEDj8Aq6a8yNYcH2
+WiAWuRNLFEqBgBV/vWnrahVs6ynHvs1Fg7Z7DTAYiqlSrkEFT3um4zaGxY+xhsm94YyOSljRLPa
qQiCglnZjrlotITBn/P/p3fTNEfjjZenazv9VkhNo/wM9YLzPjBN/xSe8NvELp5Kc/YHdimhx24m
m2QAyU2xhsPsySa8RtT4w23cxL7HfWIX2cHhX73Dj4tdk+XlH0WmGGUBO/Fnld5XVJc2u1fqRWAn
poa8RwfQ5awqxneaODT4zsHemYVOTqSWgqGNKmQD2Zp4XU94p7omRgH+FIX9RIbAFpLRXlotaPVa
zZ/leI3zlIBIhG0GCro3+KJ/aP5RXWLmBtmgJObd+150SRN/dGGU0qpbI99rVGAMKw3Rfd/u5oNp
s/zG1Rc0i1kgYbPStY3FpV215M0jzK383MQfO++kB6g2aJu6HODL1pzYISgPZPyy1iKAs13Wn5Ja
i2IUiJTKfq7ycWl789oMn5qbhkiZk06OU1tl9xJptbM0g9nEHPZfoAI/PNyEm3M4Psx808vY4Xw0
hNim1M+3D8eGqJNAzTHhhc9C8nbx73y/YZ1ViwcJNe+mgZG+p1fewFu4hvUH9DM9s+GANgEFdZhd
jScFH8e/Gkx0eEaq6I1o2NkdZ/hrk5jOryNiD5erNZfQzSgCUWF+bX7UyK0RQ8KEzpVnzZl86GZY
NZHL9zjMEE4BqY6KS3txz8+WYJf0UlaZp/a7/PaFEa8POezEEkWKjakJV6a33ngIL4h7fne6bjce
0gHpER8z643NqaEWquYEkvBRpKRI1UQJEWrDVhNiQms7cGf9jUguwelGA7EKFnJfSjo6ZEXOAjXd
qJcieeSyr3CeHkQVRUvmPyUo+M//28pzUYzRriql0jEJ+yW1vybMAQVv4Ms/xi/ZoTQdi3Fzg9R+
ttTrw0Pq/DKS8ZLvVKvowxZc1oav7rcHgkMtlsIlqAtbdL3pp3JwHogz5Et2X1KpQBpiRCkd3j2l
ofvePSMlP8tHCQLNtLlD9Zm6fDahETe39nQbb9fkyFozaSsN3yQ1dSU7dd7piw8me8UIYMlIXnA1
if5aYYtT6/oARqxdb4RpgAwRx+nvItDylsnvXJRvL/yy5CYPm6FfcLtBDirwSPN+omb/wv+Pd78X
3Nth119O/0j7UijOuK77C4BnoiSHEkoOte011jNAs+bknL9psUfeZG+7eQdbO/aTIiN8fM68VIjg
bSarsXZnTdlxQ1+1la52FjQSETYGcUsCHiiiLsVH9gGdWsuYt8W9KaZ5iVyMHYcPAW6k4+ulIJnK
8/37ejWUW4ty4IZ3yLvECUV+oShqxHs5f8suX1KIS1u4mz2/ILq0oPkXMI7SvLSpWvMBiDFL2kw6
Cws9LPE2hrwstwkt2IC6k9yuxqwqkNONdTjox6LuxkeEtxod2od6gRm9nKwQMMUT46YVyUeYrpnP
24Uw1MTOGTsqt50Z4dOxb+x5S/R6ARLdb0C7lnJAjSq76o5bJvzmkSBdhmHW1pBt40vUeKKOsjsW
MWLM4xH40gXELopR1Me4e3w3WugBZ2gpSHW7FwRXm86PXTcPi0JaZxK6Klbch2cT/BizSkEVRf5G
a0qwm2Yo/VdVet3tbQ+Ii+cHWC2DWW5BiUXplsJPKH7U+b+SzpX5xwsMah1uYu/ttYPwGJIaWeL4
MyvfAIZmbGb38Y8iYi0DS2Rnp06QkpIt9WkH6WWYkkMYls10HtBce1Gp3r7xI5qRW2vDyl+Da6o2
fmxcTloOBpV/HoNzo0uDXPMgjLZPV21M2Q7HqstJfCGwqcwyEUjkIppp18ypupPuReYzm9djzBGX
FmRp4ZWbZGNIMzxpKjUEiAMW4+jk3P7sdyWqaZCQaqf5yflpJJ13IYGu/ZuNyVkxjBP0rmCqhSNH
relwhDtmFADhdCFW/jdtozcHAk7tTrDg7OAIEJ/p5JbCzGSk80R9B7tmRQmMrgV3/B8nUflct3vs
dM69XK3wH590LIyRv1yggaqJG8Ld+QxGvfV9Q622LfYdjyPNpJqbfhgolRwGKRzAtZP7YamFuNiW
HVrrj3P9i4BIo3lckwGeggRWUE+VMSqJP1H1Fm21wBUE9Ra6jEGqx4ziSj6FiJklrIXsfSigDKY1
rMQw1u6aQrG/cdgr/iy8cOEVTwCSoBu0ZjfnJANPVretfUqdQHeTLzA77H8eaww5+WPrl8JhiHXK
STbok0gE2UfEyhVH2RGKsfj6lfUimGMDejD1iBkvNBNOPxfCvpCEVoT/bZSN/6jD9cVGbUFP1JLI
bReA4N2O8NEd0MY1TCHlCZB/LOvpLvn0yuolmsRSmR5QhybRg5d0scXUbTOd6xxbP/vWIAF3hOYr
rj3TZr7HvdpEmRCk7awET4rHSA9iKyR6KVN8P/cseiEWJSRd8KEneRxkBWzQ1iAYW9FXv3JDcxfs
jtEiPgtQsZhlYJpBR03GmfryUDUZRYmyIBkVjTbMKizG3JegowbLWYT6AunsXR8v8kaM2jr6iqyd
pDrhyJ3ijsFlZ0rov8mGV6lKmNoedO6UWd1nUVN7Hh1OJqBDJZMH/DdWUCl7HVStZDvo3H33jRh/
mmaD0a3AbJAZJz7TISBh89eq2FMlGDwRuuU9657qslx+Yrf56da0JKpEjRAfPcsoLzsvmMQXWsYK
RIl9C4EJcCnsbmsF5z+pgKm1jCYVEwoemjYwkRbMu9KAG/SlR94b+/G39aeGsr7CY+wXiHjOccPW
DGcLhVw9tfOL4q3zx6WW9MPHcV1yQ0gInw+kho7/IWCFFmaRYvhaSK3nniBAMCaV5HiXXgjKBabU
WIlErtvTcmAZG1j2gPbF7IGA0NQJ1yF3BDbvA3ybXNs8Y/fhoM7pahhx3V4Z2zLa/o7vSobvh7HV
HlAT17D6yr/CycnKtM2T0ezUJc/gx26e3tjV1QDKnZOAfCbdaEK/zo++lDEEOXmFk5GpHsGrazV/
j/i9cP+JxV+OjhQodBkDKn0LDij3weJkUBtFWQB9uo3oaI2BnppK6LUgvtbdbYZqB7tQgnkd9sLC
Y0t6ksSHXbxriDCVAdsmMMYcz/aP/y3vtEiFXyiGBo4mHyBRWNCYch8KFNdRN26as/Q3luv59F/u
7o6JukjydDoCgpQl8jqd6pvBRsqp6HrBJd6rmUGbmy7mL9ZkjKTMGSEuf495qSRiJPOuHyBY+QN8
ltTs/W0zwn11l+hqiRT6ZqIJ92vFVKa1SGlY9q/aLiZbEB6KScJBf71q8U2uoKWpDQvJVibh536w
OOBzFTKiISw4q9dt9yVv0C2eXpF2w+ygEbGC2GJyVHrOUaqKeRWABCQH/+1qGtuJcbhEWK+I+0JK
Zuyw7rw/th0AeQJmSPLR19qmcXYE9Fl9o65Yv3pZJURsjx9UCgWp5HjdQbxWtlV4rodJ50ebSRbB
YhjbdtQ0Gnv7T4Zrb7VrBeRkj7tpWN6PKz+Yf5QtbirfhMe5694QIopqfJe2V3MSbdJVU7o6QbF8
cQ0EPc9fKd2P5Cv8o732kzFNu/XQPzFF3j1fT5GvTC13qDeXFD8flswNbV1oDT3pbHM7VM7FASsJ
ir5Um0goVRt87XlmMoxW34k8jXqyNAMifSOCXcSa8QSVhZAOcZKE5xAjlWiNA3iCiltuUJ12Sb6c
lpOU5dLmDX32TVPADGFceH/3Qj0UH8zok0V6bGU1dzzaeA0k6xDjyMX/75O5RUYZUFWW+eUouF2f
ccnV3l20yXsT9LB6Oc0RfhtueYA1A1E97pMRExqiZvqbv6Xkv557s23C12VOoFtBv9r1vI8uG7aw
KLkB/l5ds+DJbI/f/YPDf5h/CCEKmxWTL4lEwLZ6miXhI40Qa7TwX2jyPrtTcVsMV6eZv1F3tZkR
SkYQC8QM2MFfwM8JHH38VaRphMn9OsCghlsY3av+LzZ0NNq8cwBGb80rK1jNmtii2th35u8cfqVq
MclslS6lf1kA1+W2uEDMEoFVzus7N6bMuu72TLDKnth32t114ucygkd/82Vx4EaOrl4dLJTuPJCh
fy04Q3NmyAoj/c1Zz6D1B3x0m6LEO4Gucq5sw+ezkobXlgO9NPfNJgcKAl9TeuOnqOiEJnN/6JJs
sL4uYnzrW/uWqaHR6cs0jui02bsofh7hI6mvgFhM3dkQdKCa2I/UHrZPUpz87L5fbVMWUY0d6XKD
7CEroOJNsH3JunZ8Hqx1L8xdDfkU5tAxkXCrnH7313wYNvlWEhQwfhTtI9KP8B/+la/9+mabOom8
W7NGB3Zisb6OkxHnLnC5csr1uwuXOi9EtkPc80X2TkDNgFMtwh/ze+16iwR33z70TfL2jGeBeTUS
ki3yqr69wSWn5mo6Wcs4UfJmzFV4MOS2/WX9JJrFSRYWMHBpLGwVkAGZWwQIKJZTcv7BzyXmXvI3
HQKutlJImTRY7OWIvsmzcpbNRTehezJI5WbDm9cmS7Lyt9FvZeVto2sh0j+t8rODGpVootiEjsjL
0daXp/jLk/JpxtDqywuJKa8VS7l13OK2x7lXL67k++By+GdZ2+MRrDKVhPMimh3xPl5VXzv01dQu
OhdaoR2m0uO3J3Y3HxeNhLyqfgzG68GRZZLi8hSg0xAMwXp6h6BO/FsIOH5PjZTBC+9WjNMv+g2S
2iz8M9wQP9UNMTv2vtaKWBokFSFe64Rccj8WUts2bAP7nUa/BT59cpiRNGxIJvuCruNNJdrrnw1x
PfjSO4O8iiHeSG221VwiuV1pUXyCYOaE5SZ0X1ENiAA0qnus5SzKQ/epigqF2WacXaBnlZGvkn3U
XwbRopmFHqDC5j2PFfFRXSsLP7jcGp6FmzdrkTZ7QgiiEfKOxSyeukPCFHkRkgR1Z+efyk9PhjlE
FT9KbGMqIzm1WauMb7b08J1yMh5LvIwUvET8A9wxulMZq/f+wvh/01E10n60PCq7V42paEKY3wEJ
uGmfKzeSxIErNPwp3sFJBnOKsB+eWFrPVttsBtoVGVPrLKDJmFwmmLEPGiFW8ehPlZ4+Uj1NFVKc
tLdN1BMU0QAMnAWLYEzQCBDPqD25U4LyAaNY0dARDwyN8UfTb/vnYh5+tmhskIWMkb+m8R1sRukR
626c4f8IUKz6mORLDmqL1tEOX1n7GOcGKyGRgpMw9rXO3/WETCOT2N+nlmrKaYHGmiTeYSxv7EJy
bfk8R9C6XgyMWIyELJknpoJNgQfUIGlSOiQ8odMmev+VVx6oVi2XbjksPQnAZmYu0wMRoZ/EzW38
zsy0AIIOzECY6soZZLDSYKAdlT3xgbfN/kYetfIsOenmpdF6345l23fn3c3/lARlF/d+ygVmuz0k
DG5JVfV0AEeIbfCCAErUEhad3X2nP6Dh4oT97kb5pLctQIzGnfxLChKLRfYn6GQWD5k5ZGczQmrw
VfxMwGgBfhMYYt8Lo8knV5X/5grSJK5kWnVveGZgF4KTFVY3l9wswLYUVbkg+lkadHaEhxSfjp1c
zMXCE52fE6Rb8GZFsj8yk+3PcAsu8pSE8Ig5DJkTfSVQBahJx3C5Eq1sAfS7q4+YGStF+GzHPAKW
eG6G26HC8r7W+balO4dWP8wIE2RdEcgubxttZ9C+ubAvIYkq9WRIGzkPmEeJ/S5BY3SwCBem7Dfg
37aPwnd+SOK8DSx4OJeNGyjRNl3RBLK27jTyXTWo8QsxClvo4LzRsxtszZfjuJ+R7eN7F2+TzriY
EUtQBmzSRz1kRQngjS7JfIv8yEKTthqCCgfPoYFhTQ4ykMhspINRW8nBgeLj7qXIhDAEYyR2eUVz
w9xYHdjzLSKOLV9YfKztRULq52/BGuuLvCakg9ddUYmam8Ww6JJy4Md1dDQwDjwoXJj0RAHBPsnn
dFEEXkfdKku38nq3Rc5HxWcVcCUBUpRiW9dJwYgs/CuWhmysi2PouYzOSByDjampmdKs7R+C3aLI
8aojo3jNDNXNEsX9OUtxPmRCyvY14zZMwxOgMExstghsXmABPoo1BgFMIJDp3Bo7Dh0bsMpLg2iM
qcgzqvuNJmyg6lhQk7ixJLTBofvkJLnTkmeg979K6/MR+gFvZh3RxNZKXQPpn/h55voZA1dFL6az
jaw1SawakAxNubbsHFJhEmlqLdA3bBcEIgQItp2Vpo5HWT11y/QzyL8FS4MWa3oYRq5/O+SGonU7
8kb2R1/BKZIA/YdL/M58X4EWV72Xq8q7knL3rPFP/c4Ne5QfozMWUOYNYUNe9LyKEdO0LbljhFGb
m2yFWcfZV3GgnSHjpK+dvdE4VWGx2DI+AbEpPRes2nODcBHFcNJnGxXm/+p3jmsVRHCXTjxXH/xZ
1H2CuTW2FLC7Tc7ACLu92dq6yG7XTGE+3+LQKGHrP39jhdRXF8oujo8FK+a6guei7m5GQ2OjfgEP
ona+feRl1kESK51/WSzaLdEZ9cL+VIFp4JQFfy9v/KBVRX18X9EOEBlqJkvmTlgaPF1BmM45uIgp
7oGst/Xihgl+AlOYEn2LsaDRZSGUXJEMWFEuT9K3JGeEqEf0Kr1CROur+OoQSehdlUHOodizjmMO
o+Xm9d7N0QUS2YB1Crc4rRfpfrjruHx7JYIEQFdsME+f4JIZE51YAMQaILiOR6ib3sE0xG9b2Atu
3NG/ocZtOpmD9WOtXZ330WFGBUoU0e5Ev+TFtY54YJb4SF2QY1i/u8H3kv7f0vGw76vULaPtlHzP
NmIbmBala3KPQ6cZvsU7FPF6dfK8X2v985CzzKXXU5XsZFpgpul9IVYnPI7arhVYnvRhCf9vS6bk
Apq4+49dOJKvVCyNBe0wscB+ICt/JjKJ80ftN54pzRelMJecLly/n6X88kQrm6NEipVuj66soSIe
x6hdzS+sTIya6LB8ve4h6GYW9ML9LBPUPDZzjrjPq2UiP56MndhC1b2kpHyM1EarnyZB8lBtF2LM
svu51wAEu1MSmQ/+zrHgFPaU8SoxHCPgy/93N19S6h8TGW/RyLkV5ILNYaRchvztrJuBX8CJ9gTo
nM+PKSpqfQLV5hdGFmdPw/KL/5/+yBNwmvRgcJC1QXqK2ngxHDYTNawqMHINcDpUX1Vop4gH8N/e
d2cKT+v+O2qeVt/45+QLiQxqQ+NkX6ekpQfIjkUM7RYzucBS7aq7j30EMgtgicfXFpQneksja/BS
zUqGApFLLSkO8OfGt4LnqtM4Ty/W0SF0wZAuMP0NilLhZDPwuYNnf5RMfZ36gImuHNkWHOlEAGoo
J/cuiNkg/xAaL4igJWVWpVG5ZzTmNHXyz3QQ3eKISX45nYv+PZIhkFTrM3VEVrZtf/SqGjadiVZg
qSBDkMK1gJXRHKtC1YqiLZlOfVfvvtviEqoJOgpr8B576Gw1zfIBjFgj0OKHM87yYm8ZQqmlY4tB
oQNG9yFO7MpWR8fNnblP4VUYbUedcs80mA==
`protect end_protected
