`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
8ySVXBCFASnK0jewLYFws01fvIsjuPbpMxby5l5DSUDbGCiJGTjnmr5eXehjr1ouO1DqyxsSy5Et
n5xpHL7TTI/KLhMropiRCsgtUd74MsV5upPIaVYzw4vpTziBdBgujwXCeihTfiEUBAb5bdaKvqCP
ibbKYeF8qY9bUOuRK+sNSoNttxYmWms+7ZxC2xu2130cy05S1l3n+tn8AQk2Gtxox+PldqM3zHEG
KX13mLY0dWJ3uUrXdYFpAmL2eCWxCPEGL7UR2LW2lg/eKZhd4a7bkm5/aRd6jxNCESQ1OzQDpu13
pv0mbAW1fuO9nexnt0qI7tGlqLT5WzF/2czHWW0s7/a/SXuY8eC2pG5SOLY7seDT2c6e1MmVC+9c
pVciIZXLRlgjKEK57vn8xraHB7nhzMnjkgXqKRoeVOxV/42a/pmsYDxmz6x5Lzfp9RRbe7qKv2dr
nopc5tqv68vkV2MM99yBtwhIV2bexki9WqF7DV8KhJqeDm0+ozRa6QUoWi4zt4q3lZTTZlYH2zus
3PMMglq81M/0UMxX5wfOA/yvhO2yQMtqgL7cy4v+e9QNSwpatsi67u11U37lsM7Qkv+Nu6Bf+ngW
cwKSsk0ZDxTDoRf2Zl1a3TfON8xqr2VylYCYbrC1QFNXxyjILjDKl2/IVOSGXRO2oN49qOVKmXAF
As87/VgtzLwTCLh4LEfoOLmjXvl980gb5aT16IswzpCbfE8e1Pd2YOMxRnlEgeQPGAw+CM1mjyrr
OH1+jtetY60DdA9gqrbQmK/xJgAJb2KaZ14EdSaLwKicEo37uExO+mh0V3P7VAS5ivbkQFbE8fyx
3/mtTM/Aahe33gzow84hD3fcRwud94thRniB56/yKJ9APyvc5RQvy9Y+abB/yRp+t4JyZQfvBq6E
alpeDZuUW1nYepfvpx6azI7uhJDwHt1gr4lfsIcvJL2Jh5lwZlgJieWAH2cZqcY52i2+iXO09Srv
Xb3/Z9C6/mqmYyypmlQBwhrP6kI8S36boiqE4lHzGrLE8h38ezu5daNqomsUIGUeKO+8gDMrRqwO
WnJ+4dPw1DTt40P/P3HT9mDkf6yvfu4PBcPT1kt4Dvftf4/vQq07KgK5qqxr5L3jDrds4YkWp0T8
8IS8wIGk1Me8NruLZZ8dQfSEusaQ7r2NoxouzNxOYIiMx3CpkQoWPSc6EEHo3nNAy8CFVy71ugO4
aBjo0cuIDam56LBYPy+tSdk/58Ka49sY05g/S95iHuNfaKp7TrV3EY9uJ1W8zZcvIENdS8Bfq+6j
Tq5qghrPT9mwdbM299dffpK8FNgmyzJcLpLJLTYNYM2XOMq17EI0HEcERaInKWTeHWHTrWwrAvoG
MaA0VXChZPXmDU0SAMoszc+24V1jN4LdgVOnR/rjGFcYq7Pe6bvGlZMYa6uTmxn6PrsmD/6/pRbx
Ukp0js7DIv7nRsaMWa0b18/yhKiwjjnlTWG5Vi+T2B19mE/vEkuReviQqDJxndPoQZXZJ+qPGegx
U03L/TLEiRiHYqZBIB0MaYzmpiGVzVusU8xf6y1PmEztQGBPLuL1RQgUe/ECljH2E2osTkQo7SM+
SaRQpYO29vFf3DpJdX9Y50cQuHDRtI0MegMMsjlk2l21fdH1xVkJ2Qs0+MKiuokci5rzbzXpe5jf
Fcez+b+979cMXxW8Kel1VHlea3cSem+KHmzUWCYCW0W1BGf6bO9sL5/akwMK4VBdgcDDwcbzdlzS
yYERnFiij+16KIH6OPc9jtKBlGd7FWtPeTVObtL7v6tnDSYPW2MWRu2QB2mJ8UXh5RY+0ek9bVDL
zIJ+t6XZn3U3SaExRrXX5zPQfY8I648dxaFCpV2SvPtOTjRtb3o8PkToycB7KYE2v84j3T0oBVjB
P2wAuIFadBLh7ZaTbu08gmOzexUX3/aC7xMnNNScjzRjMbjJiJl2DuiVM6oldxwgKvfjwhTzmwnT
/kH2ct8LQnaxtwDN8U4qYJfr78srQdi/APUFhVBwlyBwasdpvtn9kLOhNKysNgSaI7wshiBKpDOE
781wvy7VoYl/d86gMRC5Z/6jfPt18kRoYOafG4Mm+gHj2mV1zdZ5UdaS2Scx
`protect end_protected
