XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���u����d�� ��g�o�`@�*m5��f��X)Y�7�R�6�н�*S���<��Q��J?,F��%�45o�qt"���9�t��w�jX��\1�1�0A�a��<�;2Q %�8Maf͵�E_b -a��t�zc��9��A�n�ު`�wbͦ�H�}��_=���,R�q��7�8ڳ�9o�7a��)��U�21;3�Wz5Y���Ɋv�uƤOs�>�7�!i��K�a��M�3�1�%��d�\�%$�C����$����p2Q�c)� b�R$�Y0F��|?~�)T�4Ԯ��%*j�]�^v����,�6�ι8ƚA-��8v���m�W0��W��1��ʐ��|�(r0=�<����z�&��.���uM�h�=o��4J�S�9�&����������,�7�~W���ܜ=A�S��K��uz���^�\5.e��X��M�%|d�o����p��[L���=��Dw��xY�61E�­h������ڮ0�2Ww�'z̮�M-�&�f�V��5ڲ����������='i��T��w�DcN�	���v�H!<��Z� ����1�o	w���g�����%v������ӂF��:/�~"�L5��g]1���T�}���.�o1�&��@d:��O��١R(��O$/1X�;L�������$�_�M��:�"�I�̻�5���Xd=��W�}���	Iv�4������'-����� ����,��Z�PXlxVHYEB     400     1a0ũ�C���^�Ë��t�д%5<[����=�,��vn�y�	zWUy?��D6���e��|�9/����A��|�g��+�A�h#�����@��f�Ō7�n�n.f�2z��N�6�IR����7L.F�ւ�e��ae���,|)����"�A�#�~ӫ�>�0�:9���bQ�$�����*f���am4`bp �=/�/�|�W��?_��H��m]���5Y�����N^ꟓ"� �
�a���e��@�K�k3LUx�a�7c8��כ�M?6J�J��ɺ�8�9��a����N\��N�I�^��B���XLG`Y���"xk�hM
���(ic[h��^+G)�C)���f��n�wR���>���Fm0�Q�i�~��6@���l!�.��$����0F0��$�Y07=i��XlxVHYEB     400     150��Z
���)��k5��ò#���`���.�*�����ĭ�K����xe����E�+��tv�+p�հ��s�+���K��{�H-�YӮ�fK�U+�����؍c�a����xR�^����N��yw� �U���W��B���I�LN�1� �{���(T��eʁ�W�0�H�!�U�9Q��E<�ý9�k�����40���j�J�{m�}Cs�7}s�6t�R�e�
�#U��WY�
�3|t���ˊ-���V�����A
��U��� �V����H�PO�)H�w8��Y�qD9�_��z˕�Y(�@	 @��P���}�A�[�ٚXlxVHYEB     400     190�L�{|������ы��<�K�W2PP}��փr+ �9<��ywZ�>E�z�9EUYˍ\�^z��B|��Ҋ^:�f��I�k���7E+EKx�b�l��v'���$��kۓmi]T���J�8�mh~�{�ࡶԣ����_~˥7�?��"���.�va?)-dt �.��Z�k��;��!�<n�%4�Ia2��n���&��a�|<࢘G�掘ي~����;4��z�s����$b�	Z�k�t��q\� ���������zɜW�u`�Ob8�:�A�)	҉�gH�ot�^��@�Kd˨�d������_R����U��-<^Ä��/�r�k�.��,�7�q�2(�?O�֓c���e<Eͱf�c�^�Q�e���F+���5XlxVHYEB     400      f0���M��%P�=L�҄���P�E��؅lX���O���I��M�v�$׮�t$TdK����ן��)��3�h1�P[Ӛ+>gR�2EMk)�����7,��H�r����������mlZ���T�)� �ĳ��"���F�|қ�&QOJ�]L� k�|��߁"�~�UK���4�0��|#<I%�3|]���Ն}J9o}%�eӄ�Uɂe�ӧ�"&������ql�XlxVHYEB     400     120����}W��r����̎�Sǡ��E���c�wcA����H����?[�wJM��;��ɘ?lTr�U�዆�sǃv���)�A�	�� �b'��1OBU�렄�s䙰��u*�ڒ�� gy��TY��r��Z�X�K
5	������`�`���p!-��Q����մ���-d#�}��m�4��	�sM�n�$��I)���^ ��*�3����.	r��,p�/&jK��a��܃����\-v����X�� +�ݯU�ںsQĦN���f��丰J��XlxVHYEB     400     150����k��i/�7�C�d���K=�T_�``�z*PQs�o�@��qt��.O�
�f�_	��=`z�ׁJ��kquD'�v�r�V��AF�Z�(c�	��>�X�*Iu�Īk��tK$�_�����lG>�4)��2�Z��ja�sL�d60���_�X{�o�#���N�"
8������4��ݙ�g>*�8ghl.Bg�l+��Ϸ1,����S�=���q����ϣ�e�w��F������ס��O��f�����Z[�����LL$ �RڦK���r�`��<+��%�謶1��>_u�K����ʐ�wY���>k/j��4}�)�Gݍ�VO�X��K��VXlxVHYEB      ee      70`g, "~���N�g21G�,A>�� �g�H�ST*zr�`E��~�Z�xa� �W�L\���$D-�*�|$���E}[��������K��u���jY�9Վ�!۵��j���