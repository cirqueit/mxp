XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D��	��glg�.��C�I4ܐV�}ʄ���� _�]Ӗ5��"'�z�rN���v6��.r��Un�.���Ď�#�����p�u���Zo�ʋ��ɵӧ��*z�NSM��F��e�߾����.��aٲ�H׾�9��=�Wb���e����M���� Om�X�8U���O�9T�A�%2$8T����6hX��m3r��L"zd�d�A�C��o�̔s_)�Q<�mj�������K�2aE�D#�GR��������<�xlhT�hΰJi���d��6î^<��՗7�-���Qs�)Z*?#�U����0>3�Ÿ����j��[3�t�,o	��ún�~���u7��e;&e�I�!����3�u�S8-)��DD�y2o���/�Ĉ���g����%)w��}�`흴])W,Q�-e�ŅR,�!��#�`'�4{ř�����kvt]+������H#��I��6���!����~̝l�6v3�puSy��X�ݪ�h CjJ��h����"�eQb�7w��C��Z��������h�9%�VF�m���k&��Ѣ>Q�~U����R)�J�e��uY�v��ҷOb�EY+��"6_�j���}(��N�M�(5����4
,Ɔ��sH��K|,�o_��}}��PL���us/��-�M�yO�}ƍb�bo�|?���)Ojl����F�� ����LOS/�Krʧ���A(�e��Շ9�H�twY���D� C���r�?F|��|�߯>m��e<���F�����XlxVHYEB     400     190A�x-q��p^O)R,�T��lE�����Ov�ڇSA-�힓�b�����\b_e�w�N�@�PȊ&X����1>��ֶ��Hx஗�������B��#�_�#52��O���B�3��TE���Y(�"�M�>��T���ͻª�cv�jDU|-y�V�3I���M����Ω��OE���7�z��u���1�gKd�T�G��K`̮�f�nG��wNW�;�H��K��[����V:3�xQ�Ո���Y��(�6k]�CCl��d�W��c�T�H�3J?��(^Is>���֒F��l��Ɣ���2e
cG!
n���y�h�8s���On}�)���4p�}Y���kamG�������'��7�?�5w�3��
pW�_��)�C�4�XlxVHYEB     400     180u���x���9��ߊ�B���>G�d,ͅ
��z�Ι<-,�8�eNF���WN�*>�T'�D�&�
���~�[v��P���:u�^�tc�L��h���%Ṁu��s@���R
QQ�,�?0%[��{��	2���]RN�a�hC�����['�֭�z���)sQ/Lq��s��T]�Dq�=���y��R��A}��j�J9ۯ�����0��:�Kؾr>���dOٌ����E��hI3��@EZfJ�N1�,� .���
��Ǎ	��
����"z�a@��QbqjU(�Q޹�����}�.�3��Z�L��v*�g�4'�� 6t�AՉU��;�`~��y��S��F��J�vW���('F�	���E6�*���~*�}XlxVHYEB     400      b0��S�#��')�|�t���::�mƝP�H��L�%�V���1���<�.�c�Y�N�Ē�|:�����$��s�si:��.U*��5��7��	Zk,�q�@|�z��1��^�^�c�F���l%���_���g_X{����)���2'Ոʿw2v.�q/���U��t[�t�����XlxVHYEB     400     170wir"�@h�7C�*�����) ٙ���<"�um �|;����vf"t�v�⴪�����Y�4�n���y;ll��dBM�w��&���z�(�E-ńn��\���N����lTBv3�lg�����-d����-�/P��:�Mފw��"�FD�Q�;2���q���.U,��.���	휁G��0H��	�FXI�I���Q��m��?�I��?W��t!�j\�_I�m��J���%�f����0�i7v�XBuv�A
U��
���� �	�X5�w)݅�M�&8� 3�Pn�_�@�����p�?�����1��8�|$r�;���s?V�q�S�����L�����ᦨ�,�� ��XlxVHYEB     400      90/����%A�]{����c!:�)웶.��w�_8�F/�h�~ ��Τ�.{V�o-d��dM����E�)����BrE�v�K]�����ͳ=���;�n"��v8	Ñu��^�z��=��Xc��5�*\�C��v�[�yC�XlxVHYEB     400      90 bͤ���A��2mz�n�n���x�4V���/o���q��L#��ꔼ��C�L����7���9���]g!Pu9�iG�k(e�"�Vc֠���'��esK�L���$�D>Ĺk6A����xG¾7Hd�1�n&H'o[XlxVHYEB     400      90�uY����8a)�����Oq��f��)��sU]o��u"����rjn�p]D��am*��\��h��Ԣ˞b,��:� T�j�Bv	������w�񀙁������t&�� �EM%`w�U��4 �mO�Vڠ{#�� �$c*~.XlxVHYEB     11d      50�/I>�i(J�)5��,�9f��p?1|9�0�,zGx��3؈ [�j��/�Aj����/�N���ɔ���m�ܺ��X����vD