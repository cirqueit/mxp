XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���<;���~x�2'�3�����xN�ú�
���=F�]Xا7z�z�Ҫ -F.o!Ʊ*�@dO�6^�˘�7Z\]�m �s�TA"u�� 1´"/��t���$Gjb%�'JY���؊z�a�mi�s@���54z1�m3�����3�}��ă�Lݠ��F%�e9gI�zwJ<�a0n7s���X~{�ϖ���p՗Y/"�x^%S�X�a�$x$��'��ܧ�˾t�t|k�*@�D+?2u�3aA�P�F�x�B��/ÇX��f���y~l�$.}k	�?8�t@Qyv����VF!o�r��/i��4}����]�Z2��ɕے�߫���K�(@�Br���6e����,�!�	B�NJ��bHҰ0��"b̗C��A���okR���듍;��&���^���"�5���٦g_�?\���-���6*.þC�D��+-u�˥t|W��iYsjRZ��)öo���#n�	�T�U�=���kqȇ�@���=��=��l���g-��n������.BI�V���r�g
�N�n�%��;>&^1��n~�����h�s([��1o,lG}�
ϛ���\�k��`�����8���r���; ��*���[�#	���գK,{)z��+���iט`߀�]���.�s���,_�J���2�ݏ�u���cG�3ɳ�ǢQ�'꿯"��^���A��]ज़�g���b�H��Z�1�uaN�/��h�.�c���Q*LK�1��0gW�e��[�XlxVHYEB     400     230���z�U�����(�Ht�2¹"ҋP!�۬O:��b>���6��[ƵSZO�5�>׳�Ct�B�s�������}\����L���6��|AadNF�^o�ꏤti�,���tM��s�	�i��U�fc�XJt�l"s:+�$=Kq�q���
Z� 2($��{�f��c^ښk��Z��Y�%
ǽ��]Ns�
WRM����w�I�؇�_�n#�+)��`��1��#�#�٪qd��^	oi�+�ik5���N�MqA
w���59}�p��a2��C=���bX*�7I���rr��d�P��b��[�����*I՛���%�wZ�a�-	8��S�DKYW�ٮ�hҬ��A��	E�L������$"6ɰ ��12�f�k�8_"Y}@����Vs��Cz+Uv�}�ߞ}���b) �m}N�����	axΧ������31�����G��W�n":£���\S�_b����/xj��E#4ă5*�bяP���:�֫od�э���1		��w-��{���'�`׆U�i	��sY-H��Ɔ��A��XlxVHYEB     400     1f0n��-�<�2������`�lŸV�$r��kɾ����}�'מ���%��F�1�K�Q�����h���Y��b��" 4�	���-ܠV��f�Fi�)� }f�=%<�M�">��8�7,h+�_�J�a��Yo�M*��}����y�����h�Y5���F��V�U�����Wh��Z�Nb/σ֏�1*�EBNo��8��`2ub~��[�f�g�U���9��Z� j�HU�Q��#�?�_�)��w��t��'�#A�|y#1���$�6�m|ۃ������f�eZ9_����,`8$D|��0����Jtd�u�tRv-��%�d�M��i�nR��.Z
�	�3p�Y�4�9�{�Ty,P���9V]�R	���W/m��<�J薜�LQ�zgXfrx�-�An��� ���ⲳeZ�R��a���*�r�=��4�"
��C���3SI���m7u � Ë��X�Ne^��M+���Z�XlxVHYEB     400     1b0���N�b�y���@���ڀb���B��r��5�]� c�1��|_�dHEcY`��O<���|��s�{�5�2G�|�$a��E��<���kaaE��.f�4��\C�d}���(^+�l)!�i2A{�j0�S߿�����%��Hj��@�we#_Yw��3{
,��y��YЭ�9�SpOS��߶Ѣ弾�_���pw�Щ¶��x`pDd߶}�jf�rԯ�G%�W��,�,!qf�dC9��O�c%��aR�i\aG�c�	RL�a���7���t�
a7�������t�TwKۿ=LbyT���X�z��ic��CgC�6�Nv �L5�
V�č:2iE��,R�H�q�=+Wl���2Z�"�s�.�v���8�n��I�tCo��c[ ��ٜ���z�9��s��[�! �U�(�I�XlxVHYEB     186      b0��+�΀%+DY '�L�����~�YѺ۝�yU[�!/���q'�xǥ{Fф՞cU��%:�Ȕ��v�L������8�� ���rC�%���B������'с��P�yit*�у�Yc~��6�Ӆ,73 ���pOO�T�_��/7&� ��N���x��