XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����j��qc(�>�U�6�ה��3nHwy�NY{){q�,�
ͺ[ψ�M�K3����y�,Z�Ҥ�jp��i�oD�&=:Ш2+<�OH}��xr�ϕ��y����B=�Y�]�=*�{��V��c���
�U����ʽ���:�!�5]�ƹ�?��i��R����VO�n�l�&�d&?m�z�& �Z|�@}EK]sc�i�"��J�9c�&ǁM�a���+���g�\�V�����d�K�vQ4���BJmп��K۶�����������v?���LA2g�E�;j��*W�����^Lj�oE8�Wo����o4�2��ΘG�|����^�N�$��H�5�M�Z��9���K��N{�jk0a������������X̴K[H#�Mbi��v��<A6Ȑ�f�hz���7�A���w4�uR���Ǆ��%k,��9"�������v�
^8�[b�]ƿ�~-��`i���!����}��\:�>� w��Y1���{��*ĕ���w�lI8��Y�8m�b�5dD6���dB����ukɊY���䕔��vn�����}\�DB?
�xi��(���!�6[N�2�����WO�qp�3r�H��h�r3�����Z��j��C�fB���B��h�u� y�;Y�YkǑ
Ma(
�iB����l �>�}%a�_$���j���6PiR�\i��`>�EI������{���a�
���Ɯ�0<m�^�hJ��7�a���A4~E`w/�cT�c\�9LiXlxVHYEB     400     1d0��Փ�A"��ً+BB�G�=�!�o���a�I��C"��+Ҟe�?�y�Si�����`�C	x�w�)��_OY��F�#Z.1�>d�dG6������ק��hVg4�4��K�	��(&�E)��I:)Nq_�Ƽӱ����Pq�)i�.r��[���f�`��X��I�H��7�@+k�}9��M����by��Y��r���pH������Lw��� �s�׆w+]�!��<��9��-r�/m���&-�f�3E�f옴�m�2l�*>J��B�л2��"(�hjZ�02�<*��"�<C$�"lf_m��,7�b�W�أ���>��v�tf�&��l�P�}���~�l!���%�SŋoPi}���H~F2���P�^�E��B´:7��s���R�5�Ah൛MB]4G���w:�Cg� ~���F�N �]�c��(�W�k��Txf8���+�}�pXlxVHYEB     400     160覝�be�g��.�	w�}T�[�jz��iMզΨ�����4�_�$�]��JM���n���X����;�qY,�
#�V�ss�?*���"�X�<zC�5�Ny$E�t0�}1��]�4�_-���oI��h�
��p֯��*<�]L��L�@��o�ӯ�t�}��6��&�V6�����K<������{��w
^�������%ʍ����f��ǭ�����	�z%ro�,+iv�w�̢VCK[Z�_Iu{&wڈ��I!�42��4��3?���N Ψ/���I�|aQ18���c��&�E��S��B�P
�1)�`�f��fB+���v?xǑ��XlxVHYEB     400     110�u*f-A���z{���\��o!c�ߗxq<�E���B�/��w��C�_oxs���ĂTA���$-4U��A ��l���*¶��<���`2�喃w!e:�3K�
��͜��D�O�@�@��wص��1d�K���yR�qa�qN�#x��HR��P��f�Z��y��Ͷ��w�E����3��+��uL[�=�������f�l�a�����S��> =k�Ht	T���������_�!a̕Y��,v;ؑzd=f�w�%h#�XlxVHYEB     400     110G̃d	�բ���:�w���&�e��㠯��������
!��ŌN���۔��*i{Ez(F^���!i=@�����3��ҹXA�����ڤ�����ʐQN�o������ߢ���FT�a��q&�5�EQJ]�Cr4bV.R-G�wx:�bQ[��T'�\�Z���3V%6T��
��5�+�,v�׻l�*Ci��s�e�9!/':B�Dp��h}ׅ�bI��`)��D��x��ěP���|p��π*(ϨS�XlxVHYEB     400     150�c�8�M�p�T�7h������5���!o���`ғT��[r$}b��W���oDy�+�ȴ�a���K����m*��{kM@9�@���j�tLZ/mJ#jkZ�!�۳J��cs�T�݁���8I�\J��#lsVK'λt]����U�E��F$ʖ�BJ�ni���z���<A	z�*yp�i�$��8d�kIVm�:^a/S?�KJ�H���7�R�l��gp�&������&�G�ظu7������L���e�4������Q�iǷ(��z�l�'ķi�"�Rغ���#Z�wϔ���A�L��q��������J�k\���+H�]md�p�?��SXlxVHYEB     400     190ky�����:���s�H�F�͟H�}���l��p��n�\*A*��[ iG/$M_�W��]�ІS�i�#P��yg����ђ �R4y.�@��]ʳ�P��>RP :�~t9���c ����ٙGF�N�4eꔲd�c�GuѪ��/4�a$�F`|IL�1��[f�l��{�C�Vm�+zO��5�zo����2:�l�ee~fG�
�������m��75�-���e�)Wp������V�g�� N�9��x���TmM�:l,��Pf��X�t���5�~��Y�YeN �y�ߗ�w�'(�`��o�������uN�,�������Iܭt��鍟��%y�yM�?��H��ȓ�����b�'��Y��6ĶS@�>�Sa�ڹ����U�Y9�|��q�XlxVHYEB     400     150�2T�n=��i�󥤤�o����J�?�r�î@`�e��j�=��Jv�
K�7�g,U����W�u�i�rE��6�Tz�1CWTC�� �����Y�K�D��E�!H�쳢�ɘ�����-L�0���ygJ��T���8�7��Ņx�H�� �[�7`\Y��kB%���2��*���Y�f�9L&]2���Y"���c��o��
�f�L����W�o �̶:��B��Z���bvk���_d�	�~������tI��j��c!d��~����_k���8�\(�taAO ����~��8Ƈ?CiҟL>u�����j�d�l"C݌Bd�GK9�Ql�%���m/�XlxVHYEB     400     160���NAyO�ծ�MJo�>�	��otQ��<��44"�h��p����G_� h?)o�f��%�����ջ5����l��oR�/���3���ZM�L���~FF��"���<���>N��x�r���x��+���Ƒ�|q2�XQɏ-�H���Y��!P�f#�w�U-v�I��}�l�^g�_o�Z��Pq	�zj�K�4�)R�q+�� �^ 'hP��q�5�� ۖ�s��T�7�à5�P q7;��"R��H�*ah��*^R#O[�_Y`�2&���yh� �$1���]i"c�\�L�nwR�"�>d�d��T�<+I <�x�}]I�L���fE��^SXlxVHYEB     400     120.�(e�A�P��O��1m���,���G�3���Q�L���	o�h��i|a^�(��lg��Ԛe�7���3�e<�������n,Y����`j���\�_	�%���z���_����q�� �t2i���Nڣ�L8߲kVm�*��+�i��ʢ�q޶�zzյ�w�`�f���QY�2⬇��`d�h��7F;vK��5�cJS�<�*�MI��"�h-т��	�-0]g:<��m	�Ժ\	�-^b/Гr׎�i�ؠ����G���kk���'B����gXlxVHYEB     400     1b0���
��G1:6cw��R8�I|,�Fg�}�s)ַ�-l����\�Q��j�U?��,i��[\=�_�غz��+���檌$Ɨ,Lm�Zg;��XA���-���N~�s���C���m��*����qd��j�g"*�<�@��>���X�������"%�e
�"����:���F$/�-c��q�t����ÏA�zK����;q&����B�5�!�z�W�v4�V�1B�E� ����s�gi��#�YG����'P��l��!�܎v�ڭ�õ�����1����XD�Nm��/�"S�f�0%��FW50�ئh���꾊�ᬖѲ���:����	�ókj�X1�4���h�������`�{�G�Go��EQ���g='-��˹�V�j��oB���6 !�G��؀A���
_C���XlxVHYEB     400     1b0��ei���>�S�̙,L�� �!����߬���k��<�].�2��q���pY�u�xz��V[ct����H�w�pyA�$�`���X0���Rg	�"�%��Q��_	�
3+2�W��r|0�mK{�xTaܡ�M��:�bPƒST�w1�лNK�U7yٶc��A\��s o���4d>&��ဲp�^�DIh:ܭ0	���s�(ܴ�,Y7��X���m1�����>=Q�3�������2vI��u��b(Z���[���f�x���{J��.����ܞ��Id��9J�R�j�8x.�1�R��w�u�S�c�q�K�-D�)��)�>T���h����7{ʽ{vfb������! T�6����+1Ġ),��V?1PǬ�S���Bzͣ�_#��P�o�!+�Tϻ��P�>(|XlxVHYEB     400     180t=
j��'R�� ����k���yK��Z�� u���fd�!���������㳅�ӣV�5B嚊�9_��˺nur��i��n�e���d�Z#fp�E�R7�<�͗Т�=�Fo�
pd1���.�b�]e��I-���1Q��ɂ�T��S����e]�� ����3��$Wmp�R_J`�T��_�/�a�#�oL(��V7U�)�y��x�5��6����K����PH9��ˬͧOȇ��'̿������s8��X�,�C�i%��e���lDL5�K�z5�N����_P�@�׮��/䉭Y%��Ң��E�'�m{�':�s������ �=}Ρ>����
P���I�7Zp�bFU��"O&>(�y�:�zG(<lXlxVHYEB     400     170��ZZ5�(:���}�yv���M���9�Ju_^��\p�O~-Bq�z>��t�q�
p�An6���"5΁���Abm��;+2�3p�Ɨi���hY�q=�W{���T،�Q���h�ء�����:>%W܍�5�X�a`�_��S�=���
-h�����zd7�Q�D�)������B���>��$���@�H�F�T�^T���-�\����.Z-VG@�ǖk�G�s�YMi�u(�?����u�Q�؆�y�|��bg�\pB{?E}1HgO9F#��m	���PӅO9��g�
�.0��e����hN\���h_2���[������*=R����J�����RA��ӔL��$UG����XlxVHYEB     243     100��]pY|;�P�F�M�V�m�҇vſ�fj��Q��[��cXY�Zǀ��{�����s#��>�Ẁ��3�k0��|s��لՀ������\�x�u��`��U��>A`9��q��\5�IZr����7���[��O�h��1�p�sBԬ������\$��:)<U�g�_��O,����R1˘j�g��҅�D>)��߁���8W�p�*q%Y��yux�%�?3�X|Ov�+�[��W%y�+{}z