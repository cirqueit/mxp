��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���:��1.f��k(���zp��'��FL���s���n}ŝl�+6<xޱ�t(�  ��۸э�#��Q���/��Q�}AlM���������-$4�߂�Xpx�����RԷ��p���r8I^͹~��F�C)�bC����R���S;~��׶�q��A�ڋ��؁,٦��:���T��$�Wm���Ջ�m	������<@욉+.�k!7��?jv9���xF�TY�)�M��(����i�2��;V���B~����ߨ����C�����^�߿&�<
���ײ��w���E ��Ӄ�q5=c��`��ڧ�ޘ���aO�%�ӽwC�-��gZ���)���-�Z�~��2e���!A��[�foI �!y���=�s��1����}��ַB�>�
N�D-�����SƗ?����@Fsa�b��#m�fTV4��phix�
>OH�H^ᾅ��3\�,)Jm���Q��`�È e��!��dM�u��D�#aֵ���>~2*D���)w��w7�_�U�`�!T?�+�lĳ߿ۥ����R��w��5�����^�.� ���L�N!��k/U�C��+��Y�8U�L���Ng�@�މ&�r}Z�ޛ��'� ���F�U���I�jq�;2i���5G��/n�]$ �nʮ�אTy����tPl�Q$b7R��yJk`�SO����-}�e.)v8��/�l�O�zo:}왠�:H�l��:�Zxu|U1<U'����x��4�{�p��j�>�di�ZN%��蝵�o�C�Xg��#�[y��̠�B�%���T�]WC�4g���k����vs�W�lA���?�~�����FF�k'���}�թV�6��jrt|�aW7z�G�yb���薥N�֡���Q��8VL�$! ��i[�h�q�'�m�F'R��,�	����=.�l��Q�LR�PM��փ��\~�E>+��U�J��7�V���z�G��n�a���J�*�H�d����Տ��V�p�l{D�v���S�'�u*�9��z7��N�X����-asg���X�"��H��ן��31p�\ �3�B�H9����g����XK�_ �	����n�P�]@������|85���&�d�����@�k8B�;�X]e���IR�ŭH
���?l��T���tY!˵L�����7틭��
��"��4�ʊ�O��|f��\��7�ޅVy1<�Ʀ6�],\��q�kh�	��d��oƹ_x@�z�/�[Ǥ�O[�mu]�;9�#[����-*�f��r SZ �I ����'5=�-w���o��N��	�tx{�e��t�!�C�f��z�����h�����h/����m����v�a��p3/�W�be��J��)a��W%��T���j���f�ٙ��plE�c]^��<��4j��K蘍�_��Oa%Zs��A���Y.�?r��;r䂷r��^��=���j�9`��u�`�t�Mb��q]�[���� ��J��G�:�_h�ݣ0~@LKw�Tg���F�%�v�S��j]:@w8IG��L�x����K��r�),�-�4�F��0�y��u��gn��"�ȿ@����D���%K�m���#K�@���ʗ���ZV_�M�6z x�q`'|�F�ÿ����>R�X�X��n�n�)J���'���RYO�8�tZ�'F�K�ª�!��D���&��f	ɱ͛�K�>��<ԟ�w���	�;��`p�v�}���k�,������9�N}����w�fV��Q�����5}s�����	Fk]cZj���?�0�LY�c��.��d��Jr#W�B:�}�}�OF_��05u�5M�ď�s�Y�z��+'z�B��ɹ�b�^t�.u:�A��Me���ڐt�Fz'�`j!�3(�C�S�	�q;2�(_�)��G�	��,�q�|�;�,y̰d| HƄ0�r+I����)Z�>;��_��i�l�k���7�n�:��Q)م���Y��F��Ѽ�ó��S�]>($���R�_1��l�
�!.i�6є+���3�D�bbM��4�{Ya�Q�t�����K<�\*S���%�B�R 
҄7�˽�t
 `w����D*�%s�4�3��CWG)F=;._�ܑ�Hd�zw�IM��c81�B����d��r<>�apm�6�wX�M�C��'��}���7��8�-��\��o�Y:�؆5�n+8Y��lD^�,�#m��)�w;�A�o�q^ͤ��Ȑf\y�v]疾@�;c;��HK�5�f��@K�O��]cKuP���ӟ�MK^Л:⹙sѕ+5�咽�u�ӝ:����W0�݂�� y�D�(b�o��r��V�0�X�i���"�&��*�k�c��j!�ˣ���E ~�D���lC�t��_%�}�G%�E�gj�n���A;8��f��1��!�"�K���&��x�o�C�����x�a�'D�$м�$Y;�g)n;O����6CF���W��R��A����'��\�Y���i4r�3�Bj#�+AEҢFj�9�y>�`s64"x�IRAk1��%�Po+��7��/x��FS���C�8G.�k��� 	{p��+�7�d�^	�<�]}�k"�2@�κ�h����÷�Țر�Ŋ}g��L[��įؠ��RX�HqYٜ�f�h��.}tE�k��PŮBu:����C��&� ;?r%�3&{�}܍x[`��"�"�	Wa(&P+}�����ı�L�iMte�/���ZS����8�'V�7���x�r��v�h`����i�>�e��.Z��<�eil�����Ӭ���?49a���+sC��S6�u4�c(���ޑBnc�4r�i��/�[��]��uř����w��jJ�;1��s�k�%Ε|X��m��і]Z�����iI��Bq�r�N���C@�iq/"�҈��Y�l���X�4Z�������5���C��n��)զ	)����%|\���;l���$?i[�ϤI���V�������q_�'�j�y�!.��Y?:9�j~jp�?i�f�!2�pI�5� �k�y��"��V��.�Ɔ�P裂S~d[����l�Iv��v����d��	�6팱+
������_-T�и�E��s�c�YT��{�r����) �>�O�����i֘�����p�-��W��jꕿ�R��)6W3l���{���o&��w�G��b�� ���:X��C<[��Q&zA�} ��ڭY��~��a9���z9�nu��`�"�RzB��r�Zb3�c���~�8�t�	US��郯��)ݑ���A�Fx���]�����rd�G�x�j�y$�8����`��گ�f!���E���n�>�� M���4��-p���ē��9C���I|J�2)��`��L�	��2P[��32>��F����_7G��Nf%GJ�e��9�S�-~g#u+Db*�f��eAv>��w.���+��b �7��_�P�u)'��T �վ�]B窓�
�2��7�a�yR$��}J+��Ç��p;�� e̲�h>h���ܸ�x��xa��J��YV�v!" �~�~�^��Z��`=)�/*aρ�r��;�Ă��NDÇy�)Lg%z��nb^8��#y2GX�G��y �MP�������,.`&����b ��g��x�}�z�uXu▿j:�\q�SP���I3Ӏ+^�'i�%�x�x*�e<e�xw�ȍcM�3��"�5�hZ�`P�45���:��j�KNA LpC9˧��kVċ*t�RW��;ct?H
<���:޲�1�
��5:J��ag���[0NZ�dJ+D�VTzX1&2v<[̹�y��C�W�T�v���vǮ���V���t��j{��/��R��a;����0���VU� ���Wܠ��/�A/|���j`H�i��DB�r-����p�s����1P��.�s�?��l����\C>�n�-�e$�T���~�1��=�B~��V�mB��u�y���y�~DV�H�,\�JQҘh(~��]J[V�����2ޅTZ��%�$2
�����pjp��;����� <3ި�$l}2��b�A�ѝ��i-��y��}b�ycW�b����d�|���\�|��k#%n���f��2�[�{	[Χ�]=˱�q�ުl�4��mH�LHH��1�x��	��;[���P�|z�#��F�<gռAT��_�l�mܨPJ�g�E��fɼ���ϰ���'��AƋ@�;5��_�u�S4R5:�z�.J:.�*��,��$te���jMƗoꭝ���/�QMƇ��ZU�d����=
���wW��ҝKpID�R�fÓ�e}7����y�=�m7Q�c�/\��!�x��6g���5Ӭ*�GFsn��Ȯ���7��!�LQ{�Z�^�yY���l���l���M�S�)�����D�
K��R�UH��~D�sIs��7l5:�FD�1��܌qy�2[@���Q�y�(��ss��j�D!�.�51[dK�꾷8�>ݳ�7y��)KϿ�Y�\��H�����x��IC���lBOX�B:�~��4�\���֛Jx�ɷ�B��v�A��tUy��R���f�zsA��$Ĭ�U|T�q~P8�@��;�g�4p�۸C�w 
@7�"}��uM�i��Ο��<P,Hcg쳉�Qd8�\ז��z^����s0Q_Q��0���fН��tl����ݚ㵭Q�Y
�]`uf(��~c��SE���%�]P�S닭N��"L�/Z��sYM�*(-Z�cG-���0XA�u����<��W����ʭ!a���ӴJ�:���υ2 L�I�	'b�5e(�T��\��T>��<�i� /������Q��[H!|^mW��8_����)��a�c	yp�`�*Z+^T ����?�rW���)�9����:֐�7�uՇ*nR�\Y�9fs��b�� !��"�scE�n�Yԑ0�-���v�y�˨����
������!:F����wK�d(�����$	��`��3�t ���r^�I����eD�\oE�����<cN6�e�XAs��k�+z	>Kךo����1��k����o��T�Y=+�,������f:Rʩ�!Q�d.	������"�,k�ٯ8�L��G��=N�����8� ��Ҷz���d���2I��՟�Һ�L��v%m���h�����%2W��h��Ⱥ�`	)p��hض��ƺ�l�i$���f���}�o�0�=^��a�����6,��@�B��h�Y	E�eNn�	?��;��ErNP* �
uvӳ����ts&P^6?��G��\���|��^��<�L|_�.aL��~�x���ݦ��m���N�+<lH�Gcݫ�F�!������d�.v[�3�T�G7t�n�*|-�T/�N��5ݿs�[��
t�{cK`M�K$|KQAa��ڗ�>{��s}�:.��)4�-�c?I��ű/D8uˢ�l��V5ߞk9�«g��-nY�Cې���4Z)�{�|���e�~���3��M����`^p" ��d�m'Zq��D��h�K?���ҵ�cIXh9Ȇp��fc���oaZ�(�#G���(KL�s�q�F�sJs��Փp���a��0?�7�=L�]Xӄ?���gq�����d.i臊�x�`�)���Q$��.�oCGƹ<����֕���VHbK;�O�
��JJn��'�_%R�5��nt�ZJ�Ny�C����K:O�V����c퉯,��o���0#R⮿b���o�>���92K/�}c~4��~ȴ�7�7ݻ\��+ʗ�0���"Ʉ'eJ΍R�#	����WU�]�M*�K,�<�pΑ>�#��]�ֱ�23N�/�}��7���3F5���,�ˊ�w^՝O�٧KL��ϖr�<����	�����V���a���G=0���$爏9Zg�	z��?��f1Ԟ/�j�*���l�dQ��n�Q[�Ŧ0az�L=�q$��Hk�gQ+Iq6�I)�P�v"��-OoY���f7��}|]wҴ��d� ��愗$����e�r�쳬e�7�}]*H�n��ϭ��8��T.zQ�����a��vOW����(*q+*�h�)E���0�f�z3XO�?�f��E�л&*s��~)M��G�4���ܦ�<������X��67�t��Z���u�tB|��K���(����I%�=��7��e�b{擼]�]f�l,��ѱ�3vO򏢺,(S���p�G�_j�.��P3]x6��\���
z2SJí��xA�G�ńn�PbE �M2�i̘ˎЫ̷�y��A��	�/?��Z�C%�I�v2�"�XE��!u�����*9SF0'w������FV�C��]��w�����7��=�.|_�FJ!�u=�q�>���>����_a���&�.��z���w�?���]Q�
�<
C�+X�r�k�o-�I��M�g�����T��#I��X��>r���ڴ�ҲKZ�	7��/��Q�Q�L�[�e����|%|jR	����臿�xG@��8FD������f�ݒ���w���O�:���X9��Z_ŗ} �I�pɮ/V�R�V���T@AD�H�D�7�n)cS�o��4|l�^�*��ϋ䭢�|C����W�k�'֎V#>����N�L������¹	���c�5ʿ�~��ܤ�!�06�8;
N�X�?/�~FȪL{4��ta'p�K������g���\ڳ贝��F�Ӷ�N�.�uw.�D�ZO,�M7e�kW>�[2N��o��/t)+V��a^?~x�/�'~�˵ǃ7�'��o���qӃ^��ܓ�$��m�8}�,��rl��&�k�yC�ֹk$PE��`)G;�{7���X���U���y�X����׃�`e�p�'*\Mh��Q��)�oT�������e�<q�W�ʫ���!������K.W�%%�~\��<�Y!����E q �t*��s �P��;�sT%*ro�	p羹SAw��8�z��ty(@���,2b��׾��Y�)��ۗ���e���A�T�����9H��?M�C+ ,�yp"Lp˩V�4|�ɉ���o�"�B{f9,Lx
��¿}��Mc���Q���B�Д�$����Q�0MKB�Y��1� %c`> �V[�wG*.��X�</���t�Ϝ�~� B��
UM��D&�2O�8(�*��K2����Q�N��U��m�q_lKO��p��#���,+f��ף���o�Dے�?��5��A��/�MGSb-�T�j���.Q��I�ou�&��/�����}�!��&}s�ҵ�5gp��fvJ;e�X��Jx��Y'���º���zfC���-%r1��h�6^��qrR2�����8� T���z��i�;�/�+��T+�ڴ΢�'C�~�;==�xw]����%��!����F��:O߶�(���O&M�f�K25�5�H^����9w
�D*��:�#W�Eq�	4tm�3�(e���FM�l���r\b�'��+%i����2L��������os�����Y,|�����������;�����Z�\Q�ᘘ.o�(��kD0����[W�iMKx�,_�'i������1<��8�(=Pc<���Lo->��J�*�)�5�e6���Cmm٫t��k�Op�^~�Y�oU��5���k�>(�n�y�y"�C����]�T0��i�����׺���5!]@��������?x�����75j�P�k�T�A��.}����Q�5l�UCNl�(�v\V�R�� �M��L4`\�ЋݮKE��%�na]���th�X��
�2����!��t~��7��7Df��u�I��O_��N�����5�����EQI�s�E�<�C�e�_�r)N��:�6�YJ��L��H���{KD��*ӮNpA`�|��C�.�EI{���԰@�M�b��/p�{�D�$#웖��+����EM�M�B~D�V��IKD��h��"�n9�p��V��|������9��!��J�{m�}��a=��v�����- �ř��%F~�@��M�������t����͙����c��_�x����I���s����QA���L��E�[�Q�O�R/�ޠ�����oͷM�њ]�S�Ě1��axdA"�^k^:���C�I�|�.��Z��ͼ����!{��=^�8�0�{���U>����6r
�j��h�~Q��	�G�[ʒk
��dr_�h�);/[V�b���z[;<��W*P�u�M^" כ(j���~ �2�kMOA��� [���w��cԲFT����,��c�+^��ys];pu ��:H�3eE�����)& -��꒺�N%��o�U�#�n��r�"�#-"c[X�� ׫���T<kj'�Q\��׮}�����tu�iS��9u��Nn8FT�e�f֎�����=�<eq�%0�7�Y�哔�hX���O��R#�����<����N]�Ȯ�\��vE���F8T�U�ZΤc�'����,˃ՄZ��G�J �yMnV@7"����,�C�������C�%ƕ�b��3|��?���~Yl�$��ע�򈴋ic ��ɝM�W�<��%���$���stOԈ/�$|P�q��e<BPӹ�A�3u���$S��=<�'nj��ı��P𾘢]�$d��vK�HAl��IQ w�\U��@��x܌�!1�[�6�U��n��=�oM����� ^,�FG�We�*-�ˊ�IM�
Tpy!Vf_�\K��<4��z�|�0:ԁ*`�7�k^Gk�dC!���m�tQm�W��i��|��q�kL�#	w-��Me���A8�]���8�UOb��6(MJ�l;i�u������6��W�������kw��`!G��pe絗��z�ǲ�?���an��F����#����(̣H�e6&�w�-���e�ͪ��c��Њ�5�����rĕ1Sc�LQ�`	Ԧԃ��>�	0С��ke#�E��b�Q����������=V}pĥ�!�!����ms�+�ЬK�5&�6��7
��;���R�u��|�P�O��z�8k� 6?����C��J�%���d>�ɫN�^W��1�;�ѽaا�7 A���6�����8+��ΩǑ�Z8_|C��B�\L�,be�GK֋V�o`�����;e���0��|���k�Dv�IL��Ny������MOGfA�x����nҌ���'O��%4�#�H��Uz�g8d6�$�R�GZp��K%���H[
���,^�B6���2�����o1����Zm��M]5��������mZ�(Ώ�KLJ��X۔7~���90{ Z������x��Q���׫%h2�q�˙�m者 ��}�jTb ��*Vag���oQ��Ӻ|��� P��\�.j�_Wq�q¿Ct�p�O��[�G3�Z���
X��%�g��M�\}�٠�G��zD��v`�$�(馔=Kf��QU/�3q��W��̤`�ߤ�@$��\Ԯ�/�ûqꗢ]�z�r?�N��k�_xed��!�6m5h�Y�ݰ ��e6�ԁ�V�/R���b7�o=�ms@�j.�Nޘu�G���\�#�H�K*~="/�������&��y��c����f�o}��2P��3�#���{�kb��}ߔH�b!��=�ݞ��wG*ݶ�演�5�ó��c�L�#*q� �Q��?Xh����PkH%zi.���y��R�C�W5�`��&�=`�o�J�%����U>n��w	^A���W��}`Zՙ('a �L�����L���J�N��3N��;����7��b�T�H�{9��ɰ^��!:M���4��^R<��������ϯ�Ww�l�q��>!UT������� ���s�e_����:6�N��t��I"�Q��g��l$.vQV�H�N��[�x�OWf	d6~	����b���Ki�^ ,b��ՙ���ꃾAmU�O��r��Y)'��h�L�h�P����ب��K��] 9J15Ri�g�6r�t��Bcm@�f$"�˜!�GY �����[�I�3�OM>��5��ᔐU���7�}�����q����m������&�,�R�J@�)ܘ���H��m'}f��g0�Q�`|H��sd&/g+�����F~�}ԗ�=?'b��Ey>�żI���x[�p��`�������Q�;U��-~gX#H�0��-�]��d����A%2@��������M�ۚ�d���}�����T�23?��4���7�X��Y}����+*����hu
��(b���;t��V b�����������t�i����X~
v���.�F�l)�#�j�}�J�ϸ0>r��*A��4�'Ň���3���O���:KuH���Dv������s��H�.cC��7G�6�@��!�=�:��c���|_
:��w�Fз�d��am
��]�*,m�)H}(��a\��Ͳ�e�[r8_3u�	�3��;TEq��bmTd<4�Ţ����g����5�aR�����4��v���yz���?�!��ǒ��򎶰-y���{ �6�S�`G)�v B���c!�a�j|����q��O�7I��ѼU��Y�l.���q�ۓO��h*�ڹ�Z0P�<w�Qe���}ɼ��D����$`�O�=��~h��aߖ�HΔ�X���V���SU(XF�z��8�p������K����l��-��B��[�����b+\�繛v��9�X�����f��D��\�����mO�+�w�y4s���,C�����}Z#ts��G	�2��ڋTn��\�?��Vq*ʢ~ g�c�P�˜�_J��S��O:/q_u�!�[�L�̣XFlwK���w�u�;X:�0F��Ф4�]�.Sh�g�}�Y2Mk���%��4�m�R�L4����*��X����+D��OȒ�	��S�>����PSWc�b�`%��BI9	*���筆D{óTDK�K(D�W3��H�����M*u��G(�����a�8WFv�8Mr�h⁍vVX��Џ>�5m�(c~����l��3�'�������O��c}^�:d�K�8�B��;�D��H�7)�zc�S����$8w�4�Z�T�d��.�Ûu%U�W4;mWņz�a�De��L��.n���I%;t8]Up��3J�%K�aZ���u���E,UP]gn‍w��P�i�����J��*�Y���g�ﲱS�;�ʬ��?�0��zEs�z����k[A=�^�eX�Jd������R�[A,����,�9�ٖ�mLL%x��PL��p6��K���">9��s�XO"@�:����n1*^��V۱v;�xs�g�$��Z��㚩a�4�fr�Q�x!U�FB��WÈ`G���~S#�\W�D'�����8ns����B�4{�'޵�7ᒷ���I����YST�D�RCW�����.���+�/��� �ܢ�1Y����"��1��WĹ�9�`X���P��J���k��a�aC��:_�Xܑ����0�g���wKS��
Ќ�S<��Qp��zH?$#X��nsu�;��F�G�W����ʉU�+�{������5W����D�o���h�Û��O|�R�o�pr	�.{�pQ���U�%H5aJ�r�����p�sT��%��nE�F팂����GP}�QKXI�G�4��g��g���4�p���\�0X䉞��`GSp
,N�����O)�:��P�iWc�>7�ي��8^/��O�a�o�[�f�a������E	ϼ�u�i�.z�D�r�v��j����;��S�C$0^���cֽ_٢�Z��y4`7�ى���E� ��{�s�﫫E�2�"�S�|C�����C�^g�';?�9�bJ�!R����{1�[� �QE�:e5l1WJ��I��!�XjIh��j�.u��T ��GE6�G3X�aT#q` 0�-S�9��Hg�BAf�	C�������븖i{v��w�I�9/���j�j����Y}�3���-�,`��H��!��z�`R���~��d���C��2��'!�����`�Mk��Fߌ!��=xV?��V$_:v{T>�rhc�s�JcP��r�g��*E�2���<n�H��?g���J$;U�aK70u�z�{]9񭡕&��H	�*���z:!^��+���=����SJG�zFқk�w:tO�Ժ��O|�T�竹�g?����(��"vc��;;�&��9�ר��I����a�\h92�m�F��]n��J�.�������n�4n�Sd��ƣ5t�~$����~L��&�{4�=��F��(NJ�f��5���s�Y��P?���NV��_�z�c^>>}�}�����	���e�Y�K����d����И^[.v\S�����`����2I� IZD�E�]ݹ���%h�ڼ����l\�&�5�C�����f��~{�T��/�s� �~)��i2fw��i����3���;�m*$���֟+U!��g�L�:&�[���A�nmERK��"�42�߼�閍�1�L~�r���W��o�q�Be��n���W|��"�9���W���)�����II�#����*�F���"e2Kĥ�&�꺎$���&\�v����|#���Cz�t��+n�7�j%mFy�%upǱ�<��{K��*G��Q�x��s!+��8M�挨��2�	�H�@ʉIE8�~L�+ �q��n�������W�+{�]���86
�H�cS*�����*QTw^�޼J	 �GǱ����?�J��5t�Dl z'���]مsT�l#MY�IUx�l ��
/�>�Q����z��	u���(���/�d����4ȁ0�wQ7�\7����A�[�u�$�$�JKh<�6������ �y]�R��忖��e��ǲ-&����Ny�� ���Q����C��^ccҜ�.�,�j�uФ
�c|t�$qi�)Vst�o�4�%5��M�L��˒1l��`�+����QA��*�-,̷1��Z�c�y��#�'���F%�|W*g�`��g��w�ֱ��"D�1���-�lX�����f�Z�lP'x���-�5�����S�zN�v�\U-Bq�<�*o[�9.l#Tn@�[���Yx�hrI�)��Y=2�t2m�E�AOE�+39[���G�c"�D�$�0K�h��W����mh���v7<O�R9���$pC붋��%�=��Ax��#�/M=���Y��5���&bV�4�!���Fງ�]1q��.�Ց�&�����	�ɩI*p�v&.��`��J�?��輅Í��2�1��?�$郷��WQ�0#h5��"��Y]�1)��7�UF�
�����-�,*Q��	�����%���T��x�3�<�h�SN>V$����)����(n�&z᳆�5����H݂��<�>e �5�>�3,�}
���+�fi.�:��<K�L�߈�e���\:+)S3�e7Y�}/�f�b9�|��}���t/Y�[M�O�&l�r��/�����@h<���Uin �{6�.��搩�v�M� |W1��jc������{�h�s�h-x%���/2��^6vZ��2��bl�+�<��9�|�[�&�CDFP��O�q�A��V�?���(�`c��9�7����m�,�C]�׃��n̩hzع\c47Y�7�2����JΨD�0��J��5��R�����rOj�ӣ�����վq���,�c ж���]�1^~6HT +���?�Aq�F�x�:4F��A��h����¬��Slǫ��f�6f��Έ�hiB=}��.�c��z�b�;|��w��*"
�yB��4�����q�d&�/az^�����]e�r���P�F\�,�s��*�%���vG�R��`��=�b'���K�c1�d���+ɒH�l�u�n	6l�ބZbwi�ƒ�Bf�~�b�uq�oRl���*�1�LKw��ގk��m@�}��C�eq4���*�Qmq <�hD�+ Q���L�:3��Q��t�&�6����/R�:�옹�6�a��»�;_?����cs	��d78��W1�u��f����ӹ��D��(����J���/���H����jx��+*ŁrЩ��!������o3JdJ{^�rZ(j�\(�?˩�9�����h����5��T�V�W>"�K� -ک����!���N�gZ�ؕ�&��<Y$<s�V]_䦍��T���<e��`�涇�mn�D�c*s�xD1��s��0���&=�vÞR�U'�P��T3/U1/����6P��P�x��)쉠K[W��v"��)٦���0�w�s�~E�&���J����/��PϘݧ�>���bf��p��8�Ӂ�?u
 �¤@��7�Sлc>��%�|V���,�D�މ���e�g=��GG�~p��Bޡ��4�����sCI�_��"�7�ZM��-g��k��`7��:�X�����Q?�9Д��ھW��X�C*fN>-�(�
Lg��ג��S�c�vd��b��׬3���T�rc:
-+o(����"1�+�Ҩ��A��	�ؖ¼iħ�$��ӽ��A�q�B�	�V�*�4�(Ed�g��a��e�J$ZG0�#�c]�V�33K�`�r��,���/'fEڹV�@q�.�R�R\Ii�.�_�cW�{��Ɏ���x+	Z)(�S:A�I���_���j�5@4ĩs��\���+�C�S˩�2O֝�ј�A���U㤠[����j��gz��G =���z01]*80\�/�z�\1�T�q��i��-J���(��v����Gw._���'�+̽��Tϔn�Fa��s�켎�P��{\8h�;w��ҟ�� ��7�����=խ�"�#,�U#�`D��
�bF|���.��D�`)%���o��V0�r��ĩCd��}F���	zd(�q/:nF�1���KA��L�p�L���Gqp�	�N5J��괴�����4�+S�F����4GW&\��o�˻�u��?@�ǄnJ�B�� ɿ�.J�*�������r����]��{F�`=�����󞌌���oM�N�/�rZ\������������i;%D����q�@�&��Z/�w眃��Q�TVM����
Jfy(�-k#T�1 :�;>�|��_ $�2^��������	�
T����I�O6y�r|���� �.�վ=]��!bE�<q��]s�������Hn��/�X�[\������(o��3i��g�ՆZ��L"h�5jGt��#��ldt��8�/�Ifm�:�N�� GC�I��GyrUۢ�9YC���v�@���#��*Z�z4q�<C[�^<� L�Ҫ7�u�!#�9���.�\��R��ZѸ����u��nq`,A�ђ?\K20�.��m���G���kQ��h�O�'\�L�)��$([��`fЎ��F�=IA�a����l���{u k���M����I?�;����l��L��|&�R��#O�||A[9��z�;px*
�}�:��S�;�و��QbA/�5\�,�q#C�C�C�s%�7�OqWW�j0d�9O�1�{�s���%�N��U20ob��O�v�O�S{�n֝,�1jΉ�A��A��ӵZ�K����Jp��A�G�a�+f-"��� Q'�nZ�Bv-�锫�]]6o
8?*{M�HCZ�F_�N���n
�m�jI���1�Ld��|��_h�ڨW:}A���-���(W;�9(��?xm�B<�:��H����ן�r"�inT�b���F!�^a�x ����.���	��$N��'H M�����[��v�f�Y� ��̟�:�x	�q׉�r&s<'���SqH�gf�=��k�z/ǃ�1ߋu�:�j=������G�U��5�lf�t�,8Aӂk��`�tY$�5T�@���vXi��+�G�_�-co���Z)���3��~Fߊ�����Q��SYY�g#�$�����U4�x�+���W&L�X	���tjxX�H�d������̚��)$x=r(�����P��Z��
Ha'ߺ�1������S
����ڶµ��� �`˥�M�����]�rg
KTX Ccs
��WFnV�����g���=h��~�R���Tn�����T������j"�T����*�^��T������)�F��+{X�\��)�e�%�9������Nu���Cͨ�i�9W�J���LL�B1X����3;p(.�*�ޖJ����i�ify䑪c{��VqZ��S��)q�E�
�h�`XC �Mr�Pj`Z������Q�������Lk��M��_�W��=ѦHq�I��S=�:��}��d����[$qpK���ˮZ:7�M�#�*&�s���2�q��0F�YgI��hy�W	��?�`�܏c
hr8˼�^���&q��*�h 0� E354,�����2�����`�$�O�\��^Qj�cd��Щ�؈�]�rNgSY3�Yϔ��,-Ԍ��$ �2��45��9Kg^��a_n���T[?��v+�3��D��_X�$6_kƫ��G�U������ob���cϗ���C�Je�Ϣ#'�u��^o!3�C���0���y?�k��ۛłH��3�>�3��M�e� t�7���y�QZW��l�	@QM��.%��< r�
z	7��죱p_K�l�nI�<P�朶��8{hm��͕c�T@��l"���
t�.(�I�s\�c���jҕ��S�FI������x$�>���֔|�kl�p=-I�#�Z��+���c��c,H�T��R2�oO�Č�Q�.0�����{NT��"��L��o��~g�z��k��T"@9ʓɏ�6B��V��'I��
�<3`��X��s-��S��]
��r�:lR��c"$-3J� ��1�	�&ե�	77�׽cL��8-$���*��Z��)#��{f��u�W%�ͻ3�+����QE�LD2�.4�]�N�QC��xb��(�ӡ��UzO��;z�֖GN�VFB��<u�7���/3w�>�=EGy�B?����NА"#s�=�׿���=��hb9h8�o9?/�H�2峞-ڦ�&����JL®��`z	Du4Q��=���'I�N�ϰS�6@��c��]+�"D�L@���_�yv����'A��H��>����f���N�v|��@QWXĵ�sx��$QO�i�z�0���ɿ9�����c>Q=JM���>C3w�G�NA4�
�B��͡�
����㦉���H/{4�5J:�/�N�T�V�+����x^!�F��־o����xC����獈7�G!/�I!os�%y`�����4Ո�b6,���"�Ll;{�=N7c��k�qqD�[l�җeQur*�bT{D-��A2֟h>�Ɠ�F��L�ɻ�1��lT�wem����0SyzX�:{��� �\q6wY���7.y��R�~wh�k����b�o��7�[}��O��$n{���=#��m��~��k�<��3<:y��c�BS�K�I�gv��doC)T�`8���zd��h$�%�J��rڨ � ��P���P&{� �WK���6�Z��(�ZPÃ�1�*��ޙ:���`|�f��Ψ@椚��J�+�5bŻ�(5�hGM�pI;?�"�j�#D��*�gR'�g�!IJ��SP�g[B�ԙ�j��;p�w]�a0�71�܈1�Fc��3
M)���ҥ�Is�IX/�/�p�yM�'0=���rX�"�/�8�M�uG�T�vr�z�z2�FK5ׯ�&�w����ő~S��ft5Fr���2�o�;�ٜ��Xd�B}[�brWk�'K�
��7��)*��Q¤&��3����9�R풎��D�AݞU+T�)Iv+�=Е�
v��|��rl8���x��������@��C�Yn�Ùqƍڂh���̐�[�.JV���OHx���V٨pug'5��A��|\��@�c�� ��9�Q�"&�k��,!�B�rP|n�sɱ��OU����J�3u�}d�Z�	�6���fv� ^u�X�^	4��Rq�O3j�5���Q��L�%=���ߓײ��y +K.���Cž�fjP�ƫ����uWJ7��ò,#�����o��^��F��V}*i����%u����FL����CzH�[Ǔ���J�I���Oqr2�
�dNf:9H�o_1�*���P�;b�Bx�j���J�OEeq��K�;������pjcg^5�R�(�����)�J�W�#�O��oΌk,֫�tj�Er�$�{)�cn�x)�ߦ2��X���p���(�-��1�L���q*����������"&�dm�S��@�r� ��\�.!9�\=A���~k��[KYj�=��@�<��m�:�냂��	��[�o��������p^U덥bZ�����[��z���5�.�`�t�[����ѨQ�f۠�Z���6���y⧩��3�X�l�kp���Y��A)'w�,�Xm,7����Y)�M�.%g�K}3}��,7��_3d lkL;?�fy�mW�>+g^���G=Z��M�`4���r��Q��ԺǱ��y�P~:���
r���C]�N���۰#�X���s��@=h�N8����j]_=�
n�m�S�8��V��V(��}�)?�I��5��6�j�4��(Ҩ�����mluFϖ�
����Ľ콉W�ڿA���2F��rT��WH>.�&D�Ĝ|ܼ�FOu��f����Z�:q��J�<�d���`<'mn��@��;��%i�����v�>��#
$�֭<~�R��]�3�#���9�'�[X3��8�<̰'l�X{E=��3��?�}_F��Ya'7>WV'ru7���h���5��"���b���T�Gꬫ�*�B�؈�;�$�D쾂��t�x��}+�v}��:>�P���;����\V�:9�\���ߓSB���VJp�!s�kn�R<�Y��d=>Ib:��t���S P_%(LY:-XXi�����w97��(�������yRl@����\���P5`9;9#��J]��Q�#=�6����A�݁�۩
4��:j~/"��y��ﾍ���T�
�gq��8Ѿec��+|-͂҆�yG�S\p��F��Hp�a�B1�О]��c���sq������I�D�/-��7D~a��=@A?�+h	"'{�j��(N���y��"n*�
J�Ib��G�Z�c�{'�-K�L����T�-��Ώ��E5��v�V��%�,�7|Tj5I�T7�0:�H/�oI]yP3׬����ǼƼ<a0&���{`�sɒk��P�������Ѓ<q�7?���|^�4vшh��HE}�,i�8��8�[Ѷ���}�H��"fZ���
��	�߅x߃�o'���T6��{�Wu欄���Ff�@䲂>i:(��FX�&��	Q�m����-����3���v��+G��ܜ�����)I`�A?���;�Z�w���j֒����@���r�6D��A'Q�F.�	����vu_tM*<<W�6���>��c��/Zg\:��暚u�����e<���;�j@�������dm�B��f��� ����w{d�1R����ӶL��T�2��!}F�i�"<�o@)y ��m-�e��l��I���dN��g����x��"�>�?�������1��=�d,!m�AE7���@����>O���J��[�k���*k����� �Q�Jki~�~�:�'�k�@#�yfD�959�o��8���~�ȸ|r�(�0�L��2u�gsp�흞��sq�8�A�yk߄�.������`�r�\��t%�����ct41԰��]���-I��lV�=>�J�GQ99�s����¨k���bUH5 I[���G����M����Ź�X�C�h�����%�Gh�O�6���D���(���l��f�A����i��V��F�-3�毛��e����
E�螤qc2u�M�ĩ���ƨ�������{
�^�@��K�Wb�nD���ծ3�D���o�9���S���"���d���9���t�%`C�K�O/��$��0����g~8��"��PN��$K%:�B��'�V�|����qVk\(s� �Tr��#.z]U.=�o���'w\��/�j"K^�ň܎~ioy��{S��U�o�����+˹�m�˝>���Z�U��-[�Uq���(�b,��z�-/wFNgW馣�MU��lˬ`�%$9IkP#g�BD�l �2$P�q$2&?C���=i�"�!�����8@�*gB'��t1_��|CQ���B;ϥ�����o�[���ܹx��^b�~|e�"��)E��J�T`�@�!� G��A����eg ����w��O�(S?N�e9�v�l�3|��`�w��&�"��)��r�w[c����y�Z��C6����_�U�p�V�V�2���%S@=��65۬ѩ���?k_�=	�����.J2&7��m5��'��0����BN��3�+h"�s�[Knh0vs3�÷���_�޹����;�t[���9�O��J����J:�#]&���M�~<YLȮE��:�o^#�S�b��}L�7(�����閩��Q<9 �3�y/�0�n��Z:n����%�f��aڊ�^�-?�V��QS��s?�yx�������9WWG%��R�����3���l�ѫ鼲Kw	���}9{H�vt��P��/�k�������W�Re�����>H����tsOe4�ӑ#)�[�C�H&��&�4
�zXp����F�f�g�\���i�jE��^��)�@����]����~��˞�м�B� ��:Ҹ���Ƹ:�{wZ3��$C�>̵��s�p�z�u>��V]�D�|hc���ݧ.�g�5�t�R�/��01��T?Q	�x^t�U���ɦ��n�w����>�j8`O&Ѝ�Kd�|��fXe��u'L��&��Y(v��>�&M<�;s�ޅf���i�#�F$�<��"҈��>��W�/iW�9QW�A�(>���+����0Q�e*U����Ih�,�C��,l�4
��(�����F�qf�,zi��Lk�v�b��狧���:�kAn~=���|�I�hv)d=���-�-�>�����)�bUp�j4Zy��WSFf�-���3ȴ����Q�6l�D�x������r��| t�3��s;K�I����+31f@P� `�
�����F(q{���Z���68�NX"L��B���DtA�z���C%ҿ����Z�x������Z'LbW}|�!�8_Mi��cK�YJ��2�/�������}��H������!�æ�f��n)���I�I�l�z����XVB'�V��]b�^�i��U���H�����<L�6EO�|��<�M���bz熅��O���{�0:0߾��)�=���@(
�^'�+!<4��`����Dy�;�$f�'�����(��I�oKs�z��`eC߳������)�:E1�I�lh��[�.�6�,i5�\~�݂W�lS��}�WS�]�ʮ�w�ӕ���qx��v̋�h����� `��lĹO7���)�h����e�>���������pRiL}	)
�Q�tF#�狱!��ln;����,�*���gW�?�zY��a����ǧ�Xl�nD @��-|$�,��(1����7OeS���� '/�o2�h����*2���ԓЬjӗ�)��U��y�O���4�$$����`��ބ�3����՚�9g�tTX݀���$U��&dO��µ���6o¹� �]4���A��b��jH�\���"4f����K��÷5'�٥,���HRt����e a�Ū�*�я:Y1�`��)Yq��"ǣj��2��Գ��$�.	��#��٭� =s��l:��ZP�ܮ��)�S��y�U�]S\;�"2�+�����P�
��<�6��i �'q��:�Q\tŸ&V#�	 �ͯ<��_cD�2k���	�o�0H2"胢ĽA��޹�� ���O7�j����E`!n��APB�;���N�e��p����a��s��F��!��4�58���������'�%�?!K?d����n��RZ_y�)&�>�_OeW� ��Ȭ1�������=
�*I�C/1)C`��� ���&3d�`J��U��I�A�Cy�(CY?� jm��&]oR�����ϱM��� ��&��S*L(�UNs'�2�?��I�"���c����^�D�Ŏ'�p�A��N�Ύ��h@-���e���:��YZ�����K�& �5���X�H�{�J`?FsAJv���U5�@]��m�8�Ks)"�<;,�$�Ό<����\�.(mڙJ���to����s@��
�Վv�����Ջ�.���v~2wq'����_tv��^�Y�SO"\�kU�LT�4�[r�|���/.���b�o?H�u��VP���[X�ӗ��$~u�h�r
�u3���>�����L���<��(*�T��kҘ�q�& f}�-s*��Z0�#.XO)����5�W.�����\a�pv�z`J{�`�c���vȫ�:�2��B'�IG�%���;�]�c��I0 ���&/5��d����2�}%0�[緇�s�}2t�r_/%�x���obbQ,NN'![�O��+cg�qL2XM�; �������$Svh?�>:��tm�OWJ��8v�8���,� Zm}Tt5���ѐ��j��,��(
�֖�Kϼ��T�&��C�s��%��_�\u�:����c�GZKԙ���M�]�Tu$�{��3��6��A4 &
�ӂ�q@F�;8�+}h���.Q�h`}c����8�����Q��G�^��F=�#��_u}L$���ޙi�Bn'W�F7�9#6��i1���"��ѾsK-E�b�1U}����p^+V&���f q�=���)9��S� �A��' ��&b-X�()��Hy7߆��*ɫl��S48eB�"I'���q�(B�8���8R�rL [�m��TY6�Q�"Xh7X�ܛ����	�l�7o*�:�}k�c��ļ�g>I�E�U��{G�0��fG�EL�Q=��r�F/���jٹ$��S��R̿���oh��+�� ����#��m���#�8U1��D�ޘc'i2���Os�ʂr���dT�N޹>D&����!Dӡ�}��C�y9���������'O�+�w�/-:�w���w>�ZK6��M��-��ă��UDa\?=�bOG �m6��9��=��g/��V|�,�R��������:i��_���r8�ߡ�t9���I9�	�7�ϾV[+�g�bʐ/�~��:��M�D�+�����U^�Q��mB �[W�c;'6U�)�L(n�;�������_n)"$ӟ�6�w U`Ut�o�DA�ñ ��C�g�����R=\q�n���w=i��z[��*�i*߉3�1�4w��i�HI��E��̑ul:�06�)����܏�qLj��:#;kr8q�#d�(�ݓe�@�Jz����/;=c..���i���d��<�řO�A&�Q^�u0Cm��(���罬�o��'vރ_�G�.bL�Ԇ�Je�5�y��X����s�."3���fd�4m����*|dvˑ��O��ņ\$�P�D]ZFڟ5�o�m!QG�V��~���'Q��!m��=�@Q.$h3�[�O	���f�y1 ��6�r����c���L4��B��������46L8�^�P�ष�����?�jn63չ��h�,�8��8�����,gg](��1]��5Bm
+w�����op^+���D��Z/m��r��/|O�zv��V+S�Y�㡈u�Y�9���&�S G�C!�7z��j��G*�J0+�ǅf�����j��/�\ l�Sm��/%M��ĥ+(�Sj�Sd�ԥ8k��Ey=�^'�
�X�& ����z8�*�ɞ��K�Uw�|�=R8<1)qr��
/��}������n������j�x�դX��(���P��(9���F��tcG�l�b�����N�?������/�<�5}��t��ɨ��?��qmP��Usb8F3�	劅���ﶈp����^q����Lb���\�
�~ۯ 9����ñ��)W��M	�=�Ɵ ĢW�@�yѪ�@<'Վ�U/�Ǜ����[࿒yJ4���F� ���Z�%g7s��X�qk��jꋜz͈�s#$-�ՂN���;�Iǔ��#�ූt(Dn�߼�^����V�-Na���J�E�M���>�%h�gw_����AΈ�2��z>�� �&J�ͻó@�j:�{u�,A@]�S�f��#��/z|�H�����!.���(64 ngΙr�^TE�pev�$�%�:���D�p8�>c�_��lQ/�42?x�۝�']LPqA�x��qGO`� 4�J����M3�FO"�4<�)���4mHӾ]�$��p9�F��
�k �%zײ�E3�+nt���5(Md��bYt_��-��+9C��`�Mm���pe�,�1cs�o-����'���}�O�/詌ȵ���[A+�6l�PP��R�E���SR�N��Z��CN�G|h�OSeև-S�
1Xk���UM�ʣ�j�-�M �P�a�X�$�^���T�BL�-dR[i�	:�����u��q�:�7Į�Gn��ېx�4�\�i��3~��)ˌ����P�;�"�Iؾ|ْ�~��T��ܖo�=�#�֍E/XaB��s"�6]�P�'�<,a
�w/˶��i�K�겇͵ �0���5�z&��&�*�	&�pD���v�f��V?�eD'ԑ~��<��|�c�Ѣ��m�tE�aJg3�(���T6ܽ��5Q���?SF�<ֳZ�{�A�b�a�v1��7��Ѝ����G鶹�#�Ѳ�J����ѢV"��m;� m�~Ԋ�ܣE�OsUM}UFU_��&f�=�H��Ri���acZ�C&$`=eu)Ҏ�e�x�5I���k�y�i{F7{��.]�I��;��d�"�����%I�6�V�ĭ`Ld�8���RhOm�x��m����o��Dv���a?��sh>RV����Uu���[�U��_�̎�|,\��{Ύ�������������>���ӲX�ZN*�.V����b��&�Ѣ�8���
G�]��ězk��o���{K?��3�v��<^�S��*М�%��
J;�����/��Ҋ]�7���z7��<3�N�`�ҵ��q�����p����#e�� �Q������/!A���u�s�>�V�	��Q�_Ն��I]M�B�ai�F�����T�;f���� X��ҫFHWJA���)0���Z`
��4�H<8,lv+]p~��X��9�fS�9�ݼ�	/��u	I���:,�mO��E0�a9�jΕ��ՠU�$Y���ZÝ�R�cg��ܤ��|��[2Dv�o#���W�����^��Xpg�9!��h�C�k�qEj�p��T�US�m�/��G�?9���H���%�M-]����,^x��pR�@m<"�h���$�zzcDkg�?��\ԟ]�t�q �7�	��������s��%Ν��� 0���}G��v�-��5X�����G-����6Be�s�������d��*#0u��$ �v����B�Ԃ�
3�=�a�&���lT0TS~:��!b/X�����X������蕇xZ�f�	�D=�_�=NDB�$2�ȕ�\��,V�,��9/M�6e1{�y�U��89^M�|+}OQ�l�+b��'�Lx��	ug�@��'�o�B�1�T��w��)��"e�@�p���w��95����Z�4��0l����)�;'S���h%W~��W�y��SiОXK|�<��g%��Z��f��k��	��	��S1��ۈ��'V�%7��@2PYv ]��׃�=ɝ�Uo19�W�Oê%%���+g�N]�
�/�*^����B_b3z��7��� �:�l�~|ԓ��]�s�tT�K�y%��Ai�_N��m��$�*���ze��P��z̧�(�?���G��`O_-M��Y6�'�bGz,W �G�#����e�L8�Vκ���a',�FH^(�|�m''p�z#�k�k�Z�Y�Sl�X�%�����3��VW�l��S�E!&�D��6�@ٷiU7��I�l��^4�ƭ0��Q�s��츟t���HS�OQV�nI��.��˿Y�)��d���v�H��rߗ@�f����T�����KI�H�e/ ���L� �+R|��|���HȿIxZ!-�����.�o��+�����T�s"D3�J���\�t�N8l��M��˵�7�wʊڭ�����3&O>e�;�Q�uPiJj�Sx��6>b"H�AX���1O'�d #�N�3-����|c�K����+3i-
�:9�^(V�^�KR�q� ��������M(�<�`�_N�S�	j�!�	�����^�.Q`Ds[��t�>�b藅����BD%@b+w�KJ�ǅH�KH;H@����4��i����@�c�4fU�0z}��.,��-
�n �ʘ�%�s԰=��屎�N^�~Mg��cA�[2=]sNAw�G	����M��Kn|��^�M�~v���^���4|�_��t=X�fM�*ץ��~�.T4���:�����0�p�P<�&���A0�e�1U t�$D_���؀r5w$ �ٛ��CV��$űq��X�X��w3Z��P�pFz>k���c�4�"�DR&����?+�gy2����=r��V��#,w���0d1P�kBWL]�o�X,�z~�����Z�Zt�I��VHF������K���B����5ct����)K@Q\���� ��������k�Ⱏ �#�����#��g��;<b�ޕ�D?o��gkk�Y�����e1sj���ޘnF��"�C��	���=A�`�I���5~_��'{�r�W�9#�0I!-`T����]��V��U�ڤ��P��`�IHb��\�!.��b�ʉU}^���}t��=S�S��5��=Ug�s��3#j��	���젓�KC|s���'xZL�Rw�(�]�_���[�8�/�f�!29TuN���`Fѽ�<��{yx��i�F���i�8�uX�.a�R�Śz�Q�Fn���%����|Irj��1��ŵ�%.��Vj�=iGF��C�^"��c�<_hg��gWUE����׎�<�u7
���'��!AU�QD��<��T�`:P(O������7���ݢ��-1���'��w����B��&diW��� %4R��'��hC��t�C�JS!wPZK�s�e{4�x'�KY�l7�<#)�B���q�87������&n�OA�������v$����^��8��G���oz&a\�p*b5�XM�/}]���c�bߨ��*ݯ2��s�ikt	��"[XI@j��W)*	E�өӉ(>�%oUc�@�:H������ ��WO�=D"=vU�b�ڋ��Q3�������e��Ak1��e>�w<�H�/�����1��*Q����t�Ѐ|�sG��2�tY�L���d1i��g�>��Π����,� ��@O'��zl�9e��߁}�,�f㙯1�u`<V}���n�N%��Q�{��ګb��+��K�j(��T}r�p9��Үl������wO�y"�!�w�&y*B��d�+uT�H�
����"*\m���1a�0'���<���z�1MT	��LL)ИA��Ul����TύH[^�J���3}�]��̺�e���*����?���*�*�Z�1�e�Q�{�OO����>Bn�My�q�
9���s��fy�G6�������P#����A�����]-m�d�5V��@�{т�H�=L;=�-[U��HO�V__[d�A4s��4�c�=�0��	��s�θu�0�t�J�9����M�-�!��	�Y.�S�G��
[�}s�]"e{%�*<�du��<u�'+�q\l�'��&�B�>>��$0�?�H�[�aOྍ�/A��'&o?�P�ON��s���.X���5�o���_�hL<�ױ=�iW��EM��A ��H�C&��ޙܒ��!��a<�t�lx�ľ����]V6[��P���}+��-�o��De�� D�"9��C9�J��2z|��*f��>P��O�5��K&�t�߽{`�U\�Ĭ�_~F����((���K��7�~z�]�0��Ҟ�K�.<����D�ȷ�{p"�۾+g����S=����r�,E�7=��u
ٯ�%���������5L�R�ف׌��t�oÕ��.�M��� ��Ȟ��0B�_��~��9�{���@ŷ4:��%YD͸�-��Gk��e �.�t)��0���H)��o2�T�/86�x�f�\�fG�?�ɿ�w̨F��Z޿�>b�c�EG:.1�1^� b~����:q�=������+�������xݜu�Mx���Z�����n�Nֈ`&Rt:�����TӍ���TF�̬�lQnX��2=�y��_pז�RиK<Ӛ�~���6�U����&붦@J�Y�n�G�ˮ���� �+��6ʪ"�x$�t��"k֊<�!�댷�Us(��.c�7<�	&X��rpw��	K��7uRI�:ļ�{c>�K
j��Jx�޳%��m�<k����~�֌��g��I���4&?+��	�FD-����V��p��=���뺨���4���ɦD� =�Sf��t+\g����U�G߽�O�+X:�%������( i��yo�������e+���Q�2&��Q��]����f�/]���oW0�ڇ�?I(�mn�`������D�/�a�G� ��ڭ���@�[��G�ƹ�GKn��t��Z�z��>c��ȏw����t���H$���7���[�#�*��
��tJ��s�&��5 �/^����n��cp�{�O_D��>�"�۷ϒ���Vy����4�-EU��_�J՞+�ҡUO����fNY ���n�b��^�Q>����'h��2l����A��J���ۓ��5��	&km������X'ҲAI)n_�Hȭ鳑~�̾!�;<���I���Ȓk<��)�A~C���P��Su�GS��=���`��nc������P�wq�=p)������ɪ
���J̘[��HK� *	���tj�S�<�K�ES�P��d��gȋ=Qx;�]�\4����O�����!�4�yt�6YMLÀV��q8�u~=���6#��Uv!cKRg̺��h�X��B��;1��Z�����t?�L���?����L�T!�����W�����˗e�?0���{>��G_ݥ��k�p�#�
px�F#mJ2C��(�-�-6��9�,6�^84���G}o|fV��	�W��h��j�+I��ζG���h�lY��篳)�����Q��S�Y��=����ڂ���eq�v���=x���Q�l�/�Ca)#�����kx�.T�7#$�L@y���� �M���^�.�5�خ6a��{d3�Q��s����cP���Gi��S�F��k1�XxOJ�D����r_�Y�6+�B �d�֨f�T~�b�a/Be:	p�i���;��~��;�ه�}w��T��a�~�TF���5��Q�W�QU=`dܩ9$��7�C�,h+������ɠM�tN��Cſ�w
���L�^*)�:��ul��y��`����m�fw�D
�`��ص�h̢��I2g6 K�Ѱ%�W i^��y��v'oi`�E0�6W���S}��t*�N�MǨ,�`��+p�vC�ʌ� �Rͱ�?c���;~͎[�����I�1i�%���_]|�D��H��ԓ"v�����>�~l;鯥1�t���"�g,�vt��jtTᔑ:-��4 �ْ,�0���+��{�vW2��r��(�'�`_�r�p�4�?�{���5�bI��3�+2��T����?�1�;��x*�Mҗ-*��^��N���ʫ��A�e��?�)zTH%�cNҝz�4�h�LG���\����n�Q�VyQ"'H��jF����ӈ)���?�� =���XUJ?��� q��{�{L�{ׁ�9{�2`��}��f�b���6o�g2�E5����̖T��I�8�f(f��o��v) ���_0�&�Hd�O �jON9BS"k�
������9*N}ӑ�N��	`�Gh��=e�*��<p��M9;	�g� ���~T��=t9��,9CDJ�j�a���4��t�*n���"�'��^&��;}~yur�y�G�ֳ5��tYg�X����B0)c��Sb��T�����]x��(�	6�A&��L���<(It���N}pX���"Q+�7�h�N޼��*�98c�ʸ��HaM�@$~��G��2��e�8��H�q��ײe��#�b{�����ZU���{=�xn-����1�X��֞�Z��n�+��E��pm�aI��Κ� J�Uڜ[�����nh4V@���/���1w_��E�=��}�*u(�RP��Q��J�M����r�9A�3���R�!BV��"(o7���f(ġ:I�Y��#�\�f眄/t����6��♯
�E����O���2�X7��v"P�]�f2���#^���ΝF�IN0�*\�K�!$=�mvFC[���pc� ���~���N��_?�SS�8�Mܢ�rH�h��\o+������y��{��o���Bt[�����Ib�<��x�O�C�L�(�d�Q��`Gv��]��'���l��8Y�?�Ԏm�p#�i�&�$��<�����-�u$��D��v��[-�V0����+Ta�B�� #��L_�Aم��~ց��h^�/-Ԫ%�Ɏ�k��=���|j�ˬ�F�;����t9�͆���4�u��ɧ%�T{�����mKW>av={��ɢl�CR�)mr=����PHN��GE�/��Ћ�zNJ��m��O71S�T�q2��(t����`���	`<o�m�NW��:*h-�>��Uċ�6'.	�8%CG'ׇ�.��c�LFe�Hs���?I,��Bs���@�ʒ��b<3�J�T��MDd�yo�~c��m�nS�_tp.���L����ߦ (�j_��"��Ŀ��& ��p�zZ�j�T���t�]��Jc T=R����n��\'�V\��D��zH�R8�$�դ�9�+���7���DQ�p/�a&�ҬE�=���5��@�`st�.����b.콴�p�5/>�OVv=���n*�`�T�u�p�+w&q�]�5�������S�f	�'�k��!J1wH�<�Bq�o|�䮙r�PN�IJ�����ͧv��/�v�]��ԉ�V������<�w�Hi�8ʌ�o�� ��#����I��ʤK�R����\iG^��Q����M�@�nx��t���a��Π��ۂ�}0+U���T���s�!�4U�6�Zx�s���@��(p�'32ZI�W����4ޭ�{g��4��a��G�y�*ĥ�0�~�U�Pio%j?�F�b���rZt�M�I�	�S4@���l���k�ʅL	��`E�*D^sK��b����!�����V�ߢxŵ������)�؛}͌y����(��[�*1.d�d��)�l,�,(��o@;F�Hq�V�'!˞fc�S4j�8�A�(*����
�=�`_>nK��/ԯ��Gњ9hj��^�v'��'C+[��Y�lҽ]�f�j^I��obt�{\ѠHNz��#[*֦��=;��;;5m�ԇB�$�p�dQ{Z-P\ʙm�ĵ���q�:�r� �'m&I�6/��tiODc����X�ǵK�"�L}4�rb �U�����3੫�$�k�Nڦ�Gԁ@��ј������w����|c��b�����j�W�]��u���G��0Z);ubT���(�PB�3�]
�"�[�{�4'O�.jm����'u��cz�1_�ҵ���o����ܻ폾��F1u��t��5��.~��t�
���# y��cH�q��b��D�d����2R���\4�8'��02޳�b����?�p d�%_R>� YH���v3���q}n:c�#t	�\`��H~X^۞oa��3*�F>"�4	�)�ll��bM1_^������D��>DD|ˣ	С�v�ŋN�eZٛ�Ad&�N��´�?�����90Oj����}6�������r����E��f���mX}�u�+N&dl�KS�*9�)r�Z����~ke�s����*6[ǃ��o1^^��c��A"�XMhO7ݳ�Z��ጚ|H�����I��CYd��>�p�O>���x�b?se��R�D����U�
�t'~��V�!��~47���w`�y�~�����tG��y�(��Bge�\ݯ[OY��s���I�����=[ 'h�q���Qߘ��0��b*��d87?�%B|�5(�}&S��"�t�4��h!��{�8�y!MW��a7�ӂ��CR�{f5�_��RΗTj�����������U�lEՅ�}�@x�f����С��ы?+;�]�;9��1���'�u�4��όo�$���
�us%�L[��y��MO7�ğo%�-6�űę�T�,ZE
0�Ѹ������žԶ$�Eq�s�{�z�`�w�L�L����@�:�3��p���",N�@lO=+gQ��ȟ�MB�u�S�+/�,��Ҥ$?�.ºrl�wg,�"���y����D	��]�}�CJ��?_	=<�jN^��T���2^!����X;b?��l��U�+�cɁ�.^�>K�_)� �J�c{�����=h��Eo_-K����%Q�Ym�D�]��e��p2x�U�1��<���C_�����qt���k�Oy&׆L%a��VmpB�t�>�7�-
�O<z���@v5&d�q�N�߀�;�A��Ѳ�� ݾ�
1��	���c�Ǜ�%�t|�Ѱ0�QVo���V�r$�I��XD.���+�� ���H���V%�l�Q�-������=��ST�Q^��,G��CE�[��%]]������f�V����R-ʚ+
����z*�6��['����,K����Sg��HUiK?9у�$�rc��c�|H��|���\� ��OsO�G�?.�@�o��,;�P=��3�R�|c�4��x��!sq0��PUP��8𐳍��o��D�[�ҋ[�������XP��\������b��1����'�+��>@��YIN��]�Aaݍ��CE��
�č�p�]��]NuM��yu�*����w�˘�4�)[}1�}�P��*!Yz|����O����d@Ņ[`Q��g����k��E�f��.��Uv{��1�'s"|�N��;5��]cY�;�̵�%�P �}}3��uN&3�L��}����>�i�)�:̑���:^������O'����h۽8���=�ݮ��k�e'&��n¥�Db_��V��h5͇H/����vc}X*�#������e\_h@&А~T��;H+��H�!�����.}�:�O�+�\=��(�N	$�������?��h�-B��H�}}��z0��UE���\vo�f��Ap6�g� �d��·�Z��h���'eqj0��
˿,��2^��}�2�{�Y����d��f�$���J�,�A��m�?�bx�>�8�y~�VBal-��߉tå�;�NI�{��P�|J@�E9s�������`	����=R6'>�t��`ðO���2���)6 �tyV�+�=܋.d�P��X��"䏡����ݔ�ˋG$��=+��~�!}{4�fIA��,U��k�gH��CZɦ6!�A�����;J��z$A=T5��5ˑ�z����Bz��Dy�����.������s��*
F0��ۣ��|2*G��O�03��%�7A?���lS�SJ�T��3�Jk;DE��x�z6��*țn��3jUI���F�=>i�3#��񫗷�G�%��}��g��6��j��i��Z[pn8���=Q���h�J@z�1GH��T����᳭�����aH�M4�ZY�}�䔅�Ŏ�&l��D���-Z�vɆ
�7�;^~T��B�A���T������' ��Hi+R���w�d_����x"u5�)۶��ǵ>X*��,D?�|�JȾ�Md�QӐ�=��m�U{>KIYe�����Ѝs��c-��v�i��'P�qL���y��{�:��[ɵ��9A_ن�{m�3��.��/3EHY7�Xf-�-u.\ؘr��:\�+�*���1���ݥ�`A �M/�Nʞh�X��>S�̗d�4QX�J�a�O��캒f�,D4 �uM���]`��EY-o�i��u�����8Ж�}�F���BK���H$��Q�Z�}���ɌE��#dYƻV�0,a�X����K�:tV�'��	]���(���}��U���վ��,qsV���'��B�`����*z\mj��.dR�����c����,B���`�
�	0U1+�dV ��eC���)��BN��zN��i�^,C�C������|�%/���z�$��G2{M��Oj��5�;ͽ�:���zqm�ӽ�M�'����J�(�;R��mg�UZ6���m�Rzy9	8��ET�b�T N�����U�n���$>��c��)��8�{J�<`.��0���k�X!�^��Ku/�xD����s�גP��{B�|+iI�$Q�?�e&]�|�}:�Vv8�&,+x촸��1�Y��:edǫ"-O����!�P͞�T~7\�cn����w��~~��'���j��B�	��V�����ܴ�,w���G籏�s��&���z���z2�~ty"��M_G!
W!z���^!�Lv+z`��ý� �
b�:�5z��3�N��k+@��3^�y�mH���*���}�۽KT�7�����i�%x��Qړ���r82�'��`ݴ���S�s<X�b�Jƻ��%�m�y��F��y���`��b0��H^-�Ub�5�-�F��ȭ�\K'��Ilu��HZ�p�9��*c-}Փ�֣�(=��R���q5zԬ薅2S�������r�y��;��ڲa��v?0�u�L_R�|'aGhxf%34��u	�r�0��ƄA�/融�e��:��<S�M�����-�׻;\~:x�\�N�IH�i��Qň]Q�~�)�`3�`1����P#�k�_�J�'����i|G�E��J@�	3,cWw�D_Z�B�D �m�����?ch�-���D!`/��&C� ����p���I������QC�B3�1���$�����7��:Q|��߀u�.�-r	�$���5v��ۅ}�FV�=���B�ocywr�Ih U�D������0-�T�Z���)r����ӋfĬ�E��b%�t�@�=��wր���Y;Z��2��$��[mH��2�pf���Ζ�E/�يg�w��޻Iˆ|hÛu3f�B7����ycŴ�B$��1G-�{�Rl����yp}Ի�E���08��Ra�T�-g���A���ʑ]����᫥���hx�i��.�BD"tu�	�y)�!�{C�!��Ԣ�jI�_��3��B���9ͫ�f�����fC�͓�m�%��@^@�p�$����nQ[x>�ȏr)�q����P�<�@����-5Ί��c��J�����������|	s̔��MO�ͨ��f�ϒ�%�}�M������KÖH-w xg6�$���P�z�2/��5��7�_>G0�CןiI�/��i�m�t�J��۔L��834k�f�Sh@��7���3��9o0r��},�CN�YFV��t�r�'�M3�*�i��eB�����/
܊AeU����������#�+���i��d��{���=�2	�+F�����J�[�,l#��Vp��]�3j5g��V�_L~�zğ:6�����K�-s~%����N�$W���S#��(�l:�険@��µiH�(OA?t-���jF�,Kf���q۷x	��; �R�)E��,����/ �kg��L�g�^�t�4�3�x�����A�Ȭӷx}�z���T���=�AN����6%�\m�d�����ϩ�ڀ�F>��f�z�7�z��V.y�H����I�/W)���04]�v���2u��'J��Օ�cu�a!��W��*�Dq�ɂ��ܐJ�O���GW��iuhC��w�{t ������%������� �=6���˸���}�h�k�cr[YA����q���aB�J%�2s�U��5��b��%�s	�KG�lIX%��O�G.ۮ�7D�B�ܛ���Hw�N�e �oi��'ʆ��'9)w���ت��8�<���R:��77�|��0���n��f�^{�p}՞�,{�՞����A�n�����][�6%��T���:�C���o��$'�� �����6�`���8�^�`y����׫d0�|�L~e"�pɠK�xi�t)R�����͘�Bt�])�	Zm&�꭭�z�b�tI�xr�ϑ�����K�`���d4_�Aٸ�-�y�?�_�jD4���j�:�ꙧ�I\�C�Q�%+�K�1L� �K'�?.�X�ǛT�.Z7�k�Y�( f]���Wnv�-s2D���(}犪��z�����[QʑqY����6th�ޅ[:Wќ� ��ƙN���-f��K���T�ڊ<Z�J���PmWF���l�Y��iR�*:߷ `T�%Զ1��ѡ��Ō�f�W��ej� x&����\)���p�`�U#�%��l�!Cw6B���N��D~�*����i�F1:}f��!�;�]��<?�å��\Cڠ"Z�~�&(I�)b����g�I�mpK>X�wg��iks��ӡ�C��q�;{3# T���2�a���6�f������	ߎ��9ra�ҏ��E㻏�����a�J���N���M�IT��K&�2�^�n�0�_ˍp�6`a'�#�{�Gm2������$�ݧ�'P��0	�UuK��P̭�t�}`I�[r��(Զ�iU~�zɓ�^��w����E췲�>y;"_��i����v�rg��������O�dh$t�B���GY����{}���<������ȿ���K�8v�I���ԥe���E�a �c:*SD�Ż.��'P���|,6������믌��t,p��7�[�[���<��
�\G	�M�ڦ��K��S�5D�ܓ�O'׉��TJ�s"��[��ѲN@��[_Ӆ��00�a� �E�єN�Bxz/¹y��� ']��\�+�`'s�0�?��]��&���8��L���x���e�p2���`h���yW$�|:S���K��<�(1��:��a�	|ȼ�V屔��;&���zd��@��d�R�"��ߞlI�F��ז��u.��D� =�dU����3���O_��~-�hz�E$� Lf6Q���>����ؑX��f�����J�@�f�-p�:&��N�<���`(���؋Vb��!W���rӹ���E��Ay�K.���[.��U�a,���2+#����:/w�<�tߴ��]��oi�9W�Q�K���A!$$&$��W��r�7ztGw��țb>}B�r^{�Y�+��3��I��'�x����)������ByC��#9�a= �U��
8�I��8�H�?����\����] g�n8El[aKN����W@H��y�I��"/d.ڢC��=k�\D�9��U>?�H�;$b��.}ڡE�)U76�Y>ܦk	�L�0�.��W�{��l�X��c�%[�/��ٯ=r�b���$:�ِ�M��@/��1��aG8Ox������7~U���Yy�*���^9�(�,��_ ��� ����j����ȵ2��sp$L��p�?���C�w�:�=��G!���x EڇN�k���,?�X�t��g�E7�~�k�B�C�O�GnTR��.o��Op6�� [���$1F�!�/:7zPرw���f��}��[�n�҆�ҏ�OSɅC�%KU�k��7��&Vx_��gFSg��A�Ӛ�=�H��\�}Ʈ�fuv<��1��T�ot��#=Y�r�e���/	����lz		�}T�fS��[o��o�x�4`���`5ٽNH=&a^�� ���U�4)�����v�6e�F�|�J�K��Z��u�����@@�*|���T^ߤ@�:0�Yu����y�W���V��,P���9��&�eE�zm�T��	2�����+1��u�����]W����J6>ob��IU����3H=� �����m�t�$!5 ���C���<n,�yB���g�n]��	b?<���$�Q��=�!m�owl$��y)y��lch\��W8�	�̣����`�S3'O3�7o��h�n�٬��16�3&1�����G���⎜��N/MQ�TƐ#�50U��ԥ���	;r���6
����X��U�_?gt͢���~��j�!���kkr��vj�k�K.:�����*dD�3��#Z=f#QK��MAI���<�n�,1���a2�K���ǎ jE���ct�4�]�g��Q�ȼ�5��)�\��<��`��vI�ઃ�{֒��S/����o6�6��Y�z(c���=��!�A�K["���߆���lm�gASݔ��\����d���vR�֒>�ؓe�)�P��{��B(y�KY��ϢP�?�P���)�0'�.��P�A�|��R���!������~��W���몑W��}��nk�U=���+ �ֵ/]���ج�$e�갘 ��"E��M��Ui�ߵM}����puD��H�20^��a���iZ���7ź��e`} )g��8�҄�ÀA�%G�}Y�$���������� Q�٨&@Bu���3.Df�)�����u��Ȼ-����I��`	���'4ܒd2<��ƕK�0���a��wa�#�22��Ǐ`;{���bo��Z�:i�Kd���J�'���UF��!�x�^�����45l��E\��[�&�t�G���#t�>�~��V��x����܎k݌	z�Ú@kQ�S"��ȝ�P��;��sli�dɋm7��N����D��Žp:�Ly�ƿ��B�t�S���:�ӱ2�FXZ8о6��+��P�M�!�ʗ��<����:�ZeP��߱*IƢ�z���TP��c����A��e�u��ՠ�f,��Dnz7�w<mHXl�D$����W�3��߽ �T��V�u}sY���r��|<$nG?�20�z��h2�]W��#�^D�E\>ӵ=��e|�>^��-�\��9��@=��pۿ?�(bo�}��D�6�a���7�	��9φ$US�}I����p�jvZ"�=(�J8{��zY��#��5W�*�̌M@���lY���9!}�VW�W��ËqU@�27ʧ\w"E�]�j>��^��(��Ȑ$�ݡ�_x����[�	���?pX��$�Fp yP��I�*���_��\����W�0�9tٕQ��"�[f�Z��1x�|���� ��k���������ʳ�I�����ᗣo�?�U�*�[�\{�>Q�I�f7黲U��X��B���C�zs�Q�eN�H
"�_m�d&6/��KW��"���8/%�_��5�'W���LIs.��%wS��dV�H�!^�uM�eS��ؘ��rC[�c=�X�����*�2��ȓ{�z�=@�MNA�����P��
���Ɂ��l��Ѽo�岄����{���%S1G[�<jA��E�����-[�b�u8��٤1EA�cT����ʚwC���V�v����`�AZ�͘6C�t�f=^L�.��#���olR�&�2�j�̮H6�����Qѹ��dI�f.L���Dw�a��N���yw��
o斻�R���PB��:�jn���c�3w�%Y����t���Z������=��}�5#��27�E���a{���A^�Ħ<k}�_���/�1-ۛ7�rP�8KZ�`T�tf ����w+���Ѯp��H�	�t8x{���O��n���ѯ�3OE�ܫ��m<8�Hu���PpGy�8ZX�q�"q�Θ�6%u9"\�$�u�x���J0��	&u���_��6Яn:i����>��@�*N�jɈ����E��W�F�����f����&1�5�/&N�5��U�kmO���N�o'�4��xg���?"��)l_��p>	9=�̻U����y�f$I����~�%�3���K�G�}��>;���/5�T�#퉭�\����?�C�� �����H_��+�8�
Q &Ȏ�����'��o��P�E����&1�CYW��0+�R!�w3��ߗt�d}Èl�*�MT�iuw�<��l�=��Pvgл�Z�a����g��a�z'Y�_Z#b����4I��m���H�B�"wQ���w '���p�{r\nv��$�ſm�}��O���"��< P��@b����[����
�a�M��y���Y�5��d�߸��H3�F�3��Ƿ����9��+f��ę�q}�T!��tuyR��� ���#���*�p�oA��6iw�ެM�d��D?�y`�+����f�y_J�ǎ�NC�Mi�c}�5[�(̵`4i����-�j3� �Ʈ2G�[���V!�����Y#BȎ ����2s33/�5�Lk}
�23g`2�RA�$�j�f�@p�2���0�9s�����  �ꪱ��80bN�7q���t���P;�Q�/?�ˀ��j-5�8�+6٨�]�4����	���І��-c�U�"2���~�K��s�$"h�m�X+-�"u����'V�� ���n�Miz; JC�=,����АZ���y(�ͺ=c���t_d�nu����1�����kƼb�e���cʢ��k�sa��̦5��Y��x�(��*!�j`�O��҃�1#Z���|���.k-{�P!����a�|oW�'���D��+����7�Z��,�MCxd�qgx�:�3�ȭ��G��������
����ip�F����e�h]hC�����S��o����y.�:�Ś�����c1�H@-�HC{S.K���3C�8$��"�?���+��7T;��~�N�{2�/��d<,W����*�9�B�n�$��K�oM3����FҞr�P���0��ߎ2��(W$Y6C"k^ ��G7Ϛ����"��~~�9���	�s^��FW���^��,n��T�z.�M"��V��˨����X[{cC���� �+�~�"����8(:�Y4SiU�c������IP�ӜҮ��OHYd�]���Q�"_D�&�O�$�7x���q�47t�a[}͗]X�S�#��Z�"�	�o=9z�Rm��Hbk'2�CU�N���ڨx���؝�`0Q�eT��=�FS�E�5���{��8��^`�
.a��G�G�)[����]<aC���O硑��C��S| ��J\j���QK����a a g����+�{����w�>�G���^��������A8�	G�`���dK��o��� ��n�P�X]xӤlӉ���U��h:6m�|�����#(UB�b�w"_OL�L��Ŷ�
`c�w1������V[J�}���;O*�'�|�{}��]v�lS�%T��r���̏�0�Ȝh!p��[� c4�Ͳ��hօP��?���m��e1z�bu��5�jH����	r��;���Ji���o�2Y�No��.R�RB�����!*"H[	�a�5l�.8��^�蠒b�#����Lf�{8^�uu��lGv����8$�#��`�N��=�S�":��i�r��mPG"�l��$l���]���"DQ�G�>�/iS�%��p��l�c��W֋{n w�oYj��-_�m����'i#,��p�u8A'Q������i��ؚ��S��t�b�rA�w�M����.Q�=:"ێ��V\���<^�Z�#'�В*�I�������A�E��I������L?�t�)珨|����ˇ���}0��QkU��o`ƶ{���qU N��dek��<wb��aVP�h`̘O�%�5�F4��I~�W�'|2[�i����K�^��Oeg=ǌ�i:�Ժ�:bPR��Ч\=���ls�v�Jn4(4���h�Le1���CBOU��ؾ�5����ȁ~���F��
Y@��t3�d�����9l��Pz�Q56��e	�0�KI~,���W�<�[��ds����}�W$�:�kJ�7�۠7��s2s�9)�³o9���R'�à��P��-1�:ZqFP�2������\�a7pT�)0A�)��gg_��Ɓ���d�3(�T����ߺHt�����J�x��iQ�R<��8@Ƞf���m*����o�t㼟8#*8M ��tQ�c��\h3���Ωh�*ڤs�lܮ[�aM;\�̎�Yo�g��AA����] q�g�,����(���R?�ӆ�����}�m��&c�����}��M��s1�zwc��;�й��W�Е�O�"��oJ}�Xlb뒪l��"^�(�vh��0��e����]z->Rfc C��>�?�F���A�Jj�b�H,���C1B��x���S�iW�g� (���+�{m�S���۾�`��%tҗDt\�j�2��4#)5�j��B+4��:��[��O�-7��x���>����ژ嵖���j�  ��x��&�cT��3�N�R�jV����A�� �ٕi4�5��"(�兖lc5r���?nlK�TFT�˄|�X[c>��@�ɉ]�8�nK��g}s�(��K���X�wp�vF��&s藗��qK_i=u@*����E[֦F,3��PfT�"�:�uK��R]�il���i��p"�L[�XO���<����/�	�Fj�P�	`�t~�g�A�7�7Ɇ�2�%|�u\��w�s���]��E�{Q�:Ҟ�d���%�"Q��h��W���d��)��x��P�& �����2�29�����&j����-��#�S�kI�a���o�ȇ�YV��%������W�����&F�8R���%d�����L/���H>EF�����)���ݷO�����_lM�b}1�)K�5�ߍS^׿��P��������
���Qf1w�^�P���Йd-Þ�^"�u��C!���}l9!#7�̐�OZ?��ɜw��0��ֱ��z��zm*�%�mʗ�펣}m��i�� y�4�R �n!�k>�a~���k���1��;*F^����Yt|+��[c�gl��3��^��3lƟY؈�A!��C��K�"9= �O�ThGIR�,;�0�en)|��r� ��<����$�¤�;���^m�{v�i3�!l*�Y�m+C3�J
����a	?,
��zuQ��� �>���sO8�p9(�������l�z��`���*;�~y�^�<��
��k�Vz�
�*���d���yt4g
�=���s&[h0����oJ>Ǽ�xh�c���Xk�B����@�(\�Wl���L[no0E劣�b�9B	�N�]8��T�uʠ�֩�nYR%Pi;��#J�0a�R�nd�~�f_C])V��"�1�@=!�kJ���Z��[x�N�ߊ��ӧo��9�+8�A��Jp�O+F���X�m�k8�v7^5�~h�^K܈S�UWne�<Va��m�j�P<9^�.����T��n��ۿ�<@Ė���+V���8��{d������9�ja�q��m�D��!�PQ0p�	�"�1���̃t:�!K	�x�N�GU%hF����2=7b����fIMw��V�N{����Lo
�^���G��ǟ\�|�
ѪU��b3����h�t��_:"���9��:4u8��L�؅��2:np\�݆n�Ɣ�pp��ΒH��t����|}����%�,�ŷ����W���$^PH�G<��:����KL� ����I��4�@�k�������0\G!D�r��P^��W�l�Ua����� ȇmy2a�˖y��k;Y$�C)A8O�	`y�B`5��U��tw��غ���r�%Yb�C�:��z�1$\J���dI�R�M{��������vծ��n ��WW?�+��Z�E�$UIfz�x����iG��n��"s�k�W�=��N#����10vC50�L�G����g�#�4_�;���Z�D�B0fdɈxn`�o�#��ǡ���ፌC�^�WJ��B��n�T6�f��}Վ��
=>�Ӹ�^	oe_-x�2��@����-o%3��=�)��8��a���O�-JB�"�����C�i���j���9�^	���e/��-B?��@fU �+,�{��%�,����|_�ڎ%^�o�Si��?GJPj�$c�7"FDg��DC�P��>�$��P��b�g2�E�FR��i&�e!��\�@TJ�s�x:�"b:w�Au�8)ܓȓ#h^W��d:n�xȞ�������f"SQ�C� �ݫ��#�I�:��32Q%��U��<2z��ތ 'ZD�d�J�#�UdJ�N}�U{��a�*���k�Ba��>�'Z�}��fދ��A�6i;��B���*\���#���d<�j��j۞�I
+2A��)��R��v*�ػ!�g ���7�O��'����`di⬕��$�G��.�6 Շ�������S�;4r�P�/�Y��h'W�����EQ}��,r�e:aX;�y�ġQ��w)��tt��]�T$�s���?8��+�N�
^Gq�|mؖ��&�~��	�ng���J��\�_�2���dE��x�Mڀ�NN��*NB����'���65"H�8QSm���r1J;���5��3|�Ԅ��C/�������I���ٜN��`eީ�'�`������
�t�_��x4,-�q�Y���r��,�zU�m�o�h��#�W��-�?u�NH��x���,ٯ��+��œmncLQ���Z��_oW�Ւ�Ԡuw������v���R����OX�4��	�]�1b����t6y���wM��R_1Lpe61����2��7���*sD����]o菎Fm� �[V��k?���q�e�(�\��)Cr ꀱ�p4�C>�(���5���A)�/b�N�;R����d��|Zdr�wV�K�˞�e�3��Dc�,�~�[��0,M$�v�5G��x�[�>=�G�s;��?}�8W�d��鑲�1�C���S�hь;�jʙ��> v���e���PaC\�S��g=*Q�c��I�Η�rÆ��L�Uj��K=�u��6Ж~L�ԅ���$v,1���� �ԭ��*X� �p��0���X�:Tm}�'ܧ�E%����=,�!����X^�id%�}c�Y砺F�:���Ϗ0F㼲�?��~�YI�zf�*�OT�j�<��o(:���V�h���ab�R��j~��n�r��0Gj>�/��)Ī|3����j��E��^ApUܡ�!2G�5z�F�X���$ǀ�J�`�Z��Ѽ�։�J(���!��Ja � $Fc/ॱ=�$Z�����j����X��u#7{��*'Y�#ȃ�I���,.���ɴՐ��4�Z9��459�/SY"=|i&[T�e0M]8̜��Y��W>��Q]��p�v�z�r�IDK�B�6e���籠_q��3�f��9���F͍�O+Y�o���d[�&�_F���� ���[?bT;�W��\���.vG���-�r�
��Y�ġX�@L㿍^Q7
:;���cqO��TB`!��5*�%�@-�X���%�O����Ơ'�W���Q�C1��_��ł�W|�NZhm��7DP�݊9_�en��P`HTy�i�<�jr6�X����������.L_�':�,�z����}�939�j-q�f�4�[GV�FRh��u�z'��V
�}
,]����Z4V����ζX��S��F�ң?]Z N�6s��Sb��-o�Rr�����5<<�����ȁ�6����F�$M4h^d�8���vSl<H/�
��jw�I�28Xa�}]4̩��a��������b��t�m�� RD;ޭ�7�f�ť-�٭K)U�m7���i\�V��m�-�|�=/�C%�Q�C�������39����@QJ��������XF\��2�Z�X�e>�L�O��%c��O����]��d��of�w���X��V��M�M�b�\���j�G�XuWeD'?h�j�#�V+B`�o�#��+?�l�p�?}tw�x5�$���d���q7�r)G��M*��5y��5@���~���d��O�h�$��Ӌ��"4�WO����'�y8^
�{��-��F���jNo�z[�Yq�,�x���kK��}}��:o� B4X���X2�t�+��Cg�X�G����<h�������/�̱�h�6�7�	��-�	�ܴ�#� ��<�Xϩ����wޭۈInP���<km�Suʜ�Q!��`?+g�� 8��@W�W��U{/S��Qg��tܸ U]�f��N+����~�خ�����^]�C�r��7T�}�����W
m?g�J)�1eG�F��i8���9�����`�BX8-�� �����v�nQ9u�Kp���z��pwT��1^$d�DF�7a�x�Fa��Bq�n{F����w�L���]oy�-)�1��i�U$)~��z���w�C���z�\f��
�����TE�U>n)��5��3s�\�I 9�"HU�L7��g�j5���Z(HTeM�MRPP�uZZ�M`��Z��-�B�x����]���b�B���.6�)-�C� �3����1��n���N�8j���v�e9��3p.�P�-��;i�Űq�	��������K�Ic�2�_bVXU����Q��W�!+W%v�Ғ6rc������_i��T3*��̇�I3)o�{+��F��p�OS=$c��O�h/;Tݟ�qwԳE�`ݸ9T���G}�R��2
����;\�6�����	��7��w��1�ՂC�=/����Q�hA�pE�FN�Ǳ!��N�0f99�Y��Ƿ
��I��z+r�7���9
sŊ�.��ݐ;��*N�5b=���p��Q� 0�f�x����x���O5�7���%*zq�eЧ�ܝq�SB�)��n������e��q�#�z���P&A���Ä'Xv�5�	rmP�⏵�+MK����>��,H�h�*�R�<V�a��d�6������lC3�$��5��Oj����T�����S�7Q�6# $'۸"��f2ܡ��݀�ťB�E`c��fg�d�xt�?}p���Q��bn��R����mͲ�7��{ɍ�
��k����tT�%ӛ�7��Qp��1tM��L��ߟK��Lz=G�*������բ��<�F{S:�|7�������	u
��Y��3u�����
"�؄
%}Q��2Zd7W�=fv�w����`��-,F��Da��L�1`��b�l(�=�N]d���AtĴ@7�F�@Y��R
�b�F[��G-���$囙5��m�X�5#X7?Y�؏���TG�e�Ej[����|59�#V�/�EYcE����s˯�(꜒8I:'�
�U�ʙ7&2zW��S��^��䣠\��ڮg��7��:�I��+m\��p���T
%��;��н�9X�GS���(� ҧ�|�ѻEG��>b�������9z:>�j�w�*���w�1u?7�[ �@�ɴJ����	��t4���~v�>Ňbd��n�$'������8зi	V���éѢ(������yLi&)V��d�g�I ����ɲ�L)÷��<!� ��_��1і��3[���������xZB�ʖJ<O���e������k��]�D2B�*S��W���E��h�u�H=S��%d"dcv��-8���3O���be�D�ӿM��C����}����`���c���f�(B�X�kD`��p����J����2Ş��Ь��E*�{��m�}�9G����¿��i*S\~߶ᔷA��X���L�n_�e5P��@����֌UT�[������4�+�uzJ�9�:��������3�	�~� ����0���2g =Z��8̉V�wMD������Ę��');���8��{�;&yNq���E��0��4�4)7���Lg���}m������s""�OD�����i��/��� Z4�\O�k�0͍�2��q�Y�d!����,Q�!'��l���Piw�qH�G�&9M�����jSz�����:+�`��N���C����7nAH �79�U�� � �thQ����y-�h� �	�A�4Ǝ�Ϊ���&Y�����݃�_����S����x����#DN\�ɯ����������ty�޷o�޳�9Ex���ѝ@�H�ڝ�W�9�ֱ�ʺ�Ċ�*o��v=����1�S5���.mf}���F����
2��`Km�9����^�����6�)��CYB4��L�&��)7ﮈLA5��]���)�+:�	��&��*,M0s\C�dNJ��2�P��y����@���Sh���A�\6����f��=���t�"��raUk녿��đG�*8�!ة�e=>xb�2!e�����h���%�Q���/��	wҬ��lD쎯��t����(WZ2�=�-��G~P��eE���9nC4\��{SJ��%�N���h��Lyg�"N�ܭ{˸�����b٘ݠ��#�?n�!y:�*{��ao��3�29S˕<J�����\�d?F	t�T7���.b I6�n%����?����M�z��ne��Co�!K�F�F�[{�u����$�:�T9����C�m�J��'���̭xd��~�\� NSE����8pG�Ѡ�^~�}�Ǯ�JQ���\�5:�,{܌�-��椱���q�폶��no�Ç��� ���fo�^+Vf(�݉��;Dsx�x�V���P&�_���$�>i�k����eY��W�h 
��K��� �����.d�k[�v�ռY��M���>3
�{z�X���ؽ�穄�	��������r���RG� b���Wk�U�R㏵9�M�q�>[ #�>�OB�7���u�oҜS���o�
�g��/�ґ"I!�������{�}��%�i�� �ftz����٨L	8�;,9�/�ꨣ��%03�*}���&��b%�
gq�i7*=�xa8�xŝ��`���TM��"1�
��Or�W�?�r/�v-?�q��2K[���lm�Cy����B��;�Q5D̏��jm���s���T1�@+\�X�Zf<����(���j�DV�o�Z𦁹�
���]/DΨ�vܮ��n�����z��6:G���8��X�%`�2���7�~�L���,w&5lΕ	 ��D�3�{"*w5�Xs<����^U"�*�X�gj�����1���|�EX-�#�-�oM�c�"C$��
��~*�r7��U.�V-���<�ӽQǇ����؄���亃,�@�ѿ�B}9�v��)�_Ϸ#���&��݂��&������*}'9��G$��E/� {���	����fB��@(��U��Ƽ�؄^%q��L�(���S�c����/lc��[��L?	���^��:d�3f>��}�D�j՘5��BG0��0A�ٓ �{R��cz�5�y�#�W��t(����;q�r5�&��x�b1�x�)ぞ��G�i��0(���	�}�=0��3{$��I�/���4���J\���n!N O7�VHW��r�����t�Yg7Ο�8�}%����vynyP��k㶒����9O�.2��\%��rN3ٴM�T
ˆ=�2Ɔ� �"aO({���[����:l�[\NOb`��NM��´ E8�%KQ�`�-���XY�n6Ǉ�f��mD/�����:���s`}��aӄx��M ����
[x�);�"s�������0~?j��<���̰��J�ջ�7�:�Fx�;`N�+�d�/5;�r�rM�k�'�+���w�br�a#���exFL��X���@���/b7{ɠ!4!���*�n!E�.w}!�Uki������r$�1�7����+U7�^��;��.����>J:��W����de��a�(˖r_�_��Ȉ�q��6m-"Z ����X+	i@�'��t��ՠ�JJ`���`@܂�q�6�<� @=�ص">�y�$��4�GOC<',�������`(��� {�ꙥڭբ��������O�~I��Zk���pgB���JP8��S���o���aMپP�|������08���JK�Δ�d��9�{���m���"���{��k疪�)�8d�U��V��E2�,���E�?��MB��!8n�?-B�a��ኰK|�_�h�&��+�
�:a↝7k>��C�z�\����l�D$��Ы�t�+W�w^��%gw�a����YE��7��f�7>7��.>3�כ]�c�s#g���*D5�R�Q>�V���iq7 ��΂���PD�~CT]Y���(�Frخ�~%l�u�1q��ۙt�rQZ6@���ԉ��_"����1��epjA���G� ďd���l<u��N�pk0��`:K�7��Ȝ�âx$N����eo�� ��	�����6p�sJ�`6�(XR��
���1��X�[[�N,^���6�MS3���8}��5�Ԇ �r5�;�":�����OVYO����d���R�X8�R��[ '��!H�_�G��j\�Ļy�ݮ�33!n��h��5��IV^�b���:�Ê��q7砥6/���J]�爵��ƕ��U�%	��SR�X����o�J��ǉ�(���o(4�D;���Ge��C�8)��W6���z)�o�AB���X�}:0��L���pR<�J_H�Cp?�&� ���K�KaH�E��p8{ �e�j]WܹX�ڥL�+P����Z���4��K,���.�_"�Q$p�T�^N3;d�-qfC�E:u��6�q�Y����(��fS�a��މ���|�f5*��@��m�z�X���&��s�e0���^����)NAj��^ā0����Z���!�]�햌����bn���x��̞�����{$ UC
	��Aզ�s�� �X��y��O�|l�Ob�ҏ��n��QN�rqN0���I��1�
^H]�c�)�;���l:{�8�R����?�cơ�˨B��(�Ʒ.a�N8�x�l!L�)`��Ah�&�}r\����`I����1��O�����?0�Ir� ݄�jwО���9��φ�'���$������/��}V����x��|h���4��:�>g��h�Upzz�z9
�©l\�p~�����t�e�&��ߋ��-g5��5�"7�W�}$,_�l�Ϥo� U� ��������\=�#��x�[ɗ��yi�A���:�c��K�)
�!���1���Z�ʊ��zd�n��[��4���>
1k��$�s�s�^"�O�#NL����0	�S�����n��]���,�I�B�e3XV��02%T�KP �ʁ�~ +Ǐ&�9X��DJ�x��qf�қ�ڼ����^��\�� �^2�ѳj*I�>�"9�B�O�D>���ʛ1HDr68u�]d�@6-�eZ]{�	����/�	�'���LkdQ�����2T)�ϸ�q5�G`�B�w=ek�G�x�>9���)ab6�@��0��I���鸼�n�/ٶ �������Vc^�{1���dy`�Gm�
�c��3���Os�)��cSU{�%Ü=`�5k*�5{P�S�}%s�.�� �0(�lmBu�y����"X7e��CU�)���),�	E�0j��������$e>ܕ�����3��@��.˛�+^?�� �_0��a�3�Uڱ���hG��1;�I@����XGHE�!=,,:0xIN)@