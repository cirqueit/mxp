XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[3�e��A��X�,sC��8mg��8�;x��乡)�̿�p;��]��,��n�\"�h�%h�#N����� �'�:��(A�y����u� 2�=�wΜ8��:���EC��j+6�/�!;aFg��g^E�*���N'�.��N��O�w���A�}6����ds�P��S�|�Z�j9�8.(6�U~UcR�Vjp��k��X��c��>�o�-����jxʂKL�����Mi0��ůM�>�����Q*�|��ث4<�9���<s:�tc?��J.H��t0Z=��̍�?KS@�",���F�sW[���I[�B�#�Q'��?H��UB�8
���!j��,�:Q����L�
����!�e2
ع��;�r�m�@�����1{`�B�����<�#�)��U5�AJ�by�Ȗs]4��;��	���{�ꓔ�������8� ��rEL��,C2�xj��N�����c�ѽ�U�J��Q$����3�O����ߞ&߉���|vv_�]3A���Vv�(�05�>N��qWT��V�e1@��O%&�:�d!��,�@F,?eA�y�[]���=�v���K_^�����y(gT�W�[>A`Y-��G��M�y#��8�l ��kx�i����kDo-���b�]d~��(Ӛ!����U�uP��[��b����D#���>x��{t�o�#��+�y������i O��,5�� �Sb�8|C3|��'�~�.�k7蔝�*�2_r�.�hT�qz�j=����_���g'Ƒt�|wpXlxVHYEB     400     1b0�w�M����X�C%�C8���בr�`�OR	-��c��9||��6x�.�W�e�0O�E�so���3��f�v�9_1�؎������!��~�om��Έ�0����~�:��krp �5SH��v�<jQH ��=��8�b���@#�����p𤻒���`��1�'�^��=?�Ꟙu�[�����pm}"(;h�Ƭ�;�g{�
��s!��{x~�&�gј��C��'"0�!������(g$��$|~8y�@�n�yM��W�M�D�痒w��?*���Pl����J���-��|K.�=m�C�Ъt��p��o�@X�a�.�����'�X-U ʋ;ǌ��fE�4j��o�y7Lp�0���������XH4�Ph���N��ͥ��~\}��©���s�1e=X�N��a��*UB6Eu�XlxVHYEB     400     170#�����x
Y��9ԔҤ�6�Z�D� ��?�c�� Q��~�n��	,�ӃR9|n&y
y�.6B���	��S�c�Q����1W�9Þ���J�c�? ]�������Tn1Hإ�S��*)뫬3@w�Om�.	��L�&ШIm���\����/������k;���H4d��;�~cD:�ӝi9�ܩ��]V��L�����uJ���B�y�.�tTުƐ���>S,d����n�����Ƿ�O ��<	*FJ���+��/�:���o��iT���*`R��R�Ku^)#�{��8����0����0��R��,a���"P�r�0j��B��G��I	`��D�Q�Z��g�����7�t�XX��XlxVHYEB     17b      f0��Qcڜϡs@E-���w���敝�_ /�����o �Q'k�B��E���i��1����+���v� k�asp{�񭪹{�^���4���>��U���I��R�l؜�BrN)0�6����Ԡ�5A�j��fSvC?W���C�Z7�M�I�_Ӱ73xY���l~�0�"�:ߤ_*�|�v8���h�;֕����e��irp�DJ�A��/w&�\#�%9��<������