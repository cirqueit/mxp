��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Ї@+����:"�� �g*�j����$zqB��`}��F;: ��N�m��v����~��ɝ�}��吻?W��y�\��4�,��� :8a&a�"d�����KA׆Q���\�W�U"�h�<�@<���-uĺ�oZ7N󝈺�����xnU��������5��g�$�Õ�����ϫ���dP�����</���G���"Ca1oM��t��t�6y��Dƫ�vO��"1aڅ������Bʀٹ���=� B.��֘\��;�3���!V�1���BB��e��c+�\=���lgƎ��*τIGSYK�ԶҠ�9T� @6��U{I�r�7��_���M�-�������$r�Sx ���"Ul(��J�+O�"��+õgJʅ )�����A;� �%S�^I� �4���}�3M! � �.Z3%�ղk�XR"�ʦ�B譼�>׶H��]z�o��Cu:�ñ���؇��ǆc��j7��S�o4u���,im#�cP<<��@Bx�U�r���>#)�n ����X��#܏̣ � x|�B��U;��!�)����Kݵ�{7A$)���kB�����l�Wq+yV��ż�	�~����iA$'��uG�
��3���_S��Þ*JR �ǟ�h֊��ax�@��x�-����1�q���4&nC�}Vu��5���|ӄ��H�I(�̓���C�0��5�90#<P�%8�6��n�R���ɪ~(�63�:m���x'�Y�@���V�e�B}��@��b�����w�r��Q�z�t�t8W-����GvE�%Fv]Z� }+�Qx�w`q��+i�ľօ�C��W��^�AȰ��G�xTI��O�]a�|JEI\<�!]�e�.�f����oϘ�ٵ�^"�Ri��B����v|�Y��s�ފ����C��]WL���ެ�v�Ύ\(���G�����"#�D!�&��}T5�t��zh*4�j\_���U8���Q�-	�UR��c�p��ջ��)���r
��.8�[/���,O�.I�����=o;4����.�"��
�����?_��Q�����}k�^� s$H��fж���'|�W$�]mWrj��+�_v*���oI�t�$d���c�h����ΈC��v�{�[@�t}��۫c��?�d������HAT��--���>mg��69�8��w_�+9�A�2���/s�*�TL�A,�S���D�#f�g�e&M}eg��R|�/I֐�%v����܌s�zx�5b���m�x|dp6m'�^�����S���FPK���._���"('��!��+��QL�u�a@�t�.�[X!, x���)�� k�f��*|����]Z"aDc����崔�s�'�����b��F��ޙՊ��֞�}�<��:yd��M*6��wA�gx�#ے�b�Y$`������h3@�;�
gIF���a�\A�av�@��er)\D�W 3!��̸m�>㼖vyo^�q� ��S���=�ak�ήOzwB����HZQ�idN��wWTU��(I�*��_���\T���H97H2��E�t�����T��&��J��U�nbc�<��ڢ	�_�L��k��<��1b� 7w�7�ӎ(�_p��(Q ��ġ�� /3;����p���uXK�y�UlPv3R���p#�Y6���F'M������i��j� d�>n�����}��'�rn�L(�B�&�s��QR�	���C�u�ɌĶ�:X��]���rt����q�F(UG{��j��'m�8} (���V������5�V��a�U�q <��{td�]�R�u`�Q�i�X�N�
�����mq��Qr�Js,���Y�Z�^މT6G���0��'�Eߏ��4`p�d�����P� �5�Yom�d�Ek��'e���P�/#��&���6��2{��C���%�,�[���ܴ�LT�g���*��b4o?Z:h���'�#��&�3�h>O27���վ�f"x�M�f�78H�-��`���F	Y����<`�"��p��YVK���!v7%����0�V��G�DJGiq�������$��m'�Z����WECfs����V�, kz.�~!�棗�yf��:2m������“�g�=+����xS�y�j�tJv��e���:`mp���&Z��ǻ���au]nӐ�xU��5!q�5��F��q�
�p�y���@�)ا/Q��sZ��CU�-Zީ����Z�D��Ή~�m��("EВo~���k��Oiu	���n��:���a�п:b�`;I�o�a�[�W�rZ�y`.�XfA�b�M�_����/Ψ�\�l4ܑ�z*�'�2ښ�{��b{�3vߌ���.�`��Z+d���9�?#�ٞ41���e `C��M��l�\�E�yNT�,��C��CL�*���N)fM��p�ɀ��X���4N'MR�9\َ�? 0Ph�c����D��Y�f~���ٶ�[9{b��m� s���FD�T�I�u���XWgx[|v�@)��͓5i-�?��k�J�����O��xWê�EKD}C��޻r~o���P��u���|��mHU�F�}������'�CXTn���1"�kv[ N/u�Z�+u��Εҳ�
�W�Ú����PXv��j7\��|
'��u�mZa`�h+TE�&�����ж���_p�5��� ]���Ҽ�"c�~�!�\����=ܤT���e�Cw�-YbC����,Y�J�o��z�So��Y�G<������s��;���(���7���2=�4M(��^aP�<(�㵆��;��G'0�i����P=�%�G����_|j�]G�Z8�f ���*y�����@�5)a��V��>X"�x��"j�g����]�.�6�n�, ���6(�"��Q��A�S_�$�%��/�	���1<lg��� ��M,��Dm�W�\tQ�
��Xw�sD�ge�8�
��M�!�1����*�{R�X�%u3"(4>j���=�O�h6�=����#G�!���,`�ݵ�u�98ۄe|P�k1��{\U~���#��WV�[)�,�I$P�4 2e�B~�m���@��{$̜�����l�R�� X7-$]K�2�d����iy��L���&�E�+�ß�G��wմy ��b�Or��g8�@(D�������U���`a�wѧ�J�1�M6�ą�X0��'^�Q�uf��?�n�"+R7ݹ?^��1r�͈9����<S�Cl�?�w��=I@ײFT\�~%;XU�QVч��d��Z�5*�����F��j�i3���A�x�2S��#���N�I���i]�wy�!�A
ּ{8)�q�e~�Q�^JYO-^V�P�x_��dt�O��ϮSC���1�)�S�x\�����S�Kp pi6cvRkA'k���|��L"<rU��)�����.�@϶q_P���W��l�WD� N�^U޳���\?�����*�qQ��+� �W�<	��o�m`�7u�}'�v�-Ζ������\���&����F�WQ�-��Ѽ��}D��*"g�,G�>Ҫz]�ʣ_.T*�[�J��zD��BZ��'���e:�q�Xs
 7��K ��;�N���1W��'$��͔�VY���~*R�O�I;��js�6��}���+��0������?�q˦�)����rbXB�C*�
��0��6G�
U�҅p�L��Ng��ڎy��-�w1��H�����$_b�AM�hE}#��Q9���]�|���mN���$��I���1
(&�o#����}~h�qd^�Go�����L�h�%1��sI@���GW���U���Ҡ'�o���
��"���e ��C�������Jn!/����9�d݋��>�{?�_X�WL�l6�8
�P��/5�,bY��d�����y6�ղ(���	n�(���誢P��2���
��Lx�:%� �ġ�f,�����hs�6��_�9�|�9��it�u���4;�l��k��v����w>��)�\Ȱ'�0!B��ynG�hS��NX�.����o���ꩁ@a�?���a-�&U_��*�}�����}�bL!��𔖵k	�.���遴�}��#s~;�{��&���ip��l�2$�Osk�/a���1\a�ۓ���Q������^�r�������Rr���S&]g;A�96�BEL�֚�o�X�e`O`�]�4�J�������
Hy !�f��M��H�.�sڞx
��ձ�����ԁ�<j�}.3�eB9�R&�%�ukcn��.om��;��ᯊ����G!���M7v'=�*�������k/c��g�3&O��Qmډs�����}4�[Rp��ZS�꿶gm�!� H�1�T���^ɬ�^\e\��!��)�i�֙ܭEi!2H�	뙦@ :�����rP�ʭ���H�>�f��I�@�ܙ�*ӳţ�[��Dz���5p�r�l�yN��q�0\��~��G�w�(FG�X?-�w�Kڎ��Tz�W�>��ApZaI��CJ��Q����� ^0ߥo]��,>��ԯ���i��B}�"}-`Y�%����D�z�;���w��D3(�Ӳ�q�^�D�"1�	�����v^I�\Fv̋���?Q]�rVW�RNv�-z!�6�8��R�C�W^�"*��Eً��������+� �^t�5B�]ӹ'�|�wH3�X��5`�Ժ��cV��Ah�?E�����ބF~�8O����*�����g��gZK^ڎ�	�#�-lz���9�~<Zi��#eCS�����i�흮�	�aּ�n;��s�B��}s5��f9I����<v�֢}�𐡧��������r�7�Xp��5͸�?s�&�u��&fᅝO/j� ��O�i�"I!��D�oTzF��(�?W6��d�^����'Lc�!1�g{A2"�g#{ ���P�}�,�����(�2*�T����t��R�M�;�%3�v�Z�Ul3aEݕ^�68"F��)#0�Z�v�lC�T�|@�ź"S�h��o�+�W����A��2�ψO�{�r�p���g���}^)�dJ��lT�{=�/�q7[�������t����A?|H���r�7�֊�k�Ƞ��[	�ƞs���1:l��
�G���E��(DfT��*?�6�����4ϰ�.X:���'�x��W0�o���,߯��e�O�_ߌ}��NV���"�s_&��	�E��r<B��o���Ƨ"���7��#&�y��i�:"��"6�T=������l���� o���YTd?;-nь"�9��DrJ�P*:٥��HH-���Ω�\�)	7��99�Ru`�l����l��Z�"�8�%���R�Tg�T[�)F�d�pok-���	9f���H�I\�M~.%�qd�~~�#���6>�gD��#a� Rt4�q-A��Qy��U�P<�yH@�O��.0�ӢͶ�T��?��Rk/2ЩN��R���	φ�D���tLV�.r���t�Ͼ���ڑ\$�Y���enJT�=�����Y�����K&�-��R}���B�#�]��wD��dO4��ֈ1���KwN��'DQ��֝���@��������R�Ң����D��F�8��@<\ЩA�
�^=�a��zT��U3�����i�?��&���"�C�T�/+u�$���6bT���J����v�L�_Ø^B�8x�1��|���ΏG�l��$���"ēg��a���N|�ɘ�׃�`�������ʫ5{�6Gw�rz9�	G�C��G���}�/���c�
F�Xn��&��?))�Mc�!����<Ekm�h������"	]eL�>.� �R�
fX���,�4Y�&K�B42C� �`p.�5b���V]ҟ��'#���� �����~D���}ޡ��6?�K���l��e�ĥZ�Д�HH�����C��i~�>Q�jk��y�)�˸v}�Ʃ3p�� ���a"�CU���e8�19�
���9f,W��'��.Ζ��ZZ4�
�ſUv�C��ǰO�[ڞ�ȹ�I�8��z���at ���ZI�
�+a����g�DZpX��� 5�����s�O�5SX��F����W�$���oMF~�M�{6�d�l�e1��\wϧX����zF#>GW�?F��V�/��M��6Iz����Bq��9��o�>�C`b�"�^��v3������&�*�p�����-�nf>�7�ʘľ�eh�&ں�\�����溾�,� �I��k�68�����I����cF-�m�1��5Xq�N��!�|ȗ���i�� x���7mAe���Y�,��֪x9XX̇�]ݕ�M�G�z�l��ȃ�w��Pl�M���Tk��Fߔ�)s�$�&� �K!+��3��;�Ĝ%w��ɖ����[�d8�㳌�A���&��fJ������ ,�����_�h|�B�J{rd+�4\�^�A�Ұ���rSP�V����N8,F�4������}�=�����P�A�$@-�.Y1e,���=�ܰ�07*�7�}�fxկ����͂�H1�H���c?%~H�w_�B��5{�)(�W����r�=�3��w�=
��c�(b�	$h�g6�����4���y�)�93;�q��EE�B�1.�����Q�ڪQ��W�R�`�j���͕e���Z���/ث�]��F؇jX�.s��7H�8ဂzv�R�6ʆ�7���揰z��N|���C����_g��2�&!ٖ�蝐~�##�"t��Wΐ��b�e\�x�|[��V���oh3��/�bT#��L�X.�� �!4�G�=�aF�]��x8�::����O��?�~C�K����w���9}��E��\�Ey�t��7#JLIb>��m-#���b8"QT�0��?zRM��2?���>;���i��ҕ}_a=���m��k�~.��HP��y��zo/O��O���q.|U�3��,\�d�`'Z�p�}s��|����%����-<�@:O����K�I�\M5E�>	�RTE� *{�!,ǳ�Wv�'	~*|��{�6�c�6N�>t��8�а�g�5h:c���H?bt�@���e�Ϻ_9��Z� NP8��� 9���N��X�_����4A��7��BZ�4n���)��_\Y���`Nv�
���c����k�w���9�6hi���D"�eq��	R0֭�ּs���r{AA2@�9Q�B����;�����K����5[����t��_sc*��=�ؚS�F%^�Ҁ�,��bG:`��)��6�_%K��ɿ��&g*\��}h����^�t!/��J������0
�I6�˘�q%��b�ܘN�AF�-T�bC� W�+�F�	�����q<a���_����m˪����ke����� ��r3q{��Y_�<khaԧ��^��ոϞϔ�jQ���a8
i�&M�]���g�O��n�K��Р@���|�׀�Q
�e;��ɔ���!��	�NTKx#���#L�����zn4�V�����Xf��ќ�������3������Ɛ�#y�A�?;"�EN��Ϧ��+z�����	��#̝B]�q*fh��zgq/��w����^d��agB�����ů��bP�C���J_�^����'kP��г�;%�<�QcF�ށtX���j�b�����x�:�����c�gTO��{���"� ��I�#�n��ZC����M�(n6Dec�S�t��p(6��Yp4���<h�_%�c[�LM���(&���C�q�X$_~�����=�_E��(�wF��ݕAʵ�ƅ�JV4��iuH�͒��|�5
P���,;�����[�0�E��,�*+�/�,��d]3���%��jO�V�z��:Yu���(���������i|�05���-�-�&	T�O8��T�����}�L�l���.�Q�V�=��*�+�[Ė�*�fwڝ3~�P,��o�g%���=�I]28?E7��l2o�"�^�^�?1�]�-�<�kT�2�����ř�-��T�B^�.�e�H�X�`�U��h�!�4��v�S$��� 0 ��zCT��|Iu�����cs��@�πn,녘�6(����p)�l�~�1��%5�xL
1}ɐ�7�W�h��gG�1\F-���N�Hp�as��;�^
6s�E��#�)�"\[ڏ<^7$�r���"��j��o�,�mT�잧	�W��xb���/8�`�қ�ҩý��qg�	a������!���C��o���q�����9�Z���j+��I~a__��祈��$?�v��9��<�5q64��4�ٚ\�u�V�{�D��'2�(���_+�d�YI�K�b��qU��f��c�5����	MG#��3a0�4��M8l/	%�s	�6���2�u%����:�yq��;a"�4��݈cߡ�S�����9��<�Tڲ��Ӏ�&.���:�dIX�IE�l�n�Q���C���Ny���F�]�aQ�>pV�����Ъ'�mU�+,���!�?Ң���p�g!�趯UTo�nd|	� ��*�f$!˰zM��4!.�O�յJ�6,L
{���SZ�j#Q�� ��:�୸m~,�[�ہ�u@��!L�`Nv��X[�6"c�yL��_��mFPKv(�C��]chd��_��_^#T��a䯛hm��5Վ�B�`q�b��JW?���S�bg�o�躟�3Y5��W�#�+azy�Gu�4ō}��<ϼ�Er�t(���ʊ�g�+%y�D���O��Ƽ���%qL��qFQs��ߞ��h��R��x�M�}}���>���g̩��p^'mխ��Zb�y�fù�w�*�%k��'�Q(CQX�-�~�|A��j�z�M���L|��:uc���ᱩ�s���4����l���(�7���ˉ0ϣ��h�?�C� ��1�Dr�z�ƛ�t`�������;�Y?]+� 1p�4Ŗ��+:�D9#�%�=V�UB�U����XJ��S���Ap�RLٺL,�;;%ŠD�{c^�LJ#Mt&�n)iЇ>��X>1�"�(J�o��ػ���!��͵�	�����D�Y6'i-|�r�c�J�ɉ(ٵ
CNk^�5�*ze���-Sϟd�%Yō�Yo����ϟ9��;R�ϻGӭ�������x��.ġ2�ڶ���~�,�xՏ�4�  ���̩P%��q�B���$����,�[��1C��V�j��\����뮳�Гq:x����6�����/�7�C,x�
�^4V
s#�n^�V�"�<�fhQ��� .�(+�v��u�Ӌ"�<����p�}�aT2�3ґ��� |~��)��ANG���Ɋ���!��Zw�̺�ED��$J��KI�������E�s�}j�]+Ԏ����E��~��J�`��qZV%���rj�j��bޣҪ�Jr���O�H��PE� RG�����\��u����os1�\{�\dRCq_��;	�Q��y
�r�Uǥ|m�Ҭޒ���nn4p�ő���5��O��#,e�=��D����4��n�V�������q�EC^�"�lXO��H�&p9����u\���(\ڐ��&q�;�/W<�7���kBF�BVk{'Ā�&����zh��^��>��M/m�@���^R6aY�8�4R���Ve�c���'��QfA���=e'��	r�+�w\��n�L�g��O���p�L�7���g������_��+�&��<�)-�p�U_Æ�V�W��,g��G=�ܟ�gtHm*ȶͤg�{��a�Ɨ������UP9E��[�#2Ez�F�8�wO�|a/����֭��l=�����7p��Ё
r�n��\M Ux-�V��!��C��9�Ͻ�����*����} ������F��m�����Hw�DDO��D؎PKD鏓��u�O
3%�|ZV���(�.��>�C�z鷅�!��i$��fxK�_K�Y�x�?M��n=+�{JV�d�� >c��5��(8��O�>*���nۍW'49�PP�;�;O�
3Y�a�ĉy����{��leu����>=��ឺ��eu�����	�L&k�M�]8�܎s�xL�~,���3��<P-jj�~�|��o�]��f>����`6��3�Vw��7|�S?��P;��꩙�i)R]��a�J�N�6{}�h$������-j�V=_���\ʹ���G�5}Ǣ����]�u�<��	� "��I֖'�C�mq��1����Ͻ�kG�f<�L���B�ƲX���W-��p�P�&�E��T)mn����i��P�sok&5׶X�����m.���}H�ə�X(!���j�����\�|�M��?�x�Ax-/����8�CSe�B򜓽~<-���7�������rk���{�n��l�-p;S���I�>�ڗ�A<b�Kx��aG��Trv2��? ��.�'�	]Djo�䁒�s�HV{�}l:�#��W�2�`>�a��JK`������ap�(�K`	x����X�Ӈ�_I�ȫ�$@ne��ľ�+��IK�G[�����k؛ݤ��f��  �����v~���忳.�	�腀_�>�쭑�|���i�����?QAQ���%V��bQ}$����@ ~0F�a)pD�)k�a���[�
��|��VH��� mNm9�����6Z�!�GB_��)͂�}��95S0Fצ��D:�铎A2}����4�·sX37X��o��tݓ-�V]k�>�෧(�8d���Ɏ�WBy������D�+2��ބWxgn��r��,��7o��Ώ�?����
5��z�"�0�GAJ���nj�*��զ����K��� �m
�����Dq.�¤/b�d�����Ԑ#�4�p��1��#�[�߮� 3sT}I��$�QA��f�_��Qz�������c$���uX"�����څ{�Pa��j���2�����G/��g��!&�4��R6�&�L�2(�g�M�=�ˎ�2���M��HQ�:t� �}��gv�k ��j W�_#IۖA؆b^��h�NpF��Ŗ�%L]�¾���6I�)�5�/�Ђ?�J�2^7�Wͻ>��$�F��˂0��v��W�1.�*�[U��l!c��F�3+��+qH�\V� m����TH�c#LbBЅ.	���43��]�D�w�vN�4"g��j+�ԚK���V�/�P�f���mg��ћ���
YbH�2��Ȧ��:1Z:r�P��%���^*����<������b&f� ~ظ{��ވ�2�o�Ֆc��7�����
p��̗`��6�D�\�m�?h!a}I����V|R�#�y���+
 �W����q�βEӼ/�
�m7����B߂�D���9��=��䄍cG��v��~��}�X�.�D�q�l��g�*�.�%P�h�o��`����ab�)���.S�1�����}2QP�t�e��/}3o�^�ǿ�v��`2��Aw$���MY�(�f6��՝A���ޥ�L��a)�ώϢ�*��YfJ�RD�?��c�
D�3*����}&T�8t�kntE[��V�b�ӭ]�)�A($��Əj��b��$K]����D5GW�:?�j]��*c�ƞ���@�i��T]���b�%�3�8@6m�ea:�l<,9D��M(�ޏui��X����PV������phY$ftB�c�g��_����I㢾���@�U6)�Q�A�}c[���z#8��p4�f�+;�+��k�Zr�`��qL-�QXm�`����brm�����v���4�^�:�8)'�"U�0�@%I�:&��wjɪ��s��ٳ��řt��O$ꙮ�݆Zv�#W���CR]5�y�X�%�6�&��f-1j���;���e��
u�O���%�*�{�CBjI�u$��PeI�������3��u��h]�jZ"�P{��%~*|mx�ۺ�'���'׈T#H
ڋ�V������ ���?K���?sb��̥�}�ev/�ꠦ���v���.p@`��C�!'��[-U�0H�#���!���g�᜶����g�RzR�:V�:a��P��^m�_���� �qӅV$��A��^�=��AG�B��:��5Di���k��Ņ�J�M���w@^U��	ѿL�nT���ӵS��x�ܺu>�<s�.�hY8�����N_�]�-��9rAo9˗;�m+��G�w[��<D�mE��M�,�ָ(J��ד;)��[�JzE������CP�|���l8���F���sQ���S��u���1�[٠|��}4Ugs|8�_~�v��j�p����
�hB�g0w���y�۬'�e�a�ܶ�e��#����\T�gJ�8c�s5%6_D�?��}�b��v�,Ƙ��KI(ٶvL�)��O�WR��g�ϔ3�M�Ph�U7����λ/X ��o�����P.Y��=4�@J�a1���J�(g'�����sR�э�Z��[b���o"t�6!ʸݰ��������S�^v�h�0 ��m��;���]z���0���"���g~��e��Jth�w�1�b��E��U�N�������mY��P's)�1!�"x��"�X�k���O[�v��NB2����I�<��W���î�ТcO�?���`��5� ����UK�Ɔ]t����[8��r��d��ʳ�o	ʦcI�}7JQ��/P�	N2��r� ]'T�H���Xc���[�5��%��8���4V�V��l]��{����d�y/2���Fc֞S�H�V��l:;�Z��c�0F́n�0M%�Y��H@�٫H�\ �nd��R�k�j�8!G8k������l�U�����i`󄀘�P�J�w0�9
:]in������"�W�Ҹ)���`�?�a�"�^
j���-~�����n���R�;�ys�+�/����t�r����K��'Tȕ��:�����0��
H�f�#.�d����TY������L����b/+�gU@��b7'zfmD��Uh<	��:diH�&Y��M��c��N�#ƺ1�BW��p�{���p���п���֘�%�c���b�aH�.����(���ir�./K$�Է��ؐI�:G�
�c���K��Hxn�'{��b�Q��,%�.�V�d�V�g|Ǡ�8��I��'��� �r�WO[%\:ҪiSGV�{b!ľ�F�K"���ӆ�[������q�X�|J�m#�:y'�(K�5��,Ǹ.��x��M;�@��<.�40x��嬆�j.
�H0�'d��X��T��ւ���C�11rښJ�#w����N����p�Q���/UTp���L�8��������v3���%���P�Ux���?��QZ���ɧ&$U.�ˑ=���){�]��U5�`Ќ�i0(]�`�\o�-~MV�D(rc�A#�����og@
�.5���S�T;F���<�A�ۿ���h������&Qj�5�X;n�����\/���G��ڨ_��~P| �7�O�E03;aE��x��L�
_�t�>���3�̡M@8�b>U���gL�x-W��! 9=���fV�.��a����l�'��n�
�$�̒�����7
��KI2C:~�5o�M����5�κ�K�!�`Vl>���:S������~��P�:���sW/C�U����_qMT�$e��R7e/t%����%�hh����{�o�OP���O�G_Dw��LD�R|��2��'D�`_T^�1ۑ[����1��	�v�s|� T0D�b���eTZ�x��g�Ei1��Z^> �	{�U�x��[4D�vt� (htQ���g���U)׎IZ����m&&2�� ��V��ҟZX�y){+����3�':�_� ��y���~����~�{#��,�;M��bURd�3,j� uv#���r���4K����w�3r4�7"�o�����<u�	y�>s}>(�T�����aӓ��?���X�֝��d�s�Q�Z�v��ӳ"��ӿ�O�)v�Yf�s�m���d"P�k�@��ȫ�x�ߡ��k��W�W4ѹdPg��	W�v�Q%��-&�x8���,!ŗ~"�$Kǥ2Z0�iދ�&)H\��B��@��z���y��/Y�?5���)��m.�s])l)����@�����\X�:s�~�j$�7'T#�Zڳ[1�0�-���м�%���*�Ej�s�"�DК��LE�h&0w��xA#��@��O��2�XPL�#2UeF�G��X^�q_(mb��C���u/�V>��M�p�i��,23���/�-6��'|��c��ߐ�
�Vy��DM� �R���!Oӻ?���>+x�;�$N�CB?ȓp�yFm%�FCb�2nnc�m6�<X����JzA��X��r&���K����k˫L׳��H�X�f��+Gg˫��v �kU��l��j:{V8��y�Jm�ɣT��^�{(���y֟���3�){ ���K�8o��m|V�z�X��l��i�/.J�Q����T6�gn��@QU3ϒ�:o+6����Ym��Ƽ܋����z\�R��:�����E��~i�BY��s4sc7�!Es'.�h�G���D��dL+���b/\/�㱋),t�!�4,���@�s�SR��G7�\I�_��/Ѝ mK���G6M����c��z?N�=��j�O����Y����}����T��?Û���o�pxg�82>�C��X�E~J� 0˻���|���![��C7�٩�o3^��ߙD���#*�R ��}��q&����#�~Ū�jYP����"yS\)���}=�f?A�)ư�y
whW��w~�P�*���8�&�v�0����jRfq���|BC����;'aU<M۾	�D���h�̓ �q���,��)�":����"8��Y0^�m3b���M�U����cT�(`aI��*�&�t����^F�*Ul���ɷ�N�*�DMO�*&U��χ��ܞ�-�����d�K�&�,���#���1!BR]�x�*O_7���ּ���; i��[���t�{A��^�̯�s�3�u?ؓf�o�YU�5?L��-.�����i0fp�����OE%���@[�m��l�j������m���LI]g5\y���Y&�<�5��]�s��vE�M�u�Ȇ�)PƆ�L�<�*N=�ޯ^��i䞂]�����T���O�$2Id�rn��2�S��7o��� Ü�#R�"y�v8��H�E@��Jɝ
j�&�H�w0.��U�  �q�hS��TG,�.�&�����Ǵ�w�oA!�uN�շ�!�SBz�v��H?]�N|S*������ع���r�T����!��ZG�P��>3�-��5�v�j����8��J\,�z���W���9RZ�"�q��sg5/��N��*2�1^�B���"1<5����x0��ŝ]�!���2��C����R�fd��V���Ǻ:0������! ,(k�X_�.BQ3��`��f���,LM��()Y�A4[���O��(�G^����l�W+�ZO<�,�3������ٴܩcX�w�NSV�k )����)���̈�*Q�}H���ժcn |�!�Q>L��^e��E�A2�(_���QPA�V`/]�[]~[s ����a�!\
�gPJ4��;\C�Z��:[R�>1W�8Ed�/<�t��$u���ƴ�5����6ә?�x��ᡵ�#nS��M� $05���r,�2
���	U�o�Z"��K����ro̖|^Y/
����i7$Z+1ޙͶU�d�"��1f�g��#+�v����D�������!���׮v�K"+��'*lŚC4&d���G@��1��@�����o^G(���<�4��6;O��c[u�qB�f�u6�:���묋�nE{˩���z&z�F�{%ꌭ7����P�6�ޣ�G�u���q��g�u��[���RV!�w��\�������%�?O����G���
h�l_���m'<`�c�4�/�7).�2XJ�U$�a�#�k�X�̽���>A_�l!����!��:5���lT�6t�/GG��e���_O�r��#���SY딕u�ŗ�ߞ���!� D9�?WU+N�A�����Ej�����h��w=�3�&��v ~�4O������Q�*
d��O��L�>�wxǪ�9F��E/��9���@ '5�٦u{�-H��Rd�K]?��>��/%�qڐ֟z��������コH��$�h9� �m�7R�8��5���I�C���<i���s�D����������Àꎫy�?��vXB`�p�l?�N�a6Q��iԂ�J\�Ք2��h�oN���V� ��R���C;� �TKUh
��e.08L������s�S�P��}_�ս�YL��7��G���&s���԰��U��=N���l	�k�^	���>��S3~���{˾��1�0��t�+bV�e��{E���H�dδfEI1����x�����Gu��<�	���H������(d���z�-:�u#����_�b�q9�ulK'��ܛyj��sԽ��8��A�����E���،<&�8�/�A��