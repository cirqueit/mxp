XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����c���3�ֆ�\��^�D{�94�A�1(�oP{8�$�DH��$^�ٙ�-k_��/,Qy���� ��4T�U�w�������J��PY��uI�*�|�8�}��-y�C��2��B�{�,̊A��Y��EB~.�g������<���{b�8>��vR}f�mK�f�*n6,��\�����ZQ�VZ+��԰ʖ��Ԡ���>~袃N�m�H��:
���h��x�?�0鳠@�/�֙}Z�GPE;a(&rTz��g��������WY�6Q6���0����8�E���c$?��Oz�}�m�}�J!��z#���[H��lI�6�9Af�ەuV�O�i��:��2.g�֬F8���;R�D��Y�/���D��}�w~m����n�/�̋n!��Ρ� 4���v�'2����D���O%/e�}wFw�V*1V�g@�8<�s�C����6�k���-Y��}^���P��:���>(���z�Kf�ƚ�{cS��dQ����c�.�Uzs��8�vܚ�XJ��_�B������LO6wQ\��Ѝ6榢FƐ
8#៲m�kb��֯����u
�xe9����%�TmV��ZMQ>�D��$���-�K��kn�&�|�,�p�1hJ�,����Kw(�<�I�}_^��lխv-�!rz�{���]8KF�@>��!�N�q����6MH�oocI[���O�뒢.�g64�;����'@�|��Ί�]f�6�"�#XlxVHYEB     389     180"��E�@�zQ�@��\�;A� �`�
+y�w�Δ`�\���������(j_1�[k��C+U��%��QKn�و���߯o	v�Y�Y����j��&Y}ZWG�́f�Sc���#�G-.��*�����͉(+D-��f7�{��^�@�;�ԅx'�Pdk����r#�[��B�T��H�t���)�N\����{Z�����>3�j��cu����	
���`衷7*��9��������[%#�c9/�	u��︃c99��-U�-`�{��ɻWӆ�.[鿏h��H�����k�k�J]�D����y7�=�	I=�g���)R���G�_��M��?b�#��m���@F{2�Yr�PG����8��+ϘڝIje