`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12192)
`protect data_block
5W+q4EGLpYPhvmORkA+vRcEilLVoeVD/t0XJQKTma3bClR/6ad1TRqm+r9DHJQZQd5DEaQJ1C2G7
WYOIfJ1zRnYHwsc2eYcM7ooezCrQU0QqQwL2bWeAdQ04FZM60NgPHzc1hQ34mQhHKJfJswVHQG5C
ANDXDn+3lZNxBG4idU3yAwp+5lQlxdfFqtiqpPVZ0iZWrY2w4EylfZrKju4pS8fbL+gJXq6fTC0k
XUUeUnwMSH0z4/hXbEjyIshXJpeDCGyQqf7Q30SdOoLWd8O2sBc6pyTq3rrvfvDSr+6XS43/A82V
Yo4DUdV2hjH+tMAcN92/fUF/raksooeJ38I/rw7mKE2kF9Tn3qPdG12x1iS+NVL5Qe9UDybCHNCB
Dif4svjYeiBwtGO4orb8q41YEOw1Xsz2VtfKlCKd87VZhHeiNQMdi+9IPN9u1DxeohVouHr6XfLZ
2/UtZXgtGVhJhEKPJBGm1OdafWYndxdn/qgTc51KgM5Ql5tuIzGeXjol3d9uM6y21d/z6X38GdUw
G+SwMGlcbeX2parPoe+GohOCqCL83OH4LJqDVUWajwm+IZ7gUO2mk8D5f1JfiOr9dKQ2upbGZOeq
XTveT84QDMuXqoMczmWO187DGig4Dz6PNTa8ha397wcOfHMiTZE6KqYoqD71lkKPnmOJdiWwMNHI
TvdJQ8IJduULKD7s4hrfdFArMfJ5azCsak6N1g6h4fgVowlzyfsJ8oo1+tLFu/plngQ66JQYYVrJ
wCkzGLKzO1ZFM3shb2KPBRyAze537hs0LeI+g2b02yDFSMq6IpBGfxaC7fyr9FWfj4UBlvBEvjRp
IfuNO3S+JEN57XlCbAUYIwBh8gb8FHYU5PtyBbzOPsGpp0Kus/jtnD0A/7fSa9y+ExZ8V099TksV
dUEik7eW9Et79ujE6ivxG5xst0km/W7cFtiBllGBMg+tGTjr08epyAhc2BYBy7m8QepAb5t5sSlF
OiOHjq3KZViRn3V39T9RGtIcucjcaGcBOZ16ij+fht6GiXWSv1TeI7o99AiV3m0dpmiD2hWgnhkp
nGrotMTd3yCib3DaRVFTKkJdHtVSUcyc787zjZ2wV4yGZ3NJwHB4Iy3gx8sYi8PRQc/1zIN8jLIk
zDn905BpyVNTdYXnlN/Wfrv4T1l4AdoHOCCbIA3x16gXZhOaZuMFJiDf6oLWP7m9ATxteE4eQuYv
8y0Is0tF9xDc75YZpZsCQQITmgDL/AgL4wiK4g2/t5i7WJkGvKKUei969ATyVwrdtVtiwY77nHyF
RiFBbFS9ozwA1XV/YSkSG3npQW/TgZA1YnrjynBEPQ3VVdHVV4XyQn9kAsrzYo0BFFH7NT4r8H7D
ddVHQ9+qH5/VVAs997AQkzFENe31ErLILYOgFIhIgf7+jFJDAw+CfBF3dYiBOL6+3ycogne6ZP8N
uuTJPIL+wO9Db4B/Xtf4Md4/ZzdMRvMFPkVPEJ6HwpSxDprDYiphYeEgU+GHl8Dj2X/Z1t7CTWI7
WiJp3AMhf8vowmgzqIjO1yW67B1cH4N4oO/FU7Vov0IHoBxIoXWsL7jKtXBA1Pe6CdURQcxet0yx
yt7jEGmKy+7zC2u6rF8R7v7jY38Y0CIUz8Mq6V5bLSKghLlObI5gdLxK03yog3XXH3753ItT4Iaz
sKOO9L/5MnaqQAO1YYfgMdTXsY79FIMozr44EiYUeQTPKzwQNc/FfIOjUmlOyy+NIZusfi1h91FF
mXWbA/BTF2hJJdeDYcANvptBoiZfydO5QLyEmVLPMqTXp9dwUZltTo7IpbEQyERC9X8dXNACaCRd
ntzNt5cEZgfAO49b3VxcnouMonYJwh7iLEQRKEhooDDrqig9FZ07v3U9vx9lj++idvh/oWC5wEKH
RzQUlByc239yWkiqTqa+RNjbKFLDGS/YSP7LgJ8V5kA3iuq0F3jE+rgiv/YIM8sfoUibEIv3/kkK
Zn+4NGLXQF04Lw5jk0P/NSXqNkP6o9v5zfTmUJhi9wT7jOSGyh0LpEvnIQ5CeeisNSQBIgUZdmOA
U8j09y1n3JIt+Gg5L6W4fgMlSIhilHyRICK5PuSKNMWLv6oWfpKo9Mj9XsQ9yIdP5ColwJfI+avQ
+JVLvQEhrdnssQrfqywf3AsUAIjOz+yqdmyMvIg3nz3EzXcpwqI7wD7bAkYOM/qQ1jcPHN7WwHKU
AJ0PQl68Joqc9j6JQ+VYJ7D45tO3z0TJyhWqjtv5mpXTjTd+3su03Q3xePOq0g0cRA4usDzkWO4N
KRZOsF4y61WOIYBw5jZOuBO2H8e3C+QK299LXemmLsFUVOfDxwISsKhnRYKrvRGpryW/PdkFR3LA
XLcBMz7W8y8GnbYWKfnV1wVE7qyVbJ7qcRpuOsydmR4JMo5/juJSOPALpFtMA80M3NFUNECC6yyN
Bncr07pYssROnlcxiseScMLBgsXzHEiaVD67bIKiBziYflGVGU6U27styExCGQu12pa7n1CdKIKv
yb0UwtoRZFpxxZqURWNHXnuKkee2ES+WU6Gch7HJ5hhYc0salnvockXD9cfUUOMFr9DqNZu+3m3x
vzf/AqXy79b8sYHre47wZkcBeO8RAS1tBzHHopOuLSdzmJBaUrki7dus186hn3jM1QRmscGxra3N
Cy6TMspT1TC93HVKT2Uoqux9l9EYgT9MInfPYC+n5RIlIIY2YaPg9wubUIRrJitKymBCsSiwUnt7
vKXz1moFS0lxylsjnceKr8/lHR1FDbOLZqoc+dwtNFENYjcVhd/jVjZ+H5cKv/PSjzRTeG1Xyug5
jiicbIv6JL08reGvVFgpuHYoZguWtxH0jk7IEnuiTwiXI3PRFxDQhkY7Hj2IBxgHjFX6GJzZwYdk
nIeWAk7D2cIfJZ32oGtiaZR/hlGVEHo9jmYKx7bgaQG9Q8crFr1tEU3c92jtiM9auN/lCJuPwUEG
hZ6smfGPByAONmt/QKT4guyTzm3gmesJGLVrEW87P7GIKgo+mUZGijtUTaHdYn04n2/pBwp3njLR
bEQ5kXuOrKDuZXznlPBrNGKr3rCb3rgQ7HAxr6VhIosUuCG5WPU31qPTBn11QVk0WydOp5J3rcUq
bJlAdK4lu9jvLEVhbbkeVjYh3EvUY2HpxEXDDF9A+BBmIftq4bZD63+8prBr8z+VeeFzFm/cTrv1
VTiI4v+lsIWFEg1ULdvQG5KRmC2h5GX3RNDDlSPyBZnvAKReD9y019qm5x7bjW+QMpO1eGYBZ0Aq
P7HAojjnDmcEXAb/lApl3v2aCHsJYRJ/LSsJ7fHPZdtsfP60TGsCmYBahY4RLBECYXuImCGnUXLz
AznAkTyABl+wkycFZC+l37iL/fuvHy0TnHT+zls5LH6xqh3dHLhIyAwJwD40eDSXfVt2odf4A5ry
0mggVtsijQJ4EEDhvDxYSWy8qbQzZVkKawo4f5tTFqke4siFYyWHL6HLiwLTiOrbbgqZHW+0kdrU
NOmCk0PIDfW+MCwJApQq7R8c3G8x9eYBgbq6OUydpjKfdqE+UWogCmCrDSHgKCn7wC1TMoru7BeJ
Gg7IZl1nFVcdJSMoHgN/o7lt8WJ+t4RpBkZIoJC32lYj7TLtVrFYtHZrB3NeNlIcczE6BK2UnWcY
+b0z5ETx05ty/vQ2GTdAX7Vqm007X9R2npazeoQNgP2iin11JkReqOGQQKP6rObGWyaWm6OkIli7
QN3407t9APMpXw5aasZ1ezI4/NbZ2PIjoFTMSAVKZUy7Bru3mP8Y160Pzx4JLi/cekf6Pg3pTCrn
NOoNSV99Knf8Mj3Qk3dgyxgTNI5CdVK1C084OMsXkA98Icu0BfmUN2RQUK27DceTFoRLxYOzYfop
QwGQsKyUM7bIVy3V8b8jQUKAnW25LnIz0A/UJqA6mqQHsCBxtirdF81RXrhYp3cXBC52BRe4kCfk
rQixplmwrWEj/TLSiZcmvtJiixPk96Bk/lFlWVEQ2GwTnn8t84FzG4TP/e77P0GKpiqqlgsFBDuz
+3l6w1AYdAHsiJXpv38lrs8ADsbPstmlvY6T1KyTsLpnUCHnRJgFE113XuoaNkOtkZ/T9iBo0VBe
H/zev8FMdbYNSZYRNTaVE9AIDv0OOub0ODWXNkU+r0SrkGr7lChjrdipjc5pG4z4k5Nh7E35eI18
22J3rmMmGrSXZXYtUbfY63znLbyTtaORP1Y0aZUwGBy3NpjVApeJ0edldXcBb1a2/6pNLg1pb7vx
GysCukAyiunmMD9tng+ey3lpqnkBYbj74W2lB/1E8jRRH895wKX+uctpJVLvUEOp5HK8kM/TqzmG
iblbRn5asW3DKlYG3SdqiKYH2lulDZKc2tHa3UtQKTyM+FKHsMSWIiucOXSalrJ/t5nUAd1gCBRj
1wOZ3rPljnevavfnFNdt1g4tAvPEjkwFQzA1z7W0AhR3EAn2r7mPeHoSKcjElIEjVMB+UzaYoF/+
b2zgkxcAhK1AZ6DK4Zgll79CSpWsoaIlak9trgsRIplQ5cro9Ias3WwPug7hm3oeLmFNKLBX5lDR
/vsq57usuiqGuyuVNUXk0pAtqZtg3z3F862kHU/vtzzelxz1EgWBqb5Q/Jv95HItv6i4IXVDLOo9
35Qb+IsFuuE9USQIRSv34+Mq0aA/GB1B9fmpqOrGFBI5Hb7ZsazHpkOlLiQfJwdc+xzW9n1uhXNE
OLfRLHU0FdK7CB3yWXI1hwNvnKst7ViPk2a3jWEvh1PpqGIPrIVQJ1M7hgCu4wWCDPxUmpR8rPX3
99oXlP9NGEyWnpWHlCq2Lo17n6PIhKJPdsFARgc44Lr1dPtMMK8NDhpgdg01SgX0j+ieqrzYLD+P
ZtWhctQjKx19+EvHN9lg3cewRC4YpJAUXMPBNqQVR2d7XzRoMvk3B8ijSEt525VQ1/GNELCs5GVv
cKxLV4nAiTlcjqyOO221aPTcUEfG2BcyVbYAzACX4r477g3A5T6k2REwIzOaityN50WPrlRtoGlX
H0nOr/sPzsL/wbJ9qUIaDHu2skShPaHLNLm55/UrkVK5nFzOfLurMeUQXvDjVxXqDChSnhWqSSVb
CvFcOjX5ovaM+k6awI7radPGin7WhuZgolioSvYSOyDPwVZzwciG+Gq1UoAKiwaQ2ejoXVi42Y4B
sjGK9+Ft+XljJ6R2Hk3KPhgupS0GQa1gJiE/KZiXIsPqK1SMoDAAVMx/34FVCWvzGbDEFi2Oar6F
8j8NNWtNrbz4mpwikiqm1L2VqeN2SJ3B4/7uAgSwmuyhzU2J7QYf9+nnTIkqppV7dAWiGexXR7Oy
86QsqhqHJ1+W2/mNhhsjT7C1jyxH3F8yOTcvN85DaKfynkVlcrW20eWZaTizlPcAw5wrMpDH+LES
nrkwtgaH94okWFNbrvtYPthHS/CdVKZCN/LL4HHgrhy5k5pcgotVNq/2B3kZbnwNdm6Hh4R6lrzo
ZUw8yzJH/gtipAaYdYrNFoCyRwbn4kFbnhGf/+e19Njm8Dc6/vwK4fTGgsmbCrMCRWWOpuNxAmAZ
mgktyhyY0L3a8Wy5rI9FqGgwgPLTCgLiYMpyO5BEBDvDaWpbORZta81QF3Q/fhk+phYJPS3SpU7E
ZJbrpXSbRg/bsndg9mPV7OdmhBvgPFWtufND0NLJTkxBEEzNfKSyNSnsMweG7bhFmEIc0URVnSSw
mW/3+/+XUk6vI+h41K6h5kdiHB6U9Qn8iQDuxD/Bgu2Lyj01az8mliaHhJ5VIxEojqjBC5FCSGWC
frlBeezsJg8r/CLiDK/oTwDtkkSY9G8K/gjdeJC7IJR+laAXuv3WSxTO6B8ovkpbXf1J+Aefhpdh
WvPqNH/kAirDnAqlRkDHGK1YGnsoZ/U4ek/kb8IPe9hQ9ErKG13oIvfEf2oBd3ky1nDKO47mUWlf
5m6k9WEOJDaGXzAUh4DvpF93g4O0r4ZEAA0zNsezE/g4aK1t5AFngFCNpKf8nDhd/6dx0s6oUpku
OZuTb7uIS8NtMcgnavKt2Zd6xeNGY9K5t5V3DGB9fzem8a8DeE2a1Zw8LdMCvyMocZjCaXYXMcHs
M+4AQSjjivcidsP14HZCq97vzHEzVM0CQfkBJVf6liWkmBGdBTQnDqa8OyomRZ6S+NLkw4k6rjig
vdXF7wyJbV0NSH2WkRU2zIeZlRaC37H24EyW1HJ0YaW4KVz6Z4B9KNlIc/efX1UuUNKO7PeXwupn
IW0Bj3z3vn0CWvk6Pqga4DqDaRWayKziLCY6YUeAJQc2/TjYF6E4c1g27t51dLSzHQGTRuJwsBSj
Knib5Qit+o+TtsfJ7r/mS03Ww2h9PSw6sMBvox3eOzrtTS6sXL/DSaSniqvumn1XStGVer876Ya4
ZGc8MivmB0sUZ/otjatKRyh4vsIoKaiqZz5sL68anT72MtyplliDG1hk0EicxGbjgEt88YTJO7KJ
WY+LUyzDdb94paOsO3+tRXHBwbJRZbi/crJEMEiOoyUSZiUiJRekySi/9+85RtojntsKEcsrrVla
UoPSKTbdYfxRZloYVsnvGiWU7LP4VIngYplSJlZxTQp8bPt/m/rUdp10w4EjbzkgZ4XayyKXxZ4I
GO1gzm129efvd7o+3JXU9r+DAi20mkVJY5Vo8U4vBcY7sQ28etVz67zrgI/X6QPqV5uOymEhRuet
dtmOBlFBd6vrY3bm9AtyXP/FHqTLhROMwzol5GHuBudsvpzscvHfhsD7qeqQV3Hl4svSLH2ot3r6
DPPFifcTCRmNo7GUSeLn7NFyjQkE7Pw5JMUHEsueHHy7AAPPnn9VbC/Un0uKcXHYHQaTHSeQoXsH
KXQiEFiQDaurRzQs7AjL7Mwdsf6XQw1wU8ouYk9W/T0DKVyrtzmukIfC9C6ITv3ZuVWud4Pw0tkt
5grInUZjz6+8SdUImbKyjcAo7bRLRTuOjBl1OvuvMlb3QEo5sLBBDa5bgXS5UrqdQRqGAKJsVrFO
p0eg+egtSM3XBzL1+XV/54FbZMA9yu2XSJUmhBVcfBBvrQ/MsfcGfLd1Yvf2ilH9supA0QIHe2L9
woj1CxqlhE2CpA2pHqVvSaf27ND7glGqS17l33kLccYHj/Mt64Jd7iD/Rq1vNA20zN6F+nslKAKm
oHgf6Ptp1ViveNITu/kI0QkGi7ZMJQ/06rZ2XT4zDQ/uOCDYsb6Q/DcEnRlGVEmI686ItytnOEVG
pgM6pW2kcBWJPuH0kAFCjbdHV4Pzutn//7eA011c0cPiuw7cjWRlHccEzjPQoBLOchrG2z111Q6Q
uBf7fGE7wkmNbxwFapVv5Ezf25Pbs8fnBhm3LG8yUv85ZKyuyeINJo6rUOhf0Yc0Fk8CRIgtwhfL
VTB9GHxX6veEr5Xl9q3jZRks4+sqpgZYB88J3qjfyo/46HB45T867yL6iR4JcxPQNJw6Evij39yu
r4K1Pphf6ZFcEbed6/gpbhtHAAUmZZdTeq7OqMjmvdlylhXsCtk+bD2uXwfWEjiNbJw4egCId3+z
sp6ROqqmN831wG12wpWQ7o74vs9WeSkGw2STrT+pzEKWm9HBUZl5uA4/L4w5LjcMjq7DZd7XPl5T
rQgCx63Jv60YVlbWR11RDonC4aCa0lYoFs5YPEEPCU2tdaxsupwPQDWpljVktpYxmfAlurlJCY1M
8XjQ0KmFqRZg7GldBmjm71ciPZFuVVLZOwVXBwkxdAf56D+Ob37hHn/y9faZjuTk/NlzySj7p/VE
Q1QKNi4l32BnzunZribRMsff3hm5QXyr9m1w0UG4doj2q9uf+zbLeiF+0OakIBcfCwCvMCxBOqBk
4cDRLAbSG59a0+EjdSWgwh3xNsvVY/c9wysPKjw96FDh0kDA6vBjNdIGNzsn27YwRm9ji2iXoaMD
KROGHepsoHeD/qjX2pB0wPeBLCRN/Ti0dKFHtNHwmSkPZQcB3SZ+R43UHCHjaSxxofK2diIS536P
0ZEEwwX14uTRJQZrv5m/c/8OXS8nT2PE1Hs3k6VThtRFq4oA+Fl+ptGWh32RsyPhcs+HrXhXyQCr
Lj3k1nXgd+k+ySEfTeJMxcQqttjvL96Xxb29qYmGLyy0YJg57dxuHBJ2Y0HLLNBO38cdkXytq4Fu
2fXmixY2m7n+clAgFwgxagH9Pji/sdsQaL1Ilp70etPEFzMF1V5aanPtS17QNet8AE5Ko+ifMgtL
2vUy8WGSyeZpiqoSGWuc+tOq8NvZnTvvGdBE0uFHkqjWfJXe3KynO2kdkjABwjSNPmbNAqTRPaUl
iq+iru+6xUZBCzCXAk5wuLsjsGsNgx0OQAlZ7XRmQLGp0MUh1S0TPR4QvuU2okkK5w2iayP+Vx9F
jTbVYKu034BatMf0UWhv+23t6zWp0V8BKWoYAEOtU1eUqecxUkXkA/1809RnvxiB37y/I9UOQOrW
Y6te32iOYtYdRHdfOT5Z3nV5Xt5dVzCzO6qN0hivgc6qHZFoGgn8N9Gs//mtyEX57DCWhDE1PcvZ
C5kRDHykNTZxbJEwALuoVZOmEXUfXJm7d3D7Nn9XDUZR7IuxqntDOOLQeBmzo1yAM1988LCyodZE
2LoCXxZM1ZlWg4j4C3KGl0Z1hjEdVnYRuXS8yd2dI/t7u68pL8vb69VYCj5bRQv/vy8uajrIo6S/
Rihr1lozZUaDA1XdDDKM3FJ40zeHvtq4UUVPvMi1uBTMzuX/wvOdE74mrNALkgLkHfKxRF1oXYNj
loVCEsHGepquBq6ZIzOM1FVJNSh1y/kQXCd53Mf9NzFbp2O+SAsBP35Xs4zDGuS3h1PzQ+kKsbI0
LIg4KoHDlHBnweuPsX98Bx40uqKXDY4pq1vAxPOooIr5xNA1aAaa8Xmosub194w7JcNONE9C5ieO
830Vh5R5d+ANZD0Yu7M33nQ6gxvwYL1xYsX2Z70qnWGN+xjMDslXDTC/gojI4Q4PaUTsPLdhFt4I
8uMwpY0Gn6ScgbxxyEQ83MsMmhIttfQVspB4XqbnHLeYEE5sUdzPxVwaZWAzNcH5PSSG1B5i3UnX
ZNiOOe0ZIX8QQpdHo5XL9y1pqqohs95+RhBQ/7B3xigm4VGGM6qBvC1ZKHD2YvWTzQdY/fLYIzvy
t6Fo5C+1CvtXwh32uAAsUIy/kUB7+dkFjBTwAu2Z1KQmmLUv9q7Y/tzJ7VYqqffl8r6eSjw4vVD4
RNUnPv/F8RZS/W9gsBh9FFl6d7Dy7PZQ1KhIwsQczVg6drB7U8/k+06MzJnkQCXEnNnbYAhE/7OY
4OsOyY71S0DuncQ5nvedIxRVfmrMFPu7bI37MQZm98Ci2RZpruq/Lnb9OSGMJccSxVyZLLhFEHmX
Q5aUVKSBPUkPI7K1ZDg28G8wttTbWMnUpKf+1z8z+y9yeUvcoSB2q2ah43Zynx+P2dN0T9pioGHF
e7KCVliuu3JJrNZ2fp0cIqGyLx0K4RBAyXsVb8O03UyZn/PekoVdg2uz60mv3IBUFgoQaIxsK1FT
ujsbrTCpTQZ5OPNj3O6LKm63wH0OpbvT9w3BCr/AvUHfcMeDxrfejV0XUPW/rIo18enQqcDQNl4Y
xeV+m/KTDcfXfyygTP5Zi6Akn6CZIxyiy5xcw/UDXa/MUBZg5eKSvhmCCPzXAtDcAjEl3EVxnQjU
c/3NxDsCjWn0y/Jv3cbo8ROP4udRSonXGS53BZrPoSuXk+u844DPcl1wPxebg1Dam0WLw/VxerMY
SW5IH2nUy+fqB+5QzwPdm5Y5f+S6DYnIegnNMSV2SYFRLdcB6nYpQ9EQS6NsbP9n0xwW0Zb3TYsA
WtMWgELiuiZmxQYgd2AhPzygaZVPWjvkqSNJS3rrTuW6nYi19Oqy7NFUhTdU6/0zuo+3PQDnmRBX
kvaXMx7kW+pESYJWQb0H/fyM0cDmcMpjCcokuP67ttsX1AHTfDaun5lftRkvwmHqZGjiQZ3SalwW
62jJwKQLjvQw5EmmAmiYU0Tey0z+mFcXgqlJhAhzSE2t8pIs/Li0RVIdHsJhihYsIcviwpfV/Dit
C3tTcjOgS1jS3LIm96QwSA19tJRSWzaqNdFillUAJfPP1aZ6Mf704xYTcKkKa8qdj4EW63Kg/q8U
hSvfTUYrc0Mz0C2yoGRkrTedmQ5M/zx2TqqRvvAxISuHdXXSXhXDAKqfCYdGJxuTCSz31aAch1U7
rD5Zf3f4qJsbvDjmeUBYTdnolJIUxB+ehWiCG9qPWyR7BO3EHZXEswJ68ElIW/WZwKrFd1WoAoGW
j1Y1yVq5WxUZDhlGP/es4VR/JD7mOiZ8GRDIk5uM6e284CDtj+tcrJGmhDH8fozAPcxqEo1ETWHz
S0gGhsMjaWMK8odTL4AUnfdHf3orL+PrYgEXT9MvQxMPV3FlXh+rZXN3/UL1duqVXMuuFqy20EJW
6gfR0ITlBA4XNvHNgLJ2FADLek17p42j/kdBDQH3pXNMg2dqOG0uwaygpQvI7zoJuQhabn/gDjNX
QTIPv0n2Vaz+LMN2EijXFYu6y47qsP57FG3M7SINxSuznacT5fEy7NMHrALdcLhNV7EolthGepI2
1YCQ42Uvf82GiGUc5xeoYSxoUo7Zso4GEVo8LrGCLw1Un3U9rFy/kOS142gdXev4s5neDA6jktvk
BVlIFyea8Tc+vyb1Pg7hhKioaM6ov/gBSDG57ZADFXIx33a0XhhsYnLDkuaXc2f1q61l+YItbroL
lKd5S7yU1KgPPBiyN8t0zpeeZ0m4J8L+LoiAIT0/mJGoCDtBKVP3SXIP+jYfVpzMffBC8YuqW9ey
AHgfNLM8NWl1AoeqIAS2uNHOH4N5tQcsSMazs/eMQ4aG7OF1ayQLZBV8SYCB5pug7oWn5M+MyqNw
8pZG0PzWBVoya3fy/ZtmEdxaLyaL4xTjiWQoVJfKEP+zctNJAmTQU9W6otqxMmKHYGaCSePbl5Qe
33QU5H+Bq+QoyQHmTKMQ9OfblbUBuClsvhe/Qdt3YBgZMrv9214MhyxFMqDtRyvhCna2F6ouhXxz
o7C1gPAltqhW8Bbj6mpwys1PoiYAmTPR5VlKTvGonG97aMUT85nk+fCvrZGlY8l7Dm30RT/OVn6F
N37x2MYl01xIps8vWM7jNKJkjl9M+/s9VDm+HtYKBAAiMU3gj9WtwBjvCieg/INcZezDv+Q2LGN7
SnORZ8Wx1Ah4iqmk8RWnCCZZ4RnVRw3PJue4e6x/krRQxrmvNZPM44B15zvEdAI4YSFkkVPZMjGS
b8xohRQu5ckmQeMUp3Op9w5tiDMGLTWhmifQoZbBwZvati202o4bh2NYHLuOaE5WufaLXA/H3QuA
aGN7H45udrZGH6g1hHJK/FR01xKRq0NM/zyoiLQ7UEhveDloND90DzpwcAp/TFaIzrubsvkdv77U
FNf3Fo93jvCyNftqRn2/Oe1Gyu5bWNqDTCShwAaPqBNze/mrvzfWsGsVBYfaraWojjMaokZBSfaD
SHxe9Zf+ry+YMLTm+JAOO0E6x4oKZcicDjsaABo5n2ZgIy7ihY2/qYZvlRqgx0hSAAFx/IOX7Y0/
zC1BNfVrNcrG+KR2IiUKJfmu6awEkrKmNU6mXsWSMnceaKmMjyHqN+LZD/n58LstFPBzzeaf/jSm
/8DqACUJwkphM+oq1B36tsgzErAsWhybnwlrMt5ccMDQVIkLy8/35EiDwzSkV5EmErS8U1V0XAlU
MdzfKJ3pTAf7R8V5w7AJSgn4lNf+TUNhkB9NyzIz9rO+bpdRzmBlmdvwSrzUCYZbkAsvSHkB5sws
TlG8QLx6Bd3atWjsKwzORTwnq2SeZKFhuzeQhKHflfKnvu9+FXFOEwkYV6cko8NRhEYLHelsj44V
oauv+Tk8wKerpSf0DdaeWUXsGh0sCi1NKum0+PkS2frs99zT1iTmNc90i86rJEetlos1Gg1q3/XH
oc4NrDk9AH3Lf6mjD/UY1xSNwF0v9r2y7Hb+BineSvz9AuMJZMp8QxKCBSCiWSd6uKk9eYJVSnwe
x77TBGPfui07SVEsBAnzmR5IcCKVys2qblLxm0MwgryCz3PIXrMII5VZvRDD2SWzvXXegX/dyHwY
wCGOUAHI6IfDD6ikNR6wh9wNrZn3ntLYfqvLsJl/Fnu9ALUbWx2gdglyPLKdPC9J4sF+l44AYdWY
93PsAL2nVYDIhmnus+YXB5QHIXKbSanfUWDhlfQPrkZV9Lc42tZl2mf5W8uIA74jgPa4AjSgT+3E
OSEBBMElhqpoGLjLpuzTpyo3SZCPw4jwrlL0sazzXcRStOd6XSdTzGWtPTPIWmbZ0vRUgpdvHVV0
nkHjiTw9qkRIMEpmz9b0WeUT6k/OX8syVKdYk+u+FZ9hbFLd6RRp9nwiekCCttc7VVvHhndNF3qV
WdrlFwrMaeYPwIbZLj/gsGr6ufT4DbRe3k52I1dIQaOMJb95M76vijUmb1n/SgcBNOARjM3yutGw
KQXHiO4sZMuzmTez0iOASTbOnb+iTCsMKPVI99QSL51kCpL8uI/up2N1Yg62vQHBg83DlKzBWQOz
4+5TI+E19KNzy9sinXpbrpBqvOk4xeJgz1vsEcdxcg/0itwN8CGIx9ynIB2wroSlok3IY8eSuXM/
5H7hm5ownBtgWSPTSHYtWTcVTc5RyN6NxPrQxv+rsW6ct9sXDIojPLpe2rYvRSilVOre7dFXy8MX
B2fGvJMgpqL/uVin3nDyIsUzyI89xzvaVOJ9ESLPkr4OE8zGdgepWNkybMSkVi73cB2uqDAX0YvN
zILmpRtYWF57GLuqUZQiOXAkrO9zIboCvw9TsM6mINpvmmBKn7Nmhq72PQMyTGVo7PxYj3PrXykl
GGiMD0G3ZcQzRAR3m9BAePbIayIHYQ5z8/e5N5/IN9XFU7hNxtCkGtYcv0dQyz1fPoZl5szu8LBl
c9oFsbXhdQDNa5fofZsxTv1qXpw9iJfpuGn+w0+6+O1DDCgzxEpjax0rf71BwGinu4djLkGl7Wzn
FH3vuFuL3kDc572iN+twmBQllnvusZj/MAK+kg/qwgnyhjPJizJwHsxAMdLL6xyuD/GdBfo/Qxjz
zflb0dMgTzS2IRhrpUirz5UTw+hALpNp2jdZQaIjd2yvHaPysFhZM7uNqN3Pb+0Mk1+g+nVD8hZ5
h3DU44AehZtOzNQMzNCnIugm+kBBvtPu+HKA+XBpNRJnGLNPG6TPt/5yMgOZWe9erdKxkGkb9Vq8
BV9MnxnKbycqIrE0Ilf+AHGcSdwLh68HWvYRxIBaPcKKsaxbHJRTd+IO+EP1uL5r64EfvQz4BNCT
v+NTCxEPRw6RTkn4RfAYSs8lKWaNZvpVDSJe8PN1z5Ul64p1bhsX2KK8PMPd6Hxl9jpAO8QAwvqF
UTFczJied+RIKln1YK+r5cm6KKBGMW9BcsDnYNHb27vP5mJ+0Rekx34mb2HpGTN1UDghCJO4x6s9
MJBDEGFywZ8Ky76XL4S8dPTyRFOpn1AIjowgacnzP3ipOn006znul6XYQr+bTdpHTl5Z31WEMbs/
2cZYj6eduFglB/Q9jjsado0tjIgzsa7ieL80EzjvKQ06ZNYPCJ6+Rgo+L+4GZPrvQjbHgvfuOdn4
PbiSCJWqCRIs4jz3NCv0Rsg5CXLu9tTZKY3Si12VrWLpn0Z422Ij6ef3yiKZuktEYcZ//gtXcW5h
nTmH0VGpVbaBx3fzEJgpvJExLAaRh8XYh+fIJIEI/sQB1JcZA2unq+qKLmiz3WlBwE39XAsEGOyS
n3V3E4xMkDfijjWFzloZVxtWZOrV/Hto2j9mDb3tYYdZSrzVFtadka4Xlff0UDHQ8zYoB25u36g+
fQmzmf9AnDYRvroNH7tcWNUVxVw1psVI6DWCaamN4UWheb3ehaam/Db2e23vUF/YDel/i1lGYhyF
RMdRxY1VMdBwaMOOoXM9bZ/0F+rkuoQpzvhJ9IDDxZz8ny4hFNjB0BT/In7NfymIBrqUeEvH8nH3
7oGuB/BZabnjRk0DwQIW26vDKn818hf4FaZyDCmznIjeBZAIhTBVaZ689GYCZbuTn2NMNDtd9LhV
el2syubU/zeVl0REc57U5M6RF5YL8jVFWQ298MgZWQ3e67oUsz5Bbfecy6/EZwjMlo0XM5JqoFZB
3KOf6ztjjp7MOvdKz8bQ4vNUm+t2CwRi9jxS7TY4rMozu8qGeRh89ae0y7/AVlsXlWu+H7pNR8cO
qrCXf4kHPqmOxEszRy9j74brHUoA0X2R3QoYSOiXHC5zWgEt2qh5JXjCvavsxmnshgDW3yoT/x6q
NiJX/oyIJKksgTIgrMO5C928ILnIxU4gVCo28U9RhTMV4Ye//bkPQ1FENZankZf5GVCHNsTey82t
xiCadHUx6TDuJgAupmXyhI44Lajui+eDA46KL8ORfY06Q+WzR9TOvX2eIwAnw79W17kEpJtUKlt7
qMc0t/mYEET+mBAWiV+WZvUJvcc+FBTD9rKJ7aLm2Pjt0uWLMZt36ASwx2C4mCdnanWPcsjZZnTU
iJFSvDoC+E3jJESv6zsZbn35ctgmn1KdgzHWHeDBq8eKPwMWKMc9FTLl1tvD4WUXdV8Zre8lQjgn
GeDDTv5V6Ilwc5yDGrhNPJVIgBhvSvvil7qG3FApjahM3hJLRnnJojbT7o0iEBzpaGxpTHJIb7WH
4MPyzYjtlcdGUBoPGF4Lm/BDaoSn6cxN1tRs4FFD1qfgp4aqUFFZ8VfEaO5w/zP0sP5u5lnV8vEE
LTB4mvRJoWQlUq7ogXlmNqvcz854StmkCLGCg37qsxtQhQOov/TommxPUXXfvo9q+RtpXY65MUYo
l88tfBhcBMwDIC8Y9+qHoO550XuN088R0BZPPR50vxKbeiocpO5xpFQX4FPggnPr9ijznWM63Ng+
NwGvEllCDbdMiCHTU21zh/i4f1U1Pr2zANH4dpf44e7t3kpBfkFquFJ9bDJRFn3GoJD7I40wZmMv
WldDf4lI+STC4F47nQOzlNHO42HIbGO8c9tbReyqyZ0F2io9/9Ma8QmZejbdSfBhGSCyL0o7mIdQ
kBjOWS6hEg5Db0dj6AdvDzL6xPGFGk+hAiIDHL7HtQh5/nl2vKVCqPNYyeJ73syiv10lzImYLYj8
QvrulhFW9e9QsnkHSgFUk3Lrq1QIZcTVNkq/k9K/evRZTWnV4Khz3ntLSWQ50sQ9wgTUU7VNPQqU
vPq0wopDnM08vPUi6mAebLfp9woHMG3syZe3zQxA97rCUqdRPFQvE3Ahgf1ved3D/EsrZJRnTDh9
j7ulTG52O+lJDsvZYZAzjcT+XGA2s5BVkQ2t9vUIrv+7mqfgCQmznSiyIVKmr25pthDz3LXjsNEl
bmmm9DyPxC80WD2Hp55Pe8IMduEED5FiCgaJKf6HDKZq6IRO0ND7pi6ujJD7tS21jkOw0N4S9sGY
PyYiqAJwQX5Wu6SQXxPFRfBPirGy6FFSA+4EZLtYTi7BtYV2yNNbYEqMXTDRYcYrCix22WEk9O24
zw+jqK+tq8Zii3wvjZOA+DXmCID3rBuQ7PePZyX+iAFTB7nXtN25ckuv37CP+uqBfP6ZjoCHcCRz
x74ag+ivkTAgh9oTqsUYEr+oaSKHHmh6u4I7J4Lg88DUgJdt3HmuuMdLOs8qjvuVXQlBmPPYX7K5
zO02g2XSoqYHOJcx0jhJque3fb7grYU9uDbbPGYJzEyEMmN5sYRiaVgzyyJeJgj94Uyjc9dy+xzF
Sk5DJxT2wvZk8BQ6DzJuLh3E+8j1uM9Y3XXOwsl5beDO/bj28hYg3ajCcFvB99pBwg7g/kfdmiY9
j5z3kEzWk9vll2rByQ1Aa0G+RpxZw4AXzxriRlBm/g0H00ddnPwlXvXb3zByrjdqXD7bG2Fzv0rc
obZ8BigREDmKPwe5wiqi9hkMXiwFXpbOrsbmemkrdVC90uLsv4LoiS2l4gduSkYeTGGzOz6EHKAf
MUVCJc/Qdt1RCZ7IdNezgFRWwHRpWgyVUAQt5/gAtOoHXmr7G07vubMYb38vWhK8FTsHK7tD1wqZ
Fx48xYkJFDc7AnBKVl67zvllg8tcgbZ/6ddAgBsgSMr2qfpn2VSz955xMRSfh/EP9GpxdqpXqKnX
4WZGwaFCJW1qGuqVv53iDjqg2X2ha28GDwijkDyPCGeWxWt0YtLRB2SLtKRz/NrTtoms8nIxU+wH
tfMnXOv6dW6mzdygPB0goQEV3c4dNo0UfpM2O6G8RiDa4f/2u9d186aJ7xZ3OsyuZYC6
`protect end_protected
