`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
E9CgCl1bJxuMuzmr4ii3ifsdYpjz5ZmByfaOmLG4B//G8cVOSMd7aME9vByg17bGe6Cv+UAFwlpx
KI7HKVD+pQFdsc6tCEfYtRKAjQJdIhN053qdBomMvdhRwwWtWw6TqS2Ca7xEhtSKqfmzhmszhGcV
xvsCM8hhVWg1HE6oV21rqPtCQet3JPDkWCpTqZvEbB00/3Mjkqcdsa86tcRtqKgr6/p6MxuTW1mX
oKoQG9EaaAMjmo5yO6yeV2LGWyLdb8t2utra8NrsVYUts3gtDCRnfs7c4769jRbSIdHYpggiTtEK
SJyAAvZOpqDe2FujnllUssPg4ezj5B+qGkK2ifGt9i82nKIl3geGo6+VDY/3Z0oZdPNF7kbuUSfo
HCR1FzMPy6AzTgf6vnezVAxQ9soncu/C3buL0ynCbWe1CueJd61unACWDNRbWmcWaogNMNcHFOTZ
jrgSJnnvHwWqgBzD1evn9TufW9ZgBMh7jGBLbKaQtkpIPBK+T7eTy5J2QPdxOZBGjXZNydjuMxiy
3AcG+zQUBjxz9dyjUQgkM6x4gXtYXLdfMPoRjyufFTayEx7m8Pk25+2hvjH4zN6BYO0Du3xEhKYu
4nde9FyU0CCUunDKKoAq1K4EC/q0DcZHHzso/wAn/Mxip5ooFtaov20jCBQarYXAHgW84OQW283U
p0qJeeN/+UkmcnBGLtvz9mscZBl+jYo7iUP9i214Lk4G9P9ZicUPEcPFhESxG9G6QycflsRriNJI
y5LCFenAli68JnrwAduWERKLTkiORMw3xEUqlUVqbRidwZIS0pLhDlBWHfYajr282r/CtJCUagmw
k4z0YGut1ismGh92vNKCs9+SpgdMY3UxwSdqL1iJKm1KkpthuMD7D+MHgNfbTfBtBl+YclRz8Eyf
WBWh42mssUxKMzPwLdWBnPJFIZQweo9FYIUCE8ukcqZRn9+LA5mpbN4ndEdnM3fQNku+MTrs3wRB
0X91BU++K4l8aNWbdH/uiZf87bl0x61ajzMD81m2BXZ7LtVpXmSAXgmAnkgvwLtvGWMD4e3fcvQz
L9G4vp9ElwmLnTtkMbg2WdJhr6Vet3Dszy5sRaZALN3NJ3tbdgW8O7CKB8LVABRtMkfOwpJWxxJD
/BlPpmJX+PEtgenhnurGC9oMOp+c6VOag9K4Lrwt8O0sVzMp0ySkgbJWxxkkTpBLwAG6nGsCqv4l
GGtBoug1bDClk5ogJe8VPNOcmj61uUyAExGM0Zwo+Ogw5dgtUN5RNcXUmMgZ219y4i8ZZobU7n0w
ygqLkEWJN0cwxscqw19DH0VVp3MVhNYg/Ztcr4OebN7/mmwbSRAiKR1vnGohHL3b62tn9AlzydbZ
/CXE1UjtLKP05PkQSX9aSLAZQl9VIQGW98fB5N3nYtpSfTBPLjVg8t8/lXL7S/A0ulocQ2ujTo7k
jIvTzL5pQ5r7R8GWW4ulMj5ngYXfD14rtw8mSGZ0C0g4zjp3r9TkG4i6lql/OHPXHtF1xRxVxq9k
nB1Kl7gJ+eaY5BuVdpsLkRK/BM8YgLZhL9jBN4t+dL59dUpWSqFNSu7xwrc0GCy8zYMQLPoOMjG0
HZmdpheN4I4H3StV9MIlZKrSAJTFljqMqwI7GJt4mmp9mgFh5NvmBMVeWCwFFGIFXDWiUXUuTCoR
0UqVmjn2D8mwM7ETlmqUEqpuI0LqtiCMuDqUyAawhs0M/m09+xnkNG/M21qHdFrNijjCHKD42KYa
N5DWhr87SZAqhDOgMj/eAZMR2lkUtO7n1z2kECZu3Kwp/9OKeYby/9YlhJw/uWzCKb2pbDIARvXL
0XDfnlo/8IebJ2MRqRMHwgx3xAPsVjNXrfBggU2HkYE9Do6mUhbxHw2eP8E10VsYoNl5HUR6WVo8
ISwT/nmVEQpENvU7fBg7+MKf+eTgSq6mBIxnOA9AK9ZooODOWUkKEG/8lByl8BvGvGHZKWvPaAf1
XWDhFkT4LkzxbjqOhXTk775pVFtlKyID89Y4L0n/ynTtKU+RETYNTQBJKXcp2Y5yA5D/UfotCH99
eP45MqBiu6qk25Dmit28uRow6SedIB8dX+G4QdFhRMtEDVZywmVCfFKhJhBF1xapVYtM3cqnrzRH
lZ9/H3RHnKn3Q9cJYphHeFHGYeVAYJHdGS5PzdSg37dnsBRreTTNWl7Rz6BaVLFmGI/YGGCEQuny
mxB+VVUaIOfdBRdtobuX7cVwnAB42RSD/M1O6lEtRfveq6JEj9eYeheOWW8+LbrgUhSR2/ua3mhr
nniMNLbXlg83RLFWXlTJFQNrjEKmwayBOPH0xw13TGhQNamu744MeqHx8gjnazmZdKCH1Ioaj9Nk
zMji/ajMQybRV1lVbn2sBxsJednQbXJJPqgOvCQNqH2+9ZjgXbunYJudoneaHPNVOtsaEdED0TDx
4rOoTKaHXm6UeFqrhMn+xFoPZ5lOO/6yrpPjnCc5E3DwvhtBUx1GrHG+oX1o7TjT1k4fcGzE4kJP
zWJpVDtbBVHbGExEWciUMOV0NhpouaomNn5S26Co7Z/cvFbJycODVWe4OJ6/qhDC+Gk5oQ2fTKvH
fgxpeWe8m/tVh25Lc4PHlpwVOW7acAOLfsNFwjuUKEetv7S6qpEA5P6rlh7weYN54vWXoTp8aOuo
2m+/4GlrYBBPWBg2igCaGNDyf4o9qDEtrkAzjQ+vJacyhR7NOOIyPtB+2huEI4m8FrnbeuvLYzux
aBlhb5Ime2pVbqIXTtsR0du3Ujb441nDCdwrg09emzn1Qscg06Wp3R5KpXFqhO6T13s4kaOGCy3l
mveDlKvhTx0oLmUXnURxK2UjUqaMNHDidcm24cCxMUGTntGG6b9Lhz5w/bzmF/MlqXC6xD8eLK8p
Ark/g086MEvbNvaSU8s+sN2fNwIgYJDFqsRQSYzkkV2FWxlzRwKB+8GYWsQtvKXwpyt7Pq2E9PQQ
T62+/A3oRA214Mfsy7gw8hBEBzccthn942Ey3OsyIRl+sqQaAzLUTLHiO7W0vstxy92cNLPpSSJO
yGgAbyZ+T9bHB+1YZCZ7pWNcSsvdnDa5OCBSQ3TqnCHu0rlqY9FNBSHIh/+Kd+9TnkLki7lIbHdm
I5xnlb7S16REKNCf7L8SCdiQGhnaNF0IznBMmYjQWnObmqSEw5nZifl2Yze+qZ8+TqEQTFfhdqYt
QwwJDEDt9YuniH9PXdKzzvH+4N4ngoFCX6y909IvTDYESPELrUFkg1to6m091cHATMpH6yxH43qe
LImGHcisK2CYXYXLr37kzJFxihHGl/L82T1tXkvonLbXrLUPFOXZ3mOLiLQBt7jV7ilt88SFP617
bZUox1wpaz44ps0lcbfy931UmIw8XVEjjSD7eSX0vU7L81yMbWnsB65JDrFAjkNPOIVjAscON+6t
Pwntra8qtRBD97fPQgZ7ygV5Fyl9bSaXxUIqATTO2J8SoHocnUHNwaLqHPcU4M/nCthRBzNK8Hsc
jTIk2hE0N6/4gbJ8uzR/wp9cRTaZR4aK3lNCDsD9i/ecMPef+W0/mz9o5fUQ7LwRcq6glQqy5eB3
eUKNeJDzsjFvIZW8LCzIayaVhzlbh+FThGvhM+7VszlnuUAlpncxG2fxJxTqlYwCpZ8765wqNKA/
dyqfFEC2HeprQX/dpcHuZeZASsFT4zm5Z9/M5Vt3XaZ9yvHuSQ5f/X7xhjAwiUXHL+4BUhJpmhZ1
4Qs8BfssRbFvXPGzRWVoPedLx9PJqojU4Sn32jYe6+M+/A9e4u51j74jpvyU9o6AAmmqwFRHxrAO
M5a/D7s09LfK3Vkm2M5fct/bohf8MS3MJOwq276P993kjW0wZrQ/1SqCbp/sn0impLHoII0t16hQ
aw0dye5Sg7xPxRtIz3rv4Kfzdmq5eRgj/VUw5ao/fbekzuGBMaDZacVRULUbLzUrpTl0d3csfuE4
44+bXms9JU0RLohy2oQ451nEP22xtVEvxz5QAoDB7SzzgGuweFmqkaIVox7QW6BvHzLMEGOpdboK
82tCMFeFG6F037jT/uVY1TE4U6NvndDcO4pOXtgToKhZOsG7/IygZNIMwqWBFn0KBnuZdypqRUJk
UtkU+N0c49beHfverAb2cVeumw2otuvsVTM90TqwcsgWt9Mm8VGX0U4ATcqgVyLEg7cShi8COryR
55pa7St9h5edItKzBGSJW4DZy0bPUU36izaTKCPKUjcIeM7lPRNlW3XBddmEMaDVOlPCjb7BmX3O
FxqyeOQDmOwLw5h73+TE//7dwHqcIToyMh06RiAbz1RtbbMELinfGpjWxml3ebyf0WjJg4CobvmD
BXWgTXqsR+H9NkwowkX3z3CnxeQHlpvttAqL23WmYZQeAzrFhzKalWxkOauichuiv6DBhZK7yc2L
0PqN4cMKlaQUgiEBYrG2ZxTe4MUXCBYK1wDiDa/Joz+/uWCwxRMQM4HQigjO1LOQUh99HXtZWHeU
p6aDDC4QUFtZNzA6uo2I2dYi/bDM9MpzM/2cE2vNhY9dhEanIxMeRUyPpYDpjaFkHj8G84sXDEKr
jSoWJiE5ZsvQkRcYu8DxUdWeotrcwcEYohTaKM9/H+N2n8haR91iDyNc33REZkUVTx3qqidSex26
Z9fOzlom9CMgOaTKKybjWROoQG8fbf80VeH7WAIgU5Hn2Xad1eUVBQ/22DJiZrhFY4Y5UHdachHy
4CCdR7JCmOXDujowCnV7s3iStWPWvwdQhpBdpwroQReV7GFv17uJnxX25vIG98hbSywaOlipMgC9
pc4J8PblXfOSxx22xlu25f48RJK6rciSpwEdER37LgqqMCW6mVecUWm/jd2Ps0ehzcBgu3Z7FkpK
RCKOv/Fda3hFH4b65icQQlEEoM7wjG9as0RwrV0L63f5sAPzj1Hx+VYDWkK+8Xjm+0CGflCTGhrc
BMcnHSF2jwTb77pQANX7su7vDSO5fwPNBBL/kfiIhLMmsic0igPejvpgPTbSBInQu5v39Npte1H3
VA7C4ptCxSWnQH7xqkRAcMFx3TvCzl+Wytj7FS7utNyfqhfGhGqHrstSDYkCLAp3lRxN/V/YxhyB
+96syGRo5kPtDdK4hqFkippbP3n0ckbzkYzxcFR9K1lp4EjeYjQwo8Ws2humqE0gohPQURIfZnxi
Al8XFAXW2UDYUphEhWzh/5GBDzr/Do7aZA1z8hRMByz+0UGJRSLXQlncyqLMa4rGRehFirFFRo16
nnRWMw7ufiHnYQfO2y3HWpCNjgXi9eyur6GG9LKUyIgVipyuoFikSolg9OJE28qN7XiNl0Idkb5/
aOvmGnG5hBofUKjMx9TWL4A/Fcqrpj2zLmh5G6w0hjMJT5d3nsh1mJAMTDYwoacJ73fY+HHBNRnQ
LN0iJnL/O8LUQpKc+MABtJ9QIOmHyUUwahdU8MptJ02BqzfRfMq7syGtPo54c0t82dF2Q/0bFcJS
7/fin3Il4BAqiU5h8qIR0PEwvr5PjfBE2rfBUjD2xCouvMVWgYKS1rMef0hiwBSrKhM0Z3Lrygwq
apNUsT5YDaUiyf3CVkR7roN6WFL6C+8L4n6/Il01ULMiek9yGlIz+wixNMpY/4tZJApWSe+dEcQv
+l6pysTK5VhuIgkwchiTvHlZxVr6QAmzYjByDAQeTuK1CbtmxIKeC6INneJ/E6eseq2TjA1l+NRj
Wzj0xfxdJOPkUO9g3Ndm3d0VrxVaVIOToXTUHvGibdxCLQHmdP6cB2wXDnln43xAQaHd+KmE/nny
EokwM6KrOIYdye3YCkLZr9Su5k4Vg4eVBZlgGR6vMNFGlvXuJisw/G2qF1XdeuiFQ5Fwx2P/A/qC
ssl0GixM8Ixa5LQGMtzXz4R6a4T35xoUWxT/EP/DrnZYh9tfmODK06Rs67hjUW5jLHK6zU06kcz6
BLxPunTxbm6qwsHwGcvp+DusATzB8XYTX2a+GUp/7MsICFaQaUupOxaw6n6yNWVw6zfFUxPhYIyu
3lknnH221a5VYfetzKM2Hq2u950OMCiNtGXCIgreHBQsCsys1SoEYY0rYBiEJfi1poZV8iaSKtRs
VHJuq566oXnCfA1vEUsFDC0NnCkyAIW/uB2XzllqDWqg2nD3OqxdjJcnycZy/7vl7syhlOqOYP7R
I8UTtQyYB5EzXPqFxlWXtIKsf+SYN15YZ+xnCl1lw+76IJ8mH56kjmqH/2xFJZV9TjJfEFSO2C18
hzCNCqETu/Fm9QriYCjux92WkF1geGaoEKpCu8eIRi/SK/EzrhudggQMC/MHovVk7Rfx5YhRm6T2
QQEAsNRUKRXrFrFJogyAJ1HAc9xKNjZg7DPjpG5/tgJJxZmg2oGIWpm7nEt5VcIToag7745NWjZ8
x6VaGNwgazy4oY/pxCciYbm+yjW07Rl24JDEVasCXDGMeVNR7O4md9gG3O6affmF3GqP8Cfp4OXc
HJfjN3sRz66csHd0dOr/agzWmRmrNRL+jETtow4EMYCZqLXkfjkbKe30gTwFMmyYwgtEtvfH/1w9
yMqs8/h2ye0TvP+yf9HKgVxgRc6PlxNOG+wDVnTEyaIirvjry+qgLBvTvh/7idgCFfuRKeXaVxo4
PekxQw2/o581AEJUH7yG3o392/aeV/z42jyiY8Ob3av1VeQ/wtTJaJHpytA+MAyk3ZEx3ozKUhtH
NhQC05L/ws/r4SQCJ86n5tB/kHDHr14k8qIOJAdfPURKPtLxkMECG9iVMB7GU6Uyqru4gapL1fZT
ldz04YATaRql89CxBYbgstIcO59S1FzkjF7+65qNe0/mNdfwuiLZpAU0XNLfjcKyEUmAi3lVS8N1
UrMgtIIkzYwIcvj8iFcslWzYHTBEEMxpgxgDxAsHBBf19ZOikd+mlU69QAR9P8A0bcP6bTrMHbyF
KEySq9W3366DRlwvLj9CyBbALYw92iLBs9E/4OOejvLPI5Zr/SIqmmLOlDmqIfEMDVISH2kSmwq1
acW7QOBKTev4NHcZVXkUm8EgrlLF+4JkCgAPQl2vn6+qy6VdIM6QNf91XgmNPjAdozBnr61KDqsu
Y3G79bA3oRQrtuVTxTojpJrNSTVqGCN51R2B3t8i0s8anhXbWxVc2K28LeWtViM9TWCQD1ziJvs8
MX/Uz5U7Mjbprsi5BEBcZQv3ArVmuXcjFjeiR3+Fo8QbOd4BEVtcngCqCELya5UCFV7fh5SgN7vI
tpknVELBlhwrS9sLo5P6NsUJiYImutktI5ylhlB47QpGy9qYkMq63IEf+F1CMcCbqYRgGq0PkXoT
b0ibX7PzS1cIJ1huI+cMkX4WUmI8uI77cViNkT7lJ0SRRNnX3xnPsdM7H8T411oc3/5o/q5NbEXe
+/BaNC4Y4LVKLFwFuLes8bCalxrqPk2AU8daVp7nWp1lCY5V8xQZk9+vMmLqcHEEb8F12ctidUcV
QTFT3DxnrjvPn3F0RItfvvWLWdBpMMoo3QU1B313t/TBxnRZBTZTwFZDPYFokaq4ecU9WbkvHUj3
Mi/Dk7LUAOUwUSU8yo2edOl3a0bpaeraJnIGIhkAY6ty9uEquWBqYFWL4uUHOem+WHMd2GoQqlEu
UyEuMWa8sXABCrdiNO/9D5yFlbcCNi/ft5wEJpe1uGWMgGkD6ninUf7l6zMV+GSEgcTIMf4XFLWQ
K52SXz2jRHYIDax52ep5JDwxFIrrwWXaXSVEi3YAkyMp54aq/SQlmaZE7HdKRF1fGWgJgwffIMBm
ZEQ7IwKQD+OFvygqKQqbNT1FOiu4elVGdV3I84z9yA+SB2eEDQwoizhrIYUFNdZ9msskLWwbvr65
9+8ohhD6Siea3cXJ7W1qYbJoMQ8nhQuGAtZ/28RMzalb9OfGSWbeflORVbRKJmGJ5FdsdYwc03cC
llwf5Ej3AZWil2p2mN+cWTgqM9Yo16ubrYkk/Shg/H3Fjjc9tu831kfSgH5rKKCYIadPLPXUfunI
uktabmK2VRestNXP8d1nlHBaxUUb+TvPaVUCmxM/j0JMuiO229GPkI1GAZOMakv9SNmt5tFHdn+r
x2m/bl/dPCZmOJSg8MLXBnwlPf1e/a9AK1mt8a4ydeSOt1EJiBMgTjHRiHAysvi0BXxxMhLTnEGa
Na/cdzQ8gZPPn+N/CmwUi89dKzKTK7kuBrGwxhUvLMFZH874nV7V9b2cFC9a9Cm+G7kMtL5FlOF2
jAhIZVWFI2NEB5ndWQRPZHl8r8gJ30xTX8IpUz7jvWN8JQzviFqkqy25FjTOUnrZeLCTOEBBRnXE
hxRXt20UgR0gK/7SPmdoYuulALd6GUpCTkOcz2BCxRd2bPhlP/i7DNmAYy6uEiaIeuR5BkKru95h
IjCfLCIxF8M8uQpKNrv/1dX5MLC273dFeIYl+RL9BKQ9pgA9ZBxDslKeyzyeKD+7jPIDqRTF1lDd
bI9j5zkqTGRm07U26t3MHrtr6o9LoW49t8b/IBqVqUu35yL5tpj8JbyB4Z27cmcKq4ecTwS6T4sa
o2Tb0WLz9LrDMlYew8C5LPWTb4eWMQoOwOmZQja/VdFAogTcTS0EP2cd05cW2svdhIhwKD0rBRqf
ZI90iARng59lzDlbc2OBpAHa6zKS94IdFDcrl+EJ8KAArVeP/TQjrRc7vOVj1qfEV4rw66Aiuorz
UY033QmQPqMlsd2D3cl588VCniEHWy/F62fwgOxT753/x/TGnEGsy5/88S5qvRV9waUzgJk7ajvf
FxrzvgojLruGbjY7W7V+s4uQtgU6auBCFq275erf1ECa/MXblNBScWdtuEnAaNjJP9Z4Pymw8BV6
aCPrMAlRa7BqFH+1aYxHTqKof56z/L6fSwBFiQBF5WqjV8u1z0MoVmNc3xDVq42w83clIof6QU8N
ihVhLwTAtuwOWlhYODrbXPDxHh0nVF/mPW9/JezDypC2lO0amfCWAxHXrhW/jSQ7dcQYr2sSZn92
ox6gLZiUbHgD6jdinJ3LmJ7KbXkmlk16ziFmj+cp2BoT5BmZpzW9nLTh4Etr2kIDmAIUbQACwR89
zfHsFQRydB/c5657f+FK93ldqZeOIzNMHN4Qu1/aRq1069/zf+iv/Ck/g3+VLtWUsvPSBsdoygMA
+5QYv4aCBRTqZ6TBHbOYyit1vQjWO9b+Sq6KuQUO138PjXvpZbm9pY5virKc3yGaU5leRN7XzGCK
yHS4NROtfTakSMuJkJusZzKHQKJd5V4lvxq8JdSLlox0ezBBcgXoZbIbk57vVpa3Gb2czLUwqmbl
POlv9Ak/u3cUJKOhZ/xLSbEHp0L7xca9WAa1jE2p0ze7vJsXZ/6CRlQhH1//FRevigC9R1y5fCdH
No50xTlzmFm3PketHLyRQ+j5h5QasiqbOwwHScxgrF+bNBf105ETBIkSh8+ifTVX0Wsa0gFRp0sy
/fbV5mRntmqEX0zlY5FkcGPURDcPJB6bXLCI2lkIHmXQNkKzQlDgIR9gt1fGw5dQ5gfCsMedVce7
651l54fL31gEJIdZmebtR7+JzOVFOWSTMAg/wzz3Ho9MESlu0q0ptYM3ArsBqRIf0i6074DVhAL4
lCzwXE24Hopl0zVD2aHIRpwzYYFmwoGVh8eH8BVH4HtQo7CHr/YLtwt9/XjfAzepo63YVKnxidIE
yDTKb8ieqMdq/cFrIpv20Myub73tNdUDI5V+G4XyEHYdrpW8biHp/NGjTKFT7+53IOin0y+NfdD+
/2DdyrhcrU4iejjlYt15wzPzcGLK1QnxKxhHorjFFhhTWNjHW4V2seZ8VE30AkZbRQrBd3qWGaI+
66I3nDbB7acvEow/JXFPkrMeSpY0O0snk5ABEytdc3qdEzRk4vPEiHhWWVn//yUJuHcy+esvA76b
z9ISVhXMLIBe92PdQ11BIwFNG9acvaW8pDkSaVbpMfTaBrcdZyaiwxI3w/Z5jZJB103N3VG/blxt
HQnIw2QGkfjgfcVWrD9Jui04qkTRiMc+OvHBtmZL9d+J+dRFpTSIdX71//tFUrcsn7T2KUIY3J5u
krxb0N1i986rTGCA3/kI0m++k9I6IDeNK2OhUGoEyBUWnuxowi7bjwfUQ/0ylLLcCpNnemrUM/bO
4SG8+4QSOvOf1495StYnm+IRa0u6bL/ZVBOrC2PD9uKoXK3pKQTGPItjOrfkU6RUPX46Wd2AIkl6
pvp5oh4ZPRYticNF/YKKYKxGcESVG5A3TKzbKZbmOFFjppBfJH2L9dj+gXI6O8ZY7qni4mDllBR+
dueMS4tHJOjkOsiJUUIvVI48OQT5ilNn2pDDmrTmdujPKtZ9aMNl75cggGUy8+QYgC7x92NdoooD
3IrWVQx3NfRvb4M9rvSJLHjIPM22RT1TYLimjL2lH+cu3m2oG8SUREJ3zCEk4udEKADY04v3d9Va
Mu6jqQ6ldLg+zuxHVKytz/n9F0BhTTGSVboIGsESHuKH+yY+5mMi1XwFsjLsby0edSkC1DFJNVWx
buPOHCuo1J/g7YTmih+oHc6t5SMQzmGRg//nNTW47yTvMnQ6BoMP3Zh0XawBa4Rvdci+MJqWYILa
mDjhjDynALygyabsBBvaRx4aoiZyDASp4cRYxoKJFtGqjvNcj+Q19/AORBVASSoO3njQW5l62uep
HoUPJtbofDSmZ3fd+3z1TjnDvqubAIYvJ40RqeXCL8eSoMrX3RfWZkk+7znLN3ELty58XDNHuLhx
MWlsljHml1jCD2XGyr5J5bHFnA4qp626u5egGhfYEqVuwMBhwl8Y1x4iauMnLxJtU1UdogleF63p
/lXy1kKKowzFZ2eS8r6S1yc5ijHugFBAZf5ePJDvUKyjKzEuEnK1FkLpfhgis2r/IKCsmBz2bScf
/bjAgh11oEpQVBowO91wzdCgXEa3iUpcmtGxQhFOq46DD3oDnNeY/jrj7+j93RM0CUJbAe4uSyIH
ytixkg5FNjRo9Oh5Tl6zJPhbkZ2ivVnHvXEAMDSoENb+gnunsrXmntRxNFTaML0SKFmv4bIRJnkT
EsH1A5aOVwOmKb4rdBtiPijf93bWjTOwrLDqRfxl6HxofS7qIqBEAhwSLQW6Whu77U7bsE1LC56z
n3oMO5IPtCAriWHaWHOBFzvxXebpk0zTwRqvZQ0jEbfoFhh/r3/zpW3d73S1Fs0eZyIpfnCnhx+c
rqUKnk3YSZ+XncOO3vuE9CiH1MQmwJ/JannFbFk5C6miSHpJ0gVG+TTo6HbHy4657417ElLp8mvV
yiVhyUo9sZlb+PCB/F04fy20+EPLqWAMRGVgVtqMpgCnC7Oa0GyIVtDPT0Vf9Wp2qriKiRE9JBmN
Dj/9J26ES+AvGhmSQQk5kfW5CRU4yW58SurMhnyGWlhrRNYA7W2ouAJl5jjHD9JDy0FYKIUI4S32
GFOVC4Yam2ruu4YRVoKhgvrrOPIs+mOAgcTPXOf7zT8aUt1mVcgJpoGbo0+eu5tCYNa82CJwCkGD
DROm+To9GsEbqpMO2w6yUfic6C1yYUfLW/jSKSOqW6jxou5gaLq5upgyPp/hppb1508zFtmNpBs+
6mWZcxLZ3hsyA9dfJUFTRHtnggMPRVuQeAT6m44UrgsbZvWUYGqlz9SIq0IOHqq4IRKxoUdMq9ua
Ne5st82SOoZCEfWUDrkBq4fVQc2jhjIntk5fv9b6GxoCupfMI6qS9hO7dkEjnfty5onexvtl6SIf
PMyvo2nXl00PRxTG1gKiDcFgcp8fNlu3HWOiYZcxVX0ddpxA+XYNmih1TjcxBHjGo/3ZoHuMtONX
sxbrzeLcFEEE5ZoLHECD0fYUUnicSwD5sceqwgJ3AhlqCUQvrEP6cQ31DvMeMJCX502qnAeVcZD+
tN0Rm/7XPRBCGg2nEi/BP/XP8T1vT3yt3gLIcusswwBbg3ysBscpAHg67hpGeXxhWbVQbtL0yBCe
p3qefsNaOWjFOErZzPqFYzZsfHNnosRYTcylzMFX/G5QWYldNqtg7NFWoHd3qk4gVqefcOfFRi4Z
gV9lUyBfmbR68BxbbMWhizRyWdLm7mq91zqIHIr0o89grR6F2pgRlm0F76IZRxc8bITKho0I19T6
4CWY6bsRzCa6fUumGGTyKCfY5d4vP4qBg6A3nkdWoEVqY7N9QnlWecXJ2ake8+UiNe406Y5D3ElU
RKbLpCRzIIaIaa0cvcdcEsEVcs87dVcbd7QW9yVL/NIiJIHX3m99cLnSZbFakRfWcYKbaFGmO+S/
B41Y9nVgap2BULt6gqltQ4ZJhvuZHGgzPZIlY6neM201ynHpGqc4lsfgHaXaunmDEq1BVaTuq+4Y
o2edV5XL9TrI3PD/tFZUBqU7e5K6pJFKNK8F0Sj3HkU62MF8Z1jJdEm54SJOjbuw6HObTKxXebVh
qokc9LjKWkgaSjcwXqCTDnGleJ/YU+0uPkwn+nzMSVkSpHjQdXl6rPwCnlTyPDURqPhJAlKz2n4A
9SOXulWwfSOSCiN59N95Al0EWggCnZAZwUVmvMmYH4NsNLysKo2mfdzhYVCIJGcDg6tikQ1aRB5k
/rqhEz21e+3GdE85YGEcD7evS6tQZwoU5Iw/qSm00kxbvZSb4K4yrY1/UxKX9xcfTPrdLtAtT5FN
mQm4QOGBTlnc3CDOglMAg7hKomvC0vNL5fOQB4vNksmtieSSjPJEBOzxtJTsk8G5UIlgTj3thnXz
yoI/BrRdq2DRR0GwsxqQBlJ84zdmBCUx5c+sIFd8bCeVXPXLif79rXO09QY4P8gQTZx/KD0hhsog
Omx5vBrmSbLhGvfQy61Chk1IDmAWSDaAn02xiQCVfJWyODL9c6ood1MnFks+mSb+16Ax6HlrCkL8
PFWohRSmJzeURvDnS8YgEAC6yK4fscVwwO0i6g2GYdJE6MJALj5zElo+tKfGoLHltu2k9LV6S4EJ
VgaRoccP6pZRuu4noxlR8Uh6vrfkzAxvHhSw/2fJArJr/hFQmCjvH6uuV0RL9UF/K9ZD1JWdlIAe
oIRDXicuCpMGZ/j/YIJV+Cw9XTrBjprM9uk6talgTGyRw7X4NcuxfaVvoKZL2OgrIK3YD0TdHErX
3Vt3ppQaPAUGEmun0tCwGqGb3FAFQIb1+W043/7xOWBFWnamcPYQGtqbcek1h8Lo7RxSuoNfrOkF
ypCKrbXupCvVsoncMwWN6LPdVJ14s+39Smml0JDSQ8sj4OgE6D1RfxUnywunUxyfBzD9DN0TPQNx
E9PHHn22Xx9U8Im3zOpZ+VmXM2nT08GX6grSSTUSIv3hQVPbTK5Cb8WX06DoYD+SxP7XSCymtBLn
RpFkXlAgz4sEtxFoh+W+o5UIu6SK0cl075KXh1qKEBFnskcC4W+m74IT1O6cU99m2Is6SFeEF3Ta
KvDR51yNs3KoTFmY3qDcYa4DtGS6LPo0l36OAMvNATzXAekVPLageEQPcCVwFp2Me4A4KkdguVEU
QLS7RyNfM+QSgYcbcYsBfXNtsiX2FmXs9BkoIVFBDC2OnSDg45DkaUHdwRveIjwiSBvE4ENFamnM
YmVGkFe3HK8pWJoTeVOp1x/RJpdedUgakchZff7WG0TIZ/RkKqDr2nUYXcAFokhn5ilnbx1R9pcq
deWJCTrYTXxeC9MRkYNmW9sDpqL/A7Uo2h0WsS9SHWf2jTW3zn6i/xTi8cjHlYlX0F2zFosFyRJu
07Vp3Vj//SpYP88YK9ZaKmRXOuVZYaZdhrSyP/QR0a6y2AL32HmoNCtTdo5h7wTrM71jW5hEEvFy
kVabe0Om0sqg8OO+7JZl8JX1KyxKyS4e+Y4bEa8MnzM6+sTlVA4WCvdl3zZbXpHZLTTVcLyVRDEB
FLmV8kbff3CURtGAOWbPzl7IAJZCoYPDnMIrtMgFNsVyTeQNf4uhlqgt+0LEB6I8uIWDfHaJkzw+
fqteVV3OK5Wl7LMhQ2L5W9yfU0odYez6JifEtR8vBZ+4Usr9EayR/MQNm86bHZpSqlazBUjTGRlX
i8/bzD/o1gMqEsX15EMpWcd6wzLa2O3RoadXA8l5JCY7IN24sw9Hoh5qtA32EEVkmGwATITHEshw
yLpSHAlM9pV8pwSQkuphqQ5XwD4YY2rkk41xexV8El4eoN1Xo4+4Sld9XVHeW1XDhMi8yPvJh+PC
FlZ/qS74RbZXXhUc1ZRJevH9QTptIgc88UdbJYEzv+bzpQf1xL6Tno4pkqt2dRxpng+dadEyPfMG
EykvLCDbDjMSC5BhPJ+Kp6vYaRtlRM+hxkRV1kwacRYZJAByp4B1VFE9cR4/zWKJFJ13hxDwrXFm
pc/L1Dejv6TYwkI3BWmNxzAJX8rxJ11SvOjxXhZ/NAJjzqboTfJ6EEAqSKvd4/nxROSnnPhaLlP/
5DINmWkecI+UbAl9T1ZsV65u1xVPDgmHcl0hfqXsy3559bbqi+yweFanN3Sxn6GSnUvFYGxUOsCv
eRaMuffOVRaojxKf6s0/Lf+qsUnsgYwxFxEBs7Iu3OrrzFnQKVleahYKtBIP3Jv7E8QL2F2XYhW1
6XF+JQ2LLkl9CsEQ7oCeBbIheewYikZWvQs7Jgy3F5X5LwehossB/p22rdTmV831pQmDCOXgZXeO
LR3wHDWRlsoZUqaN1QZxCB9nkYpzibmV/orU5IE091u5hs1cmF9btrt3kBMZUx8VE992HXOXeupG
CzMWZ1QQQgc9R2FfDdfZ2DJbNcgZwxK3y56ygOzjoOLTmvQvBmcUGCHUdIF1QxgyVcI0YfLb3nBX
XcrvE+x3/N93TUITdugxIDzUtQl2oNFX19x4yuHYlXZaJWHbh65tu0klEMGc9oMzUg4maN5nTLOy
rNoAHMoYg+vYz3Ckl7V23X0WcB7QNr/MXqnFJJgGYwUZdjz3YO7riVxdZj08DEDkdKI0poH0vDkx
t0mC991DG8CxVFFNoTkocSrhnmuBUiu1SBLqDQgyG12BHCQmCB11j9Gsv/ClSdjS5aa/WMfkwXE5
b8fu9c6VjiaRJXlLgLFxN9oGUf9zgocvgiZvJV0uB7XpV9b5LdiaCTxNC+48ms8Rtbzm3abhCgBJ
94352kYSSqOe2Upt+790WCDF8qquJiCxiCV3cWiEvMAEBMqhMQJl1EZt6eSVmxylt+MxwPzA9Dpl
OYG8MGDfh/GIIqe2x9Kwce/JM4hETzqDmTxhrY/PoXhN5LHuuQQM5nvzjKdwONsc35DZql1V2W+a
qsfJY5a0lieHIovfrC5rnq+pNNOpITnMUtj8w0X0Bt+ji6AXOWS3ITWcITaI+pw9ig10jhFAZOPG
dsohUQy3587W5c/JHtHhWKsE2n77pEFacG0ppyghP6VVYGVKaUD653iP94C9fCF8w41xodKSQxra
QBnWmqvmtFbGHT4luNwTYk5ns7dIXojyvkhZFOf6M5CznfVNKJilRQT5rIXuRuAc6T75Tpj1s99s
Pk4kquMqLw7SHZn6yzxaxmwMkmU65v/Zo4pQoICTs88U/eRGkAZXSLiD/dLFd3riLQGnElsBa97J
mIgKn9EveBdO+8S4zx9i15AXLt0gydE0u4UQ5iupm2F1VdcCEjqKl9Tt2gvA+Iv9RWWMCg4NNteM
qDSiCIMVY5rC6viszVeesXagVuMna5LQ7TVzJf7NMyrvn8SagvqXjWIt6wVQev3E1KdJuC7XVvlI
F9tfftuIsVsmE7yL/LKSfehW3G6RjmiPSWSkEP+T4JkQ5PwVExuqvt4uIN06wJY6pmlZ+IIyAUiK
M8xVQaZtmhtK1YGfrOEijwzpeZlE5t9pj45PGRmkKsAkXO3QkunxJJRF86rFjYdrP+2MB3CnY8IQ
kH0HyGprBFD8FfqBn+1Dua+mIPzsHIHttCcDGJ+Ecg8B4aHNn//W9ar9HVcMqSM6x5XlQ9UYpBDc
R7cFnmq+CVGOT/u4H39PPiZAsY0GiICTh1f7uawEFGLF80UpMx3LCzaCpe3rycKRkpfvkZSJmTpO
SjY/d1lJ7jtE/+osNbXXpEBSmrWz0T6ZmZdeMnMQVF9d4ZcJJGw2xHf3A51Q04Zc1A5ZCIpZoLZf
yy2Mgam6kLi9GZup/11r1AEm9m5dbNlhTTc+z2ZdUow8RaO09p1QX/BuxlL+5WlfW4Pw19GKAtw3
xEIDVYbz9jIVJZ/GfgacyMedjn4qmeZST5pcMu9Hq1wdmcnsj8LFlbVB2dYCRHE2Ji7fkDRz10/v
HrBTjTWDogoUc6cpR9u3d2IN7dcQxsI+UkuIg4jb7f8T+FjTG41JCqeo4M6Tv1xQa8t4eND9MSvC
i3WSed3RjOSvIqATRF59WGkZAeLcRs3ryU+pCQpkRIWK9ZcIJF3ZWUEX2oToD8GTI4OMvrLTQvCQ
saODrijtIPde6XSBrwf8Id0YYhFbXM8NdpjZkQYRjrB1yqoJkUOifVWq5sr6LKwJfzEmvkx/55RT
5oI+vicQlBVmCxdMVxu1V5B6jDzu/rVXHRKK8XyTREne1vBrCvWOc1wBGN9Q3rIYR8DSUCpNs7xP
VsDtBhyscS0SUQAgixoUYq7ucrVWUhkc/gSxh99Lrqdl018rQVjd+G20BOFp6wP8TXr6nnisHZSV
GAbUb8PHxQdQaHGbQTlQmEod5Oub/SewLrKii10PtSXA06z3qpM5cc324r3e2rlnIMZrEPjB/Wg8
iR86dRPlICyJZ07fNXsyrPgGWm9OiToBBSADesNl5X+Cxza2ZRtwlBYv4zfUvymYMubX1nECdUpS
ZLgfc03tJX07cIir+HAJVJSKYR3c08ate11Tb3ioOeZGqF7u+lrH5570Wuwh8RLwnhhyta1WlxPr
NI5av5Ui98tuvJQhme2lii5sCGWxKBiH59eS/eyZkR0XUFqB/AmtmqzLwgj0Ir3La3MLMIsEO4C9
q/YMCJ961MVy30X5C7Mh1ukqLLmb2QDd8YasHkZffLcsrupWsFufkHuAUmeZf42nEimAnBgrjWgV
FGY4ugIvLx15b0R6GAT0gAvDNd20+jxsqwz3ggVLKUiL14mK/zU1uwdjQZwWOXl+smABZ9d1sU5h
hU8siH6bajAE7Yx5ybeaoKuK7osOJ3FKSPysb282E3oTZh3wRa9M4s0aEZlVgumEPZUd4bzXNLDg
GgHHOkAkzehWbZPYaqmTIMt+Sya7N4GKxHT9xbKeXkdxhFALDiw52QXV8u1AtegwvLFn6XI1E344
s5vIF6luFDVxU80YsbLmKNQQF06YDQwgC7XGRfu0ODJbT+PNOpOh/jIsQ+p5DT3XtQcILZAdX5UQ
+Z2pHHiyuniQVDqISFWRvQprunmbIoOpZ/7RBBD3tnrzAe7P5NFrW1JV012HIfKwG51Uvnc0aquR
03OzqIJkH89B4Cwjyhype221NQSLl6g+dL2DxztrSRZHaJ5kjvGIxjGERF/ETp5fS8YfOawOkV3w
d3UEARuu0eZSfn8QHVAx0gwUW4tKR1OY+Fx4IYx0fY/cP7W0+hOy1xOFJx/USDi1GJz9Vgl1/BwV
X3gRZmAwYG2KEMR1PsqQwjjjwgbCc62IMXqaYnUv7LynIaATlZtpNTngpw8T5YwdaHB0x8WweePp
Z2SV56L+B7BTzT50h1h006MQ8RO0CqfcQqqurvacXWceS7sqanxaUoWrKU6FVdheDl7jFDKfTRfC
1kC0+C+uA1EeAfOLbpLXOLAdQwreosUdJZr1GWfReo99TD1USaGg+spDY9O38IKMUzeqH34JDJFD
lVCtJmNV+Vua5NXg3d6MPI9yr+BZ9ydBRqc9gix6G+AbqVn8GAUNURPcuQk5T0NzQCOktEiEAHvC
zxC0YpE0fAZt2h+NoGeiJp12YLCGMy8OIvzifrKu777GK4Lgz0NrSXJQ/mdU0wMksyjhqcS13gMh
eMd6CixnKpuXozLBR4LI7gds164HPeeQJxKyTye3KaLzXvU0KNWx6j48K7GBp/qN9oDd1vZajZVR
ymQlbwn9r25GvAkfzO/s37TOhv3mCOAZLfrhqxCObVRlHH+Uljwu5LrrAiP+KbEUavofdGL9brp1
AjD9hDMxBOCvhokMawC3G8rUx7zwZnv041SB0q7Cvn7t7KrNVp08Vj6Px/8LIrMDWI00tbbssgxd
e5yfI1m6O+G17M3THNA2KT/VJZLGPz2yRjsIyB5jadltORw5n+1tgovhkcbKMcIKUTe5yeKmfoxy
QUSs6VAsUXk5dhJBR/2UeE+Pf7jNzMQwbnZWdgD5jBIUXhJ+XTIv27dDSCBh7LRMsDFTTQ6SiFLl
WD14hWXsXgMQPh5p+2eutvkUvXpJtlxwma5gKO78V5tls/w7SCprJlm9e9fagiH6OSGlMwgmGBNh
aJeOmpQIfTGnyuir5U2YNdXrZRQ2saHbvNcYmsOv96qXs01trzfNPwwx0VKD7NM0etzkKJCuxSr8
hH0KxeqLyY+DtI2wPX57zrYLSj7FWThLHrfr4XRSBS6QhNgN6tmDVHLmJwFikBeaPVEO6H86s8P0
Wxq8y3pa08EoAaHM1L7I3MfxX86PUE2lrTC54t/iCPAqI88/CVG50jxTW1vJRxM1luxJLlungqzv
gkXjinro6DPCiXFeuuNlsZUjTe17wOb/QPCdl39Zi1eAlvvYeDDUclsfQSn70Q+onGB9UbuSP/Wf
rl+drdwIf/M/1RFcdPI9p0dvOrfZQElhT0jiV7AsAzm6SVccAjjDlMhLjp1rEyDWrugJRDd04LCt
nOUbHrkfmd1uDlz8FCy1Rdml37PQ754e8pZawmyn3Z6RlSlwdgjSTAw9ySdlFE8DCkpCzDv/r4AP
nzIe1naYW9CX5Yo6jrbnYdSBEyls/6AVFeD6rWXsugLbkbzJ8KLT9F/6qiulrnylsHAATXkeNvYH
W7ovSpHTxMcCzlXhHqxyh9peQKIukOBFb9AIRimhw3l2n5UoRA8cugJIjykZDY5HxqAtMbhBcIxd
d+FjIkMVHaQW7Z/BP3vARMyzjsejjUhHdEBReUPLdHHgjvvxNWaLk9RxpTjBeK3RqfPPXlEglUoW
h7zcC4Q4dqYFBz7Rgix6dGgzzxmb93k3PUAESvxKdXxivVTT17NAvDEvRkDcPeLiD4NnMkdv4XMk
V0BX11kNmQMsW+oregNMZjgYGCE/uXtxkco+GrAftSA2JdZJe93iqSWJDunVzaB+kZRib34XQKl8
VMVi5q6dW7jmEMdkKXo8XyjGiiE27oLlegx+9TfUfnBQJzDh4GovByQBsEwU8Y14ryh0xpXGKgcC
qxrbQUQUm4n7VZ6F7SH2ZIA+Js4xs4uB9UHwjVLhbFjLOnW8Ch6tLZ2TwKDV79VAN1O2uErXaR5b
4Rsi394K21SRP9n+Vh2+EBSJ6YML3o2CG44ckCo+WoxNfl4awtQw13J1KNTKfAwEGvdeXE9/rNuc
MHtGleJOj1bfOest5khLHGMFv2hu48FFQMAAVr4Kzvo2vWFzwRvaA2McAEUXx/XK8J+8Z5M569uH
WhvDglKtYkZVwziz4O/k25WCVnuYQUl02isNGpTxVubjBqu/ZFS+XBB/j1k2iN8VakGewsUKlPou
vuLYfQeuUnYpJRbhGWuxkmgS/X6e7exMvo1aI6N+DHLEoStdkrDRhafyQsWxPQy8T2WiAkrGFKR3
oQ5HJuYbZO5apWijWUX+U9paKs98bx89D+lPOn1TxHYyKb37+IuDREKqeQUaa8j2fjLdIie6PMu7
QJZl3tW3jffet0/0VTGC30kME9zul/QkQCDNcylvpj1NNr3aQU27sgwEf9auGDPRcX8gHx+5TUaY
zPhzcsP+1QG8Jfs90NOZP5XV5Gjdj05Bu3YAeBvHrWghhuN8/T0Iw6dCX2c9REpNBJ7QloWRgTnc
HLSnlhVcQIr6gFSMUfA1j+0uHmdn6hzYzKnUMwsIwUZp+veBWKhBzVtEz2u7COKtBUf1bc+wEAIC
OpMtH8/AxHf2mLT3pSVC6Lg4mw6KvToCDAWlu84NizgC0UwtUxPacZ9X3AofNIftvsx/wUX2oZI4
wIv2WWLT4xPtmzNlOT0BZIicIgPVO2kbhOj7OtNlDjWO1eTY6CKOI9lzg5EFaY+RgQSoeM6hvNgI
UbmruPhg/Ttn9XR5QST6K/AiSgvbA5PuRuEmSYkjNekNpw7N7ISr9s8X5ePHbjNtAmuUb9uPutPW
L508aZEXRsZurxmGbgKXxURPy1XkfTsXirsnma1s5XL/oyAC7WRGCfv82fTmFVmcGwLMr8ZpP+vv
x9n+Mz3W+ANeaiUg8O9VVbW9dndIQRY1u/sdTaXJX59ork72GF0CywzUciJO1Blubwk60Ak2XJn9
A5wr4KV4ilkzXSSy5E5GY9nu7ZV+pUT30yfcb7pwWUxFXgkYQsZJ1uyXq9U0mTxhoYZx4LV2Hosx
frNuvFaBEAlRWSHCcEf4rAleozWTcDh44kqR62OMeoHGPqEmIKwiwmfZbl8ZBxA9a7x2pzEl6rjO
V2ea94yT1UQMBGGKCdjkQU2pNYzzvQPV+F6bcmUrkER/mZth0XBYT8UBE5AxaJ3T3jBlUy5VMHpX
VnPNl83ecc8oPGkMwcHSCZy5AdIkFYiddPJgVjajw7zDiAUmpnTuxdPnXpd0Gte3wa4SqF3PVl9O
/dFMd7yfRbnkj80PSdBxI9W+Vf9JAXQUi/q4ZLmkZBhXMn0PbIP63g+2+9sRdTkDDwh9AdKc3UOv
wyRIcnBXfVDDAWY2530UlU07V+32DA2231Jc+ZqA4RoKpY/jJJ9HUhAao0ZTwH2fkEQoE8DWv+lD
M5X+3lvC4wWAQFtv73nNBWWyWw070oXfJrSO3+p5oCJcCat6Cy8Mxuq3MCWtpKU6JBiX17gYflzn
OPQT1lSX8BJdcbjwV1HyXpSK3IFN3fJoT9wwaVFTgZSvcYqdOcjsU5FRa5wx1sTkj+127OeRirVS
6z4oAEqFGr4zI7xC39eVxFSgbE7iD8f30RJrNzPoSO4LgOwxnc71U4Qgxq7ygyXN8J/xsLQMOmyP
wUuoLIO2Y1TDiryfeXfc756v4ZarFgOlECw4uqczAT/mmpXSuryxd5gxnuKnVlxdqso0By80qMoG
KRHuox6/tnHjXViZ7wS7MdkEUoDbw5RLECJh2Y0PvOhawv45n8ojMEaH2f9HklQmaUPjRvotvXxb
RHDxYoVyzCuml/Ng6814BgvledVh/Ev+OVN9zAyrHOScegIGB4tFjsQI70NYK8ILwYgWlOtmLO9b
CRr7INDAN6Vd7xleDNnx7NR85zpFjKR4iL5jdRpQYHi/NontNRZgKZBqoiDERHtiacKx1rvCIowi
8owkEP1/12OHWWIa5iK02gJJCEwV5hyRNp5jPL/J+f6kuT1AwQNVVAgwXZbDVRDCtYcLDTIbcv1k
uQElRmJVoWgmF68DBhURHw9RaX7SnYG9aHLmsf4FbHDyhESyTFsorxC9VnW5+wSdPSeXkFZK8/jK
XTe0Ilz5X9K+Sm73yRd/xkDYR+IyIhq93Emt3KxyAJP3n6y+b7vWpuUH1svmrIp3XkrY/zLNrqMs
gjGG3vSOkVrtlRdP6WrLb1OUwcuMnVz7ZWdb465F3H2MWlUnYH/duSBLTWsTtsJ352p/lY09ZyJU
hiFPF5OdgPEUmdw7ijhTm2o18mXn94mWLI+TyqcVHaH9gdmTcaqYa9RRWqStD/KGQJK8pjKyxoSw
epy7JE/5TeJUqwmGE5krBCnuSuVTea+q/qGWLOp7rN9PzU8MHck34e9WatRYpDdUKGfLjiZ9d/QX
HdlhSf32DVf55cf4kgu4PvJDnwbLTkHhsuqulsrnvTHgZrzEmi7+v3L5bFW/YIUwk3yQl3Bpmhu8
Y7WFBl+Hnv+eE5Sh6sKqnludloDZGBy+MFLXL6Wycjf3r0dFi5CCSfNd/pC48ENQ7vHEkIDCBUjY
ni4jYdqQoSM4bHZcAbeoXFxROlOmJQvz2Qwuj444cGbNPMd22mpqpU50dLblJ9kcuVKo5lRfWSKe
lnwYspJpTwY4qSnqjjxH+fpyV/8BZJvjzzLHElEQwZBD1xDxQbSA6liF+Gg8WIwizXRuKxDKWrtp
espRIQCICDIm5MF1k6y4oaG7Ue34qj8SsaeSciVKVP5qsGTshIN3urdKofPOSEkHqP3YWGj0LjC0
i0EYZi2alY8T0kaHQ9RzYNX/SbnGzR+MJQ1CFLUPAUdVmSS67N0J0j75RJ2z+xUaGrKkD4C3M3rZ
2bk2Lq1zOjEdHJFmlsWMuUMcdidE3YquXhe7089igifhw0qHN6CeJmD5dm/szWtDJfMZZ1Mjxwj5
TOu1lahkLyJIZELlbr2jUrInTexsh9Qj0MlhtFTdDgBx0M7PYWI8A/xaE0dXuDVDJn8hBw3NtKX9
AhIDI5cQWKmD0hs/wtGPHbmGUON1zAGEvrL6FYr3ogPj8p4123hLJsGRecwZjaEHWoa2ZIdLQWn3
9BTNzsMyBQRbJtQA/kjWS3l5GpkoOtyaAmM3psoC+bnf7LLHKtqPn9mv3+i5TQCOCUvj4BE9l3Rx
1iB48adD7xsJLdCCNdKMQKRka4vEwTawp89XagLq7I6lpa/XzhmMNhZMWDhcmnYWC534yQNV/E8X
9r9tayIBvuRqtPUuG29HIzpFRm7V32qQt//RB2pwoIiXD1XOPp4q+d3s13e1+GWlXsa/DfdeHhKx
/ezIgf2FNoQrWirnf/LGCBlaXrwOi8NWInu9C79bxJOrC+Cbtoue7Qz/6G3PnQdm3Zhz5msr9bLy
J5yeEbJqJGndETzzCE7Fux64VRDAQbWcMZAm9Y9AmGZ12Gz6AoXVTVC0XuT9GrU9QVu6z1w2aLHj
H4F/+nHLMnX7rYKzzzIKUaHd+B2gf3PWYxNmvwATcFz6xBiuLxzXavfAyNaAE3ObbcAGjmckfkib
ZvVPKPTImorvETK8bPnFoXyxx89kaqtDo+0ILdfKgjgAFPwaJDrEqOILhU2HSyMxpL9nHnkDiJKp
CTNBcHNBBF5ihGdQrDpYB2lE/FAFYUDcO7pP/QQBF+FVnVLuIUREFhMdwxWZAStN4kbdXxxnnshi
wrfxFuqErDlcikkKEt75D1j7x+rzjs5IZQ76hK5yfqfRi4JTHM1A1NEcbrA2TrhywyjstZzhAyOt
wkcq9EJnxo6rLsGeAiTqggQA+MT38kQ3QpklPV3Q3cIlR/Lkd9YkaYMs/U9yRphHMuKksukH3yaU
6lqcuOsL+81YdC9T3KSvmj8PRZ7qX973myPT+SQmhQP/pF7ZcVArtqJLcSbmopmLxukDWjz2WS0F
/pvsiAmvFSOti9mtffLxlfWC7r35lGwSf5RZz+MkYfzMLOWcg3WE8RxcwWGHzwtxJntlhT7PVqW5
afvr/YGX2WCH3BI/rdIeJs35JvdgpbtIPS0pM6P1sJxTov2p8YXO1kheO49XqmYDL/9UjRH1M8C6
9/ydAh2O8NKnWSplcfEKPUPlFrk6D1bxPXtnWAUCK5PbrffY71wWYk47+93x5kX8xBM5sYwXYWT8
MHZy+17T6bBNEL3iGjSLtwWJO7+fzzDlUVzKQpTt9rg1RgOGdKolp8XGQe/zuR12KWYk1IETdMa5
YxTluSssQCgmRpxpwwsYSFuJg42FQ2Or0Ry4jY20y33qfmZzWoAPrgXVsKMraalwx+v1gKwEFZRr
BREQZ/4SaKVRj6r0oOXRRgKj4oDS1icDBsrGZJkbYFwXJwokhGldM1f4UHwmKRKCCrmlm0EPUFfe
FJmr/wGIPKkSqYjlDDOpFrMs4IM3DIxPiQWFgfvd1zae1f4H1o+upLC8UKK1fZQ0qodmDWaVLZzZ
60L4LLRM955BCV4FL0QmcRbtJLAvOzsk9HcDlBkuSm22E3/83bORR6sYOkitXSdiCJUXlFp/63sX
urT4Iq46hM1ccKnlSlJixn9zZJ+5GIcYxxRHxNq1qcQ7soORE8EmxCuhE4iv3TnG9p9nPKvZ1BlB
OGnnUwY2HTUhhgoZUVvOvJZIePLwZ5fJxxxuAFbLiBT3vwjdISWB/sSpE4nh87SiEkJ/YGwcS2Eg
DEJq1ZjW+FW2eQVsU7wAwRmFNGpZ3Phr2wh6C5GURbNKBeKr3YG2v11eTkHvo1YL+h/3WZcD2C5k
vWzKfEmRfd1eTx9RomKRa4UE97PdwcnG269rqDnvFyijAp2+xcJk17QzQuS0KlvO7mIFbWaXlj22
gjgaXf5wQ14NxbdVtyZM3BNuNaFReevT0sVAjvYfWAXMSGQLrPI7iWXDZlm/ayYu++wXni0DHqy7
yytCYvl3gC3KLHwnBsYb1GkNi0YPQp+h33+at8B/RrEGiBOEm/Hu0lL+x4PF1Ec8XkAOLk6b6h8Q
ncIEg06CPK4hwmxY8jJbKc7hW29ZrltXdB3kp6c9j2XWXCCE9iu8kgbcWIiprxs9HmqCf/J8Awm8
RmdkbyeVFZv7RAit+j/Zlle5TKjbJNbGTLv75Hdu942hgtTArGbbgokWR7EHI2/hGj0KTpJC6seR
RYLMZXOksAd/Z08kNLBTeqX5eGfo85ajy+cJ4slzPm8r+o6rXhY4olpHvSpBz0O81fArM3EIGNSE
UwCNeLfOHhaWo2pQTbZqwPnu7Jx6Ox4MT8odNKHy7v7N0qVZHr5qnSw4Ogw55EglmRJ0OuT9XYx0
eBnRtYmdGm1EC3ESaiSR+zU8vJu5K61/zhNxPWsqo/pnMr+PWAId3iWfWHv/SXJS6Z9asN2+jtQo
bggEZaHqtQnxdBuPisqEg7N+6GT7Ktr8vHya8nvHXs4+EQDh1Ybr3lJPXHNGN2/cJfl2mE7mP6iu
sHm3ZQcFl+srV441Oyn54bLbeZNjSON8mCxY2K98nbixPHUqYdH0FLaXaEfT2OC/I5LPGeO52Ed5
R0SWV6zLaahuSlFY1v62oR9Z/go1/3kmSUQqtv9zA8aBK8eeBtKg2yoo/FVZ1bUijMm/82qhY+RP
EO2bdiwb9303inme3rBv3WpmAQy5Bzbn2McEBd6qh2dkBLFttSkdaU5GuA9JVbtZvmM/+Ful1RS0
0f7ZMOghug70AQXASK64P0X9lIZWJ6YjCEP4W+FaIs2FaC2YExPBnRe/gv24h4LVJMPvTl+CDOCE
L5w5T091dajE7n9KSVWBqT9ruOwMXZ6zb6+MKECyNQuWso0kTc0VHJg4q2I9FekemyJ8mf9ourdn
folDorqJzxHXUGNEhTUYqbbQE/pMdT9EYYX30LHMtf0+cDXKcE/SkdEICQrQgyUVDF4LpUn4ZJJ6
vV+91idwzGnIC/TepDr7iwnpUmYM+6GBKgMQKbdS/ZK4NqhMi5qsEWK6k9UI0CrlzS5Kskg7wBBM
gOza0MVCWd9GfWtDcfDSxzV8JVd2yGX6ZyMU/kYkU96CF5mM+FBMtHcu5vSMEkBtMtqB19xihwYv
LOrQeIF1ru0JpevAelRYUm3d1R/wZ+Nu/aWJm1xy6iXXLcMSs7FIbANqk3rjm4m3q65XCcLr1lsR
QdrrGL6tzWifbiKWdksrZQm0RaKGGgSgyBE/4YZJa1B4dKgtKvg09UR2tmVh0xxJaL7T+CPOY9qb
j9dr7ig/xmdG/JL+/bdWZVyw2FoGqYi2UCrsMZjXgGZKeVMGx6x7fBu4dy/RTuu8slskQhaMVD6c
hAFGVJ3sEXjL/j1EXei3h2NFfBwW+GNgZ+sHENeeA7CrcYqqqBflhlViukMtbH6vHtHCSxXh2kWU
RuwTDEaJxjCHuPQAGa6WC8qkNGu2uSz7C006Pq2Jic8m8IlVg2iF2ZGVjLmgZX+QYxaKNdRYRxMd
50f54d94KD5foru5G29S7QW3i7PvP+bHoOJm3kyEk2lTbzR2QE9kt6b6lngZDj9kFgBFg3fbiWjJ
Lk4BgclOUa9iOzXmzv8l44R9FzNnZOjz/JgRYRRP4Nr8JcAK0GAbxFzP29LB/9S7vjFSf0p2Aq+6
t957jYxDHWGKXyx63LxkMys9gSgGplp7+HujbJpqCcAYcTjHvA21kI2Vwmp4uv54KPSZJIin9egE
qQ5f/yu9Ls/+/wPHKdCLCNfKnl53ywNjgJ9Eryd8yu4Ngla2SO1CwWh6gPEe10kQiZcmHsZD9+qm
kppO4IS3MkBm4P8r/S3Btn2neD0u3tBSQXSEudqZ4G1WXsW9L+3KIH0C4v/s9BLBs5Vm/j95lrgC
qz3LYLK71cttTnz2Rbk1oqjjdGCzHoleV+vYZmtDUHgQVyF05SKP56klx6h2sehkFgeovCvjVjFm
XA1D5FwjtBfyThziKGKUyXJX1Vnp8K7TxnWgINmZUogX/Pe8IbENAQ1Coeje/6JjRPcg+tIXva7I
YZAeUCV5CrclN/WvaYdMlhu8wz1JB0nezjTopmEsJStbyx+skEy/Y/7ds/20u+C9hS+NFEFOlUdO
/jxlwEnUWLt182KjXEupmXCO8CPW9VCh6yxkhV2Gtzef6PTrsoARoCperMi8s9/VnJsFk81118tS
g5P8AW5pES6UpnspOknu7etmwThhMh1l4c61gVbauoSIRu61JMhpDHxsggGyGaXMwYKxTILyadP4
zUS4M7YULTdhxgefhpG/Aw+ldr+AgKpPI2junVh7eGjPPiHAfG+Sv3BXimoWrYcawiARXDxl2vMT
fLIzTzRqn2FUXIkymtgbFvwu23aiV+5pwY9orSOXH4LHuneUnVxJ6bzMhh4INOgd5fSfV3p2Cyui
zpQRIauwkpR5XzpiTkRmB9YWvl+HodQGWQlAXid07VnbMnMv2sirRcVUIIwhbYq56wdPSrAh5lzR
w4wAJwXbjodZp8Q9bDPkUL8WVk7xOkcs0gQx1FIYdIEJmonqDAvJuUmDuMw+mA6KR3WgDWkPJ7E0
yoxH2SRWrdyoozku9Y9GK0bGP86NwHgtZ/cjRD8JGlsO4Yv65pwjCvoeZk+VUi9r7jjqvt54jRup
Jp5lUwsASo/hoeKKB5WtGI3gdDSEt05fZv9ijuZBfvb7dxWnyy/+82UaxV4gl6z1AJSkkOauURwc
iCVwV5i6dhSUMadx7cO/S+OpR0Q7is2udq0QLz+iq1ozIWbWIxE+QmeJJTKmMRUzpgnZgzfxSINv
IKCYputJTK41iPhKstZtZYSRXgA5VZ1kCH0nqwqdZt7YeVMrGDgD/Ig4Q4v4d5C7AZkEg8NWArNn
XjptB64ZTDh0UPPvnZMrogS9GhR97SU6UiCu3sfGqnV2gR8e6FEjL17VrCuThTsU69PSh/+8Jex1
1sB3VO/UXgDaIi5+PLHLzyo3UavwYqfas36MT5vAwP2yRLjLzM4aWauuliC7nleLqAf79a+ZbS0U
1dTWXIkKQDcYLr6mOgeEN6ig/L49JVrhe6pADqQ/DifF4VNZJKPb4fHfaqu2cF5OZiWumYnsTHod
PFg5QogWdntQ/zkxJDulkx0yYugeNWp6pODYM02fNjrpW6EuXZzV/phmXw4a1f9ozHiIjzpOr1Q1
47UOTsxP55ueRT8UglSf9QdqfngtqhuKFqn0964gj0wWsCzA01dMl17oT7GbE/gVDM6QEhJA5GYx
vrdl3tc2t7yCDlFy5+wo2m25Q7kZp6+Rwc0OkkUTdJPbGtRJIVkrpiZj6m4UIzmdx7yoWwz/Kl20
ZXhi1XDtBq5vH3WyGMX7CbP0liaAeSMwwgoQW5LAo4UAzqdQfczvgoNEhFGExZYZGJ5p12sUgZne
GwycOiopfpuVlK3oYhDMxgJeZ8xEkkxpvPX0iYcq02PAN+6f9NF6J4SY2LCIvc9s9r3wZWLrxc44
BptYqXFu3E86azeWDK7OprcP/lyRrL8aWb1lHE6BsocgLpd+MvQU5jzVQ0kw2I5h8vLrkM00TucO
YS9TdJcUxx1abyfC9xpEaDvrjfFvShUi1+zywTflWoCVVG56zlqN18sMYYCmuxdqGzg8pgk+xFaO
Z+u1MF3kdNTEsVjrVTIe5J/inUhz1blEEXNX6elbLE3Q6EnARbCcTo98t2NI6EY9mUtALJRjFBRD
DIxsMewRIjw64Fo+k0/t/9nEUQbcqXeUaV7xrHVTF9cTzFPWsaTz8P0fcC+DCTaJwXnPr3cs9gmF
Gz820DW+RdRVgQQ06wkX3tC8RYhmfRq7iW+jYI+bY/4WnKMxDGNed9Ll6CALIrE6p1V79OogxE5v
vIk16YUNKElUMIWFyisr7bS4PAstKIcnNDZvzlYcwxU5V3jKw7/hPDnL/qPl6gT1gRSxmCRYUTZ8
ezvSKHehz2Vkw/dojZXN0pxYFn+vox31bu9qnBfCvcrvYyzvW+7rZTNezKIY7r6OdlL+ULqzZH4k
rqDhw/ATe/Nr3HIHfpufTj5CZu3bfFdGGJB7oHK3Updzk9T4k/KTN9n5054y7uVS8NWenqXKyTWN
RotsRXuW83PTayUmKryNhQdlnbeGPTo3abFQGq8R4mcwdjX/T9Vt1SlAv0BQEQjEH4nkpU2m36lT
74FUzROmOycM/lT/VpKpe35cxOhjz2CNyPMW04XDyj42nQRt/hAKcFLHLWqWjY7t6kuexefZOok3
mdB6eNEiR5iHGQZFJURwK2695rFdJ/eobE7EDWOLvkqm8VEDWjWfJvCo44dl0tBUzDR58soblEmH
XiMar2IXCO3L+uoN7RUB5T6Sv5aF3Eim70a+mFrGjEAFp/3aetTN2zdyjgXKil5UDGLz5AU8l03c
mKqOopWiGKUns0lqf0Xb9fFn6D88DjzIAiH2YUtj7wDsNbD2f3jY9Ck0hxoRfkrtunF5mpddlRRx
aX0eUTbznLgnGqv0LHyxNMHB5hXVYCP8DULZYQW1T+CXIUNhxgWAOZ53s8oc1cXXuLB+u8Q52enp
150eypBXuhzVSShPnjHzDMEzxaC2hz9UCukYV+RTdJ8+rzeLivEPUkgn5A+5o7GaHD9gvpdcRacn
yiCsDu3z59nfN5mcWg0w3yYp3Lhtuf3HctOus16Q59IbInTW0atxXOtrFFeI9t1b6RIQJIDWLZ9f
yEQzaX9liVgnacHdYa9sowWqI0gU4tlPe6Ve15SHS/YB7yPHfnblUIYsJAKOR4bLQDKoOUhvezDv
/khss5FwUVyu0G3X1ZRPlbRmpHhYCxFWHCcOGRJm3ZobCuHSl7Slq07Oy7orDi443IeurE3nzLYc
+apS4+ejaCrQ3iUphnb6MUbZHZMhgcmRIVl5N9778q7jjuwmZJFAxnwaRhxuu7HX2LSk2VL/O9uF
07B6T0fYFXj6PVODlyXPmXis6sYOljCia5wPBJcaFMWVoy3PM34aJSGW/2cIAd74CwogzlhSxr8f
9alJpOmtLjDazr90QNQTfCriRdpTS1kFEA/Kwct0QaCc/tpKjigWTsuUlMxk5bL1LMSGb/JMixpN
5lbRSis/OGsZKRsmyxBztH19DZsa97AcJH7gF6x8DhgPULktSC/AcjZlJqQ6VfqlCT2U3xgXGIlf
io/kevxsnyBtaCVDWrP8m/cJq/MG07pGF/159JN/mJNdREdeipnZzV9+fr7drjeho70ye+ecSz0B
VzFtpWOYOfbRBXmaJwxTrKmhpCoS20CjsduLl/V4z+bbi/ArgY2puGDvqCgNU9xcFdWzG4NIRsKv
UcOQeehZ4vL0y6Ta4QGTk1BsirLDFx3ZJntVLKHt+vZXOUrC2jdP4CT6HifxLCT65gIBhYkEKVhn
5u3eDl2c6MgCLbQk7+EquRIKlu8PHgJsezlzc069XK+AaegcSxfGkQzEdHFv+bwDjslEGamgVex4
iXhaSn1ZcEieLqR6CvnsfG6whm8u1SeDoReCYPEXFXw0wK7N+/SX3J2nIwafzQbsDKcf6BjR+1OI
5neaS7ikr8HyguqXqdWVyW/x6tXrQgVoZeXAFQLugRCxHRyT9kH0irDtiPn4fOI3N3uetjQQ8dlG
g3Yu8NmD7twb+Sh+Uc6PeWllRlrR63jJwhAwd7wHxaPHzPZnG0AtBFNfZjwQA4UzxOmiAV4kX48p
iiPHAalAOIFA6cFaVqkscligCPgY8IJG3QZo7mqg8RO0AUwN/pHctSKH/n3DswzWWYKtRxDwhwCo
XzK88qpuVkcgNhD4DuQj95OEfOMsV0o/1ggaik7orMiHbaEgQ1j4RhK+4N9KvpE8HPB4YlDGc1Lo
zkKTr3fwZeUgIZvBv0uLRMFxQ01cOtzH/yaz9MoSLXXQgHoX7aJJyxcm1kGHJzWP3ICcF0VJdkqP
w44DGtaEBTEK0h2DHHUhig8l59s3ktEIyqFWi3l3WaDXwKkdgALbD8hCzFib7d2GkgL87Y/dEn1Z
ybn3C2e/QDe7mJgJHg/ulhi1QeSmgNIhvTynjKt+IjQgGjEIugqoNRVH9K0yU19QUAu9v5opEDMs
i2aKpWOisqP7LFpMUX51I06Y9RDq31mHdyC2K0XR1HmEgqrFNbMTxSoC3lSrmmhSNQo7ikAuChhj
xKJnAhsyLGnNxUOSVMSRFqUL+xBYFKvZA/6XrYH5kBRr+njrwB+UD39XobdTbXk0Dj/0V6HFiPXY
UXJrRY3azCkshWekKzu/+KQUKpVVw98BWrq1iwd2X8raTmAMmWpv9CUPen0Yl5ewFZczx6moYFXw
jhi4UkBRQ4JpqATqKPiARvjg7/l7Z91cQSVFLqhGGnx3OXqgSo5IBfJcDH3hZVwLvHnG47Vay7nc
uqBTGxMguSo3V9gEfBJohDgjzbdZhsnj/4cenxxO1AZ5+FYXsgoVrNlVaHauHR62nxdSduwmEc7W
AnUnCry/DxBcf/W6xFcoANgGUPKA6vaip6S8mcoI4ifTqGWJcIwuobVaXQW2IvyYW9EkX97HYdv9
m+4pEfkvFNPjdBHBqYK13YvpqDzUmLigRcW/zvgUMiOumhAMwp3V3ryHPU66KN9KanZjSxCUf7Y1
A3RP7BLw938WJv1GqztAD8WzeVnBXCI59zv6CFSTbZOwec/ez4eH16KuGmbk2KFwVg2lb+jp7O1z
hJiZ7vHQY3GZE6NcFKRHHK7WDY6ZV0LikK+fb6vDj7209eX5FdsFU85JnS3YKKicTu1ot85LWpeD
iPHbNDRWlPXJWMAKgtd+fdgQ3nCCU8XRunyaNsvynbZEvCrYpYRJLE7XduNQB9J5raWX6yrjKGBb
4WUnp7Ca6sztPORU3bAWqNA6W77LFSjE+7zPf3EPdvDjYOVmuRpVCEwJ4FUbFYZk7AdOwP4mq7PW
puOLUwjD6WlyXrV8gcmvz5ivO9+blE8G3AMcOl3E8PAednlkYFTBhMTq64Evr3iY5F5zB3CvUQGZ
ETCHbZWZLFmyOpsWpE/XI5aykkfyQy2UfjkfF4ynxkaVsmGgrS/15/H3wZbqJvxU2vRjG16p094o
nXZZoPV/8JcISMSWubVeLltl3gveXFsmDgwsiqQLpwa3xWt0FymIj/TC9tZzIz1tiZTi6V4pDqhi
Sd2FNHPqBuas9mKL9X03onKbfVEf00JLVArMEVB8I77v8CICke+wJ/GCbJvZMaZuDBRPjnPoy/+t
Vc+HqXW/nrw0MyAkm0cayvxsnsAgysdHbEa9evK7g7XTIVs77W1W93QyMV/vLk4eK0d5Y53utGf1
U+WBxDADUh6OcniYTEQQ+AZo4ya+5EFeyhnop1cEqEK8lguDIaSxQr7C+g+9eoJyAP5AqTgtcBVS
g5Zna2cWV0QV1w79DNBAtt15uPcQTEmV8weuEfqhtqbFAQq89ImxnzF1bN5IELOfOWlxT/Q/3F+t
sGhP92Z1GLX0Bb8qOVpschcc/EvSf5YWZ9jfl4lrWu2iorBF4+HCX2DPW2P07/EiReJTudwyAqRJ
pOKSpQp3eUbvqgVydvvvQP/vZ7HlJmj9s9wH3u3uOMb/VeZK1aybs8U0/zuXwCICxRCHjjAm4/ZY
S+VazunOaUc+cTzFyjjmNg4s3btNatMWF/T2bxVwoOK9oWRSPa2TvRPqrKLZTzAN/HKmeZW8Gnxs
t3LRpjV1CWkdnCakj1cUGkGyL80aM+94JTMNS9nUTtk45v2m+4yMTCkrCozJ2e52sgVaFUZMuEyL
02NS1jH7n/YcS9ghbUSZ/mDgqYaM79gFMDv/mvB15sgTdJEwQ4W+mYYLn6hFS8VbGFEuockdNOqr
qjC6y8lSz9CRBreXFWFW8nyHURhjHHfgdbKLNIuaYGVMBihM+HwgoylYyulRi2CQw0fOqGl3JiBD
C3NAjD7RhUrt3mJBv/beL3pxhlfpOYed4F/i9YFi59JfrqvsoHc6kitlzKM1QZN6qyE6dgIkOcme
zw/a9IdnRRzF6bExWGDSNFuLB9y7xMQ3YEO4CjcfsG4kT+Z75WaxBLrKZCAlt03btoKzq5qKb0fE
qdVqmokd2C353azR2eLfsNnn4qzmdtL8C4UGFEwqfMap9cI4PUqB3KqQxxPujB/5rw+S7el3MoZ+
BBaN4UEeaqjRPbjtJMIravPNwR561ud6K97NP+iUYSmP460gnkaettkjqaBP07bXI5AAAvJ0WcaM
5sFDWD7wQn0zJFz3ujJuKhuUy4TBpr3I9Z9q2ZgPdu/3auD03053v2DnNT/XlMsbscrNjBC76msb
+8u4COUZNypdY4dQqoHeLFM7+2ydIOXHoh0/RoyxSXeKaUdg1Kecs+e7/tQ3vfOZPWar2SVK6Ika
dtKFB04tylaeHXK88dBj51NY4CDonPtucCJVRDnXGJJf8uuXBFNFuK+7vYz9HoFPrFOudK8Fv6u4
7L+fZYfouJLeOxfQHiIVArvZXnvxabuSmKYh4otjCuHfuVD0nm4MHKJYEsk2Y6e3MduMyc9pbps8
3wHOxWF9gOUPTM+9wsbAkMFS6uFj3uHmFcgFkTGQHlgTiN/YZiHIcANqSMcZ6olhljAXkV40UXSz
m84gniChTgaW8pbtx35YvaCOIZyNrGPh1S7RC/juGhuq9RWvXE2DR1oedMXULpEUWnrDlf5nCfwW
dtyNEC690vhFrrprFrq7trk+5wo+OL/ccDBV5rwkHiaHup9JkMCsPMXL8S6pC0uvVALvH3sK7Hos
8Bzu5oada8oDX0JqI0A16VObMQOb4YX8m9v+vWaABHcLUAcN46HUr+Ew+8QNiWsFr88l4M/d/AbZ
X7dRsJ/8y5CnLuBvk1O0uI1N7jvyePLQ+fFddpD9K8a8LHb0rTD06Sa5J6pNJxhTBIlfDWrqQ+b8
UtPfIT58r9YfMRG+DpmrAcQtgv/xnYD2nNF88SAmdctdnAOFd5lDBGHkLdE0yensYLMvrFdk5zWX
B3ggvh4tRY4cKEp+yljqmV49cKoLzIYxsyX2KCcFo8bi8Phaz4ufYKhlxQkDV9ZX+3Q4LtRWcAR3
2yhm3+vwUvsMKA/KzZCC/OIwm17dgVHk4RWN2pqx40ktU9e37tNmx552FHqQUI9+WMQsfFNPAYZU
a4ztYIFiZ0yP09Ncy0Q+s4iRr0eHN6CRD0EAwVUcEoX22UL9j6QADC2F4omQWBzPrVmAXB8jVi35
lxbq7aKHjh5VUl24Zo+drJo2lsrA6IgZayQaOSS6t74hgXnD8faVPpcEuzuC8xcV4Jyt07Io2NMp
Yl330SHldtJuJDkek5cYXaJB+spIL2lUpa59s1K5d9QdZZiWVAk+evW0hvsBOZQZJc2gpIoRn8qD
RsYAOhhKTdL6BI3hXsAKnVDsSkpe91GwL93sWb2Up1Ky4QNaTG9Pp62P/RgSDo30AE5vY62Mputu
0grnoxetuOPHCeuPKzWm78miQSjqKXFfKw6MEWDlXVPevpZXrOI0V5kHcRJQhl0zwW3rDWaSEW1c
+tH5B7C0e7r4a7u1zlyCMEZTbndeTSd2UPRZtKrQVubVL37n2h2i7adTJ+evV8WKE4o0Qq8roXpz
+JD0vjiNT7rgfxpzFUJeyBovQhN3KA9YZyuEXLcNqDeMTBqmdEIO5fyNygEICYzquA3uGBtnR00+
qOiJxFFx9G3I9DHU/72poNHMi61l8IRGPYHoPRl6J1OrTyoyE5iQldXFdnuBuPJxs8af+GbRHcgI
S4ZhDFUvcYVGqOnOSBeAe8ErzgCRsD+XqPYX0Poe9BIzqTlRvE/whxGujdT8csx5VCawUcsaMNcf
Vny+rLE45Id0Ef0wiznGCIt8xQs6LYUFxuK0csqN8GVAWwkT8SKQx/rHMeimvqV2Of3pW8/bvzuU
RGk0shLRamoD0gKeZDF8oYe2vhErdZmP8Tqgl7DwyYRbWMf1tm0bgtiVtbr46BfxfjIIv7mOq82e
IbBg3lAi4dcR42SYe4s69H5v5dNm5WmXY/sAegE0G4Ly+A8zjYXbMm2wnEGn6ENNdcqZbcvxmACX
RNV0MDFOOw6kSTiywg5LSikCSWQQ2dEAa03T0t6+eDhTjbdK2LxKIIy8TujvHgh1yKsCdilIpaS3
Qi45zUz8bdsFwsSThcabI6JrtuLXhy/NTz4sQXHeqEDMUvDJMMn/75PdBX2Rl2ns+Y8bXdSJdTic
Vhc6DmTWqovaaRMi9KFUEAHxIfLfuJ7++atwONp1ejJePecrHkNoccoITjflFBqPopSOh8Tg+/q2
3x2rfeU4gFSspDsFaLkPpxuseJs8iVbsN6DQgQrCxDHf5NDFOj40Y94iMfaLeRdLKawZ/N3iks/6
TI0vAjsGGcDzIEfxQsl07WuuBnGJyO4VHmSn+OXRVdJoRqG8VyzxTuPk/BL76H4wK9XZJXg6bDkc
mKDV79pRcCalBoNJIyH6pNdoLTnDbzbJd7Cnoh+Nw2nVXmndZVVbwQy4yFJCvHOsjgF5Fi/55YAi
TQPZ8QLcep0VawUPIfddMWtidy++K06tSyfHcyTRMKVGWDdi41oE01oXxuC7Rq9bkWvC/JZdAm5j
c+JBL9OhHWth2OS9+jjDxPvN+v/abK8cxpaBZcmEn7s27BZxM+HNMHKWbZ4qqrb7yR0WtevEqap5
D5tET33bspRnXIGpV3X1etp6+UOJngZIGjv7/uKaN+za36DJXM6113xg3+rEhHveK08GsHCs8OGP
olf3OMUYpIKNu0fq/WqFWwnSJ8uVYhAeHf2+w/7kKRdZbl11ed5LxkRrScLHDDB7wpo6RrzRAUYb
hxCJ17TauHk3EfqqQtbxUr/oMdBIChv9at2LTY5n1yn/3KyRFOeur+T7kv57++kmuMSpX/csCAHZ
O7qCKT/Y6IdgQJB6VKLYKT5lbZ2Mp/V7md79AjKF1fwlK3KtohcIwYjQ3Dp9WeqrjVaOajiOzvSy
3nkNubZ1JtWXxMQyoe/pHJQy3JyiBz+cnzbOnvk8mQXCyNaosEh6kjdpmbHs9EQUOWqntlxD6RCp
LW6RQyQV8GEc8Z49aTp+ozXJSpI49w7InQLwUUVd/Om8c79h6zOCB4+Qsw0f9YO3JSnpX8mitE3e
F60tIy0HGHCwHbJbL4kSpZi+E+WgfUNcOfguPFdJ/Xuor4+jOK31cAvNgMTvxSmCN1DK8l36Nj8a
x/CE/1duWAEOLvSmhRXjI4QujbCAuBnhcQIkX5J3qiz6PFstn5efeN7VdCpDDGB8WehVQodwzbug
Xw3hmqKzX/l/uuayGIYQowjEMDpS4riuzHZfq9xBEo9JSW5jaFoYFhJCVH5CE8hIqa+BlJmDHEDN
cIrOH7FcX88YNfCPzIfmwcfgroCDd8tplvdcfbZ6niToKlIPBqE9nEngVu9h6XXMCMTyM/aP3uVT
j11keqPXAsdrb+U4AdcfhwWjfZXo4w8rc8SWxOPI5luhxz/3MJvD11W2GrqNjSAPGT/Z5rOmxV8Q
UoL4PGS9+emqed4x0rnL3J1BUMRn3UicAVLLSYjivOoyvtM9iU5jayAn1YbQB56byBmYosUxK/Kf
1yX42ixLszIiUmsnRYSxO2IdKErMHkfimLHCsndwinOvNrOBoffe7dXG2/wcHk2nY6/RgDisUxcJ
2/qehJlsMJg03nEQg9hA9Z9ns2SmRhdkD9X9udqQHMX5Ey+2rkAswLU4NyIpYnW3sConl0suR/zC
z4pwWk79qmuUCtnSeka5XBqDCu8boBYETINQmSzFHlAn5QpKe7gN0rqcZOHA/J8Zg6SEKktl/Rbk
jNTCFsRCNeLB8Z1OpIn+B2Y14wr61stxbYQVHGTM+z9ap+ybyLcnLzaO1OkiGtmR60vRyZZocI+r
wj3y/xxd56XqAbBea9PKdq9eAYXhxqZjH5+qlgsBl3ZiSla3m+kB6FXgxM3cDu3UtN6I9t+ShcVm
Z54yZUm/LtYAJwt6GkaPbY/8Sh5jiJVcR2PB7cDxGansGo/hXYdXtP2uYEknRaTifEV26ofJQfPG
rB+fCJNbAomXvZVxB9FSLZRSKzbSS+t5COSCXKE/eh/4zhR26hfd9xHq2mjSJtwJRF8WZgyJFkcv
lY40Qlyb3ps6zbR26mmhC17RKwtjCLsERm23sU5CiTNW77dp9J3XUIgKga7ioLVuWZFHbzA+z4I1
FHhitwIBSGBY6ov3Xym2rXQbGnTiyuXha338xdgO2uCiAz08ZJjk5TlbMqC8v/P/SQQvJlST/Xch
B4HEHheRFjgJqo6os4GoFvIhRJ8zzG7bTi4eT49vE1KAhfiWh5J2bex3FJ7u7cEVkk9WlxT1srC4
g5+r/tKfzpT1ixMo9cEVRGHyHBrLJQfKBfn+ctb5K3NQ7BJ5/T9iaTFmFujxdBAvwS4CwfDm1iYw
E/oAUBB7+BVe4W+TRASGExzbK2xZ2jXT000Ixi98VS50XNBwQ5qsrHpnuafRdHqFJn7Kl/V8KmV9
VEnuEPImzRi6u80k47rlIt6fxcqr10WfMi9lcXp1yFvi4xs77CaaZCiqm/bRm7w2LUmov1hv+O8h
iA2Iks34+PmUlX7Jha0av2Ip2xD0dwEAqB6iQFfCS/Sgmv07Zsv6CewOu9wIFt300sHaTAX4kNGe
qIguwXAEsJhAhUY4Y6jTKINEg1o97KVb+uscjAJjLjUwYIhGZ2o1xWJt4s2TlPu+apc0hJcqITSZ
iunxOqNCZqfOn+oMQ8eX2LZzeswoA7x51mKFQz8SummYqNhN/hDyFKCH4g6n+MIrR0GaiEdFHrr1
C/Z9YPmjaAIvEHwDN8G6SYZPTRhHwgx1sSUN2FIfuJ2dNfdnioKpA02B6hMJ4TU1YtfUa+R4mSnf
ajupvQhueOWQVjKQLJATdYInFIDAMdmZ/gxyKtCSCHw1Uc4/rH9GBpX9RrR6FayaiGTE04EpH4cw
FWHTt9eTzBKQ62wtnWlELu227hW69NjQKOGzXBw1GdkZXEvUh9gkHpmnDEa3kojUdKJVRYnEsVeW
uYtAJg3HJ8zwgJf4dGk7iGWcRDTZvmeI8p/WqLavUwp8zJu89IXzkLKsjYIBxpBN8HUir6b5vDEj
H0sOyjODa4NwhQRbLk7TFgDHfKav5MXpW7cBiQd3iW/3SUbm5yAD7ofcObjTCqDPwdVMHc3a9Rau
Ub6V2PK3wK2d+fkKnkxa37om/zsNiWTH6y0u9c56zuHdU0KNVLp+b/CyoG3M1N+1mAY6h9qoN/sg
c1/70k0+opgji58PYdAOhJV7kdZjSf1Fj/0P9CucwYPTNuMMeQufQIFu/QCcHpfrAobQe5ABaiZy
O6emAa+tX4S0NSWtU/ginTVe9gaQyANGP40WR+TecnX4H+77+kUDEmoPHyPo+sMJ/gJ6iBzWxj+u
3O193SElSYyE3jYEBTgiYeGgT+Ir9+mTIVQZVD7I15g1o8Nz3d4zpuVy7xMBWmwRTuIqdz0AD1RL
NiIyFOF2PqBOc8RaUYz77Ko7lpGAZgWuvM70OVIiMWLWKo57SJP8LHNgdNeSBALGsOjjIwnMRNX/
3bW6kPqDaom77Txyvqr+6KMJFTUIZuEqS629aiCCvGiSpWyPkM8zjq8LmQ5nqy8krvs0YVpJ5NQ9
Q2p66l54GniezszAyWJGgTOXols+sNkuuSmFy+GaY7DR+VGeKhRkfjM7vAn7QbxxZIeKlibVp+R4
Dpw231aPxNP5wAB49s2ELRl8zvZygkWyrHuUMJsJ9v735RGxotK/lqVdiuhhGRsHPfdLHWLglHdD
o5a37AO39Iy167lFmbAAObCCu14dvlfnPWeWP6PEHs3mQZ18k74tSUHu1eQU2pAgb0AKPnE/TWbe
d2f1kYtxPkW4LVSB8e+AgLJ2fJQuu9/5UrEF9pIFciW16lxP/oEUsf8KIs+kzAcgfiQSZt05HNJu
lU2sb6LM2uhMqK9FpPCYNupLRkYM6Ft7jex2uyBEy6yonOGLMF/97dLNxEsLDUIPdeW3V8HIpFLQ
8LrkMnk62HHHClbHAk123vXuYer0uiHC3ZPaUthFOCtEJwCNEvzbOZk/Wb2pnKRG0NBIlK852xAc
epragMl1LTKgoSdLIdhhTmlNNQ2hL18F2mt7tjm64FBnW586JWVmvHhxqEH767URosCSwSnRDXpB
ojLxOYw9tN4+YAwc6N3Xqq/2sxo3YzHpJm93vXSBKO0xuRi8g4NfBJ9DPI0H+nQHzGmvEA037no4
2MDMyHRkb8G76u5aJeOKNFopRId9w7rt6gCgSXFI7vmYbM6ytxDjKifoGv3cBdvDVBUIaOn055NZ
gqaRdTYhm4JSIgOXKk6uiZM3vEngVlZ6NfrVTjUDKLcI7GVKD1QL1TET4X2i7xAbDS6N9R2Kphtf
Xv8c9hKihq1MwH0PlN63NRiAajANjrbquyYrFILKJIukzvnjCEltgoQJTjYfrEHZzXyAXnCBt4ss
4AVmM6Ob/uG2gO6wCH2XmeXBdS6pQsf5DvcEcNRMrAa5WdrnIzlN56dE3k+XNpuXpYoCxAhY3SyU
V8F3eGLguaNP+ctVv+QzPFVJ02D0Jr6uyizRvW/REg4S2SnrJRLagXNJvQMNxGwHNX+sakqfu/+W
0pX/va0HSGcZ8NmetVAWxFeMWBNDoOn3zAC/MBOu4/FBiAH4IV4hcD7ejkabjYrxdDB16R6ucZti
XssP/tr0gSx4phjVVI3RHYStycvOF1dvIdWj02qHbcFF0Z05GH7BG+Wm9SWliuWCIBh5lcs+okO0
MNr/IMCDfsuaUmCNMwjDSszeY/OxNLFV9oc4EhhvFCHUZJoC2of5qMtdCnAEA3GjKasx0VBiDKtY
G3XgQr+ojVqQRHUszNPnExGRTMl6orzCuBFToB9XWuvRhI/6cFFKH5fbSKyOzKtZRVuauEr5diSC
ivkPDlULBTWiTP8hdLhQLbpY0BucN+CdQC75tL5txIaBgK1FutrQRJsMBT8rWFPxLI/odijKPDT0
dBWW1Pf2Vr2GJFzWcztmDFfU8/nTaxZZBBrvlE7Ut21yygnyK7QF1+YyY2c4Y/STYp0WZIb1STBM
ho9w2YWcG47UGLUgjPKTmUd0pDiFuofIYgDuwfZSg6cE7HhktMt1TJiZTfcAaO0GSKS2MxvQoK9A
GE5rqCX6PW7Ca8wiskZ41bJ+CyNvlNygyc1fS2PUN8GDE/DfTlnaStNFVj80an5f+diniDw3elgL
p3Yj/baIIh6dK8SyWFSJMOX91YajXu3AxDusUzmje10xxgwYi+mmR2XJOJaHxPnkW9hwChTClNsv
Fb+daeCwaeiUjsn3qDXinMs7sGlntYE9gKOezKDblXsWC/UgTSTPwyEmjSqztHcUMyLmPphjMPk+
1QU+J21C0tMWIJRhOb+7ZgXXj3GeW2oyoIe0eTvqIpZCTcTacwA0fIA+UcVES237KvthZ7v8VfWe
aDfyxyaZdprx5keO8/ObcI2npMph87RyHEfUb/se3kCuU1cWybYEHVgH3b3WyTg6pPWN1ailcLco
FDa22xCYhOlMpLOiwEXCMHIcZtvk7YEiYptuvfDyB7Y6eoZbH0WpotMrLaQ30U9sDZLlhRJ+Q/Ja
bjgiwc5+RuXZKZfRPYF9yORHYX+bgtbhp7/E3CIM+t6gbqfT3fGlNamxIXMYxi5RnzLU2iAmZBuS
WIvAB9G1pcf/HPRVkG1AENagP4Yyaft01+Vi9kTD3wR5avypl2AJe3lHcPjuudSz8rh5MYD2K/iC
2jwY2H6Gaac1zDoCNoBXz3jhwNqsrHeT+A7koL11ifEHIgzSb8Ac1AuqxuO01T7BUkS2jOWD65Gm
8Rt8sEPDC0VRQ6mV8w7gofuQOwr57N7O7gBR4CK7kgQ7IEWq+jtaE/YUCOWyz6Oond48si0BUCYL
KCcbe/RVzEilFpncYdCH6oXo8l4QvsRn5XtkbiXCVKvLBobn1wAjID4od4y7lOGJ6f5lJukYoy3d
t7fpU8WO3aFeeR+vM4Vf3R7V2rowKaoiZZWct2+Zi99+ghJiL3/32JrLS9MarBq2qZ9wu8Ib6qS/
+ZnWiQZ8yZaPo9lbqb+XQWR/it0IJSzOOey8+IUjU1di67CLa1J5ZOG0rfyoWrKBmZwEXHY8LnHd
V7w54hcIX9rU5LDLuGvDK6l4+6b2CD1Ai03BeP9fKYTp7HRuTaeHJjqz0aUjUJpHEY0zVTtCoSro
s0esmtOJM64f/AXskrVjlRanar2URNFADW5+bo5wNnpTUVtd6GkKed8ASxvxUJnSUyUWp/9Bqbp+
SU7WvwUfZiGR0bmwDU0IMDVMnc3td5ijH/+9z795/f6gp145zrF2+I1rqUEcybdyvdsIuv8+OCpa
irQ17wDReohJi3oNm34ZIg37s5/BeViEERA/ZhcWQTXUjBDS3YGYAwpTLNzm9V0s7gAc3ujM0kWN
ep34d46CPhGcGzz6REpbO+WPbSdzBcM79Kp4R/bNCbPGMT85cb6DCnRoUVka3zjoHxNw8zdSIsem
TH+2VFB6aWgB0blurrhpLZQG9tbtxCtyyPCOxssaCemiHy3vqxiDaHlawjoKc4yEu3zBfnOKCFAq
LpfwsyQNzuf6ldm7YgpG6aUzV6/gpEJLYmEVtd6pvhArHbLy9lPFt3aLsMGNWQwrvvKpvwHDLEhz
UsgOAi8d2AI439+W8pkaObSIl3FDf2SatVxi8Jaxn+lZVuU9VF0hJbTk4ILOOT+EuApCJDfgE2JB
SqjYVFYw7YItpROC5MPjfieX7K//I0DG0D0JFd7VCW0SJK/IdM0aNyrMCv2b4VnoV2EsauQFYaRl
VPfX033DJswLwYwsDZWyeD4vu9OuIBSmDR19ZD2PrQZ/mHz8TagX1i1XemTzaqOP1uyuJmrG+lFg
6o+vgm3UB9DfSTFqGjOQpQTHIQn3mtG5gqsiFD11+T7MmMh7oHOl6UJ5WJKv+hD5aYA+wn3DnrlM
YlDLbtNsd6I0jVN8JBI4nl5/93evNiGpOkpWjg8X0q+bDKwDqFsZcMD3Pxb+aFqTc6McQN7d9vYk
kyPGKJbN7aCEnzcrTDyaCXz8i5vpP5xISoukfXAJO4ucTVTUqWhIIr7zUqvruaIxAcm3MhpovE3v
GETenP+pP9gjLuygZE6ItSj66Z8aOJGLGXCnb5hklSlC8EwTdagwZ6/O1HEY6is425BSEvz582ou
BUKDPW0mEoZFUbVKs//TXpmGTMMvJgtyevPp5cNbNRJsxQoAkcNMDNSTbBXkAUGWiow0nu91pCw1
t1ddkPuO59KsBK7JNZyReCk3JMS6THUX9vQ48/tZZ49yEFsZQJ1BW1mmiDS4lJYGRdq5eIZZDnN1
gc9qlu8AxRk/FyMMXmY0XKaQsCzUQ7fXmxwio9t+9+VIGNsSuDa1sKoWPcxdqi3iVRtpzYmPNbOm
+z/pTC/98rpcuek21czGHMT8qeetmU/LzZ01teMTpoKmJusi7waDFOj/3c1N02semN8fDYbKuksI
MdLVSqj+WoObVsyZ9KxqKdjNn9BAHfqR6jN1+es3OUMg/hiSxPkJB5oCaALfANrpW9/NiBkad52v
5wF5ttP2ejJkbBzeCQxkIoIXtdaFqIRXvecA1YiVOk1smKql15dEuz4o68Ak8pDww2FWUedhgsPs
EI+UpzNLcN1UHdKVpz40d0eKRd9zeQQmPaGOujKA+y/WHB1tLXbj8cS4UkUwOOTrPoXc9L3LDSba
mO2WsuZVX7l+gOamN/NMqIh8Io0uf7P4ZnvehCGGITO0Uz/3B4Ln+njlsLd+IrzW+x361sX073nr
davMtYcPT2olp7W1n26PA1EkK5Ce24C+enqKNN6xyxr8pRpSm7pN2ENUglKbWTeATZ9ZuOJDkeOg
ygRaMHZeIIETHPqTVH1x6FoAUADT04nzlgm5FwXMz8Lrieq9WUXZYKPlME8MAMQmm6d2P4ouyql0
E92njV9bpf7eCvYsBy4k8RIL+EoAMXsf4NZV4NbIgOEfqwyqWi4/bgLlj8uP9mlHJ6TpZ/Kh4UZS
6mileXWdRfE6GBbEXc+2WH6+EKm8BpMVCCNMo2K6JpFcJDSCu8h9Fw6oAKxcUXg3U8fvmKZBAmuT
uqXV6NLxNcWSmzJlGa9cMtCpVVkLKR1D5oAPoNL7OEKhxTR34amur8s3UU4gnDJLdGDslddS2n4t
UHdxi4419c5rYVhv+0fuM+Mv8J7Az03FgWEJxRW4idNV16JIOyokEqiqBJX8qM3tDbJzXq1TKxY+
DX7lJMwGPBR/yZHLG2y16N0WL4IwoS4CO1d+VBOOM1c6OHqYM5IXiAAazltTZe4oI9UsQjOFNQ1D
JqZZpMx1cR8MaqV1O461gsdwLlj8YJMxDjNSV1tt0vYqEuCY1VaegLjcBGR+EKKpBeSRXHMKo0p1
7MegZt3/ow6Ef4zbg3zdbQPdn5HV7EjVyRL73cB8rVPNQIyuQqBdrZi8koJ/ZCbLv8IfDjqnP4mQ
EyJhp+raJIYCNdCYOXUQOboy/GgPvc/YB/zKBJ/zYzqw2xRE6e4w31Iww08T5FMcJpw3sdlzFKs2
HYzzAIueChvQt7Bg7HWB8dayKfpG7zXydC8K2ncpXbfwhv/ICylqjMbZ+IpWnLu/rs+VPbBh3Il6
G1jWVwxhfyGDwFqc3XR9P3gersiM6YkbKqMi9HnwzdPuJ6uDlwZPnM2eCYzeCMIJxquwGhkxliL4
Oaw3WwOxe8aPDVxiw/VnCuESfMN89MeiNQ2mHFgl4pjay8KOqvEa8wBTHOLkDUGFZX9uBcv+SXub
dMSxO4xr4xUmT+1NnyB6VOYbx4SADfmoB9Gg6oWEorWH+G4ReqzvLpyCAsKHKtfpD9Ceyfn9qfNz
eBxmLnl0i76C9H50hoz69r88DQS5jWaxvZS0y5gVqjIOKtDzYEe1jBTLXzaWGqt1EM87gf0Fp+1k
1rj4iccuObcmkmiM4a4ob0Wyt+IT3umvXqH3VGci9wgjSZMVsYNOFW0hTSW2yppq/se1y/0s4KpB
Zpp5IwOLKVAi35lwhtgUS3FTlSf+8+x52UGjMLw5cyZfEMJDmwZHiHxrLPJKFCEmwv0kPaBNzajo
Mp1iYwoMVrNNU6n/g6/EKzzx0jsKtCc6DxeRyxBgO04boUa+s0tdC2ldVj5LsnsW1w7kQuaJRwxa
RkoqQhq9l+b2tyEj0angCsGXBURBOyXhoYAvnryo06PkZrQdOSMITzmlDEZ9MrRmfOj0eZb9cJBJ
uT+F3xXQSkV1Bs6tVfreYHHdX5qQNFrcSSRfu10AGGm33k9bhs+yGVGHJB274Q7Mby4eRBas+bxR
oemeGrFKit0yiu0Zbjti9wTdx6t/AgKKq4TfJDXGsiGaKZZqAK5l4+Oy/F1RurbruM3TPg0bhR8N
ZL5WXfn8/VAHJXP7o558thZfThnsNBQSr2yvMByIJD9U+zyus4O3Rs8lVuBmGr/oQM+whij3X6bm
/kGw7X3ZeXrnlg++9PJzg+tl+JVxRQyTIZGwYhnj2yq6LPXR7NgkGIAoN803hnWyF03kHYBn5Pd6
SWrXAM3inxpvHahp72vO3MXrQ1YGXDuOxbtJ7nSE0TTlWNxmB6aroGCIb+l10gxikpG5jaFDTTJ4
qfkVLKgJnigfYDqoOzR0N9cpTAWWFJJruRWAnpymHOu3rHJ2ewDUt9ffXZDWawdgp9OzalKPcyYZ
HtC/FE08qAJ2Kq+J8Mym8gkD5jGdmo/VuS8x+5M0qTwBu4PrlE7B8ztSwZkRT9kkZcgrsOWDo3Ww
gLXDJnpMME8u1MjbCoI8arfd2uq4waMRDK+CQ79eQPlEW5mHnHhHKdtrFzlaDvUceVSvUcqpphvE
PaTbwE9uVwqXZyuIDaarRLVz87BqxqS5Hx5bdqyjNpbn5US4l1xiCdO5uNJLbJw7djMYHedZhD2R
n1pbrrUZfVTp8nf6iztsbo9A/CVAyo3AKlWIgHVzRZp0evhnwBsFB2R+Zz+fCQ3ko62sirZF3WQM
WpVRrjwWx/pX9YIJqiHLAu/Jzor4zVP6cc1W45/18t37y7Lh0PZo7V6CKK8jCa/vPmlX6WvS4si9
IcRodGUpwt3dGbefxu9B4bDurGrEWKaE5xSzpjK+cTe0W0SVsdSLfzOwoxzeOhvPw3Ppjo9/cDgm
Y8geDjVVoSUIueraXAwPCFu3V5ZX9dFe7A2NroqP3L4d4p6ULPBy/tqeCXqe4Ut9z5lzPUEnNlyh
gOzsecE3D5BuEYZzQhWcLNUp41OA8fHIUnI+UeXytSPWdpF6zYhAqIajIl+qh8yIOz/R+RXi4uBE
mMQf0PlhCVGoow0moxXeiuv69CcZnxjqwJFrQ72ipq2jlG/JFKUYJtwNVhObV4psOzJjlsjSChB8
FMZ18heajRvL7j94vUvrbSb8lzWaT/PtqbgCg1CKy9LQ9KAUUrXM+yIfJSrNu3sQhy/0Bh7/uk+c
ETTsXp9zjFcdM1ho0a7LremvDiqux9R37O9MTJnmFJCS/2ypof/0ddc8ERt16nrY9pjdHd5rOF43
1A5ikXJic44dBJXTGQqZoQV0BQAekX0OVegb8jmudHYWRvY/Z+Izj3Kh8wlL2egrYde8ZlFJ4YWo
xN0wnBYMuzTun7bUBkbvVY4vOp9+5rMTVUKwxEZxC7Bt8f/TfYs/geKK+2DIq/iy1l0GqHeTs8u6
we844FRdzFecpGgS2KpcOFSD6DghJ22r9i786g9iI5/l+/pbxHxLlOd65A7cWzmSc+HMHrAhUOPj
5143srXEkF89z0DvIWdM8UxGAf34FP39CIVlkjIVCM4XP5ztKDQ7uQ/uY1GN8D6WbCW6ppPVu6L4
fZSNJ9hNRonRNGeUfCWQfuQpg/Jjty/Vx9xnqFdUFfkuMFl3ytnnMdw5b9eJQ4Bxx1lJAKTO5lhw
YgH64GKiL4tJtvO3lY2flt+hpszR5rHAEMselgHpWtIKImVxueF5WLviEgV6FsHuznDUXltffFy5
kd30tIE9Rtm6Syg8FudxgSYX2MvlOM/ukffJN9iaF0OBBT9FOzgrjGIApftdj6rzmjUarVWwmc92
u2fB6iAD2LssB0dastvo90wGrsdRnUDbe0foJdbx5KUxrvxKiOu5eF+cYZRxavGMdVsPwEOsVi7M
e4P1i5eV+GKlvKY02vjoKonwH2Ues+qnfyDYUXE4I2qrfg5oNT2lXioP4EPMfhXSzaWOKllpYU23
p7mF4EMU8ikb7vPE7cS6zkTyqkXsnsMAoxb1q9947/4eeKBQEQXpTDksavJ9uSCCMeoPkB7APrSs
vbes2kbhpOt0LX9NzRtEuHASo15OnFKigEo8iYPfZe91//Npf0vXhGDNKpIHOxRJzO8PwPN1j5bc
Vo4PaQWlQC1mvUZ04izyP+ztzArxoBH6Vw0H0meWd2e0zH8TC3I4xRN5RJPLfXXLtfPqR8xc33gm
STZfJ7aZous5kzg5+3GLe1QgrU7Pyl+eNm7iJSIB6GPL3w4HotW9Tu1uIQFGlMk4nSzB8vHhqf3r
JxyET40ZRZRv99MjU6msmxcb+0U5z4WdVpRH23v1XcEZy8co6P6PvraRwKx8LwUxYpJ29dr5yRZL
iqFJA9+bXVtbxwBZTbY/hHkM+fACZyrX5jrMY/huclttZsIFmwXoKUVwRA5dMZAog4Jw2QUgpkyc
Qk9ba4UHb+YrpVKdlMkITcBcX8jMD2FzHUj7K3M7dDxzvqNo+MnsMUuAeZprh6xlZc5QPpQv6/jh
PG+ZIagXDyb2F/aZKGWKIFTJCgEuCYOqoDKE42/Osu9k9ocnUH850qtmy0Huz1EfuGGTcqTgZPtC
WZDtcqgq4PHPF6fKpo67WVoGwrub1W2R+zaZtH6DzmEkIeqMI8qBZthZXpDJcQjaCqbPGVi/KARO
HQIUnr3vCQmxqKb/uBFfqxs1MAKN92RrBDxCMZm6iQVOqsV+EQxfWmYAyPHOhETkLymPBjnasByT
N4MK7MAZi8K0yYveKuyMU8siO3t3NS+Wm1E3rmYU1LC4fnICF7I4e++MNRkmU9PzyH/G7HoTMSSQ
NOdIHbyrbJhXVno1YNYMT51k4avUcqWMX0WFcEJX+R68sboKtHg/UBALUVEjlr1YBFyh8hjJRmgb
9zXk/pCaC+xyfya9fIvhhTZjERRUxw/eDGGcU5ODcRSLskecACWtKOJDMvnR8/aviiftUqdNZjKM
czjhFbjDSDoxLsHuIz3zRa/meV4aR/9hZHq2sPHtb3w9JF3Nw3+gyuC65O34WB2g72mRyXjkRl7c
wBF35j88w6PMs8MPjNcHPv7kiYVZ3o5eNJht46HpQrGA7DzWh4VIM2ExlVMhNdoSF8GGRBHG+3+P
BURJJL7TOeZq1iOe/tYumdj24zYCZ70Q/0Tucp1LSqCodweKSXkhPuDiv8OmAOF6gyylGb8o4j87
tTKQodqyVOQjCvDUxs5MtGSUYqu144YAB+LO+ByWr8zqAItwk95teIzwasqhLocu6QGimx4DMONA
x2AxuJRCqbeKvDUpaa86CyKWDyzGdxDv7j4xvViRHPV8YQiul2CcDGvlTzYwyEfQnBppxPIuLm+D
A6KTamB6ECzOd6BRtwiJEsjs2O1G4beMXem02fkilk0roe2WbeuE6BUw99a/x2l9JB3KYl2eXDCR
ZPTQZoqH+jPM1RpyctPUdEOkzwbUoflQxCpl5Q0RuyhuG9kY1CnijrOzbYIiKRsEp9yxOL5gwn3X
uqBfc4V/Xn8xJzp3KUZiho7cozD/2E0w0rlbNLFlepf7XzdPcehElz42SZxYz3oE1BrBleegsux1
SAgvgoKnfygSk4xk/l5BTQP0NY/XvOPYliqT2pZbwuC/3oeFYu90L1m074aXRcwXmdPpEVsc3/Rv
zacm26CU90PTK3jAEXB+4NEEKISUyz75KhwL0J7cucHSJh7j5IWj0R1jEoGsJF/xZhXyteQfNT4T
LKJqQBa8EvDgmX0sanrmf0S8Gu+YnHaKKxvpmz/Osx7jM3HD+CT3aFuMmoGQqbcBcyDpXzsG1gsG
UawYqMNseq5ez+6TPhCYTxt0rSekc4PyEGABFzG/z+JxweFoQ1QnyTnvFJzSYvFJovOLsdHIqNot
J+mCzKfh38fQ4lTGJlBu7EdK6qyns1MWsGUFXSBNMERdBBJsBkgYv6i8pb2s76VY9vVKd6yA3MG6
wkuvO2rbG3FHJ83MSjirRyw6sJzD8qlK0cF+OAIUNRyszPWdGYEZeXtNBrD8q9Wr77yLEtG+qRYW
tBKbee1c9mS7YrnOopt2t8gX4SmKVL3BnucMBdcGwOR6elHRdVjZ3SfBShwZ8RmI2Ber/Sc7QdTr
zPA8IAlGwXVbcJbnUTBC/vjBr1amuIehc+3VQNtW51hYjrUYfNqoyUMwaPkX91lMykET9NFAfTBe
FdHD77J6nT0tjk5sqoI9cTCBOh9Qc2Ef0vR/lpi166KkOhGOxSmwiAWVmCnpXZqe38KI6Vxb1HtF
bXYJ4PZOq+9n2pR7IufFbyCQckdUDWL7JCBS9+BhJPZpzJ2ck2Y4A5Ljq9nq8iRxqGaR5lt+Zkr8
MbZNihD50skQfzGNNd+0Y9A99HZ7pxNB64lqh+46Dw5m0lNKLRAP3cks2F7JOEnzKSuHgKIiGS6V
S1S4nThZ8vyTpUVNGaxXq4WmLMs15XMLBf9YqPbvffglCfrwxVeGEX292PdK6wYsISvLTEBEJ0ji
AsdOmtHSifjFjGSHjHav2WTkq2AOvDsanSbF1/oq0l4+6/45jLaeHlr/F6TH4DSGw/IVwDeA08qd
jLP6AybVlkbOw5UGaQx0H7DwTgq0gXuYkYBPJMobFglA3KTRvREHfclbz7gJKcqryLeobHQVjiI+
HTbEtTMbSU4lDw01IHMP4FkRCqA65boyG/jueRueWWZhAcYjPUXCqwLQ5jMBQYsDZE8IzAk1R5p5
9R4BX0fbALGw3TqrY1Ia3pqDuFWHmY8m2GZLxeJMGcRfoPHN50I8zm8qf9695/bxAfia4+eaNImQ
pwSetLTbQN5iyZVAEu2G2o6Iz/Tu9GNwxs759XhTcahaaOMPEIQbAX5DiOj9rkEujCuBtVHNN6p1
Ix5z9rVxKPRks6HGK4CdB8rajp98uI4PROi6UYS0Whg3PLxBX8f50ePGSDFcZ7tQ0LmkvmCdeFOm
CLTfdePcAlYh5zjFcqQqTOnRBw9Iy+tpxfCIQccm9NwhaBkab30gaQEkn6TBD89HbN+xc1u/EvNY
LDLmsPM9kZVxOABEMPSymvDVMjgiY7idDII5oDoXFQPVxLyKvpZp0M6qzxHlIMNRySB4D9bOY7Uc
EAhmaWcJCs8iBmVyqfyhW2+U8+ieRAae7uI8Q+QIMUHOPvL5Mn3FY2jFIR1oJJglrDyTsA0ECJYB
Y965LMwhsEs1hruxwTaerc911M4E3amwVHXpjyCnAuFTo8aEXAD+BcMGrmdMRpKvi/0qdq4ZnwRC
ucT4Voi8YaUe55eJryBCDkszF/os9dbBuPaUwKPTHKdHW3AplBGm9+LmcMk1maS3zAYHGzLG09Vs
oJ1RcaY2WAxD/1unN+mP8+uQwsE8kdpUol4S5eecFjnpqvIkkKCR4CBq+TVX08MQp4Tcifef4xoS
R9R//Z/Vgjid0iwOfdzCnZBz2A8xxTERN1DClsiHvZ4/ANwQJQtQWIGOMOr6jR0YsW8dx/tcG6w+
CPtdrR40SEXkfn6Ul3tfk8UOvKytQzQoT/Kx3aoh6sL4yb/jGETqauSr4VlYiCmC0yR6I4jtFFkc
vx42KA4TL79ytPWXtrJGxZJy7A5srbM6fkSPQHFAmo17DUiCchAUFPVIpPoS26oyT9DupiQPmI7E
mRTcskSp052kOGVnQPOKFiv83v2vqjNK+nFgWTZI+RCOHcld/yKAckPaHAybwTQltMf90x37vZwL
NwZxwy8zaq2ELUUrOSfqcVyzvV/jBnro+zddrT6lBWpYHChbT1uE98TvZoozAoj1YO+PmAoYyxLM
jXJnJz61SBqVlaj73uiLEt/0iDAPCdvVyU4ZtcE0A7wNSf5La5NH66oY5QmBan+LmYL9b5TA/zD9
GIK+a0D2juS9gX80dqwjOiLxb8QS5Gni/XZKSL2ADc/jqRZRA5DUu8uI2QW8RKnB6DQfvCtvkbmv
g47M97rAGrKwEQz0V0P29r6ayohh3YHhNiyjkNnC5UvjubPJhkSv8kTB4i+GTI9NUM5yg1C2O0Eu
Ff3XwA3uTwTQM+CLMdLmXacvnGoKYwDr9BfNJt/NEqx5vcLAL6O8HHkbjaCYBMFfuK4Bj7KO1vNl
gBoTJmN+ibiatOxtyAqTsIzSUku6kaBcBcz1/HSpLzs58cYA3fTawZViUw/2gUS6+7W5X776Aei2
yY13LCZ7IG8C0RX7S4GfDeQqQWThxkmU31liJESygwWPTW0pdJljECkhgZ8VKU0IX/OG1FYN4BRH
zdWXy/VUiuxdpnLGjOIpIRpS/4dq/3Ax95rS9lWPGUXW5gY+qp3Cqs5owqY3YVvst+IkqVHvjg7U
YyQPun0r247diC7lFmZpR1JBBLibkGid/An4om/04+c2zSNxa5I1e4EkRdljgBWfHd7V5kiI6Wma
RGA60KNFtJ/4Uj4bfXEm0/jcx2wqrYGQybDlUGDqhqWMPZVflf0neehZuIZWVcN73nL1+hBEXY7f
5zzNp2llotzGGNDBiS0h0G6VuQ5t29uvKpQbkhxvrhooiXRvuF2J/NuhxHcaWY3X6SWay2U1EsSg
OEsYuZW1UmMmypIxavSFsULzeHWBgKqboO9TVhf+LEZw35JqTphNS/Af9ubzFc3wz78YJKrDwVfh
MnsB6DDilXxp7U5BtP2/3bIiN9e1TCu9Y0xq7l95ln6pTe/EhBx8aGWfXEzpydMiS19cYqBK3rXC
a4Tr59tVj1t68d9hecmiS2cms1KtJ0E3yWWJgL6C+LSEQrkU0DoX6D4zh8xnEsbPz9zwMwhIGUdM
G07xAcw4h7R5jB0y+u8PohtbIFFR1Algx0Rvgr+nM6c2uxF65fySvOPVbES8JIgbCE+X4wWO5v2y
bmUuMgsfPKr8ye2JvoDzmMe3InHX9IKiBsX5wnz66ZHEZ5kyax9WnR4EXiwYWwLCAggnALOVSmYQ
V6eY+5YNVIvynEWzN8bGR57EzU4Ye4o63FUF9dIPafC1bTgmjQTKtBdqGbANwhtM0rdbe+uD6lX+
9+nDU5Y/KYn5IaNFKZaonszxjI5nU5V4AlCgYmrai7re2QjReplED2L0BTehbz0g7dF5UPgfUqfB
X4omsfeBM5+XQ6/OQsGUDF7atFzHEmMnY86gjT3fmRtranuKpQiGCorNsVhoSIpdtQmzbGpeFrDW
8tSBPL8Vp3KFeM7qycrZvTmrHbmo4FQ9kzp5TMccDHNyNZSiYADZ/FBwi+WVOtXEnukIx352Uk51
wMtVJYTBkxYPFhogLwmrUEU8Q0cceKp2W6dkb28J9pzD2sXsXnGnjyanxsVf5rlVmhC2DCVflmFs
n1cQ890B/XPMc2ND3MTyJYONNhDmyOym/KEgS4o6tEZoy7pz/jFKWMPRnE/nL1NXTw6aJeG4Ddrj
NMj9PQT4JHAIULb4FpOjNnQVzGX+jGFnmM7tZ+1JjdTht+WHefmTU/AT5ir0fo8XiJW5w/zy9s5r
6xnyKq7UYqQbXrWyhm6o3X8fEucILs/W1cxQT8EJLfGBhfGFzsDh0qrF+hnxZdHFxVw74H56ucJ3
SrqXS6RSawcu+0SePhKnRDAVvLZr86vaqkrpdqO/NYkfq+wYQHwCne/SUQlJQGGGqDnY9niOfurR
3DJQCss4FQQW2Pv97XHYZW7N23ugKRqcIuvuHDNcHAlr2ztQsot7lBPKgwYFf1/k12Oz8Yj3G9FQ
HkSHW6FmzksmVgDxhWhe1OvqECMAIcYtcky2v+L1mqVFXxp+oY89cdV95e8dkdmHBHgqiJCe1MZm
n9boP6Os0euJ+JkBFl302Ay9NBqyHHsnPD/Egmvw32IC7p5Vi3yE+Z26mB/vX+SKS7CAIfSn4w4a
Pfpuia2ljfUEmQufrYSMMr4Vk0mqfPieEOLnsgucxgfgG4IS+ho52qe5lVJiS4whPfJIegec5fEu
K4IWHRAmLpSp+qA04oO6q54ESe3L0NC0fW7G0wx/QZZ6nGdNvqBWs7UKx1yXqdnPbqkD9oOGrqeY
zerdgXTY2EBW9OAlWGe50sQRdB+sftv3+SgkLQIgY0xRxZHtU+dgLVh4gyIE8xQmW+hDdVzGeO0j
c1/GMrTYQcHKFVaouNy9TkQ+HvlsPVsvKaSJnj1ZJRcua18Pi5R90U1ufeL8mMclo9SJ4bL+3mm5
w/lTQwDQ9hIfb3cwLPAYonsRGDvpARSPy2Q85GYMiNNIT5CronKVUgwPp7WLKzMXgDuF2q9wKrDn
hsTf1ICKbKSfQxbSROWi3ATljvFxz1fWGH30J5Xk/Ny5tamDmcIMQ4QOeH/3LgoB0Tx7v1heqZgw
fUlm27A8sifb7/4O0zpJ8G16/ikZITIQOPsBIpq+oO2xVBPKgfe78ASPOQrdYcuIvwtHrPuRp2Wj
0Hh4dh2dEm79kTZhmtQssFkXaGl4pK++aUZ91NqrhnOysYYJTr28/0jw24QR8bW1mJ4jKYj8aeLB
tR8AMcbyU7oGUeE1Sr2BkJ8fCVn18BNJZjsTImriCBPzxgor0cfMWm4Cl8erUT0sDaeEa8jbzNGI
QwB3Xh8JDkmP4hgkNiPFUXn/um4DB0XBi6m8Qg/NnCsmCybhX1/bJFoPpKRGQ0yNhbCnLl+eTvhQ
gUxfugCzQmMxQPCkCYHbeOmlQDncrNLPaxHYU2XXrjx7iaPJuhtOZFfIgjOr3HEPS+zYc4+3GU+M
1BhDvRtOytokWIH+Y1SRbTuj5XFOx4g8EIEQBUVsfAjHWKXLt/0UfzdZs66xiUavdfs+gazEBlF8
QeTvThXTriJM5/HNSue7I69U631vyXQahQCFt1zBI/sOjP0AzK+9cS8JcyfMFUzr7XNusxNeYXPn
8EsWx0WKMrKxDa2NGvji4ovjU3NVWWTjIoC/BB/X6baRaWcuVGLxQQSjs3NIwLmrtDv2Rt3VDhf7
f9DIoPbXg+vTKvGkCNVOjGA1GssfRaKxmFH7q/vniBJ4SaQ6WFmgt46n353Px89t+1EbtKf8aEdB
X74lfv1EgEJmswtsU39WG60WM5f9XTbwpn3fADZd3aixlhGBjVGVBOCYUvdVJvxlSqWnLZKrbOt8
/HFmlRz6fC3LDNsXNjYN9/1ft33MRdlb/mSxsNzxMXYDdKHe7VLu+jN4nXtpg1rrmmP7AgfROdHT
zhXGksiYjmWCLXjm2eTbQ8FXaFGQ9eALn9TdnZR9oYwoz3LYgviMzP1UklfYiV6XgTnuZfuugjJf
FW0Zwg74dTNFqbxhVT7rsthP98I7/OiiTARkCgT3G23UFROrtEwWzlziLt7fC9UhOxtEaY5E5rg8
F/TyXQHfcXalPu1Fs0HxtEJSMGTtAk7x93/yQucVFXRIlGwYLy8JCPkloMQ8Q7oYA7oAygS5jb86
DtN00WziJS29R7OAXyf0AnH0+0p1ZReD9Y2NFH+lM44WVZghlBu6JOuVJbeNl7AJpkJvwRV3oOcs
mfHOETESDPmh+6oIo0OEfeQqwRletY0OQXHmQ1fmCl4WtdWEwX5hedy1MBSkJ0y9POf7CnCbfFop
ZsyuAB5vdT7pA2iVTc40mXTv/NPeXa5llyOtxTo/ilHXEQjr/n9BkQDaUGm3Ra0rlXiI9NhTd6X7
DsZ52hUjyQr+odYbGswCuQpP7t4Evre+SsCfg4QBvldkSNXhhxTZiPxn/bTFy2znnzJr5u5eHdOk
JkihLcYniZ4ooxQPoSTk1VkxkncnDGFKud2HIYMpKnyzyxjiUWNn+Kagv1q96w8vhNONlbpJO3wO
ZdYAiQhWKlr2XC4xKP9FYhuHjp8K6EL75ipAq2WC+pw7i3nmfNUGKzOCzZTXNBN2w8L4H+aKmmi4
fP95WIIBSL7bem9omLalm1LYa5dIlez6dUxS5rbu/c9KEwoitMrpbuX0QfYQmtWms7sPB4bBmGBV
fB8ASCKUCVhUuJmxggCaSGUcHGEvhqBWufp7tobcnCHJC3hHdHFAHFO+6znd19frszdmm9K9YM5y
ursVvZ9YC0/oNAaKpi/deNvZnAMh7R/0ReqgVFHDQFwjvK6N+mOBfTNcCPGcl4Hfx4WhVIrUiBKE
j4rWKp96Qw7pLTBloR6P2Vu5eKf/ZWHkrJZyZ9POGiGmkawuzJMGxAd0E/iEOoUJXA6RNQ4Ky1Sj
+RiCUh0fwkiMEAl8e2ngqj80tmhtMxw7hpKSVcrTZcRktWBJZo+gJk+/vvBd98Kwi9v04QZ0HanO
ItpDgJUi+zXGFgVFKAydkTfWdW079NKCWaTPtzTjLDGfpuinnXEAdW6mUkKl0B2pccOKv9FT/gpr
xrHJ+Bfz0mPMkg5IhAOnyks52wNzpxRTHNaKua1/tQ6GQZPlowycHHstNxb2LtLnnsOAg7pdywxP
p+/4BhsX/tthHmeSLW2UH/C+fgiQckIsd1zMJEpVJ/vq+vAL4si1L1CXVLV9Tim4nDA3e4Dtukj3
uYQj2Ogzc3fhscmlIUeZeYKkWPHS+mvDubxVmw8WwKbsROTigsKOS3RHNsDU6s91NHa0MrGe6vbu
MsWmh0iGOK6Z3foLrmrA+ie9+jR00H0Bwgu0dLY6O78bcz87I1KObOIxCgXH6iN5ml6mR9ZiKYo/
x2YjaA9YFvjlIN/gdU/ZqvO/H7GjBWu6X2AFFGnxGea70gICdYNQ+55rE7443Q0DyrzJ3iQ/jLF6
t+oHLvmptJc9M6bG21HxxBuD3zTPe+w3RXn20YObRNWjdgQ6f2xFBpkcNxPIUhCgcExDkhSuBXi8
9eJrV1I9y2+mcyKAXmCvf0y0M/1226e8C4EIKkyKAB3wwkp/1KfTTUpnX5Y94SGl8xQW2ETWmOYp
znRHfftWVjCgdRZNh9TfAwrxnGXDwgcEqZ6+r6soxLHvRgMx+In8cphWz/izk60ClnN0UjVjRGxa
rpj7qhDcGfyCRckvDPV4CtWoro7ox05PcYtRn63ngDMM1hKF8UdJmi/gxw3wPdmRQMa7zJgmZoWz
thKMB1uh94kvw+MChMSARQX80210SAaZZpmH+5sOgHrDIPSKqxuzlUxkkuCWG8BCpjg8m/2tbPLR
lNNgVhvwo/YspgY34SBKU9y1pWxS33Nl24zb3TGDHao6g1b8p9KW/G0V8RasVtvEQ0hb+GXnRbKX
k+xdKC5Ohno8GRvIcZFbzOdtPpZZh0L56Azyg/fquNsr2EQs0o5MshlzDk1VrTLP9QaHbdFvXAOZ
clLSdv4s91ahq6vJJhT6fkjnfJ2ssR7wPgQrC3epjzXEStWsuimM7sdeZf/iTUYF2L7b5mRB91gq
t0vptadJZEExgJpqxRaVINQKGZqW/d9cDaChMAU9JlMEudvsJgcDyzpKUN96ur/tmirER2vwoDXG
aVdPhgPYQ7u3lBlUdkOxhmv7J8LJLXaPCoNqPfbdmTyAHctKw9D57eTLGOfeX2r1+5ElWb7bxHQB
JlaQe6U8Te+KcVB4h1VutOjBp07D9YKpSM4dI5H6a/b+KVCDCNOVrf43nMVOV+6IXAAEVvr05CgX
9Q9dbC226ilK76lfBS8ECBfOBF4OiIhBe+KOgLFZATQ0PW/Q4zXJCGvN12KXYH7PjNXal8daJm12
ssTvVHU7bxQT9cdTFMwfBiGaxDwRskbbhUgbJfBoZ/nBMFk0a1hlSbHiWELFVyKn/VcQMrewS2rX
cAB1ncVjtdjrEgY36sri2ts19lKOnoHNeODCJNHkpfZyK+EYMAwuKF3M/fdPyKTk1Uhp7GU/7k6x
vX29YI9blcxsOpRluqsZIDs9Yxoq+Somg98Swq8P0gEGdzikEvD/5YTHzGoVPespWiC3gvvrj2fW
qU9zL35nb+oRBNGPBFGK2F0af7oxfUlY+5uX/fFJL2zWf2NXBHsnIqkkItO1D+My/0FlkQSyWHmu
8JqvDNl+X6TG/D+FIo9TQ3dQ7ZrqNb3ii4PKeJteIt8Wg4Ik9kv6QjV/Nz3Iw6aQ0ViOu5+UsRfi
11AE3daxZmbgSj5fbfamG4thSOP3/ytim11mhfm2fgF17p64YSoI9tEXKdDks0gEQBO5Ha15cG8d
aZo7ckuq/zrb61YqLJ+DSqGedkJleqsup7vut+tSBsRW4b9OsqCY02UeQR6v+4tyllpN5oshg1iZ
hTPQQYBVTTDJSmLlnIHX7IYunXsrMjX2XWLH9LNfp6wHeX/TeFz3JrDs2ocLcrpFwAYwj0Op3l9o
NyTH98hR122H3lMauzol0uneWYhcUMoL/Qn1v0cOotXSrxzioglrKq8C1RKHTTcr4/CPTFeU4VxJ
24Di1vTAvKaLWGHKjUV02muDmw7+4hyzDd+WkCqTuj8WleoxSaRcI1qyezd+kqa1HC8h8aSaG/M6
6zsdvTPHrMzc7EJ3KrIadNcHpGSpPMg8BDCWyn1K7RW7jbdnKEbPPMgp3Wewe5ucPD8JXQmJki6/
p4m6q/1xRPjs4zTQD+vAa6H5cfPGF4ZljWDA3JD+GVn74li7W7oru/1Lz0uZ8lLWmqZZ7sVSN/6z
lW/sq6oaYMEzxpgKPOtJgLxxHn9FcT2ct2QiQD3HkPv/lJ1+zuRgdJ+AjY2hc+fFKifCM0hE3+7m
9FY6hAbXKFhQbTZmbnrmccZ7BJD7oS3Lz4914xapoTMlhnLc1sTutPrWKk2K9FbHFBVxxwyMBhYd
D0AYyr43ZF5D4eNR+7J4L0w+gPzoTJ/vJoqsJa7UI06TmiR9ng60NUOxeGT9mcLElrvvZ/4yuq+B
3xzniWuACWpQ7I+xXXxfBWcaufUGcVKCGxQ6sKUhG6OhU3ouySXDwH27hSf/bC/hMKu8fvjnbVBJ
mTL8DEIicp59MffxoZjwpWjdauptQL3i1HuPvMyy72pANfafIykoDIX4mJUZHMAs4UgnN/DqRA4u
4AKQVl+xJTSLSKCymgQUWhWblI0XGOBu257q88QQWx04/rZywS//wK/ivQdCOss4uJNh4Rh6LRQU
0eUPucMmI39bfpoZVgbZVvBKJc2gXNZ9dS01kI918f1QJ1f0oWNsxaFJ+67tfUD2ruOVO7M5SKrs
/LnpXQaRhYD+xActgIPUnLxajEcSOsbRn9KsxHM4sd7hGlqtp/u0nrLkrY0RDUOlm+TimSj03CIZ
RRltlMpOvQ8tT/xKLOTgre3fwwh4PC9mFRFdJ34MvZiUGnVFODFoNFWGkuJqvwsdQNrUiRKQyh57
t1UN3Hure0gwgrk5Pg9r6Q17BKQBRmhgvvM542kqY3pGZ+X0SJy62AmO41wFPMuu5A6rWL7R1pz2
852eavaxHUCx1xTTErONFIC8dAWklaJY2nFTbtcrp72z4iG2CfSonmlS14+gP/ITTljIyHqr0CWe
+iAhtRn+P0fI2XGk2IQpHiuMjfaG28B5cNHTDpNIr2DYkqFEvxd68hsh6rg8yOtZYAeW4AzUu7mM
4IsD8Lzb8SBV2LsTH22yZ3IawnYB8C84qNFfnyJXAnZOZycvB9CFn3stMFqKavxFLt9B/WHOfgbt
0SSJL/EJsoJbTT/b3eLpwNoPxk5wjgX+sGjjqpKYJh4p2NGYLhNru24OAWhmWCmpLtDFCzYkcSuQ
EdN6eEyHQK7qBnxxGfOsX7kt5jVnpNnFVpNfneKY2CYczQGDgCeYYk0T8sYusT4f8o4O2uEgkkwE
I+JlgIz3yALxpCwN5dNMwi5LRV58LehR490uXciCJfWs7Ul/I0hMbzR+le4Ubkfd/FFYKaECP7cY
qx2UWTv/IBhd09iudlwrR9QUBHttuAOwPm+7i+PS2odxOK9+v/JjdYFhSrIcXDmijNfUrT1uD0VT
Z4hPAaNc+6ys8qUvzNPA2BSeOTtzJTuxWx1bbEPkRxjheiy0Lm22g3T1+kiSnMFqrWOWgGXVL7x2
BCRHkHEaVWJyQn5+NFc5DgfDkY0D2lUAoY2AVT1T9fbaNni+jZaCBE4Zx6M/yGrwauB5G6tBqEDC
3h50NNHtpMVvEv+0ylGtWSxyRo22Tts9XwHu3yWxCbhNW+lbjv3urNdIdNNawaWXuMpTcPmz0FoC
//bbf//XtNnzlCpo2IjqOAs2PiJWchPcFbid8/l3e/bYkpuNZji0fmuu2D0jh8vc1kSy0ynculiP
B4JMUP5a/8PZ8Tgr7X1s2opGsvKt4HVkm5C4nKQjLJKMO+WWgI6qaQpjPXBkuCn3R8iQOgeGFYZ7
FvKqDKmNEWF3Dt1ebspGJl14bCZJkNB8ittecd2gjwzVVqI271JU7wPqKvuXz8ZZoxWk2SMihGcc
6UXJ5xOy2yooU53qHOf3U0yjEX7z5/wWM12pvY5J4XhQk+8gcZa/kuuzFJVt6zep6ON1qYyCvgwX
qYT7cynqoaTa0ssu4IXRZBabQchPDO5tTGizQ+jdpJVp1C2p9KFYMEgJkaGlKoaENyvvR+iE46R3
1w8sZn6ivsVG1x2DgqmwUgFvtUld6CAKVIQ7OZPz6jBSx1WcKVPb2xtdQokK66nNxyiFU0fiB1nD
b+dtRIQbyebdCZQX+cW/B6IebR3Fi/g1/64SizT+vRJtQ7e7wWOTl3ym5UUpQqzdw9ABSq1N5/gg
P24bbYD5r2AjeSySV5R8I/hw5IrjMqYAt7AwMH3c+dTfEO3B5BQoaNVoS/fla4gnOuSXPhqcuo+b
9ph5eFQ+gUMvuBxhf4ccv51KOwfYlIPHETqlcjX3iTv/yoVqHC7fG/yCuVrzvKRk7/qlAkdXnRwJ
/OBzD02X9rO3/syvzNpgR83j91AbVqmIcfrLqxZlCjiqEL52uSv63JkhYCaTT1qUmfHcRTf7voBu
+bdAiXEKrPPqxEUsFPLJpwvQChh+H4RFGu5d+DoDd+5zPmwK7I280xlgpYEp6xloDxMx3zfJ+abz
rKdiQg9TN/L4CL3FCUYPNZjcXVcz4kHSzKe0kaH8kbimhvZYND5QJAxfxAVqcc7sD7vG8G1EaTi8
aYQG75SNRI4pdX/MzBHePBWEionJA7mhLxnRUMoDGQoH/l8aQEOdcrkVujyWnr/tf+PnugkJP74T
M63lDsApQd1HTB74/azYGQwg0MWCz1A0EZQcmhJS/775b0wEGOCNy1ZVL1eAWGVfFOEdqk7/B5Pt
bDKWNIJbJ8po4crz2n/n1QK1+QG0ZwCO8OeZ9JKCk0ZpxgStpHKG7tFGTruRb9Hx0b/FjDt8/6B4
Vjg0dXxxHu6X8vPx1NxC8APT4QAqyZg4Rw6AzGOA7j/R+vr0QnGiyPPpFgcx0OY986dVAkLB10H5
PZKB65FTVzRUEkvLR0wmqkvNqPnQMf084SgAZ+X3bJqM2PU3hg5JRKgn/YpeQM5EtGBrHi47OXwf
z0reTHBpLlMvIwNOFfwObUTc49ZQZwxSG/ovmS4fxupnpetGOa5aMFGNbZTuiY71RrBJ9ELSyAhR
+drolCLvyVwCHkridMX+Qe6shoohEXVOw9hB1Ugn0OQCjBZ0Im0lib8AkoUKqQEGlGWv31j6w5tQ
btYvH2mGowqYFAgxfnYotfZVzF21a5f0/ghCDQ8Blj4U6LrpYYdQT9efF/LEOzvGG1aUV1phIbCd
Lh+sZCC8iZpv6uHO9muMAvwwuzaZeROwDVLbsrKwybEPHzh5+3H8U63jDUWnq03Qyu202mzfER8u
/otyKr5HW6kgSC0qL3UZiPLbR5roqvomcJmJILrutgaB3S2bOgqRIV2/wBDACLzP+ngaCFyI5FxE
+wP3tTTg17Z46YrvY3iYAyilvg6abrkRbh3/EpcehP12NtlKHReqr+0rHb+Wl8bZE94pgGfPX4Is
L4E6PzRnGTdENjhF5jWPaifnwJFl71eMyBgyvu5whKl4q15/nkcA5z45tw3Fdup8KmoKXp238Gz6
OEHCvKi6BZSeMjlK7IdLVM4hk2WrRX3OGYlxdhJS4G8Zk3pGBK7fv9Z2H7NIuzGzjPUhOJj1DBKp
pPSC3nm7b3NYP8EJ+XNUB9HAweWfkmumfONIpoMVQLMcF9zue4lwbfdrR40IMW0MkwxB5KPGhaDR
r+SJQzVXUr0v6HNKtMcOlci45kU6lT50krnr2WVakIoHnScQ9epgk48M5x4cnd55uOJNOkRc8OlL
WZKz9+86lRJjHNsuqvgE38iItQO/lHowmgWnWM1naPILx2aWzAPe71BGWlO0My0tu+EfXFuvrs0K
bmcqLk7Ybi0bul06HflhknkxY4wLEqWALJqlNaRXmu4qBGPeuQxvPBjNMzeLb34aytsBf6YMQp/w
2uiL0xpVGrDNVUnbpqLxg8a5ZAVOA1+jSp4fPixSlpDB7AjDqli+VX6pWo9qZbpII3HTYWTLpAuv
uk7PpQqJMlDVC9uWJ7i7eT6qSx5TDqpWFskio3B2hHYp+Qh7ty4zXEsFXwd/OmTuke2Vfyt/PbSA
ko1OWfS318zPtoMVg8NbhGhy59F6Sg0ARo0ldP+stvskjAFKMIOKbOWVeyFtIy+aOVWqfoWqkBZ4
/fl5N71PM0DvqYHlCqTfePlivIToqlq3HZ+4suXzcQaScj87rr9uQqIK3zE8a0w08gEjfTLi+ydU
xU36E+f52GMRZJgTGmRdF56Z6ZY+/6SYByl1rlp0BDje/lMx8IAwfg7czzipnGP8ZNVRpImp1wSu
RINQElOLvLBCdYgZWGzCTK5zWAq/y5MiOaBaZWKhM+3TqEOHogBWTrxMLAEKb8wcp7DMbyVLzuns
8l2quvyuUmalkYe+uyzsUx7NLUDY95RhkDdm1nJ82SLLkfadAk7Pb24hlNrwfz737bnOZzIaDQlS
v9yceNLraSTSjtKKpFSG6ULfYMaBvo3DJNhh6sO6Fy8VLamkWoffwPcAzgz3V04ELvqRZk6s/jCD
uC4zxsHoOlKnPDsTxp8pz9FwVNp4eGsoF67H6cbAonZ/+TwBGf0ROPPCIcYoTUBknwFqnuUIk1Vo
/sW7g6UM3Ua7xr9zqIAB0NdxSsPuy5Eqo/ttvM5BJFBwf7WBmPW60p5gh+BrTxun0EsBwtlTTe2h
XZq2a/3u6hJINFb0O8fQEix9UnoQWyss4pBOANi4hsTjOIxsv0LmGMYwnrjzS+OXgrow57g6BXpt
UUnwseZ5IGKeeipNaxzVVlgnGYEisQG6+p9gDN5hkBH0+nHGlYhmtdxprGyaSvLd19pS4ebvQsqH
8i7uXs2dU6iyuxPUgOZF0yPYQbjP361xULyY+ke+ZlIzcND1I264tktt6Q5AtgFmCKl3gog+Wfc8
Q2euxpoKBnGjBtysSANVxQQ/LLPsBa//uH3VvPOX39OPGP02NqyRtO0dbuUdsLa8uVwT8WUEwzBe
nKiNZpaEZjuZy8Muoplbcuu2gZYcPYEhMfWS+XniGVtPLje7vVXWgthQzDRZNIVsvDuUgLM3eKZI
hR07Lh8TgYbWHJ/Fhax7zy7GSHjbZ6xDsPTufkVvq9KackJqy4ilsv7nuGzQc+dZoeCzwe8dBiOV
j5e38in+a9s3bSIOaN7pRaA7Xz+TRmpaVflcbqx0xhAHgVHvfZ9esx0KZilIJIt17/UWxwHY9BJM
B2fxM2n6wooqd07BSC5sFpYw8TnmgaGTWyA+EmHKKGv492yr5vf+YNeileVm8bsinjhSXURI4mzU
ByUmDAXK/quKXP9b4pf/l97Cvsp75UywyXjz2Ks5Yq/AycROSfIOtSvoUz1dbLaUBG8MRnYcdEEg
XdIPz9zzOhZ1YPcLSq7nwHF2DTR1J8TION9wkImvH9ZXjaM8qCH2A8ZEImB4Zv2oJAWo4CdzNGg7
0q18PNWFtv9iFUxkBGa1xIq3leczLes5xNVRiZ5Mx4nL+8UXUdZsw4f6CWiwwcA/NVK8yAJmDxR8
An+1Q77EAkrjYDWnQLiZS3kiZd/MJBtuiPVlM6idFUfIz+EfIwDO3GbPoDzpTVaPj3GIFyU1c9FV
861h03Zp6fXeacOZB9UhQUXLbA0V0q2yf7VYCUCyT2fB1inuHcSuiKQ1MU/3vwoTt8DVbQoaDy5W
s2WS0rv4ktQhDLR3wILPn0wZvdAfXzTdGd39WeS8snj7SPcSm74ZXwd2oglyV41Noexvx6rgKPsk
jSrzmtu+urIrvrVxQZI1khj01RS5OhgFJ9e9u3bzFhPkwjN4bCvoV5hmCM4nxkwVG/uLSzlljAxK
PLqDFsu4qd+9JwdPObZv1L6JMnDOQspEAsrTP6jIZo71QTtLbhRtjzjO7j7GvY21SacMXpqNLWPZ
4J/0ApsB4STqyeFv5Q2Crip/t5PrUio/w8KvEnO5E14qt8UAwVkMBprv5EzEHRqNB3WxpnWOCL+y
UodxOfYxNfO1+k7P4ZxCAxj1ijYCLTKHUlDY/ZURRTsPQFJm5rOjqo3S8oL5i4ilrABUeJznZ2yb
CNR4WSP4LMbTG2UoabgrdLs/01cb99wajgrhXBZSEn+FtBBHCGRkCH6tm2hR6SZPOQUB7aHLCDXM
3VU3ynoddmEOSW1JeTglxjuP2APC+WgMat9YnC7jmf+IJj4RPGuMnu8Iyqj9FJQZLa4D1h/rSudF
uMKScAp18Js5PXenCTJx82mConIhASZu8IkxNZD2oOv35q1rjhpT13mZ6UoKR5ZjaOb5F5Zc+CtO
n3B7O8B6uzScFO79uGhqxcvPhyEaQqVW5Tb2aYpM4Wl/TWHT2PZBSD6sh4bVuscUZCL4C+co9eg8
a9YceKa1nOOqOw2+7E2ZChVhsFNBFwOZ25DwxfJWQOjXsN0IkTXbxqtnk0PZr7/e/UUyXPbhNfef
4hfg+HnuCcsAZikcDhD4Z7RH4Kbe80GCvF1a2laQl5imCQ5jp/TcJMGKrOMwoNPHWrv8p7Rw9NSC
chb6mvyxSXwzYCIll8Q3ugNjFw8RuBeIkW4jm112ERIPMBuktARhxoNrNX9ConB/Dfgc9QgdF+Pr
gTFK8ZE4JARb2sDcOidKwF+1fboNO6HHRrHxj+Z1ybBSVpxNXgbQT1UAYXg1ilXJlRzwOFbtgbxX
Xve2wneAWJsAh+Dm+zTMpEF1F7VUoYiJ/+zzGSJl3ZHmg0nD//kRAuAg6lqVdZhryPyfwJBd21+M
LO30fr+0KTrTIvrWCyxqVBTqScKDark2zZcWvrom7yukTBw451DqamyCTOkt0qH1LPGd3XkYJzY7
3kyWstPmhaZJY4+G8gPoyQAnsp0sAiffMQyJN1VSsVx2cG68uRaFSSHS1w5awFIufLPFe+BDZqIx
JRq4yr7Qv2O4pUvI3el88ulAbkGtOub1+oDwRWHUzWooi4tgABLSaHRgW1/+18mt3e7t5kk/s00x
AsAj7UL0ZjHprMw4ephMPjDBFAUkr/3YXGe64BTF2MFccEwNb/dm1CyaLkqYs4qDaaA+ZXkC55Fn
qfeA3ZvwZ8WkOyXoePytdO/qJ2gSz4Kgm5V0prpnxTdvRAmKlOd0j1fevim3t2lYQqxumI7WXVQa
DtC4+Iz6j6FpPyIFD7GrFBmmelPZES2stn47YiG2K+q14/F6lAgo628iLV2xhB1eZaVFgZNkP8+1
fmfT8uOQpiWti+kD+eUGSLNcNc/wh/mKMJ+xxXRF6XQ2WEcpjqF1i+Acvj59n7epL+iMOrWakcLC
68wBLGDKq/YN0aE8dm1vE4gGNMIlPpg35Hwm9OFIqxZ3FvrpM91N7y95c1aUn9dEbaGV0v1BC+v0
sGEnoSxiw5es7aAAoJoUzZnS1N0BD1LlNHTBx39QslFFrUxzlUuwz2RCMOgiShsEXbgBbYo+w1LX
GPj2RLxasAlM/+ZEkn5eX6l53NFv7YWIXS8iKYL2vCTwtyu9HkIuw8C+UYGYpxtWFN2yqeut98I8
jO7y18nSvgAV/3/Xx8WT67h9269lCRWFXyn6hskNEpAqJxbVjIgqzELNjLE0un7IquUG66eyuup9
DIiUqXWEf+xFlS82PD0okZqbdVR02wCLH9atbZECugOD0e7XK8wACBi81VIGaJD1d2bNBSFlLCOu
8HkZhnPLOczLdCnCwQq2V9l4yv2Lf6Qt/oPKUHSQ7eAn4xp+47B6cZrCN/A9h4PJuTkG4/bOeIbe
cyFLqvk/vjP+Rw4AjzVgYpXXg9opJkPg/ZgN1K3wCsS9pVwlQKj0dPyo9qwmkOksYtFLR9/v97Qy
XfqQiXS2IdyzM/gtlILKjhfEgO2szo/p9H/IuSc2VJLDujHXZLY/4p51BSz18SgnDsJVRubwrtJ8
NKeZzaIVCCeqr/H18YFyjPAi9syncH0x/PyH+RRnnMGktW1lkpCHT6ME0N5cvF/HsU1hKeRPIDoR
e66egDlaTy++BRSN6Tr+aWcz9KKBmTq7BespBOy2AdoWS648GxBYpcUnhHjIOd/ZJUNyxnvFo9rW
RDlomalxBE/X6TPXjwHTFEey9n7ADfHRr9MXhU+qgdlSOctDcYIRJTXMQOR8xx+Q03b7StF+OJiC
LoDL86CrbGsMv0aag+OK7vTJ0XDtdby1UEX0HgMVDuhRUicL+TAZ7d+b8zLG85k7ixNEA/McjRrB
h+MOJ53diou9BUSqTDAQBZU5QR47RlMV48EN04gT8gaF4jczRE+YfRgsh4q6blIC07xqvaOljYxv
IUIpVe1LogaCB8NqkRpZOcuN/ZiBl8CwPiG+wfhH7POGV01QKSyv8dPmbjBp3u6+fOkiF7+xtsuu
qumhYOWNTwuuHX1vizzLG5gJRA1c7DNeCXWFT7cxtoHNpv9AD+QYm46N8pGumNeyC8FZXUgT+Jx0
ChFiBADZ4c9cSt7IaF1iQiduEsqUpmtYUfWwY+I/ZvOs4nnGuGXVppJ5pDi2YOQAUnaYwF0ub5Rc
9/xyGmrHNJ37raadDloUiFZrNo0NgU73nI4O4963wI6WgGsFBAF1C7GVVYjhkmsHiEQFbY99zon/
7zmjFv6Zs9RXdjzR2RtL/Dhc45TRlVUjuAMdZl3aiEQhD5PvXonsgUtgtbiGKungnMpmgKJ+z7JX
paw6tSR8fpipWPYmVotDOaW7vrBZarLTG28ucuCpN5Lp4NSED/IhZoBUAMYhF4ZpPH37Lpxx92XN
0j3P02HOfEUeQ1XFY2BRv0+413/LZlEILTn8mZuBvumtkCdTEQ1+9HLFoeofBkm7Q/DmDt6qXsm/
ckKSWz207voGaHODaTEx1CTpSmb5QEfffWxX6EXq7TsA8Hot93PWU8IhuYLz7dYckUWCfM2h3947
7ZiJjGDtL1plRpBFpA6XdQqw5uvLkySNiHXcmFp7ZgFFGY1dTfpLJfhqOl1vlZGDYuCE2cXTtiKj
olhG6pdZzvvH1GRA9xAI31aPMTQoqcSE0k88gXoc+er9OUV1tPz+b3Z+OnDkFujojIQ6JbghVKQM
mCm2prEQUVG75ekutAW1HXaNpDki4yPQAyJ9PtMJv4PUfZ7lHSwPOXd6nx1fs7++M68yAenC++O2
OPXB0ZDbphQmf2S3YYEBaTf/kCW9OMj7TMrkeUy5LqcATupzWWmp76D+X65Py1e+8lKtwK0EjY5i
g8YonoBXB/gW/cz0dmXX9mbYOUC7KEje9XSdJIOknh5YT8u8JQphxn0Ni4/dQjsw/X2RFZTT5Go8
2LMGhiWQPxHQXJMK7KGa7FY5f4Pg/xZexAA7cuWSPJooclWtfbdDkf72P3/CdpNaBWzF9wzgBzuJ
91Ab4tTsBNqFVvOSyYy0tAhRfPgzWprB/xhEE6pcFu44cFFllo3/KweqVT93zMNJEmzBXM+xZuqf
cjLteBCmocuWjkrMpAFba/iUUqxvD8cwkRN/anlVOZH6eZFPO6tj0G1FuRpNVh+XqZ3XV8mFl7ZU
AuWHVtx8u687giIe40hhqI3fUMTGnbuUG2RJuykT5G2mUrJQUPT/53oKdN/xPbL8aJf2thDU02zt
ZBd4JfTtJSXM+oVAFp4Aht1cRm/lqc2cH+mPNR289WDrRM4caOPgv/qoDWi8M7+Mkn8Z/SRjwIjT
Vh3kNdXvlINeuqurqMXm19GBQbY7ktYK/1NyuPyOOe3oAYxV8nh3LqwMec3BT5S+1GkIZNMYZ7zV
nbO4AhESCCm0b+einQ2WaU+SR/Vng/b+qXjm90hsLkIbPuM28yeiJqgJdjBQX902b+uogntfl4v1
9xEFXowmEjigvsgcoDBFL+DCpW0EmKZNaaKAPvqbc2j6e5BYg7s5cJ1NlsNJwQH4rbBhZeAOelTx
SMoI4FATac6IEziCDz8wcO34WmLVnTW7z0+Ss6Uq4PpHpry6vXO5OJMxRv3cv9Qc0g+i5n50ua89
ZWfsKsaVgUIDSX0AsiBS3oGQefH3zQIKFBMm7TRg6yDC6fdxf+sA5p8G3q+c7F3QVoXIUKK6eBQy
GwEvuHRZX+noPtbBvWH51Y0FQlVE5ZSFAC3MkqFgcPcZ58BPEfGpmCN//3p43X4AO0uq9ZSTpkap
ZF5lCmqlfTlgYvR4KY3oqew88P6TbjOKn2yqOnxBsA3LtL+y7T943Iqaze2lWb1RSoAoBxqzrcEs
QBYM2cZwD2B9kbZTbGtvSLnzKtjpkNhHFpGanZrB4I+oMgDDy28jOqVOEt19X/gY2w6WCY1ZkXIK
yZQPtA3XGeBb0rlJ7N90iVYtbKGctZD5TZtXHf3bqnLbMiLxE+bMtHY0QGP60yz05U4xRN2pqiAJ
Z6u/+P4LLS/tmnZHU8/Ud6HCZ2XA7KI4obLp11Jf95bIkmxsiL+m4is22P1icB445P1NZxaNjhPi
c3CM6pN3pARNAYhC5iVMgCq+H3nRMyjeLnvEtkxH6J0ulA0kX1K4l0CJSqwlIlrfOFO/VgtYFfcq
j9/R6+6aXUYUjYGtbP1QivD9n1c8l9ALxsl0zV6StsQ4ngRivD1bXsIZl91pWrbQEnfvCds/MTX6
EDN87PRdwWA3tq4rShTa5eny+1LRz49HAQkPQ52+IEbzbO/zEA9uYYy5vt1g9j5cP1VlryPaIbC8
E4o1omkSD5DocKayn+LvvsEruENwzKuBux6qVOTRb08DYTG37Hnz2lCuafo+xbOPV+EJHok+20Af
h639VKhVCqDJBaH2zC271HK53O4jbzAFAT4s/ZGAgnGrXBF0SwRAO027VsH0i7Tp1JecdmtPFQ97
782Jp6AJkC7d+JwdPkgrXA8OATvBF5aq3rgptmmIlfP1y58DepL+QSBalTxdKFpr/mQbthio3P5W
TCUv7KSlUbZBX8adY+6nFf+i0djhsRKOEZ6+47P9DcPK3GKIYMsdbvAHIMfloyZe768yGxtK9XNG
G4Fx7wAVc18yJvq5d8/iJEjUsTM1XYOv03U9ECCN278BaXolBgMKzJz3vXQLsEewrK6kOvDvUa/M
rIsdlysUyrhShuSyLH21hE+TjyhSC7ewOk3O/lTteY2xMrxgvfKMBfcTxOkg8AXFQNnI8ursp9uj
yUDJBHHP6RO+E20fL7sRaTKbIzcEhSozykMMdQHU6sdYT7XogQRGkHueTBaG1sWZBwL9V4Kkq3LP
Z8Btp5gDX/B+y6cxuGhbx4dhfB1kPuW/HSYD8iXsi6i6mUtYvelt71kkg/O7+BGMggg/AzWkJW5w
MPhrPyKHF0jUy58JFDeqvNwhAKUVWr1gi/+Ljrmw73TIP1AmKLbN2vALJWPkOAekwmNCO+/OiPyX
k6Qcb2xln9Ul5Qcqh2p2/aJKww4zCYJzc/KNUwHatnfaiX04TOTooFCGf7idBFqYxnmeORQ3ezhk
6EPhPNgaJQgsey2mOXGCxzWoymvQEeH4fqWY7fVZ6L+zPRyGtMVHVCZT+xP1s3yQnsBc41mn1FIP
qlTh8c6ACfkPGlIuvl7qBmXQS5VxCRdfAtGSmayTizpUtyep+0SZ3pIj6+UaTS3fLRHWSfA+Tex5
oRwEm1c/zvxGxjOqCFvaTRXtE0W4xMIHF7xsYfVd+3aXH469tqRCiQ/wXyRIsoB0tkVYG6hXfdXv
NwJFw4WqlDyP5FB/PIUEnZI1iV2HM5J5fAbHC+ZUjWJPHHW8/drt7XlQc3s5eahlP7qekzqcsNc9
78SKP8pRQ+mlVwL/wnkEITXu/6F76cOB9HKnwMo714C2yniRzy+y7b2xNn64zPS24KKyjqtt3+Sf
THddJo5hnNsSZGhT6FMJohxXQpuK2+pHCun4csWOCctX0Q0lHE4c6kJnE8qrf2m9aRl7sUPKZMyq
63VDnX69ad0aT2GIj2+Vz6RffSPFWP6bFSna9fZ/7lO+Yl7QBMmXvViGIq5mybTQltj9P2mrRub2
0hkv4AQjkc0GYCzd6WayZMQgSlgU3my2m/Oq+dJtt6Ys40qxPZH9rDVIT4cpnOgJZS6CiYvzSMc7
HwT0wuY5An9bclBbAGbLPmtMCeiXylvcX+F7duGEmYxJv5UPR8avvq+nT5G4PWQ2sXWN8zRI2SMH
KUmSIcSo6plnW/n1dYQn9M7VOVLt45ufPUevxrHaV/ZJobr2wej/oqk9k29zN0wDBoXVzvzycFzd
zdPo0hQV0XVDDuM/u1DLeAwoZiiGhuj4t9ivl2ICkjSWTlWDKbFPpKiN15zWLA6eEBF8hl2pUHNm
zKTtYJQQ3vQlUr4jaTmlYcmL+Eu1Keqzsm2MoAiErr3e7LXWWsTuJZTzMYbNnvFH7BiNX6jHGkhw
n+XQbZPetpf5R1G5RJveEnWdoLoE8S21/KrCjwM6ZiVEN6wyV+5KWkxnWcOVOTYh18BlRFWR4rfe
cO+TcO7jh09v9V/L3R3VHbrVkkyZhbkdFTdIxpruKL72oeB4w3TJ3i3hOyHsVxXY805e2IIZjhbs
1AfBl5xYq9pPGahQ0aG9+NEtKzcSqsu+XhshN0L3HWec39KmBiSAvar+0NGLo8ho46YNfW3aTsz8
XNeZXbdZXctbj9nHVP3kOzS7/ja1qqPsfIz6hd3QSCVcsevC7+XUUc3QYwf8MTL5/bH+kyNv+sb0
hC1H4LoJWAf1c9rMSb/tC0NtwDwGsLVDtFbtWNKMqxsqF6QN7KtTLbsBXza2Z1l6/qsS+5iFDcps
r/cp7WHeoqoEmnsXqW+I3AAcugh6C5laBQ12hRoX7ETXLi2nx9Rq1YcI33n7EC2XYDC031+uwDhD
bghe4ImjhnUYXBhKZHzXolzBNECFtSXzk/dgamCac4S9hIWstL4L+ptnoQ+uFn0fFzS6CEk+0Nsn
nFPJaywzOyLpp40Qde8QXcG1Lq5su+Xzr9oOmmltGN+5qAr6LKH/1vbEhnjS1atnus6jpQbj+wuy
fxJDoOEXpBkM+qxHIPu2ocMg5B/i/XHmAy6/n8pFuip2IxgNLVUn7EbDwGekI5VMAfOl919ZYZKN
3Zsp5a7uRKYDbnrtGBfvy9MCEcKH0NZq9Ce6rMOZls+fSil7/JxrQkQ0c+kQBJJUMklN9/sQnis7
ZVQbjxhKY32P5Nlm3yGjvX5QWGDf0vAXgbLFELmaonjNTHjMLJmA6ccN+yPUDyPukzn9WVygVDOt
D8Zd3U8VGQZEdE91QHvzA5v+zbSDdCtCW0wwoEt5pf0xX9yHrx6pmEPaESifDEwZFwwbtn+7+psg
SM3djtB+PGGDh6UXa9uH/8bAy3RIdeOfrpeL1iUQab+EH193RpeYErs0G5qq0yMuqRb8YUbwzIzw
TYlr/YjWmEh9oyQ7iGcja67hiUrtWoLn2PwTEjHwruXPr5GzPZofc0kjpKcWt165/YFuWgujtjJX
KKaaBFgV68vUPWn9J3iTogpWnJxASbwY9qASj7TnBor84IVe13QL4hSJZp9nPk5Gv8XsJOVZ2+2V
Aovj3GcIUtWvY21/XvFrFB9/4NoMBLEFDNLSL/qrhg27JKA+zBVgNpvMQZ/2coqBme6UDMPKDRc8
GSXxIu8hUP2qjIqrvbUt8vcnJevM/G22A1M2dXFQ5HFr0vrUauCM5DzbiuILr1GZEYi5dc7Pvzbb
NzfbQBlrFoQjfnavMVoQy2sGh6F/+Zwk00BjY70tj8rX/shAXd/FtgMfW2XPs7UygEmKG7K7K0hE
uJfbTMvPRxhcc7SzU+wXoL2aw6A57HDxdO+k0T9Y2zEGXyIS1bWZFT3+yP5sAjORvcQAruiB3hJc
tTRDEUaVQaOR42dGAZD40agbnYBaHPR4NKVTeW4IP1qIOfOH/Q9xqqNKV85mXeFbcg3F9mRdGQE5
eQI2T4ewE7wjT1fiVR2Iyvqm+GT+sjGmLPJXPXOH0310RPjWOH8GvUFtJqO7xzluE8Yrzp8TG/LT
S4uR8jYiiIhi6crYZaaJxsgzEXKlfE3PvG/WyoO01B/iGzLl8mkfg8oeAqzzfCHevobF9VQjldrH
5zl5PG3v2DU8i0D4/f37RCkqTdk8T+mzqM6Hio5nHMxrT4j5pQS6nFr34WQfpiQU4J8mwF282aXz
OIE6c6WveO+QuEEBEA+9QhOx6KSA0KMQQpIA0Y+boR54hrSf8HEoCf9JgR1ezwP4IS5T/IK+BAKH
wWjub/x8y2OlXBOgItsZKcvUEELsEecYb/C9P50A432JH1vRewYIIPS/sXQ9PFzL+Yjqgja6+lRj
BtkshdVA+RQnk424RZcnq0blrbttHjwUkGA4nrqvpjNYl7jmDSfNDgTfQMU7+il43zxDYfvsxNkw
i1PDGwOExVj9iPlh+sNGtjBls/bB8SWjqDYa8cU2wnKZpjkYaH880DiwVSUGH1F3cJ5F1SoM9UmT
UP/J9H4tl/2pLRPbg0Tpkkgn/qOrXCUZ/XZ7ckTUFPCpx2CAegp4vphBmNToz9EqzODy8BAFGTbv
Qnprj+6SLbbxtzuPLz1QmRSWEH7WSwm6X1t3kDYN7rrCk12EOpHAndcqw+Nyj0H5IpCMc0I3e9Ue
nC4SToKkbrfB52azd89rBT6XGiDyUStTGAuJLfHmOLoQ8SMhe3msbtGmhe6MCmWMx3L16EtiNTOy
m7Imw97bINpl+bQBMBLYqLjL0CUn2oiLUlau96LUb/tne8gzAzOqL7GzRb3jJaf8OeLoHJuNfP5N
e6Oun4ZGvDHOF5pVJ8K/BQGWznnn/lUg6LoqfzobcVkN8xIoo9BgdVoLDxjK3VYOmV5W/YKc/klo
X4xOZptkSiwUpBwAUlsnef29wEQVRU/YYD845K0FrcjAnf8eZXclc481X8ZN6SAayE5W/9dtNs2I
VjEkcTHPK0auuyUtVFxUMT/aLjoBRyldpgaOYlGhvDHCe9APjKNH6/H3XFyDvLJvWxdTZ5NdmfPm
zADgSHE1gt1/+cmLK7yTYd3FzcN2/aBm/p4GlSglXhW4Z6uGFvr2f4a3bnsIU6Ml9F7nAswAOqyZ
59sO0LdZO3QryPmaqiX+sb0NLQsUHs0DfetfNQU30YqjbMr2HGVv3eidKo0JOxfh+BJgoVZqQifv
LOl9BvenbggJfOIl9xAuh2MzRRzFuQdCZCfZTTlZ4Q4AOGtFWYcFEhrg8aiCAM08+Mb/dsGkJjUU
S6S7WKDnfcW47UtzCINUzaWNEkdWBM7vDoqHEWD3vi7rx0z6Yy1G/vnQEHPrnqKKHLoLpZ8FtJb4
w3Z8/85wgifktLBGbNyStrX72Y7BBBvjnvvzActp2+5MMpH10wZxbwq1yQsnQCZucuVKnDMA6+AR
dr2tZf3UjdGheN3pTIP+ejCQQO+2ikmSL2zsnvpHI021cum/n42XT7VMjsffqB+hs1B2rJtfAh8o
SHK+UkyTwcoMiXulLJLzjJr3Wc+3lREuv0RDtklJy0wgrB5CpmRITwSRa8A5jBlb0rKafHrIR4BZ
9BtRUP6NDj6Ke4aCwIZ5gFJB+WDC5ddZizFw+TLytLCOC7XV+JL1/DjrOikigeNgRYVffh3mG6lw
/WAItNk1TI83AeJrP9BAR7hvzZGuw5LS/hwbZEB7+gltUv5/vjndSNxcQ74djCder/qPlwV9O/gs
71tWHKU60nOcelQBKWleTpfpstsVb8lGYOfOcF+i165TpPETFUsMy2FhZIdxiQHguDU2Ira/pB3E
lqBf7P3WS7BdsZrfkUdnw008UJM3G597/SPz8GrZ+QarXiX1i4hCZeNugA+wNBpaApK5GW67dLfa
F1i+KznUHtwHpVd7ofxz/f1ORu4B42+g/4DPBNFaJXfCdUmJyAMa9CE/yBHuegyc0shIv4NGfHw0
gsR0v9iAv5AUjk7VdmrSeWeX2T30tkRxZYjIDAUcaCCT+Ci/Ok8w1+uPAbpRqYnSeNfRORjufSyQ
dZcjr8JZvERqOgOG6AVTa5prHZaJMobb6MnT8JwG4SLJmsao0IXzIjNm2RuTj2RJBP76PggMmbc5
xlXNPXMlRTsXGRt9TvQVg9IDQkJhjxHpDMI6MV/XevA4iMiK9pyy7kMSxsw2CzqYPq4l0Nv3oN5x
e73Crkr3I3zFYCT6H2BwC+v6wS+lbLQbGX1ej4qcrOYfK++jcV2htUtl+LO8PS4ZtL+quLKEvyJv
yjaQ7zlVXFoyR3ix90fEw4I6sbDxJxIm7bwe+/mQyL5zmBW/pdjiJbfHu+DE+ZmbNhQE9TwwAtJY
Ai1TJOR914pVvgHw2etex7dzvEdMwDFAJH37gsxdwxwpyRt0kHJ5mvfc+LGb11UuoN7xULoLZSJK
T1bteGxeqLw0bVdKjnivROpTTygUbxrOcqhz1hUcTmjO+RDmBxXp0xjJa3HhrXf8ud5EvyykO5zX
SGUvb9AjbV+7x1QekHXrPJyRfex94s0tGsOOJgIRExN9BG2OxcVIrHZROtUBwirJSML+WEcXIzaf
C/jCQmwSuFpMjCBE51PPkRK5FUyadJCLyGMiI84jENAG8w4ZQCvlrEmTU0MSy+Oq9jEv2mdtbRRl
WGSn9qTCPT4cqe0e/btEfxskOt59QWJAaBhhlnUMdJ2DpOlm5Hd5pxTif4orM/FMsza2iidgjWws
zfKMh6RtYZOi8G6CYkiRfnEvAO3tFD91UKhOXhxDhgcULKfF1X2fWM6N1hPdzMvh9HnwwrupkMQR
k28o2LJn8wlhVS0MY3zJpMEbaYiEaG/7ns7OUuu9gklaQ7di9NjI8YSdaX78WIe/vh7mvUD94OLu
QqtrfnThO9mLSYZQGJ8llHv4c7HJ4rfi2KN+G/5EquwttPHXqIg9fHpbOQjyFpz4okODfbZHVgpb
4hLAVa7iCC0w5q1de/7uG85RfKmeqJJXBZR/2G8Ggcn5ZHe+k0A9GsyFIw0bXJ1L+zcsAhkpZwqJ
Pxs6DE4IXJs6QVPHcFu5/J2tXHgaNWS1c16hk+HbA/QHlV7CuEZg2doIZPR/q61tdl1/AkIZw+AI
F+grA04hvjrp5cStVRQVioHcsHhzD7DnVUazj1QsAeQhuNdRCNdd4mHYCSAxPHH/g+p1B/fmZ+BC
ACdI9Q0u08uwtTGylFYlv1C5mcls5QHa7qrgQUJVsgjgmncr6AnCsXwVAu6P4u7gH+H2pj/oA9hf
JzLnz33HHWNJAf5JBpiuGnD6vlPtYmjlV8jEfwoxrQxxQfnzLORYQ0o+J+QjPyDy79JwnFQr9i8f
0zm7C/wZc5Q5mHtQlM6J8t02EEFjNaoMlK4naA8QK86htw5+THg+2oC6uQjvGvib7MugEjzgMiKJ
f+U9L3DeVL5DNoKMpBA7INkvrgdoQlLYsec5a7/qZUBDsZvWxC+CKBiFG2gpfaSW9KfNtFwsgs4g
af5/4vO/WbxF21nxwXsY71HILYZnDTb7Uow4hPPDZFQqX+YBcg6CwByHy1HaUOzs0fu8rabnHwTe
6kri4t3Ze79LVf5UZqKdCc85SIDSQmEAqgfHebZ2Y/ohecDkHPeldjrdaCpKichFopDhJ9vXS61C
4l5JD66iw9H+5vlFNJjDBTg4oG80flXxFkBply2v5rbADWU0I62HkZdcZqkzcCMOZDJGJJP5RGfD
cipQTmgzCJiT1YvBhPfzmZe43qgm/PpWYroOFDvhZKpuCUvuxIiWh671/w+jAnYHS9F+dveXvTvF
E7/e3wUsbgPjFi+eBV4DB3uzQXTU4HM82j98MGyoBJTTBr9vogcVsThEYcqVgAyLAZf3/McZMNxE
0V94sGh3dl3GgXULcqQC2+BbRMZcA8X9OLF2YpdDbQLDb5PdyPAl2AxYrHZBYGFxyENWePU5yLeD
KYEW7N7QlX6rnttkvlvl/JMwtqK3yym6F8QbEjFXMHjyoUEGfKkItJDDo4WNW5jnxVQOOIsuRsvb
XEOke5xdCaIfalwSjPW4rsnd0AniGlz4GTpx2Tk+swaNOeLlxdthZj6I2kX8/bqtpVQNdCZ2x+Kz
ubUU77PbY2nRN80JpcePzNYre5xhFUnyAO5dzdR1E4EFrr/rzrMRI8/Jsq7QcCflYkNolkoaWJnF
KLLqOEmVkLqBMnVH9r/pjZcvodryanSPwVbzCmGeUkmXBnuLLuViMxWLXqEqzEfFcGgXmg8VKt83
ztGUcSg8Gg1Xg4wvBacWNTKEKdid9G5wDM5axVRywun5WsRuHMBk6yZ7nwUdPLOWWW14VNI4Y8Oe
DQoEyAsz4F09kI3o14pf6ckiHSavRCjBQygEYIjD2Mcl+0hXqmVoWUJ+OYQlOx+PdnuxqD56ggqe
NASHhXQoe0nLVj2HcxM0QkZYNdAnK2O1Mc670FMhpXyC5ZGJBiDVwY/wv1lmrL6GTkmCvZmqyq8b
NFAneAQuzAbATnN0dIVAnXlnWF+uzb/A2Uk1Kv4+hcA8yWgnI8o/VyyYylTAec6mWY9dN2tqC/4z
xS3n3N3ALqKQptHX7VcBBX2YHmLfaQ4IwziyRA2BOZ/yaLCUDb7eZWKQ5U5Kc5X1Lk6Rv/HHvI9L
bjmBUhr+BXwbUwuDx2+irA1eILtxTPywx0nypGV7TLQgUvhL3v+de0zTdVUcfRLq8FpqlJ0gFofP
0zD4qqICt5lAfxnrI19o3gJwpRRe3k1OohGFZn0MWOT6Zg9dGiiyPoPDdOBTYFLB2Nmxqdp6MDx3
MemQEWTrYUtDkWMBQToHZewlQb2UXQVCF7OdyKWXEmuSHwxFmBt9wqExFejJtcawKjycrC3D0+sU
dZ2tEqoHug7dl4NHEDMzZV6m2A0uDt42UHBSYAm6B8mVIDXpD23ZPu+PwgtV2pUZ+wD7AO9qz/4a
jrfJv2y84YJJ4X/zdOrDQ9542VMwgPlLvzjZKphoTrdn0wV3h4uK4BRs1tpJ4b1eeAGN4aSYHnRd
17CoRlCn32PEe++Lw44CmnFW/c7cfOLCDm2bftzo/Bc1WJvs4HsasE26VVdAmpxkgpSvmJ9pBY+6
5MICDI01P/pbPkiCF95ZTOUwRy6cuLMTSW7zBfLn3637PubPtXjNpduGqdIW/ZW1xfJXL/bNYrxv
8Hz3Zjw+ilN2ixIGLqNKjGJJ0+RHx8HxwwYlNItuLiqulrPtJcLyS25H27r2NNN0ecU5Z7+fcc6c
XUA7Hl7oP++qhppnM08XwGEY1azN26XDzK16aLejLa/ti0xoE5Y/vjyObFmpfKB5W44Y+9gZ+rEb
6a4IHaQeLeD1ltXsCUhMeZpReGPXJr4egNIEbHlWgeTB4ollOdRd3oWRH1aKo1L5T8YKd9zEyxCC
PP+9IfnRQkMaXajNefFk3L3IwxOGH1PQ9WhZjr2yOB9m6sPFYIQoyoPwvZRSOY8MA8yWyeezf9kk
Nl+07kpt4aFVPZpz90XTh8WKN0e48xIhYxXM9Yd/iMPU1gGN11lnHX4LhwIQSkBTJDEg/oB44Vg3
bmY7SDLp5Dn3y/FIQR39A1mRpBZqzSyfjMI5dfS2Q4VVMwBbGiRHup+AJwEzQ4oEDG+3GkvPimX+
JreSICh3kR9uUNbdMfvgov/oiJZUf9WdMgaiyBXvIStIeQVzObIW5sDLDhx/zeLPqOinPnAvZuVC
5z/bw+QxCHfkNhOCKfRuZWT20YNeliUD3qaQRCZWwQzQPa+MMSJs3+1DfYma3wDUp7P9guzNPCut
aHVFBWaseL8q49yBOiUdslca+6cOkb0PWxUDQcG+ZAFCM8RySWMAJN+aubmkb8J2oQU2aP3LVoe3
YKtaDUNZnHlIwwtUcNS6gSgdvdvl77T2RY44dW10ml488Jk8jxzzZ/ftEK1CwnC3L+7Bd2N8B3eW
l/ZiBj4CuXnRiHuTYLRxjEk5rtFR4kbefUbSIpXcz7uTDaRFtY39WLaM0Eeg2HgtTYd2IIgXCEdK
1NIm5+IaP/zTDnN9LF+zZsRyFMQZCt3Xfb4sLljBhSo/BGEpdpJ6vm2Jdk3fuheD+qzQuQAmRoBx
6wrLZu/n3b5HQ+3K43t+TN02AJS82uNMN4aQp5e6wVjWZb1Op8XQZBsL3pznSOnlNQa19NiTOnYZ
287IMSodhgdDwKwjzyx13ZaOofnl7V/0jVH9ufuFNCA8rdT6XJcqtBYH26jGQIZfBmqF/BvNkilW
pc+O0BWes+j2/d8yQdKa3oCgQ0VI/0BMwtHPju69HTVik5kNOfWdag7rcp/AtAwfBkoUxndcJyJP
v39D4Scuz5kqO+GnnwGmSYCx2QVl3YKUj3SGHJdO3g5WbcYC40StAD+xp1uyK/HJdT+xVhGC+l7r
mRK6uwsWk6yFcxiuEsKxWyqFM+GIqw9WHnz0Kzpq0f2PQF4548dBUacP+ktj4o0vvC80fNSViVGv
AkMZQh1CiN0kYq1EwdsyeZbalDj1K6aUxZwzbKS3ueDgZSmF4xcNAMom2+CurnP4rT+R6O94s+9f
IQ2buzNZecZPs/yeL8iUlmVr4BkjN90O6uu16WG9ZdHatpwXzcVfsGRHeCnBQgTsPXWReUIyGDrJ
ehnPzyzSBNqrGzfa2EC5Ux9GBcw0qpF0xeGdW0x3zItpFqxkO+fvQi9rdnOkFNyfIN8Pp5Xf9eqx
f1PrFUm4k8gxQhRfOoZgw8xHARuqbl4A9jVJvX21siqQF2PoGV4iifHzUfsVtrkE1ir7akmlxyeQ
09sBwWB7RglzkKUFjbqSYq0sIaEmZlozFVZvQ5Cvi9O7DWZZnfViEQEs28fatvrISsAw5OebPjWX
MToAyeWQb4xcSwUVoJVcL4Ei8+Dl2xcrL+w9rk0k/E9mJmf/kM4zLs709Ax6o3fiZxvvxkPBMCRR
kPe+IjaYmxmrTtetj467TsDIZ3P/dzCXfbCZXAofDwHxL3fKg9S8HHVRYtG7ki9LXYhNbT/4jVq7
6XQ99PJlnrOMaYLnjwZNHgdTrU8mjkvNY9SpQebkx3xnbTnWxgOPeyMUL3Zto1SSMUlmJY9LufG1
FQSz9roTX/TqfaxT7424tBQRrki/hfpGrTK+Nv0/rAYhVLfHrn1a6v/5cZr+Nv+rTNjNMQm1Ljp1
8YkVk/ogI3/MrPoAKXFN7mSbrzD5FPQKXJ4l4ygqgHYuzXe0rwnEFkMIV49qcVVFvJTJY+Jo6R2N
rpNBWkHjnxC7PbneF7ducb4FMY83Luje0V127SooAhfEuiOyQ0IpqlyOu8gn2G7NhPqyNaZsQe09
k66YpDmaq9Q5gh4p9VfX1CT74OBjRfl1B0cK/zXglHdwj3UskFUqj4PALdtASBY7ePcutabMLpoM
XZ7Fl4QKP3ehBIzoz9J2G/+eGnSESPUDm+hwt+YjdHTPeJu2BOTkkXOllyAFZAil2U0t15cD4Hfd
BQN50XCogR06rQfHHHe7qe4QcNBhsfXQTppiRmIxfEPm9jBfw7rJv9y+P+aWlBwz2zxPbhbCgyzW
ZBwtiF7aNOhV/M6OYxm/7F2AaLknL/7ZWnf5hpqxd4gxzWW8j0EQcbqDSr4kmk/l73LVvh4/+m/7
Tz/0uv8Xvbr+HHyw1ZavDq4yqfnMhocXHF+NTOAJ+aMlJq/LvVkhB0r4AEsppL6/X2NEJWiQeysx
aL2fdc+8u4XzgEwkAaq++G4hASXxsuYnAgDH8PPU3lXln3OLiqbDSFSXcNNIN04ajdGlF4pTlBNF
+64xDlXNU2UCWWL57kLUoqOOrRLsmSBMsVFRlMURaOLdMW3nR5xU7AqAornE3PeR1XG0mEaM2EnS
B6fJ0RpXYVtRp+5op+tjtW4ZbFrTa+Di2V/T5d95Ea4oKfb245oFJvfTVEg2lwl1lw6Q2EAaDfKo
zw9IdM1Nb0ivzrrIrbpbuh7nhMnbYYrQb5JUuDRjDW/I7LkngwBVDQQppPw6J6DBLilCzKwe1co9
sgjT+yL3w8i/2Kb+adfAX/M2qSFlJv2oazizPQH+3OfJSQ65uDu0DwFRDuq3gtULyLfBN7hThEkH
7+XME2mw3uqCd3UCXOo2QH1seuR/SoaAHLWUgkdMyMhMou6ruA5lhyDxS3qdEAh3aIlSq1nQ8fVx
PFMO450kqn7OKCemR7Ega2lhRtBdurVt+0W9HxCCwUzXUYWtODABDDcxD6pKfxVNI4SXiXsX1bml
l9Xwt0ZGngE2IjcA6ibjCs9qixMoSahKBenAX7ajEe35zxGDBXRlPBmluz3LZUDOy2BHPGXsu8AU
3snTHYRHszMq0yqWgjmJp+bp2cw4UGlE2ht7Gu9zruvfvtyUUWfYbABlVKDZQS8iiI5Vkzb0fHzN
gJgT4Tck7ieO+xMs9d2mZSMYPmmQBLOzro5N6ZjXnDudM+I2d8BNBCWWzUtsWrL2NIFFj2QVkf6s
DdOHutk1DrNFRVCtzLRYwRI6p6b71z9giz74nSWAaGgiyoqfnKReA5dF9OHaixX27WsR/ezBcL8r
qr5GisIkEFxQvABdAbzD/sdYwwK3hsaEoA8CVGlX0S9BGaa5A0fe+L3HFz8fQft5vt8vmoHTH6CX
j+sebOytwXrWFcyFwoR1HEO8fzIyNawtMCt/pwLyWn2rfpol7LJvEPWeZumX8GPgIS9nrUF2Eojp
xrZLIesgojy2Vww3JC5rkulgDvKpAE1IsPr7O5T4clDg4I0JFTMGnkAXPTm40SdsnVhCX+gj9pPL
l/URq7+crK0WTvrFYi/0zyQ83NTOCZY75bcusiZK4LUdC0hCTb1GJkGCzkf/LnYdqV2FtlNa7iMD
q9qJ3PN4LVVf0tu5THc+duHU97vQlpvd4hpNI4cMzGJZmVrxg3jkyzr04Zbx4hWSr7fYW8MtrZ0y
b0qbpSOYmiBh3GIIcJEzWTyeX8ZWZVqKCB6WMh8uu3HZ5WWOLoSb4JaoCZ2OaF1d2WuHchKaZzLa
6gnZdl618V3ZSfG53cJAsCVkD38WPEFVx10s0QucAlFzax0stguXKYR2rW37ooM4MaIT9jFjNlQA
tcCC5EEIjqBq/xPBFX+Xhrt/tML2nlZupFKb63V0TFiwvvss9n65fUZW+rViCgY/iM+U9DVbL/un
kdt1qqVGgKLgfZPraKWudLoIqv+OyEy/AHx0zhYjlmUAuFgswv1BJWVv88pT+ySsq7xS53GfZeoe
R8YaykWb21zSv20CKQcYFJpRi6iGcfI6rbfSuX8VTN8RNLPtFt1KEsri5ND3Pc5un/44p6XGOpzG
jdSQ8Hz0LnqQnOWeaQJi97kut4E2yOFxDmb2cHzVkqsKgzRuVtgdYphKLEx6PeKjQq7ltAv9Xx1p
FIS5gEyiLzD+7IwAiQTiIFtVN0evIJuNljvG1byYekD/HJZisc7DclHtnt25yjEg0TbGT96F6bcj
glrwFr1zPUVnutGuAte9n6CfOk9HB64kXaxHFJWrsmYcp3aOTKRphPIGDJZWCxM7wzrCk2IJA7nK
nsN+wvKTzZ6IrAFX3ndLwcUOxDWfIrPZxtX8Ersg281c+rT9mq3grt0vJ+bj1qsuuaIMOxHKwcjV
ztbCU6kvb+I1IbBeRhfO3muQosLkmoIhw9iYR5f2Y5iHtwAMIQ0JVcIJkdQuDwvmTd/+8F42Dkmx
CH4zf3UBtnSsQK1MGqZd4XnhkTsM56EtuDJrEzuSRoGQKqJhQwS4bFu0l9TBNUnnXHKi5QTiLX/h
OKppJ4qNyScmom4iUhEDXxPnKxJGmujSZRxhOmh8injdTK8UysZqol1o9zHMN+al1IuVk7PVDlPy
Exkb7GLQGnvhjSS7p373YG6QQbZA/JYKKd4RAkAx7BRqlY/T+M7br4LELLPVJCy/lQK5llGmwiwA
TV4KcR5SIl+95NVfnRyiIQESJatguRxo9fL/AE1sK2inhrf2OLwE+ZIlSIWV0HsC3SgNBej4BC/D
pyzISxR7lo28fj1lw53Sy1hJfjf9N1rp2vPv04vCojD5h5gOoRGT7IulAvsvazRFz/4oyJ6IuAr5
SSELf7x4v6gGPczYtR+pr5efopD+fpFfoGZ5/VGvVeCgo8HE6Kf3pf5SFOhfY81PvlKYBl8bFW0/
hoLqYkcIPpyBbZpSU0/Uh8iRFlOVfsAxbl0USwt70+qswmlDxYLozfOMEizFE6v4t4X/GtXSU6O0
/VFTyZn3G71rLZ0sMwJj7CNJORY5byXmzVehpYyNqqOLTYVzh8t8jX66OT5GoldLMcVnvSW/3OHx
W0qZecD0OhujiOl3yAlQ7MyZuvwHTqht+IDNEaFjB+gfc7ty2kgDM0gX/X1u2x8GDgE1DmS9TuUy
FHCrNM4MqqjX4/UutqoHqFkYeqXgGRWGRsBHC18tXkhGpKyJPLPjS7MeGpQh3hjKx2+AwzENNt6E
x5UY/8zCDpZOpuwlpHfVS3QGEaRv+1mNNkVtn/yipWTY4HzdAhL3HqnI3NPP/Xm6fbpacYElUsX7
oXuBJn3IjEtABB12zvd2sHtsbmf4w3HXlGFhg9gFTbQE5XX+aNIr5rKF1V13r5vmqE9Vi5Q8V7X/
pKBEJQiZbMmN9VugPe88qhx8a+aHXMonlwAKcZ1+MGD+ZFsw2B2gPRIaNNGNHSR0Gt6bi2EVurwm
Yo6UhbRppG+fbVIwhkP5wEvArpPBjWE3V4UU3ksGG4siAG7txYgaB3wON5VhX1mi14Ccb7EX2s31
h4oBGSEfR1hQpG2I6XrlmD4XNXE3mIX8t19vTHM/MypsQWWHW1JtZmVWPtB3AwJJbGWigQr3KKU6
AgJYdImV0ziKPsJxvg24ggizB3yJrXzMhYLrqiehJ4kCtvH6bRM23qrLmsD4oVw4CBsuV3q5RFTK
LYRVhiDCs1BIM/FQk6r0D/pbtQEZoxwPWh/O8uQKv8B1IoUo9bWv4NK7LlolAorqVR7AupkQs/1L
RL5Eup8bp3mZZKWVRVxfQ+dwl8S3WppY6v4CFFIJT86IsvyufJ6mRHqhkV+B5RHoWJpolylt/HQO
p0d9seqOo3lL1xFCrdOZXyrqJkiMKnIfzKcFYc0DLcNyDXORts10/0qcB2HgWz0T0gbaPCyK6eTO
7Ju88mMRLejOaw8prRs7M2mMSWpOOUgquC44IAhPdpjFWukoHUsA6+0TXWIcoz4O5/3cxmyMjaXG
cbH9zpA1iMUuLKyV62wxc59wjm33d3ibwN2vBXK9hgs6pSaQ/mbojfyWcULbQTAZbq7HKwJOIgTm
0akAceIKYeE9RaSlqDc59r51GoFApmNk2OhV7hZ6JCY0KCCwafl7o2OUocfb0WCJs5k7mcn4xlJW
RaK1fUotA2ho1o1+/Cozmy2Ubqt3MvPMl/1LKakEkKXztz5tX1xSDE0lKjar8PeBwKyoVoCsEdGY
WPI9V3wYYvDDsQ5FZQlgLuWdkcRoSCU037IY7li8CorM0g/zU5tkI1IuPFT/FfCQc7Is70TsPOxY
xnZ5aCm9iLDvn8vWCWxpSjbicQ7vn+omz5WY5/yn4buGfk76CKdfpJ6BqIUgunyMYmkUlKR0/Fnt
mOK4N4TNGsDqg6znhpRX/TGpJvBIz7PYhnf9nqVdbbFAcM0L2NlrUtcBnLjPKei3myDqRdpLFy3z
PnlH/VCjdR6SnSXgPOG0RTZ3Mwy+ZaHsAfh1Jtqe4ycVu0XYukevgB6a40IXLxE5lidmSgSdtNHk
njEkP7Ox21aodOwc+7at7MWFs/0/7q83m3XnU+haDtFiy1jUtiC4np+ESpOxN8il89zirBytap6b
huoXeg//G/Wki8Spyfj1ZrSK0uAo3EXm2uOQcuaToRsmYYfPFh7xXRLei3y38blWnUUCqgpLt/95
6Dt77Cn5xNXeMe4e78eQte5MQdPOdV6UgzIG1yTkN9rNRNvKBvX8rnWdz0V6hDiLgOdRGzHwUQBs
RgS7shymJtBx4k4E8AWmK/Jt4qFi9ynr57JpTAZs/VC0+R9DBinMge3AkS+MhU3S/j0S2UkjGz3X
F9FDJ/HdSTnVBIPIAyAToehr3tn08NgJjMnqa8Y6dDnYWZ2tGdQJmXKD/V8CkHGoNYw628H4YGXN
onYmWL+/OwKyxCk3/BvRIbU87ct/xZAee5jjY8rypjI0k4cRoONAoJfVOcWGnUrZF8yCEwo6sXj5
ETUBf/uRtcuhwDjMgIKaxol3ntgbSbX8URNtHorJgELFkeJl4+HW/7UGvUEqMf6ZsF8TN2fuc/5C
/unki95g2PuGblJSwIg9Gn1x30VC0F8u0yquXq/xcRJ5C6yEYSFeVCB5RhQDVO9K6Cc8MvpBdRq5
NR+GcBF/6zSG7a4iAcFchTCA4nhT5kB9/pwgD8Q4wvBrWWrVJO63Kpua2qyU90CeAadvx5Y0cQQX
WOqS2EeB4rvLbl3IsDtCGY3L8vDQyAMfMC858fiS2H0+9Y7lTiDkBIXns/BcblAK1kgK7OyIEoTi
R2h5QZy43I+OeFaSHok5eg2VeT4Mg91KXLAne+/G+N2LOZsApyDNAPIZJ8Hxt99dSCK38UBvI7Az
ByZ/XYRbzSP9g6hDST45WuQAcozazGgJM63ZG6UrzqoZrjNzU8IlUg+Iof6FHnFSQtcvABmRjOZv
Y0N8jPA5KccJzfLD/msoUOXwr+Z7oAPnfONw6sO5qk5T7lk+b7V7Ha/6xiwdwJZRA66AAkYEpmHu
g2CD97ETG/tDr3DUbbAOy4aLu7HYs+S6NDj0HvyqvrBpvX1m5RpKefZMf6/daavVGdYQy+CtzEJV
78WToPfDDukmWB2ybJeiVVCW9ZQma7UVgHPfFIXaO0EolQQweVYZGt0r1877SIGR6ZFozyb1Uqpj
9GwspMwGnrdZ5Wn7/uruittg3cGXL2Wtdh18YFtlzYBxF0seYbUFbsmo7Q5OHPPS0Tv8kH9n3oDP
oPKspTItIn2Xko6kMQoTyMfbunwq0MglD6aB8DamjWwGIVRKOUdE5TrDq1GrOjm/8Aq1hm8mHRok
SNPttLhnt12Ui4TxwKhzIUPTjtOMXlIPEqWh93gNQAmvZaiVK62UTmsvqLZT4CGxPsa+YnG/EB44
6QgFwuhmaciM2exK6eAoBLX88kXuaut7LfudZUjq1r4MjzO91iaFgmCQllsp4lenOBk1Bkyrn6LE
qt8Zh3iTBHmX+WIAO31SMre3fmmZsF3MnUey2o6rRS8rBxDA7X7VNKPv0pZNG5RcjMeaZvgr1sFX
gG3s3vsLWJjw/ucT7gp+duPgT/wx1q0YbbbS62Mppgr5xgAJSt6xrZHgoUwPg75+hJFNq1S2MqDp
aMbZnimX6SZ+ojxHNebI8VSpriGZWz8/cshfLtPtpu8W7pa2lZ8/uw7vrzIxzoekdv1CV9eXsYxE
5l5IIiAu2NvqWlidfPwDm7rAAzcpbu2hfwaAMrI2KlyV41rhz1EJRYq6W9W4osHz8iyP0nnQ+z3i
5H1x3GqkWQsBMVxTXu4T1F64mn8VQuEjW82IYNIagSF0Q/L5ho1xo7AbOPkctav6ZsPPJusrZKkb
/85+2dhh5tvhu+OtMm3VuUlLiWx9AFhEcAlWsn7M61NYKH8UE80OlkmrV6vl0CPj7Vi5Nx8PqIHJ
32NyZTQ3YqoZjVpZPfhbiX/9CgItMeWb5FKKuBBQNDPxW9CCji8JXpeOM0VLDMMMgwv2TXkQcVj9
WY/gmsSZRwaz8bTUQSE8sVOJ4eHnVNaUyR9Ps5IJ2WoSf5dI3TicFjobnEhIyl0mcogt2Nyqw5LQ
0huEkhs1q2sIqa8oaYcQZg3F7jvCMgCjCVSfvGBz80fIV9AgoUlih4QYEalFhVA2Kco/pFh+R7AX
rmyhMahRMFUqTnTMMiHdtj11KVF/tKecqizb/n9W9GZ3BNLR2O1s2SwUsX69+Evhxu++56BBvRzt
5FmDEljeoRhCs8X+XUWP/dd7ihHX0SobbdBR5klamqCpJBJCSMyouzsEwqW/Wblr8Wu5covmNnPV
PGX4KP3KV/f4LAl1x/k51uvvDs/2aceowUy4yInNDMaLE5tL4pRSmPm2YA3Xp8UPvYRMNo+mYa5T
9yDLMfYVxpci9fenrr8Nyx2omkgw4ypPTFXB6mBpXAH8ng8uMdd6dYwD6vod4UwHqA8YoJGoy1IK
L0jFqnMl1zmfJDdlM8+jh0lEcDPbhwIDJ2Ck/1t28dw6axIzWV7kVOMa5B1D3N8lk0S61tWm4aLt
4gO7zS20fGD5uxBeKnt/7XtmReRJs6TzSVBlehJfExS9NFkUKVD9qRPMmgmF97LDL5G4Bu1+BfV0
7fesW/n2Idyo8ODlhJa7V23+Azn5L0nNksQJaa+n4R8dbG9JLs83mL3MoT8liNpLWVChgD650Kum
2k3y8tjzawqFPtUkNE4Uf/gUW/0OV4clJKE1x/YzLo9yyG9+OPGHWKeyhlIdRMf6qBhNKLs6OP3C
z/G+ihwYNRPn6d+uYug785FIfVrT0eoTsrf1sf4NGwj0V/uiIMgyKfmFdVy/YgI+hJ6ZKf0DO/Vh
RCMy47AgerSOq3eCwq8TVjPNggQ/rY/remts5tsU9gF6K7VhqsopUQak1Q4bDLgjPK49nNYNtc9Y
yvM+3AUX9GNELD8vkr/n1Os98sqhEwEHqBjKN07cuNrJJW8pmgNPi8MONfEg7mIU1Fi+r3lIl+ss
Q/bdKWV55NUyoUbX+xKbQmBKiD47rprvzj+IgQrzXS4L50mAMzHD93pmDLOiS7YzG/myeQEjx1ts
0ktYOfkAVRFVixSMvCH/PyY87310+/8cZ5idbsYY5pVj2S8HXlxPKvbNf6MR7gDzQhg29gBU1CWk
EOH0O6fTQKDBlvhlj+Z62CJxLCeL7kX2Xi7J6t+jyhJSObeNOXWlAsLz95mvTXAGEyM1fOE7nO4a
9ny18uMj7IlMjhNJmRiXCBjzTt5RylxdrXr5pBtFlDMJ51avsQxPEs63D1Wxsqm4EHKERkWxjgw8
IJ50Df7ms+oIwS5zQnj73LJki/q/cE3E/Yf8snv9JYD7oaAh3kZ/XGQPIBplxGSDRAxxuSnFX/TR
m4DctFOy5i0QK97BAan5lAAJaxinVd/dWUM2pfICxnYoC+r1kBuAgZvlrBTlLAIZ/tr8nvYTMSnD
OaZWi0W+lHJm6KCFJDjxlKbIl6w4u27deodhMxpppyMrqgNfMfIxTtzQazp95HWlxN4WapH9dI00
gmkZOPMSOVOQKvHKyFs43jAtjcgEua0Utk5C7JLEmq7Xa8IUYRAtWJ6NL+uEk+yQsNUtd8zY7YDR
QE1wvwyCBnEU+qxwHtdXSod40kdReqbmhpuWh0VmTEecvS45MqBoi7vPFFMm0f4Iem7s/ILJtE2K
uTJzgUyov1b8H+c49+daoUE8N4+AFdhOem9ax83q6DdJYBDCQP63OA4pN8RJZEMcRlqa5pTyqTBp
vsVPBPsAr+LsV8KkMUVBurL4zoJKbr6EHly6X/SW5CwlRAZcvbytcoth01PZ0MrMaRPXoobqDeuy
uevjJs6vxoiCakvv2AqGAxn04QNtrl4Kywr9KCWNgREuujsNpwy+T0ZWhlntchtVdgiJDBjDF5CZ
DvFQEJ0H7ca56pw0OJZZGJ6TkutR9SeFUFHuR8DB4IaHi3wWlmPWxlUnKtrPMXFAfYw9/koL7JWY
+YFMKYfi0QEdGLa0SBpY1052F6Rxy9bzRGE0k2u/1vPC+0rp1j3xK6F6/18SWXEfHbLqpxw6AVPH
YwpMV4B6N2m0N48Ou7ghR+CSBOO0nf6ehZc7qX2bhGgywbooOqzG8dlUg3b9lnX3INvQ3N3MYPAB
TjA8d/vizwZy70pK9hgjEPY5I6WZfoMA9+4LNca6xDdeUnSlk6pi7yHsM4elU5BDpC0WidgBWBsr
5C8K0wwmJcTlxY8vmP5QVkegu878PXMYTRMfy/COadpkfckSQUA+IkYJGDMDJBQ7r6pWRGNKri/3
zt2Wq1nu/stD7T29FhgF8ej2ptADsUwWOhV+Y+5r2YwVxR3Nv0/WVkCDl1nFQqYfAsnT6FKPrlw1
uNd42dQh6pJuMu84n4ODbTbQ+5QUUjbmm1GEmeKuD3UNXK3p4VhP2hEjcBf30aI0InqJtUBo42ll
FXX7cmzKpoWiuOOYMN2UQN2vP65wRenMk0uUgsl2Ix9pdeyrJif3ExkVZyavuEynRACd8XQO8q1q
izHblFXgyspxwfMPRwJoqNmTMknThPRxL7b20rdoI75xTvy+LW2T5opOLoyNUWl8sJ6zzGx3P3Tb
SwPe4iNBiS9CXUu94Q70Rsc+eH0DZuZ6QfXBdw0cATMus9uQJ8UNO3N1/vzUtY6SW9ZeSIfWA563
NyK+ostsZs/g9LCHRuzC6SN2PJqsSzMm5N+zl/tiKwRRKr3nqp8TWxnuXuabB3q3neNcLplVMldO
1WZiRZCUIWPhfGd++B41+xZYhKagvaETUPyck99P4ZcnAeaF+29lsUlSjUbFcIgnlczBfuKCPfVP
GzPxWRe25hSkFFpEYYBNz9sr8+1jOczNpklai5MbrrVqqvtQxhBqZCNj61LcMINo+jJuDWThOEu8
X4ZdEoB9vdK2zinMSS6Psg0SdSlOuKdWV9SQQ2K12LfDXmQqGVt9gkYxH5GFOynM7eq3UW0LjCk2
WirkRLxtv5QGHikR1yE0dZyymQjj2NWPdoc5eSPA1ucfrttj6peY8xeN953P1tgct5Fq+Bq2z6NK
dxl/eE+rLEgC5ILkcQryRjwbUtY3HmLlJOQfuk4wVn9Jz4EFugfQhdnaiJ0HLnOfSvTcRYsa4+ii
s8W0sRfppqDfa1xVx6bgnfOftTO8v6Pekqho4v2/A3VXnf2LRit1ymVLdC6XDuKcka6Jy7n4nxhQ
9K9+Dia3HvcCRu2U2tw14XIhneFoeDnWhiSm7PJYTksqQHS1DKdtO3+8OtuSZzLNWTKivT2aL5cU
J9d6YpTnXOym2551K/4fTOd58/H2s7Tp4z3fyyJL3Dp7Sc1Xu3hzb7304gw4aHDttii+avxAxssl
3ZdOmrAa5C3Bo/v3TrkabOGYhoHrjdU3Aa2JKVuvbpKfO3s1XTQ7VhhYmXu0D5i97b1xWWmoiD9B
EanSPUZbgJAuXHFNgxyfgGRZlTGtod8i3Es6V0KiDVmJatKxfPG+yMC1g+rJhkll4scAnQ6JZ5wR
g1QdYDxF4TKMP9useMZUtPD6CSBVInkgiXKKKSI67ohqcl07CF4Ed3DLxpOvHjbVXnvDkABo5nP4
Acy2bOsCHV8K/mid4n2GAdF/e4COdArLWhhf4AgL+jeYqphg03WOiAe0exXqi8Pgn1NO6YH7aL7v
8fLMNd5NWl/0TigCZgW8enZUPq2UNr5lGGApEPU92s/X4hJBIqh5PYcrV5iWladInhY1AXKv1yMg
zaRO707+Ks7VQA99HZFcHldQcg02QNvDN7sQJWYBxexssLMDASo/esPIqEwOCz+Zd+gfx5uN0XCE
4AHOT0syYivP0OSBeRnsgFgYeN2fIOh89vWdb6szu+3d0e0UlUQ7FG+zydRnmDdGgOlTa8fOv2Ht
PMmY8jh6BGBQfh6SHyGImyggpcrmz3w/BByMWOv/8wVeKCCCP2DJnb8UarhfXLnAxf+LRo/b6yaD
iQH+27WpPcOplAeL7hQMyxAkpRoIk4Fg4uhO1mJs5AfPGfXgCsppSA5YVy7kngLunip+ewmrMLyV
Vec9HVIgN1x2mMgxUs4Gs9WxwX2+4894GULzzwOLVKy5SF4wAyagcucN4Bi9uVn7L9P22onTGONu
IJbxACPo7Q0iBkUukAI9OaxI5ZoFrGVJiCMYTOdKFoGy5ikQpDO5+veyYV3GtqDmHw+JUb3VdgQW
c3gsuaHpQvjNu8LDRdKHYfied2s4ecfZvpqiJz7gutqfv/cL64c6ZuzW2JADUhe8/BttR410Z8lf
ZxypC9kPkw0eDf6UQdGpELBkt8n8opH6yXB0IKEKfgRAwoYPyOofUyEPPHEy8K7Pxnz+wJfjE7Uc
55++5MQb8kZbfuLS/XFQl7hQLg58s8WvcO5+y9Ye8frTj1EQfJCntZ40BQwUDwyRJfNijWVAKcEW
CyPmJ7ZNoJzcl9sR6x5OY8KhV7oE8axsOUb6JOtgnvmeRQKPCwcKJo+d1NCBIJuPxbGuG0U1+ADo
WzYXd8pWuMbSxqkJvdCK2AWWxJtoU+x6yiJxUcKHJk1k4xQLhAV1iUIaeoHwxSmxuu+VAM/ZeH0I
GA44pbQ4WP5V4SCnJ/ENzsNse1oUxr2/Y8AqoVP2r5PIh/TX5Zhr+RtjsNw/XmfppnaIgVC/BfZX
t/T7NRTVCBY+iIERQjq6pteND+usgYjtnQHRyGRLxdKodkVftjQwnENe5FtrGFV+R+7IOU10zphq
PNYr98I1PWx/LKAjBfA+CY/jCEhlCFB8iirAyTopv0FRINZ+KTO2dyzBeqw8AlrNj1iU08sunOKi
1NQP6mDkiiJdzRJL47o4jP+Xj369BcwNQ0aCJ73t0w8xmJC9JWSsHN99byKTXG55j4m2209pC0Ip
wvaS6bPGku8B07XI9xOqZ41zyQl16UXGCc/sd9anQXXr6WHvk4heJEa2e1MbVsZHy8bXa12SVwfB
/MtX/JupbSv0BHsWzUglS88wWqMI4WQzIQAZ/sLXIGTWAFSrNlb+OHZ6CFtqtgeFZ0AgYXvqFilL
XSxJv85NtQffIeAzT3+/GYRay9Tau34WQ9TzAlvgIhNoFtEyHpB2vYLiFuOIPfWKHL4IWmMSxHsz
d0pTjpCH9UPuep8lP2kDocUD3a6OA9Z2PfnWWiWz0PY8DVcLiP4IIxNzJ74Rsgypkktm3EG7Q+My
q2+G0lVDLR/CqadTgKLiQd/Pu+1PBNTcDs4wMMwuWeEVp4F2gb/LBNbDs6DjSR2nu5Ylm3KvKuhE
rsRcICrYlV39INakb4SYcTlQ7vMohxwaHkmTyKZf2OI/7pMFa0YNZ2OD+yoiz4ToSnOn3iH9iu9C
9a8L4DDTYuaVJKvekUXuLbbukwLSXkDCsZziqKxqTxCsC2i8ZvL1xi0xJAkWtIOYXGsB0sypt2CO
ywLU0qKRbh3hKlsOiXKvwW2a62D7PG7T8bcr5orqg01Hr5e9O0MChkX/J/oF882lJRjwbpv3Jjf/
cgx+YgKcUWrKXQjMuicN5odX7GECqsyWVgH6wLdZJZ4aDfY6UefaLdregQFL+c2pWJ03XBeEV+ZM
1zgP0GchCA+tyDYtpMsPNMYUCKPoKFQfpktsAvaUtJE08XBJZEd7SXfnjlJXY7ndNDwZTVoRqars
jsw6vltKz7PWLs2MS+3JK2u1Md+suk0jCqntysJ1ITSNYCKwpbIXfzvzdhymg1dIopQ5TXN32eSu
wA8prt20JVyznqcSLVhL/4Kmq/1CqoOxHFpE8HpSMLHbUrIUtVfMRxBeTt4aXQiy2efn5mF40GiD
SlNgZEmDvWdrdEycdpB1JsGePKVNhxx2VrXdoh4/9WCGUIgr/ny88M1r1+c3Fm1HHPGZJ76ugjAI
X0/m3NFNDBkzL7fxiXVO0czEJBsNEZ7sRxNssic4iDgoNiFyAEg9YovCCn2+EvA9Z3xWC2LPB+sj
vUnHdo+epFAnlVvTpOSuXBXjQbXLFbn1VSZ0wYFjxqjSa6uQVRAyVOUiPS9VgVmh/qY6jELnqA3p
4T4jL11215cAnR0vZZj8DrM8q/b8KiGCL9+ExuU7f9zhgJdbNWIR0Tdv81pzGrbC4KwkLYKk+FC0
LR/fcLbyQ53ALvN7wQXKAn1Iq5iTm5zguzzYhiJMHejr2hkYuXLvuJejiqexz6HHcOaYzNlZQ/7T
fF4u3gV6KNIhYpZP2aGDMCcLvv3rusHXGcrTuDq/nWcqi2gYvtI9buXckaXbydhzi1GDOqCAQVLd
Gc9nfYwTwuBktNb8mMnB1o7APBKc8be55FlUB8JWSMqCYvBIwsX+/yP2e3tkrOVBubvK3kjaDTGX
6aPLcmsRHuL1AmwJdvrObJ0gl/zF/HMU+qp/YbrKCR94nPitA/CHRcQ06fQhmMvpe19Bz/SSVhPa
K08QsHgit/LEBHT6JGUJcbGZgsRPtvxCrSy9SN0I6ah5zuBVfWgWkSHKzfFV2iN6hsgezbiH/369
1QINxuRQ7tYIHMyWlhqdXofbHpj+t7cYCee3l+fF4i6UoUuuMSJ+7dQQuG2ZKbg511S2lTy9AZVx
gzDwkGhPHxQenV6MrGrBw3+FdjPXA6OvlDCR1wRvNvrfauxtICblt02fSzU9qAe/DwKEbg14jwfV
+Wc/nMrJllK1L2U3+bEUK83mcv5KS7JYfeaQFXPJS0EPo2P9E917F6FNynLKh267r8yRof9cZ7vl
dxgTalaJhdf9YUoFbJoQzUEbpv6gF3dLJYAti8wuj1VrbvvzybNgoS+8KsQ7qabWweJUL1UxvgI9
U2UaHlHcDxCdGXIliH7jLnYRAHKAi9MvJeeHPKuCDIxVawpB9AmJmUUw0x9lDAO99131tLsUyjpI
rNhVN+mYQ0G8P4TAlK1JTZ2GomWgjv5v4OTg15NwYYTWvWWD4H6SI2BxX0BUOE4cp/vIIQtYkseO
h4z3yCKPnRLfW2ErqHoHTXk6Cy6KFKydFUap4bb5efvWoHPcRlqBuIQYbJw9sUsJytN+KndzQpfR
Ov3XdWZtI67tzZkXPdPB2g0YK8FHfSvlCObi3bNFQ+nupe+rPbGctYVG/i3RC8raWBEjkA4tCPK8
rhSUjvP/JqROxJtjfToH3kCpHxIuWBbmHAg3E0xIdo+TVWOFppo1wfSloIDOklNGsBAkPO/yM1k8
YwwDQEl0ivibGnnfstMuZykUCPERoPwJSFHQ1ww1FVCp3wJHL3glC6tH1Esn8vxGRwu74sDCnFqm
i1f+EFZJQsjmY/YU5Fqz4CPsLYxvaJlPDkJ3MlITCs5NOQYvboSOmut4K1KROrsQctYVlCZ+GF4+
WgDQ48azq61dqOAWCpXpnEZVmhvQUBU6/xOY6puKtNSRLFsS8/x97QSHAP4mVosJBQ/OemouckBk
Abv2UBQ9TCxAhurYO6FRJlYqPEdcp7gFQOCAylJyvgdEq4YCnaVWPwLXY2cPYH3h2WJbKAeb9Uik
ig315Qcv3itgurvRozCnXqVsK5ltxaigkHGtYVOqDuW62AkuB/PoJp45f1pAwnk76/rDfgYJdoUD
4htXesd7LQMEyKDfLA6yWXg3AJJ2wHcMAn5chlPQp5EN/p2n4Q/+98ak3r/aohFrhQHxIXbR47ZM
xOebLxdlTaVf+USIj1A13ITmVpN6Jh3X3YxFmtldQ4YqrjZWEvVnv8c6Y1vAYpnyxy2MCKeYyS60
hzev5UwUXlSofzvRPHTkiEBF1uRyUlX+jeuwT0ClmYJeE9vY9yXOShf5mxU01QOVcGg+rm8+lMwq
DQ1gAQA2bCHi5zhqbblyandjjPTp2gKGqya2JR98Rr/SG52ZMDDXyXS3PnvCKHCLdfNC0Ed8cXdk
qEKF2VPowwHwx6DdnJbk8V1FJv2WHIbQmqWbYLltXKLygOFDrFUh008vTVZ7ixUl52nrzKJj3L+S
vvKoYb2mPFO5spZsZRlA53/oaornMMwwioJNZiRM0qAZuiCqHUKstxIrlqnANAvt/rHPmopPnKj7
9zgl01+KRJeumiUqX+tPFCwhzn4NVlLakQcmbou97JUwsTajUeIjMqmHs223WNA8aLZzOyLGRO15
MSkGqUrtHw733yUy0bjiXMl2Lz4Fj6QfccGO7keoA83z1kNhbdSgcIDxRLchdEYnSFqdTVse+WWd
tr4aTIMFa/ZADDNIWLkXFbYK8TXER82hrMp1mLc5lkyqp3YPPKb/fL2TvLu4n6omtRExFH4IfGkW
oCGbO7jmmoztBjmLJVuxt7hYU3E7RrB2Xd9f+3NsdaI+FTTZZudyt1WnAcVynBjJuYDrIgYPBDkm
z72MMi7+IU9pl9MxiitqKaXg5utFy5Om2cQzawOMDvYoais2QyZE3221FK4v706WRdYB+79nZu9H
4mYALk+8fNFRaeA5xifX/wHdvrv6HgE1oAIX8E4C0eJQmCgNIT9U22WuNuQVCW018m4yUB6vMxnq
EwGbgcMoqBxQ0lCt0YLCEVCzD/m9UY9NdJtkRrQBf7ecID80+IXQOFwKuAAKYnJzigLLKSfssmYt
1/jXFPd/J4bVYVeoy0GHP2MQuJoSRE7qwUWa6PqiGbeNUpGnyBGfheUcCoR3xFL88HeAOoNFzeEj
Bt50slEqYsddsyrfc2A29khMu2wge8FJjaDYYWvrhGjQcikEBzq6p/5m7W+26QauFLUyVF+IrPxj
rPzzHUFcKUtiaTvtldpKBuBMpQEfoCTPo5Fe3JIOQ4409BJlly03gpjIORWMIfO5OW0BdIGKfLHs
DtmCVYXLsXMvKOBKl+zAO4mvdNceVuh4LhYUuZWsOQ5f20lYmeaxP1/cWp+Po5vUVDwzwCeytYxB
POrgVFDDYwKpZpzhSd/ugXQyWagdgIErDQj4eQXkhk9LRp0xOW1rxf1H+0uAzEYeBay39kuGMRGi
9eYS6fVAvFQ3BM5vLdf+rQJBhXNfSVTpwMzi3gPa6SdIhfSiBdAhdU/O+ASZAsW+q3mbzf1fYfej
CP+12ypdEj5WwrkhKSsMWkKj9VpRiAuC8FXWD/ym8FLiPKqlyT2uI9wmixbN+3mz+ADOD9R5uavA
XBjxwZ3hPUgAbM2/wENJHHph3l31HKxZMxa5WBg8xrxpAZM8deKxifl1vKTusJ1F+Aeugd0HtE2v
M0mqkweDPnquC6YNTQ+hFrmTwCFET01Us4CsnnrjflsSQUcFK8Z3fsyENql1zU8P8lSJrXb7bZX6
ZGYgbEr1Hl3jZsgW+1yJsJaoaBrX7k9aFJHcTR91f0N/QegqYIAGEfKsYw+oPiDIf2Rxa/S2f271
oO8RylKjSKMeZ4rQdyzlf2nt9j85Rle9oohNUYmGWUSeHGUND0rXTHN2PzufYXOtFW1q9EYN/QpP
GMQG52kaVw5mS2xKp3tqROF023BqxAQbHyb3GUN7aQ/JFmaX/ARxpoPGOJRF++hoaRJYgcLR0XwW
V5xNjsu0elVimCif3aPX92sAlZF6wQ9m2Jb8KMbcHwYZuugHwTKviE08uN02XUkdBn1ZMODN+yYT
e7Erysdmrra0kGqoP4rNO1pEbGVavGO6OkBYDi2QnwrHRXeYjckFnPiiCszM0tDS6gCVPLr3poeH
POFwYWxzNV/BF6PcR8yi8TtKcE2WHhV8zEkj6G4ricnXV/xCbrj2cCy2WGmlY07HuZOiXi5L5NTt
+RAtUdHOv5jUd2bzgDjGRChZZsFxsuLb09z6pVl+u01GLCJkxYYu5BQ88ss+oIkA+E1hVG/iLZMC
rWkJiSVSCTUPVO3SJvBgtjiS/VN+vVQJcTnCbEP8EfFLCCo6wzzsilm3BIWPvBcpGWG4z1qDc6ba
qCmRZnAu8q0bX1fT9y0tjd/n2sYbKuDuaxyl+Gt6j4syW1KAbsE3aRw/OPml3t9BLhH4J/8A/YZn
SDKi0K9gFtLZctwu28l0gy8oMAPliYx+gxx2diUBt40Yd2Gsi0ACvbzxAeI1xq8bHxhsYYLeD79P
xVd2eAchE7uDk4JGKwfswIhXDBEbTmD7yVhmRUx1BBXssk/PGPZaPgyen9jgQ+E96saeCBVTcqGw
48hbH6GZuc75837VHPvq+x1ONG4h9CcD/+98a0WjyPa+H2PiYQOtWYh8ADG/xUz51mBgINwtQMbA
dpRteJxfCzpCwcAVwfYYU2at2YQZTY2g0yIGakoghyKRsaIrKSc/eycyDlF5T5Y1TW8LYz+imgyd
nMIQ6S8y9wGcoIZH5Kl9lFsQ49h+JjESS6UNC1Oy/H5oPJWRR9L9jcakXcX4wPZLbkiOPcDgfxuj
XbgCl1pb729k0cIxc0PQnlvtvJDp3CHe5tqGFyzxIlD1MJ5eFAB5r0dm7ZRhVOQKZN3cB+J9K7FS
t4mkbFzq7Ew53t9pKaCINzXThelEQJ7yqzAMo36TznfqvHc/sd9D6SORRTBcb0jHCIJSxHJAPpsi
e9zX2w14kfR3ocnT8T3Vmlh82b6TwQoWXARx+c/jJ5pHaSEX63ledkVX3t1pb/otVUPUEY7VodXy
DV4ud+tQyVnBNeJZm07iQpk7gUJIAQ8WvnvylcSsmDakMcaP6hvLGV+ZJMhG+idF7QEoDLSbqxml
tf6GNOiUdA0yFH3LBRTklUX0HjEkhlfz2IxNxOpHufBX6Ve6EpDxhhkZQuH+6zc7sjHt9fSWKvM+
xLqMHaZMMs4TzOiBwSZ2PaEdnPoJB90Hwoi+HMjtBCUNNtXumt0Hre/t1v5hgouRlOSmi04C6S5d
IInNA3Hl2/7zyD+2unQPVdALQjjOmsZP4p6lBm04NqcBrp5zk2YPlu/9+v8pBEcERQQ7PFEJjkws
f7HL+tMb84KrXcCKoNsr9ZUa9ezZKWnq6m4jt6p7h599piyZDsD3ssmDhRb5eu2g+DNxuXHn7yd6
n6+oYy81XH/EoGWDnIMafEVJNJgzju9dzg1BjzekKvebSIv/8MtZClioLRhlLhfX6p6oItaMMEs2
2J50HiexzkGXogsMjgl6SQaES6e0voop5GVu+2R3dUq9/uiyny7KqxVwD3kGolq7MUo8Fs7R7f+0
rpbrX7Qv6FLlQHttbSCZUPjJlXMEpDF1RaxmIrZWXQI8wMhpK9prmO8QckPhbGsN9voBInEEqqsM
QV6FhcqJ7wjeI+lyUuc3DbqFWWlXVzfKh8h+F2QkZWOSva3nd8YafOZRg+b+3UzDkiOGDPLXRB8k
tVe23J4E7eIcg7QV1DMsO0Jgl7TN5PfzJ3GvMYJOQNeFlzhIUxi0k7YkaxuDQ5h8VViFbgSHij4d
ZzT0CkaIoTBmwinaKnfYtLpUX7dN8XLxnGcsM2VQk1uidUoozmgUMJpOyBMlMmhAbvUhNNWxNzXE
VmIkwVflCoQzTkv74Z7YSEkqc1GQzTQEQsh57tnPcAdT1i56Jzoc0xu9NK+VRCo8JFoO6783Zg4h
G3Cp4Jj1vOphONdak5CgNj9gx8IXyPq8O0QjiD+hBfXK7Zdc894OYooLi07+bbCJWWFWBf8Y9xje
9fOWAPs7SdY+E82HzIRoPKYGjk1OXnnd7gwkIBP7j/geAwnS1IAbw//R0reKzpEKON/qyyz+Gy+x
DKyqzmyg28G9dRPgUWeYIImn4RghnFCi9kwUh920thL1ZAbsuTdmMXqYQnnuqSfZwt9raelE+JDf
w3qdC4ss4CKcSTjDEFxGPcR42HbWHoq6WoEIeNpKHxT7lnCL1ivxqAUTACMbBUWHoM/V7YOUieP4
ZfuR/k1dYoQir51xowahLhaymtSl5rfHFEEWXqmQKFW71DjHQyd7FM/3ed9KTXgj5o2Abb3ymLd6
UpWGk/Yjncq8B75GUB6hftrEVsrZ3G3EP/YCOqu3NVRF9GePZAUwCDB0kXMnlEmz0aiQxibtj7FF
BG29N7w7KJuuioRWp6vAXaepGAfiPnFcojAqjd6Vx5FC7uE6lBaBCSnpP9T0UiEw8ykt3BIxoaH/
lS5bOhrT/dlPflrg3Gl/MCONpyrNc9aXa9PgNufboZ5iNrU3RwU5WSkUSrsV6e+LqPxfu3PNANK2
CJklxHVqgdYmUNtxqXg732inFhGU6qjDmS7qo3qCNqVUM7lZ6UHok2A5sIWbTdCcDoSsLJo8OEyb
+FPLRoVht+ADo5Xf+DLUfbry//qaOjbgUVDV2/RjarjhN89hoGWh8wqotSXQfAiHlHHLFAkySoCe
RLDIhAXI08GBkFgpMYtXNHQQxuFqdu8ZFABCIH6kIYno1JOxUxMMyh6a/mvL3D3wTkAzvvJh3h3c
U+eSoyLSaL9bo8SUVt1UtY+xfAOvSoMeHds78UgynClgA034wCeP6lA+S9/t2cbk6NiEQtreqMmm
94IK4xqMkO2qCnTSz28zNxWehdMxyyRqR6pJaQCMNNvFNGJIrhqBmlk174xCbDLT/UfwPdGED5o7
ISKY36J6UQQDZmcceS4hhwVOF87dR3W0+8wzoXYjKa4sq+ho6XjdtFjhDjzJSeXbLtDSzLJ98Gfc
bFNWbG3qy8PAAhTVhdRz1gAKPh3lhq0tE6jFCeZ4nDYzcrt/AglYcDCnRHCfJ7iUnxpIKrgYRw3e
2Y5ExQVeg/VDSglicE5vubGOzwWwmmr4ZuLYTpPafafDJ9EsavBJOO3ePO9KhDLGQobUc6tpreNs
Pg2naRcKFQFP/cWLjgJzGEYft69oTTxEuwVHMLP5PUdrHs8ASmLc6Gx9PoeGXaWFgUDNGG2xKaLR
aARSdCm+nuZss2C6RLpBe7SsIzlU8dc+1Mu+D1JEZYNGUVlPb91FAvh6ZlUn/dsWkyq5lm4ux9RN
9Gw2x/qRRWGA5GFRMX2zKRD9gQBVWB8lnd04z1SMKP5iBDEvWC3Un355HmVLeYtVVULRSd1SOHpR
f+CJRJdNXoWkPy1NobQvoz8WCUgQm7HMdbsp/WVr8EuD1COvRnTA4ocdaloIwaEBqp4DTgny3E0R
h55uYv3z0WDopxqoVxSR3e2sSnkbtB8p+znOPrSl9mLF+B2HJtJobF6mOFc32s959NqaM1Jv2u1i
1KDaGGhBxt3I1El6xHUeUh8XES91gnjJYndmIT7K3tGOY1h7AH2v0B1OptFuRxl3LaaKWzpph5oH
1+cLRavvwUhlOQVdKDtqtfErg+pLjWj+zw2g7td6fEezUAJDcKVpSVGx2wu7RDVsm2skF8r8M6B/
bC7lES66vHNHBaSLXRRV5rL1E27tzyLgq/1V9DKzASpyf3JD1xYdPLPp3RVbx3ueh01xmp+ACqtl
fZwtU96Q5yM12I0NL5oavqRgpBRSHdUyEtXeakHk+KMTyLRXW0YbVUjHTrBaOUCIDtTOVk+gXq9J
7E3hcgfHkIHj7YbB4SCMJJWUOAs548WmH+Z1/x5HgvIi+tgqw5fb0UVV/vqOxwlNlvbP0EtRksyE
+AqFPkoKY/NLMTYkvC0pMaQ2mj7HsbSJkgu5E5CLuEY1aQFDQ+swwOg81jr4WAswcSBRFv6Ze4DT
aDdkZmCRAOFuypIZHF3/I+PcSK2niNXjMRb2nliUf2Tq39yq6H45x/Smh+RTjiIQqwPpxzoy4S3G
m9DqaNh9vjp6FON6AB7qZigTZGwJpXSNV61OoAF5O6TuUgTImSfgnzm3r7u6AFXe/axrzb1sWW6/
PngiqmXCbPw3L+HtoeDPq02GHuMnuyHNwIkMYwp8fCwto38Dsum/tNnu7xU1FfzY88wqRZbgKnb3
xywddVeHTgx+Wk4g7yQquS1UAc8jvAYurHH/uueqbycmsM6AxmD6aOhekI4Kpgws8Dp3/Yl89Jnc
Y2dt3JwheSDBbhh397ETTWMGCDUFwpmYyyuMwzlVR3LwR0fICDQNwwfiku+hRje4uKZr8LQFB4gy
0TMtA+vYD0O/yzeCYh2pMAKs/MiCf6yBIZMe0y13OnvYT7Fpr6NYQ5cpu2YtaLiNwSBlGZuMmWWu
9JjdgOBL39swAc9HvPHG9iII9m7Uy1MV735HtnsPG31JaAIMcWN+vE32dIqX6nIMi5Civo2Jq1l2
5BP4IEhw2+xI7b3DvV9+2OkdGIy9OfpQRC9yTOWlGPlGlrc6t+9ZzrPPev3kUlEhXMYcbXh6m7zS
cm1NgRxlM6xLmvxT6pZMgOUVfeBN7hVHcGQSj+5j57fZ+emaxG3zq9AN11sHKE007ZtDpCRZO9r/
8jJzaxoxdOFDKENhCSvLWhAS1D25cnNWJBOhOvGLAm4/seDa4RB6e2uMNWUzDaQpzwq2VlVZ0D6n
zmp53sfR8WDQt2Hp+ToWOXW8MGrROj7jGcQxFFlaHrQVprYcQ0zjjgiIeZsqxXq4c0cqMYlBI3U1
bfk5NTz4s7wo80CiuYfazxsgyDm5DPF0nnVqm5rcNkd2FQeTSykf+dnqimcpuYztyRSwRBi4Vqqk
YCjvaF8hxm23gDADGrk0hnxbHgCe6z+U4FjYujL4/h78Y3FWM+DDl/HvLoHSVNue84DntGe0238h
KnIL2Id2T3tX73EFEhS8afAUbYs33urGX+QTwU3YvEftsWa2E9t4SfV0ShJKkv10eNtXnXjYUDLL
udXFKJS4gz27r3FZSN4ER5igC2KlQrwONSr5jyy8zIhGDt+25i23dPx9KYcTrq9QsXWJxxBeQlsU
9GmGdN9tituey18fz7U+bBlsV84InAjJus6WqIoYeaZVGvbIIXV/IFtjsB5Ctqli0d/rRYU3zuI8
EnhXtuL3CR9/FcIdp3Nmq/OiPqmM3qkhmomwR2JHFi77yLoIeGTp2MseET72uzA4Q4SYxolMFwkI
5nC6fNIaIEjv2hmDgaikp3yPkWLBKbKNx3AY0Fe9IU/Hy1KSsEoPll8KMpPBGS7091gYYinRYwgE
kmjBUZsNIhSle2dR/SKKvsHiiIpBHDPCEmeSTj4VQXJmKTxX3cCjz860xqpC8BI+J6BaMVZknr2k
RXtVpPCO8nUDMTvHVM8IH/s95EFT2Zjf39gcdaRDIW1tEVh/486z4Fye4o8e9tsSo31jhM/kRoEF
0N7nImk//uhXnUERf7kfQievKZ260Ntkb/TZNcIQlwFkBGxdKn+aNYv2tdp7wqGF+eHLnON3yLZz
5j9VpxY1iRepofUveaAmYtRVhfCAHn2FAnWwc/ADStYRjqUaslsmyycbgE7p/p3x5+O4OWYGA1Bf
6mZQIp+lSwEJP6c6xdSCIZaoQxy5D5HoaosBuLJN4NxAnVeJ8dPQpyBR4MPaH09x6eJZCT6ZaoOx
zuwJnFcQ1z4acxZhfotPaG8MMoFM+aEb7pJg+6KbKAGQwvSsuKY6bVCk62leiw6J47aIZGCOtwLc
dekXN41u1Kjoz4P/cbctFMBcG8efWTK5CibK0NA0VGY=
`protect end_protected
