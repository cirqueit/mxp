`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
xcTmviRY0OUSQgXGX5U6N0qgNIRWdMu9rKgrBdzg0MADeJlZJjR6LhRHGGOOOx2IkCrGGapyo7oR
OIoY/FsPJ6sEwdigzH3ZI9eyDyLvs91TyljQQix++nAL+MJ9ig1Q9bBa1YptpH2VsAZHp7N89xEw
md50IAdamPhPE+lGwEQEeO9pu99lXb13N3CvwBW8QTy1DkPA9WNC5O6IDHhP9CpswkULTOXtQjqG
euR+FgxQvqeLlIdf1RqJwAWjizoGUK06PgWV7UKKhJ1PwVCSTyZni7XSe3Jp6zCT8wavajvRBu5z
Hgts5IGqdusErKbqniZv/uMs+xQGx7LAlNwQL9m4nmAWALodTNj8HlfgeV96X6EkGT3e6+6nkyIM
4cDen0XDQ7RV3jJOGnthGhWYMf8cY3IRgxA+VNyn0XL+URAsmNIjEmx3i6SvikLIy4CBZHnG85av
jXm2E4udrDnU/GxseVOYniv1BWOjCxvAFcDEylftXetaHqzjvvrp+G8NSSEGA+lISIjmjd9Y3zvc
mtjE4e+nu/ACj8MbBEzPwVA/NnYAEefXsyrnx/CNu4n2SuMB6oC7PVTe70iYtHrzeJeud4VRmTbw
OGDUBvjdPKNfJAHqpVcG6OcTNMDByKQHfCC1wPAMqxrRhz7nKvk1SjKT0MiAa+kkacZpgT6t7Gpm
NeV8B8ACcMcJpYoKF57jBqx8mwAM1bZE4r0KiCvcKiScC04cFRL8rEqSZ292opKO+3mBs+wC2KC3
vVRpTnboiSV45Q/+ZbGtzH9Ja8NKFy7djHHi9NRxeQw89wAjjU+Uo1TgTGjDZ4cPjY6zw8gT303D
YGUK0tXs2zjK7Kw2Eg3xXpHPsfZXmABH1xUO4XWpBa7i6Sr4L7R4LwziIvgP/DwbQFmRBjGyROjd
Ar+j/VsGh1a4Uw+Vg65mG4vw6YKiF0iTS75/SI7OySrPs2tGI3vaIp8QUNtmkjIsDbNYdJNr2E6f
mdRM6Sskdu2TirZPBKy6hzr3Cr41WqhNRUHQrvTe8rX2uod88totH4IAiFYo0iZMEmMqHD30j6Cu
6l0UQYojBy9qDUz0rnuI1DTcGs5UUBNLFJP3ZL1+QjMH+aCyfcPAhwjXkcuMkkDeAZknA01ZQ2U3
KaWLGid+S+llLo/k0CIF57+VlxIG9sOPv6DncVR35msezVC/lBfW/lWdUlCln/zDI6R7dDTpdeMa
UPdICMM/jOZhWm6oPEtCwb1pL3qCpFz1kfKOweJFCyYCN60x+dNMHSjUAxoherk37zWpbmsW99nh
auDGnvB7RoQR2eB9wWhVbIZr64Ct0wcx6oo1T49yHp1N7W9YrlFHzjbsTfz4e+FxLWmXfG6dIk9G
9DB60nG9aBgJB/BSrjLfCuMxgpQom0DZ91aMWvRVhwnfWcImuujU/Qkb1nDjA1vGErFkXKH3VOnZ
shDz1VLBvG4WTaMiOoCu9hWEjx2qLUkPA+XF+kwnMJDaGKHBXN0IOc1rgg4CE1c+iu41A4BxwPWQ
SGW5+1Z9UNvvEx+clLYA8ecgNeqSYVvVpL32hUZNR5VzXMof8OfIKUNPaOMDVoUnjolDKNRD9wlJ
ECPtHh5DMg58vwkzDOL+BP3VcAGY2IL6LBmg85S/pOzunsyEKG5UGoDqd2NvQTzODve3t0MD3jOv
FoG+rzJBXX7H5tYC1wWD2wHUV2D27iojoZfeUxrmxIJEx8WFdqgb87+ryTvBjHxbU0Sq2ZpELEau
dlAKcgpW1yatpaIldph6b/7pMzBbSrk6e99Gg/LPtIX+NwMGQlg85S0CXapMq6dL9J4cSYKzyXFV
6q+MgEon2WqUJSe0rSo70EEMPcWNgD63PUuUullodUKxFJp4VaqVk3t1uwvzcjWwJ4qKN4Y4Q96e
KpvWv6782EEXql04yTy8L+jvgx/NmMPB4wApL19ex06q8vvmIeuG108bt/KX5pjmSnAQpee82qHI
rw2dLUY9vl/0nbmzXHpBvaN9kvd7GM6e5qYnW7PbjBVtufPbaplzWeX7y5wXKYE6dGrDuNNJutI9
hNHjsLRBl/I581Rjrl/sUiQ6ig5nJXsDannEBdxAApYPaNtBL9HHcHDf7cM1
`protect end_protected
