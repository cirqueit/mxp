XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� �%t�FxY� �-�["����Iu�=�	8E����Ԙg#�x����ϫ=��Z2����e��r���m��Qp�܇D5�^�x����H�)Q�T��Z�&1�w\ ��P�a�>;�hߺ���Hi�j�
�uZ�=�ױ�g�H ��aQ2;$����� ����f�u�[�`�b�<�G@�@nR��i�����"�մt�?�{T6�R�*�v$��:�����*>��7C4��|F�FU-��������ة�CLpmo~����vR˼��=�ul�2x7�<�Iw��!��V
I���y'X	�Uk��I��i��d��K����VZ�\)ܙM���B1��
��Z�=�����߆�-�P�D3�2��PZ�T�&жf-uzS�,H8HvWJ�Q		�̺"���bڻ�C�h�c]�����S�x�U���k����96������M���`}��6N;ـgY�ժ��"^F�'K�r�@r�ӑ�Wt*t@�vَ��Kz�)j��Bv/�>���&�O?�"�`$Ǌ��_�p	h��i��V���d[=l��ҟ����Y���&��O7��`J@lX�!9�Z�x� ��Np��?�qF��&�����UhM���,JTdXM���ʁ/��;��Щ�WS.�A|�L�|S�����г�&�B>>�/�j��K@�:DI��<Ր�˒帹��������2����0cF�#�T�	_B�2�DgQs��u��8���������	@�]
@�� 	���P��dXlxVHYEB     400     1e0z�>�� w�����q�I0��W߬4��9�wZc�M�z�I��Gn������[(J�C���[�|��];(,A1ǝ��U���9QCw�I����j2�T�/��B�\�c@�0�]`&�_��R�v���^��W�V�Qq. �l=��ky�B{�kO��-I�&N_��Ai�0����1�Sَ�{=�y�o��kax���h+Nc&�)�T�y���>��i�����
�M+��� �Sk���Ek����%��24���ER���8Ȕ���:*�k�˦l�m sGj�s��E$EXkY"�KSY6f�}��LQ
�?t�c0�D����!�2ީ�_��R��d�ER-��LԵ�xn����?E�G=�s�{�3չ?��e��0�~��Y���(`j����W��!���2����V�K�O��������]մj�<���T#E����5�f.�n��XlxVHYEB     400     1a0՚ӱM�@Uޏ=�P�ɺ���r����@ᬟ��>%�mԂ�ɍ��
l�T����&a�'O�Gs��l�2y��02B#�E�m�Pm���%�&d��>34?�Ƚ�<�a�0�R�W�$,�b8�=m��K)�m��d�<H�&}�&)��Q���Ivg5��r�¿��F��1.�xY� ���^����;��뙫�v��q�u�j�q��&$�*��D���T����c:���[��h�H^Eُʀ�t�f%: �fw�xnmGD�Z�Z���|��ǨƫE�CPݴ/��w��|���$f��mf[6*�!7r��!���]�R����x���]i��yj���LWe�>k�$61JR�.~�8W�Mu�􂯲3N��p� ��}l��9�Y��ٗ��@XlxVHYEB     400     130H{u���ꡪ�`�t+cc��x�㨆������k�%-v��4���k��UB�6�\��G�옫wu8BK)�'��d�<��� ?^�oG� �Ӟ�en�>��/.��}d��{~�<ز$)1��{��ڟ��\��Ŋ���1�s޲�>߇�y� W"�c`�t�V"�JE�þ�<�@Y��\�) |��V���ͱ����~��.�>����r�ՙ/���1*}���n)M�&v} .�̅:�
�S��r<���>�'g܎�Qx�)�@ٷ�n0�ڐ��/<��I7�W�3���|i XlxVHYEB     400     150�Sx����z�[���}�Yݩ�pHl����]���uvD?���Í�|֌���s��Ao�����%l��Q����n0�ŕ��s��W�Y�_�X�s���j��A�8NӻD!�h������]9��s;����d��K�*��n_|}O>~�Y#�����o���4q�j$�Y͖s�RF�k�R�4��;�����E{L+w����r�UEy#�9�GL&^�h�n]�E��e���{��������ۃk�O�؈qƅjH�\�m9�܄ҩ3��287��EI*|)�vi���z��MJˉT���5� (�J�>�}���%�V��ù
IXlxVHYEB     400     1a00k����iiS�3o3�_"��q�2�G�>c	ǝF�]�Oэ�o��N?!Drl���T��f��ir9�e-�{^I�ҥ#�S�?�mC���t�{CWc�W�ҵji�M拉8���\S��Ʊ�s^3����R4/��|ؙ=��M�Z�<�H�Sz�#H��|��
�<|�i�p��P�ֽ<#����Xw;oP7ⳡ�&.��L_=ߊ$�OZݍ�+P�o�9(�ihRt3JK �e��@��Mų
By�B�|�����}=�&�͋���
K���Kn���ݣ�4zib��A"=�Z�=�{��݌�X|G�lQҌ����:�~�c���E�krE�L{;��nOv>�m(�cPЈV��n��,ۍL��>�����ds�=bolb,��m7ܤ.���"T�ڤ��z�j�-Q�D��laXlxVHYEB     400     180���;4zi=d�����T�ղL|���쓾�H�x�EӞ�k���0[
Pb���&xd��[�#��6}��E:��c�?�f�aރ�7�����y�]�������&ȶ�9����q��"q2	�;��ӵ�wg�A> ���'��2!	���|����m�"�s�ȜΒU�}������aI���$�B۳`;��Έk�z�삇(�1����)�D.�a(��Hq�����_�ja6E*�hh�D��"1W��l����r��Ck�����4�(TT�ɠZj�H�\�!��qƳ��{���9 k��(�D�'S��[D.�5'W�*SB�M��=��r��>�[�����x�>�k���㠞��� ;��,뷼d�a~�XlxVHYEB     3a0     1705�Ή�?X5K�C(Sno�΁�C�U��%h��tޱ[&^3-�F���լ�VF]��JAlW} ��ټ���;��{�p�=D�N�w��-"N'Ï�؊�=l�|���}7���#�b�R�=�O�+��!�aޓd�G�ؙ厺k����yܢex�ӧ^1��`-�ES��5]q?J'����[�HH7��� �w�<|���:Dt�� b���������C�+���DS")�=B�.S�����4zjB�<�Z�������n�T�W��'�Wa�L�B2�]�w��Cl2�Q�����\���	}�B�E+t��*z�M��k���6�~��g��*���Z���M�'�7b��