XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��XV���B.�~��+�T������n��v'=&.o�`l��t`�!1wV"��e�%p������m��2���93���Pw��"B�ɥ���4(��D��d���4�a�){3#�88�.�驇VZ�_���DX�t}&��ew�P?=���`@���0�=��|DUn��J�YM�<�J	�f��0���B>�|:ԕ<$�E�Hs�=��IS��S~�7@N��u�6 (Ѓ�Y����k�fch.n%��C�_(�FuD�S�{D�|3���Һ/c֓�wb���f��,�I��>�]"���k���PۼX�~�ȟ�|C�9̚�!�C�0�Y����E �tm��	��^i���Iͬͯ��O�Ĥ ��[�?]�_����ѧ�@�M��tӷ�U})�y�g�hP�U�K0��7��(��꾑f-�dp���D�,B���*h8��E]i��f�^����%�o/��]�A�=�,�PP���*�x��҅� ���D�m�R`��r0�̢N��h����<�	�V���)s�!���
a� &������\�pEx�O{rˆ�v%2>�oq���+�G���&�뭡���`
`��F�^�~u����I��"�u����
b6�#������ـJp��P�0M��NB�F�%�G	w�9H���$hM��z3I�Q�6r�}/)�u"L�w��+]~\��s߶�r9�E�iz<�)ם�$���$ߚ]WV`-3�ai�h�r�|��$��'��ʯ��*�=I�XlxVHYEB     400     1e0桧?�Ŧy+��Zt�â���H�V�V�4xV'�ZDq�B:�m�w�u�V<^��aE�_b"��T��;��6�Ga�~#�)�<����G'�z"�aX�1����T!fz�%����8�5��,o3���a����dH�R�3���o<�$1���|b�����j�q�Pᠿ�m�g�(��MC��α�,ֵ�9>��d���p휁����^�U�Ԅ�v�0.�����k[�rw��p�;�kH�����>�ZR�r˙ſy��|<|�A���yus'[��ZC�q%�Ya�I,%P�v��˽_Ώ�zf��}��6�D{,�7��є�u�X`R��w��ė[�!rcV�&:�XD�d���Cwi��Q��l%8�Y�#lc��
͈f�/|��x� <(���Y�/c]��ξ!-��-�1��g3�e]�C,tN�C������:#���a��e9u榶�~�5�eXlxVHYEB     400     160�_BF	A��6�����Z�hH�H�!�}��蛞9?F̫|2�o�':�t��_�>�_�nK;y��b��R�%����*!#�֝���a���Ll�z��U��\�b;�	74�Չ�f��({����l���	%Ʀ���h9�YngW��hM���H�t���c@�vؘ^�W��{�D!s3@�S�H��ǂ��sƛ@�.Iv/���O�E9��7�R��Ҩ�>�]�U���n[8��u��g���]����tN?2����,��E1ĭ��MmEVU=U�Y!���0NH��F�F�P�Y����r˫��:�\�%i��e�1�*f�A�ָ)�(���:��:��XlxVHYEB      50      50�k���̳krԓ�?�(2R�5��<.Ni���b5�O�g�1\Y��hФ��$y��}aLl�n񛔈��H�q30�����£