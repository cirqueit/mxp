`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
FmBXbcqBUv2jbgQu902w9asEZ8wmfDWErnRFGliab6t/JZYC0bztEneGNb/kIe19LXNu85GrTQy8
LCcT6iWltyXnb5Tj1IPJuruYzQsUlJX6SwShrit2IYveJ+x5cNa6XoeuT2SWW0sy1EqLIKHlYVcj
SZZQ/jXjdo22AeM0MVvdKICJnBWBb9ImOLZLlKFv+LV+RdNTikzEZ3Sny8Q/LML8FnJsoIvNxtyi
BWeDnrz9UoK8PGBANTadHOEpAaN8GnFiw16mxFGDg5Pu9rVBgjlWkBMMkTs0O+xJDrjbI3FAR5K3
ymchmwU3cuX5plgTw7EOrUYQSMQRTEJOjkDUUDErNv2xsFT5VLn7iPJLTI/P98gCnN69ygrKzCDR
kv3h7mrfZKDNSDRDDAfo8YmKBi0U4ho1almb04YlmfN3IoMxEuhiQFAb45W8iQSlLI2CWetzL2U4
eNO/ILWDmHmUFD/0d0wKqRikrYnp6KkqKXv5cVt2/QgmnkwTb3dWKx3MyXgKVRYpqy7u6JMIXs+O
Ya3PfF5J+rbfyHUoLhjmHbHUSuJPebbo/zuKofLzHGjJVnK5PR35vlNLkHkVxT6FJgTuLeFsSITm
OFSRInQjYnVkHCzbNKnQfAiv/akB5jHyyExO2OuAec2nZLs9Galip3GUFk2zGMU8t68Mfod6/Ckn
Vka78StgwLnaJsXTFE4lTXwdxmNqGq1TcOA5XVnBYYiKHp2UBaFhzQ1Azgso0UfI3+gaMk33B2na
epwqJVEG7oPODMBkVQ7yxC5xCFhezzwFGWL2ktrX8ZrKqOzbvMZlaBWabWsKyRdpr+vsbboPEcW7
VyOcacvj4eRKyjcWrPQ8qv3udJDkdt02VYnSzLzEtX27zyR7xYKPxiapMYm66OY+Y3yfpKBhhzBR
au2K2oMx6X909a4TcEY7rsVA70abv56nP09WcbADfepjpOoSYNvNDZ9AP+mSGLYG6ulOl/nWDn8O
U3uFb1bIO+b+r/jlm9LkFyrgtuv1SFHGittRl004DVfS1d8+IoHD57m8DCh/dTHy0kmpaKNLfve2
FnILNCRxB3kjArskiUITjPFBHjNJgK0r3dwjlaav9RVaXRYN9rFrhPW8nLuFp0qxaQpaEAfjiany
Txq/rQej4r1rKo7OCh/yZrKL7hjSW+jpBkqODFoyb6DfKYd9q+/4wntAQ0ePrySd022DHxZTZ1h9
nyf6AVdYhL9pMVl2SHXR7rhAZsiwv2vDF7DmEeZLsfNjD1I1I6dgNqJVtPHpfJjSiktyFsMGXhN+
DX51uc5XKeDovUtWz2FvoGzpWo6qpFtwdAN989MdxrIWN9Hyn20wFkdBksGLfLrETvyj6MBsHusG
iFyzPWo9CcrAXbEAAkCij643wXShWhSK9/s/ccDhjWqp//uwrdPX0fnncaXYpwkbxa4m2pyVluqM
6Szmw2VPZ8MmakeChfYtxR4GB6BlE4TWo5JakMTZHt2ZKPKaQyjbL+sL0J0CFA7bE0Q5KQ/CT/mu
hE8NKpQkEY+elkdS7qXpTdVTzMHBXUP1SV44GwY/qAGp+HJ3HAJ/+jnxtPbBIoMp1QbGqDEsbfGb
Q6VfysThAaedNgJWGHVXhOJtYvIzGenj6OZZxeP+zqOLE2vSPoRddUhmp0RMyqKvl75FwEBrNeyl
Ypkq5iNERzGhXM1scMu9FjArMx1YQsyEeC4D5SV4tqUEiLj5ucoV7QzyOassyL0RM/TUciPYo8nm
bCrMDtNkOQE1NpcPYNV6FeyIXjJ6KfwsQsTV462ktAwSLWbSs9gB2u3sG9GyUPTYtnal21yENQH/
wCrrytRUhjqbNLMqONRVlvfjLJ5J4K5zFBRtsexnRwrGFY7vfnMEChKpdTkZ8kaK2MEHSLI8v6k+
NiN88yMSSlLuLfUmsN2nqdJLOKqTZwoNiuIoqgMXxhk5dQTYdqRm3YPvLLwN9sOqh+VrwBaY+/HW
QKjaK83qztm08ixtP3TmboYIR6BstMa2Kb04lPxJ6Qgz9tM9pdtqXJVcJ0vKjsMNVCwghmOZ2Skx
vsuM6tagOOsMs5/X+5Zvw7q6KOVj2QkOnZXdYw9tJKKEQktbG/dUp6uDciug
`protect end_protected
