`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17056)
`protect data_block
Z2UWY7qjw+S+e3vxNhb379eORD6OCLUieFdbCSZmmY3bWy1pbUEzvJNCAtAZ1W3zO3qO3wjdCBd5
8V6kq38ZKQA1jyAwAszV2tElEiju+rJrh/KM+Grc7uNha1lAdOOGCJNv/Fe2N7aXTmZoZJjvkUcC
rqTg5Hl1y0cwjjitP4FW/uNYEfPJ+0zqG1qVJGAbfP9dB0zf31Bd4ybtjbGn1tMAqjveod0DafNi
5AgEROjiSUYVgk716z62pBqDk1a5xDDLoHFLaHNx38AD+tRdU7IVJGJKARifEjxgn3VFv6uq28Zk
FY1yLRaFnyuAGF8Hcgx0McbCbaAPE1oJQMILo7aXRKErNBUoUByUgmD/yX+pebOphcEVw0ZxTxmG
xNYMTXn5hfW4gnU/++6216XqoKxfvJRwXOvperojAyGda1yMiIMfCT1zmdeBTEjmq2SboihaWA4n
TFXTM6pJ8n/5mclmDbFxZOYVsWOESO8CGKQCtTjKFzH7J4V7kC8AQIv2FPuN/YDaGjLkaDxprR//
G/4wJoMfaEzxLkVwlw9Dyp9wWszBcg4jik3fvHcTTd+6hyUp3pfl3LrH4ElaREfCexWhtXi+CI2R
C76Cp9fhvnveOl/tEhI9ZzmOawrLwTSyt/0+hyC2odmf+u7DpRTK5hwqVX90HnnmmBeav6Lozsxg
ebHiK/g392lYUc0v7CpsmvifsEmzPBW0gEZmo6erGdugnHqSHhwb35Px8a4g7uySXHPZS89crjXm
9sN0kYKMta1+ygfScBQfiFAFOLtr4781Y4quTm4SUIfRgF4p/fFnYBQTKluHCt1Nc8M6jClHevAb
cuN5hbjaqGUeKyhKQBiWfjxi4NJI2jF4Na6HQgPFjFGbn3TjCCq9TaMu84B95GJ0SYEPLkavYZJ3
M4xARXRi+bjT8CS9/vYP7VDxIBvt+Sos2VuLK3w6UQiNwF/gn7j41Hqazf667dR0UuRaRm+cWKVE
VYMM1+zwB/gN4FL6dr2SEQIWGHjncm4W+hsWPhCGwQZN+GmIsq+I1lkeu3PfJgUXN293X4ecTrkh
pmlv8XDxZaiiR+TZbajNH2T3Nt31kOjfgzQQ40EL81mFJSe/mXUj07FbhOIoMPje5Nnxtz2TKigq
cpfVUgWvU3B2bglcaUvHPVmy04Dy0oYP67/V4H1COeoe6CxZhfBv0vuKg+5Q2M4vIbo+uIwSBHHT
HnfveqnDvFlZ1uBGIKlH+IywBhPyGKbQ/uKPhFtELS5GNbAudKH84Pi6btnvW1zT3ob1Cg9LDHCd
j+JINT1Y7SbdOaWEHwRx0939m4DT7cD+M3f3Fyv+UHpbgXke+zLu3Jl/fR2h7kNwrcckRXbJqm3M
Gj+pf1pcGKMH6cZ00TVOgjDLTnYlW7kURQDMzioPyMFmghEr9tIlv4E/EtmwLP4tZXYWv5ykpovm
aOsNjeiMLujGHMT5SSs3QrdOWroKzJ1LB9rUN2uFlfnfSD8wFm7ve3aKQrvLthd24xNAXWYFK/EK
6s6RnyTzQzb0HxoByH2RUK8A7lNqt48nMcI0oKlVxa9v6rLk/ECwqhDiiVQWAQ97O65UG49+G9K1
I8A0Q4EZH7qIeJ3hOnr43OopPrF+63qNLW5ZGIthf9Mbt3Y8Si7+NJRtflEAG2Ind4at083geGkB
ivp/brF+CXNFDX55tYL5Ceco4ONmq5VWAQz+ZXdldZYF91a9ir2YawvjTegG+qvQJc/8izbFoqkB
DFPuGm8+KcCmoqaiO2UgBWmcvIAknOKR8wVcA9gsvXUVQGDDRDxfzOMhUqTQZoA/PCO3lvKoDc1F
DASoWMRI9ZqyM3OV9602D+UvELa91tM5ecwE0iklDCRnbUjFFFkP+0UTPlimHeu5d7Nd44ixd4K7
9JWnPwWn/wgyMnG0x0PxqGjoV4Bji9GsirFAmpOm2qWBGfFUOs0rvB6PUKyyq314jrgMbn19TA6w
LKp/ICSePF93TlvQ06X5/JuuTBDB5T5aNdrhUJGoFpWHX2Qh1fu/H7Z++xKkPIj4IbiPtTP9Hzw5
WACEGBStVH3Dqk+AHdO70MpoDi4W71KSdNTgBTrq8JyAy0yVhcFJlK1MFEIE6eKs7/SI8GlJ8yxj
fu8NVuQ9fLbzGmQbYQzHng9myWQMrscq//OF/csoT5ov0cOxYHTO9Y/Mfy4WfJb8yIw3mRR00hgh
4f+RarGgIYbVozNjecNBbHaYjETUEmrWxw6Ph8W++d7xs2NgO84G68r+YEEbb1q2segnmPAwBuUL
rEgWch7LwQ0Qs6LWHLFsy1UwC1j2QGUEsE3rFFyg1MqiPghziDqdvnfk75fEV6s1OHhfSoPENcUP
2C2pzxr/dCk8FlafjKUZAiZy3ShDGU6/72g4CIvM3A+Ala6KmRSyxsjx6cVNKoAiy3c/MMEfvTR4
JQsDb1wWUqEzRzDlAu8ZVia0+1t6jx64NxT2NvNFnRpa+zzGN+zReQXdpvTynhW23xsG9MpJ4tBW
tH83CRPQ1lqg2quqy6vd4PWVdqq6/4GZIvzM2/0BjwsywKFxhYFBJ/+yY1WDLepuF071KrC7vI7A
CLDCowNw+XuxpnLQ23pJNI8ZagBieMQXWR4ZvCMTG0eE7eOvS5Wy6GWKJ14N2X7o2NEYQctgOmSp
Etmz6s18+XPz3dMvtf9hahz6AZIhKt2h2uCdvFbW7H4Mg/KB6q/FwPcm4NTJJjyWqcWVeesRlUd9
hUA6B2nSLUD/sH/RyIHLCjAUKgl0d2gs0noa6+zTx7ft+DRfi656Uj0SPbYRaKf0NUJAv6DZMyVS
QUYxRcHn4b7xS5hSK6YGy34yXVzzn9lmNVbxE3+iUH06ACsfOGbv8frB5XrYHP3aJLdDmr5ZpMsu
XcC+AJ+3flv48yXCo77KJHqS2KTGfy/+gWTDa6z29D4uFP8I7IDGMzVOGFlfmn7s7o8Q85XuqaIN
eSOWeBBZsxahTmZJRdeg8c2RMYrZKAe6RA8VOjts0wFFJ1P4K6uADVJm/j/hxk7TYyOesdxV5gv6
4H99oLpQ7ketMwdf/euntbZpNqFUIRGjpOMGBuZHlT/vol6dpZQIZnIlsORt10CRfqcwCcKB+qaC
mNE8YhPEXbyuAW8jD+sDw3KQPgPrYe24lREgIQEXMiurwMYkXlfk2oH8x6BEZPBBbeVVm0yoVB/2
Mowk6EXnA9NVbPveCVgqLE7Z8u0DfPrXrO7vIpEHkF0I/taYqOjfcdnumG3JannVljCjD/qaJIFE
YEpfcSVNbtEbKkS+18lKoCe1wEFgXrCmPZfsqpozS/i0A/3f7lW6zku+WR4qZhqDjtaDIbo61paL
hSnyaE6gJJDrumAp6j47WihAUPf+7LXj6/z5NlwnUDuw+nJP2f2YiqWASq6iBSLFpxeo/jZGyUTp
WJc3J+IvPMzPyNVvI3j81IQYCV1sNBVWjlgRykuFcO6r5MoqTgcDg4pqo7dlC/MrgDHMVXSGX0d9
jXS5CLMYrPr4PRwJPyScyWb6QM4CBAFC8l7xVZq1PRIJ5HwMURcFzKCxNZVKf1oJ4tO6j07I+Z9J
alyucnF9PZhlOKAxZG7yzGAwcL36VEuZsJUarHAIlZCvVQ6Eh9N0wISxWJ9Y6WhrjXrabplA0cXw
EdOMF1wRTCv/f7r8FHzgLdDWH9G/mtLIWlnnkmin6dJX6UwITfCI3fvwmgPTeNaEF0/LG20mNSGp
uJR2khuNhplL+Cyd+MTrY438VXmyoEOCa0dh+FjDfIarT1oR4gYxgSddGt09OxNpZLvWEXdYD1BJ
6xLny3xWmcfFFe5WXORC1uzG7vkxP0QyLtkoQ8RswooiG7vwH08KkKiKaRZDAXsaHyxl1Sd7xAlG
d104muvirzbw0QtRGVG8LpHqQnMLJ54N7rDFovrMV3a1riSc5Tv37thyvY7sK31i8h1+DlraSf6z
QVArA9WsXEr+mXkc8+fTV0Kp3I2LAWooSNRHkf9dNAHOhGWQaacjfM5RNoslB/5l/0IJNwrnRVKj
v1/pN6xM4zR++5oj80sDVPMZTjF3R6b2CGQXHQPVcVfzuYG3oEPcnL5c2lGkfkVUEWDLCsaWj1zf
rfwRqegI0vVuDK5Pv7Bk9Q6w79oivzLPPsIjmGl2JGTm7ORlhLz4s3cgqiCBCn1chN3hAjgP9+Yp
1S4IkegGJpnTJEzL2O0IZcas0VwjMKZFJkOw9Qhs1I0+hxLKWXXgeuA8wvMrFTeJmPW11HefC18s
9r3HRpBAKNz2WbWJ+111Tp2nf4tTPST+RNif3Z1Gqwiwm0+x9IGh0wtwCtk0jgw2YxYhh2V2GNy+
IjYr8VQGtbdFLKQrYwVm5AcyB7FIi8WOpulNYeDsSgRoLbuoaMxk+TPT66HeuBp/VjAalurn8q5T
crT/0LORAmaHyMbDIncOyTQCwouxkp1ncojRt3lU+f8HZRkPX9XpuTytVHokzQ01lIFpB6E/Ybgv
XRP7hvkny7cc/ZLixPMPJhzj/VcbErKsgcn+jYTl5puP5pLCoJlnHZsYgLBF/8JpLqzfsamwQSVF
TVBR/FWF3rMAUjmWS0z8aRgew+opk50WTvXAH6kHRJ0QeNztal3GkPA5snnaSI7zC5mBkLlz3ppD
KzofDGsK+jXZ5agpZ/MXWdH1k9m/AETOPwoeAKYlWncRzylguxu84l9pP7i8lD2NSgQNsnP0wCqJ
L0vKRTsdeWAltnErl3vrX3mXzdE7TBN1TLDq9IJzKFQ7pdo1Wyp7YAoaImVT7EMH0113ezW0JpKy
GtSc0KI1RzENzdFL1PKB+gA8rBVc9q3P8Hb4C3TFiFXophLpyEiH9ArvU5SLFIgHcSWflY6czMtz
tscS6VtArtkEp/kOUObi9bkVbBdFd1/94SThRT+Boo2KRs0MeUpc3wblDlP3dDq0KEIE3GpbYN5e
/lP9Ttj4/BWRCQW+FOQUQdv+easOyk+Yt9OK869OvTR13b74qaJHIladO9xaY3/cGHEz5EWuS+tC
PSw5BqQW0G/8pJu8v1/emBzq55hky9EuI5eHHribmg5X0JZkdV0aemzbF+kTI8WtePCgL0Sb61/r
88rwfFN+pGs6l1w3Qn2fkBQGMH34cxCfAuiwzisB02ynIcnDYOGk3rqnTEjJLRBm7VzyS8RjMdDZ
T8IJA2LpreQEIuivhwYAD+8SOLolAFQZlzC/WPFACsKpDU8IQ/w3BY4cIIUolcdD5590fV/VEaDP
Apk2hmeDW8LTlZM2zui2wX2eU28fB4DJ7XdL6bg9OQoSlUcSVLRwBaMz9OqjRrC7Wo8RNqqI/AKI
pnHUayMJGYQYUUbo7jsIc1GE+YTCJoca+F3q/4jVPTrPESkkJawUgBwl5x14k/UEsqQv8hN8vbL2
V1K/A0P58dDBufzHteO74FVq8vMr+WsXsI+kyEWosKVqflMCiZMZnzhnd/p9IIH3TvJawpEsz0Zd
X5Bq/0yoH59wus/BrPMxGJU8/UIgALA73AvDyeMZkcGzvBrJ4GDlZl/WrL8Fi4NMd6O7dHGCyutf
d3jhfWZ/3KNmmq22OJR2f73UR96VSSRm9T/V8vpvbOK+tq+J7j8XrwfR5ufkn92UC3HnJGabMf+6
DhHhxXtrkTi/D1H+myUFYoM7JbBMw/MFRPbg2Au143P/xvO6ba7shdSWffbRovSdIeHIooOr3I+k
JGHQ1LQKJsEXJw8c8zhS5UXe11az/P40KHV97rfWiJ1RMNKLeB1ZlT8YSgIiMThJpvKACOD5JeFX
+76gS1vxnwP4O5VqDU3FOojwkZY/f36/BhIyipvjgCSQc+WV0lahmaySMF0C3l0hq5x5sVr+iOwz
MA/pMIygd5AdqrZETzHxq9W1SsIyFKh+y6v8WMXzlopzcIx0sZhNcl+HMn/lKAcjcxL8dzaeK/TA
ieugzqjV8HVeo+iG9hIlmJ9OGklrvoV03d2TZgm3VpdOZJuxiTXtVRink7o6b2r2MrC73iqqPrNT
wimEQQbzITs5vjYngLEKWP9zQngaimkiBeCRlygwJUQ3LXUwR8AiXPW0DOLAbASFcyMwKvM3bgK9
G5LocXSRf71aOUtK3lnO9qbS/FBotRuFkpmH88fRhNH1U8yAsK5+tmlhQYnqr7ZotL4RuRg4X+PI
l5qPHYgunmR5v38uYZIyJPg8vdaeWCYk9GreVUJQgdyf4xqOi2QwV+wM0SIsaOlmUX0U3ez2INta
/C35P7Euie5ELi2hZgrZgEa2u9J/tyBDVf79d6+o5q0jelgikyONDXdBBdTI4ra02/XDVbUlnyoA
UNz+yyOjXOg7rPSMMV0qVY0K8Th3mHWYjmWYFTr60yh5eRRv4DZ24ihxztRZkzaMQQmc/WUz+iT+
lyHlo7d8pdaIJHRZ41IjRKDSjSQjzIQaX4XMsF2g61Tkpyq33MlEqgnFM5naH399ji7bWM74H75o
pblNNmU34RSPnJwXdnxYmJ5VOAjd7aSxcrZhkOgfCKU2hHkc9bibPTv2jrG2cv6mAfJSdGRqkxLc
UAfLBLWGOvp2/W2xAxISyQXzAaERaOQXWDykU4fYuS346ZcGBipiZKeBtZVFzqmCGRQj/bF7UMi3
UCt9OFV7g6iaHz8kxqAOAUJW0+xy9ljtV+b6cu9UBvF8dWF4r1jky8cqIGMYWRTWoqHfsJuZfVEK
qMxTzTavZfrchESRXTtBhg2Jz+gPnmb6qnSf2oFKH2oygEBpXlJyLVsV/Ov/+qfxAFsE4v5PQx6Q
tjuFOGiPTbz/wQGsWHAzDOaJqwdcWurdF/TxpH8ot2eGLNjXbxuIjjofTBULyhfa4+1YFrFqUaqo
8hYdRReZw6/Cjens+TN7SGUOQ6ONLHPxUVy22uOxW+7QhAJE5VbOMJLdVT622vuDHrSgh8aFqgDi
+XwsH+m4dCktMfYvCga9/8BgtKfocKWgSG7Fz8gNXUoYQdZAjmE5srGWpehQpp2Rgw9BqWF5TgR8
cjzAMkUJ7cn3fdOJ0gqzd3AZUc0OQcKjbmKzeG8oUk9xR78/RAZvjlFHsisJ5FWduB5/RJ5SRaQZ
C11+leXpYqgy1SCDIrp8v9gIRkrb+CF5xoXhJIVtXKbn12qHgLpaW0c3pISJTu+/qE7uvq98tprU
gaxyba/cUBcRPLcMIPbGUyjdee5XBDyrvWsWen1cF3hdJcQXyvMDYoOfhlldFo2g6MOVrh8p4DzO
ylkX7pFYCG3142a9y/1phRnJ16YT3sm1JC5qt9vbya+03cGx2Vh/NymbFa40TXUs8Cjdhv0jKQrK
GsDuj+zX7Kc8b/duRFf4sjNuhrIMLhTgeqYiiu1QXSoB4QqN7oQGEIBGo5VJAEsX28GG6+5RhV7M
v1Y6nN+u5MBIk7pfJwbarL5G86x4+nBP1djFvVvjsg6CBH2TtM55nAsQVWCKNQOE1BncjwBlsHdz
AGTwDrLr99xLmhGIZ6MP9npp31ASB2cRPSL6tt7xE9NaAKYygxcjp+dk08cuFhUhrW/Yme7E0ps9
WwXUsarIUSbgw/Ur8GZscvuvcYPqFxvwfMVicKAHRMhaWfbXkoE8JGpGGv49xVmBESc2R8zt4ALT
Teb6LWbqdhCGb9LzGFYMSUbvUmh/xiQkUJ0QA8EWDBDOp7S0US3K/cWCsWa7sSrKkv8Wlb51F/pU
zuXfi2ErdtwnrQbT9OVtYhFV/UYdocTbXvHBJm0kHgHnjfDEnJwz9broOSwOiiWfAUreVwhdeZAo
5eioa0+RWbZ15Pe9PpWu6fQ/eqTSEJRCEcVxoCSozv74mEPn7c6w4sT0FHN7avD8wBUi4GBMD6gq
+GeIp4YZnE/ljQOJYXZyCZAI7tyxgCvWf3lLrBWLBnI+b6ZZCEN46ELE+NTXqbEDCfvqFAcfsKJP
YZ0LvWVZvGSmttqC3V2N3TCiqeuUZAi7d3kUhwUSfrIhPeKiRnSUDEOjTRdRhIo2DdQ5dkWgYanf
i6xJZbEY7GNkd4oKZtmY+4pAknbFAhrqzOkIq+u/12WIu1Ljj2xlyBVq8gtIOHxFO1bnSrOTIHO5
8mhgRgJgBzQhKZbF/vB/b2DEVBNYfmR1LurXg/cmGELPDJGI3EfTpZZjifSmD0jo6AYzU3/D9ejx
6ionxq4wOaAnucFeCkUjHeyFiHOtGEXGZhfznhVsBUWvaFeA6alus5/v+DvCrhjoWrVN5fzcntsy
Y606AJvq2jaziCrR5/3lykvrzZcp1qkJ3m9aOv67H1E1qes6frPn84oos5j+bKwCv7KDwqSBJiGd
8ZLeOD/xjCXiQ/PYCnYUN/1nA7C32ALEiF38H0SIPIXWn4krDMzCZO6oLhGQQdXaFETsgAzafKkS
Z2basWMW04LxUt3Sk55UBa/cJLIsF6oKByQNAzlc/FQMJVrnxPfU2y7pxzI7Wnj/w6n54JoEVhRt
lY+P8iE0aZolQ4NYY+/vrc5u9f2rD9qR+JL80WHl42WKjru0EDhDYI0GoT4HLC9xZvd7vDLdbugK
0Oy2B3f2dXosYDcAJE4sHGVS3TFUi9UjjHegEAHgL/d8VxbWHqh1bhxZh+6d2xcjyrquNuI1dNlt
L4Ivpbk+btB2Y5h9A/oSBwewXlhynQ2MRBoHoVKhAki4Rg9Z6evAZvar2u5WYDw5+URNgRwDXICi
PoMrbY5v+VUqFW6bwgozhF7mhdUAZODQh5XlmkFHKj9zEGP3dMkAvFMNHATS1dIR8lZw8ops+oSf
wPKxZTNBe13E1zoIEqv5oZVCePDS1zR3qxXwJ/JkZA/Z46S/MKtaPP8IAeLu+r0C5ms9XTsYWPdG
VA6yYOS9+2KzkhRLSj6oXxplqoon30JTjsAPOAa+iMeiDSL0iAwbJ47/RD43fRi+TB43f1XeCILO
NX3a99uSvtwsyuf2O2CkjKF70P1dsC7MrIml1se4Qw8uML+9ftXGPx19PZk9T8eERrOpPazaeIy+
8YINxfiwgdZtv1DeWh/COqcPLW+1qF6jKxVDy180HKszMCMLhPX8M8GkR7nJFalJMjcowvMAGtqW
bcqdoE4xv/5R//fjW73WZYBFhaO0ueII4n4bluIUorgmjGKmP+7m+P2vnSoGu5dSUdS0W5Zbbnje
2MIBCp8PRZaKqaYeosdEUeSyl7sU47v/ASnhsha9Fhlrou6mNTOn36jiMp6E92PUuUn4DZ6wgZ4l
ytv1s4Yg8DmwoaEubW+qwG4PRjY9I+lbqiZxWihgy8YgDokJZUgsy7hpRGHP+TqaQlGuy6OM/GXG
tM9Fubn9Qc/V+ErtHgK9OMUSJ/C5oXVWyHG1HEQmm6bU6fz4Bg4PhSX6sRxsd/2bD7e4zJlnQicv
26sOvCNmjl+D3gHq4dUm3CWxgWyDrIo+L3NfbVc5+dZBq6YB0PtGkvBmKFSfDNa56JX8C/y71IIQ
UUOOcXGzid1ZPrVHwyVS8sjmCDVPIvDssJ2TeegYWy0gpr/tTOBY1Q/BOJ3JpEpMFYMeNAlknPdX
S7vS0Txz+VvTDyTL9OgOJAgDVwxjJ+03DsIFT/fmPqqJTeE50MSAHZY6L9HewA7vpOHPCSiMhORn
CXinQnZob8rY6Jg0o7hWoVpiqCfAmgpIZk9CuWeM7fRquE/3NhZKj0PrJMxi2Ni0PrNKQIMtZT9o
kZ6JYokc1rhUnRwTw1aafrmRK73FaEV+kImtTMvgUyXXcbaIsttdF/ycSaQp3S7zLhU2qrIbBqNY
aB7/zsIOCsuHg6N+eDwyAdVAdkobdr8O1nmn0yfwnGZMzexzARKJILMQsbHeDYW+DIZzbqL48F+U
dtI61BtUwmsY5pB0/PSvOYZkbsO5OeMyD9xj+UpHB/zL1aOv7nHHUDKMtLE5zPIPntd4BeDEVWhA
w5bvNV330UjbDDqe7Dk0qS1hl2xC3ZVoLOZsAZOP3RSeFrsk5oh02yo0f08fExcbIlq45HS6aqcm
i+FKqE2OG9LWlvd18r7K3S5+TnTD89ARNvxEUiH2dDSHQCZntT5+0uWw2QD4o153H1DB3XaUegLn
p6byGiAiLV80zJoyVIik5PthS03jZIbjOHk0/DK14Rpn2wKQNdXSh+yJM/s9ogoNyAP5cHMD/xyW
RvqcSLGUlh2LGasE9wtcIYiX45nu1ossyy79qLlNyBl6TawfpKLt0iPOl4mhXI9I9cgeOZ1gNVrg
szKBp8ehvYpuyqT8v4TA0XtdHKgU6sfWgwxr3Gru+5WI/526Debc4/Q85N0USOuXq/FBuxzrmVN9
iqsN66TMrsHrW0p6IGnp6rkC2JAIHXn5Af9MA5WZjq8puqlV5TY2kwU64HQomYb1bDMlH/pk/YHj
khrOxBFIRZm4UdgF1mybWbXXYnHbLWzBSGG+9rSSZ+XT+4e4d/AAVD+n9gEQ+WFliaIuIzsvPIC8
FD/dHTVheZXgEmQyVErvCNZ/o3b2udbpJIYx50zlhmeTngJPGraNOixzHHvGlopTPeycRZ+JN5pb
rYOulqTVpGlE5g+jvmWevnbA8rS+xRs8jfa+IWi0X3vhce2yDQRHFAoS0fYNM+ZTRecLKX2GZnQO
Sd/4dTBkThdPb9Tw0DfTx24fSJm4lqIEEptJkkF+fVoG+i5glrJbKisYPueuvqfHmFYgWI5Qeb+z
zocLFKB11YzjyNYu288j448fpG1fdamS+1OOfMHL8pYqwk287Kac6DJmc0Jh6uEHk689WW+PVrpx
bzgeSeoJE9UzYAM195SX3ZfRHI8uoiKVniR4oERb5pYhtOi1askj0vL/2dWe6cH6rt9cmEm3Xrea
MkWnaX8RFWhpvYfmmnTMS6SsEqm4sBXMwF0W+rRFtgMAjJ+98VMJ+x7EWHMxkG87akFr2ENSNegl
Uov6g0s2Ftid+B8vYC8rkdQw3uX3wN0Ld92RUP5UbVSoqsdQusRm/vNjyiuYedZh8GH4mtBhXHfZ
KZMHHRd57RGd13IQHbqURIMS1MntG28VSY/tWo+oeFw4fvzaqhdh+XEuwxAELIyazAOMOdf2F6kf
PXjUdWTJCKJDPH7Rc3hdu0Lb5cthld3D7ce6+SaKbqoy6zP5mFfy1YWIJO+sOW9xv4l7pNPZo8df
8Ua3XkFJ7ZXXGDe3u0LOGohyFL+n7NbjBsVkx5ssv/FNrMGhrZfUb1DE3vXcKZ80QXlW9AKlwmvg
vmdVQNIcywLLEu4KdQFyw9TjJL/me1OoyqKupVLB59lZd6BWfEnPezUpLUmJISAlWA+WSlTrxIcW
XS7l4NrZI7d4htuRHHVhvOHuB0l3b59Rd8JwOjz0+drShhC/e4elOaVPSiEmxeO9c/4/bOfcDRF1
PSfYWQn9oluY+N6Had0I4k0P+WX9+/D+0pb7Jp85Yvy+oC2Bb3LJ82e4ndNCNB7nwytZYTnlIvWM
jyYKTPxn/ePZm+hOr8ghrBRl0srpqFZg+Q/cVwwAn0QsUNti2g4TJYGa5FndZlYOSsMPqONOJI6L
UquJ2VSQ8aNSgVLU+iEjt7Ps6sF8gqCdkhGh+ea1UjLyay2+7HNW5PBlP+AyzAQXRhHr1rWJLi+f
mCybKgp1qyHq2vGvuLpvh1POH0ga/sqPtan9RkzyI8yXYlQpbDhoNiKwXkE5A74a9Y96ex266yW5
Yz/TcAnFW3RFOrVaYvrtZQGrCqHIh4rFdBFvT6d741Vku5tEP97lMFFEqWArCcLehrzV6sU6FAK8
iIU8ND7fc5gi0EBjjrtQ9yXm4jk4a21n5mEsTx6S/W8rMvVD43WxydcbBnJGGMvP2CVfqTBp1uJ5
qVUvhZtU+S0Tgb0ytt1F4JdV9U62nc/zUnrEP41XpHZQ23a23IZWpSKLPMdcl41a3A0svd/BL2Q9
yEIZJWMgoWSJTQADKhjTR2ukHXBPo/zoCHSLOSGPnjdJzqeTljU7T9l471t+sK30Zimaw0EmvRiM
knPQDGRt2bFCCwXl52wBHqyiO48sOCgGPJu1rWfUzagzgApJ1oC/q+2DvSKC6p/gTXz7njsZ24xY
djHkOdT6rqL7RwezqTwbaleaj4jfSz85yCGyZryGOls7o5d9mhLfuQk9VfjUhk4wysiKHD5XMSPZ
NpnCtKwCvXyD3EEoQ5vTuwqiRchrlf7sUae4UvXRVXYUgtdYZDycOhwYuTxPcOy/H391pvRs66Kc
m4FSlC/uHBZG0JqrqiL0oCP4qYoSlycIitYiCODv6Oj+3MgWNZsWfYVPJm6caktgwgp+zR5Ri7jo
hA64xsJd7ctzyGOcVa83Q6EtqIscyHpeIiNc89kRaqVa1oZ2wQDMwDNAgF1UUUXzOEEMluVSa5zX
6NAngzftFZiK6WaAN7/PYGvahc5aYs/ljhRUun8CtZaS1jeO8Ui+DQiYHctHAbv3Z/N1KOUIrHYs
KTKNpjKkfJIPYMD0jtJXbrpph0XarUiR9bTGUCMAetWE81L8AoQv4c+3PJuPnEbw+pyJ46CiHvsi
9om2GR6jzUrQloVRw7o07sKOUzN0mlwqbA5cJHjbF9xdpg7BNJpGRf6Jquh62Q+wzb+tcvYgaZSC
amiDhmrqKMENztThLVUR+b1iZvfd2vx/N0Nn69b1Nvwhy5rIjmbyT4ulr5bFxhPntaLtZFySn0YT
VRI5VXCIpyBIZF/EkrLBIFwj7StbxihNc3nvHCk+DowDsw8Dzk0DEw4L3yiVmFuVsgz35rJCWyuB
AE8mRt+rtpgNaV7TztZNgqbwzowog95WYGcKMivHLXUqB1jh9UaGmotuO7Wsot4PfkWjkru0SAK4
0HnMW944HRXLNcVn55aSDt2kU3Izv22RMQ1EaCNKAeqhCXWwtWgMrmYUKgc3t1Zw14expxo29nrY
5oKjsWzAHaW8a4iLfy6sNT1GAZPvGWTuX5/3aUv6+0BAqox9o3MxauM6Xdlv1HBRJuQserOHNr5t
6gNitpMyiVcxOAZ4oVjl3voCqZQdtG29Sf72vJvBP7v8ajDZNNr1dgYXSS/rBoE0+6fLbYDW3HmZ
UDwKEmjdsfoQzIr0haGvIfPKUWH93RO1rNoqJJ7XgnOtmV74Yqty4Ltlzp1O7H3H6a8/EcMOdLXC
2sW5bt63eUXTcBskitX7xgBJZTzLRZ8uJgVJUhStvk2acxIqW4FIL2MBwm10KH4zmDfW0D3JM74s
Q572oGZbcB1npnyS0XfL1MsJASyI9oZhX8z9qxECQ/NIi4NwhNBtbsf8tYiYOG8IAjMwgQMrTU+B
3pmoCgLylDVaiBNG2zOShsZqlv0Ce4VjhbVc4OcAm9wKqNF9dBkHXgumhqwZcdMzF59HxntGRwNT
BZHuKksHCEMXaFpnNA2lqsCNEMPb66/Z79BnmYSlfVWJA6DVPsEszuFMqhB2+FWm+elKn6X8k8sR
jKdf9kFKECMsqBteFdPCF+vrFYc35OSzRC8my+HcsrawKIhhiwLyodkLnBNYqUWpqZ/z/AHlS6+e
7VQbtwkp2vtiyZr1i/j1DawriOgMtQOxhgRVFijNd4d3jP8Zlnph/XgQTReQzxRu59LV5h2fN68j
UNcpD9Oy6t4YjoRoyRVBouZuSOgcuG+8QyES2uTplx4WP3Y4snl1kCDcyHWutmTLFeLWlHVGcaCa
0aXgtaUCmOw98+b0QAzXVdFEX4V9lAyZqNZMqmwohsCzMZZt2UL3U6T3NtyRK0hf6JsA1F80UxB6
dXdnqBD7dDOYba0fXNYf9RcY66Q7Xfh/Cy/9dUGpBqCyqKnZ+zqwYrlVyOTdudJNjou+AJ9OlnOZ
T+eNRsqp+VwLtHLNscrC0WafA5UnmbwbDMwneFkEaOhGdlWVK968k1NBx2BHccLgAu0Cg02ksGoD
G+PveQmHC7fioYNSvwjTXBQtoaxnd1eHU16IKQy0QwA/15CXTYMuWlQi/3Xpcg9lSqpiV6D+ggh3
txd4Yb7ZoNeeQyg57Nk0Zbldw0XHRqVs+VZJs6UG6NuuoFHEcSOm4700DuTFBH9ByVhU1dsCN4zi
Zxb5RTzvp3FtthJu9Oa3Rm0CPwGroLF970EmffJbaJ50KGSuwZk9TVzfaQ0HA41shv2RGUqOfDKk
WDvxuQCiN3xGTxW8DYMlT0T2bYJlRbYX4KbCrHEGwxbex4JNPNKU9QhYilFC44XR3nhC4uDQmSj2
egRfIGlqYGNIfAyJDsgPr4OOjE3dnCEJbCXdWlPI5m58U4Sy2ws8nPz2ZHgnUqF/qDmq4b7Ywj56
9vCMT4g6DQsVdwVY2xvsxh6mTNfxjSwEhZbNmQOI8ANOc/wEwctNq5guXikiXRGsSmCEoI6IMkkx
b2JjiLOwuhv0tA6+ClKSGqpWTBkk1tbjhmNt4Icjbv3efM3nQKNgXP4XWjx4iaUvyQlbKS9QtXE6
9SwQIJ66WTRDv7fsPyHFUhMsoM6ZvB+SQFJWFjGFSjD5f1mLR2MI7xeoF/nTuv3Vw4/v4M1e5Yhh
fKd2gOwe1ZR91Y12HRy8SKUDMUkuT3i/KNYINdr6bSDv96KK+u/4USe2dI7IFracgCxjjFb1kalH
VnLPxAvmGrePTekulaa8YRcYCB2Bfqte+rKvgrQs9DAnugEKy8iqcVyJ/AS2FeDNdzK2x33VyLbe
An6BMza6HQY36s8CWcfCXmQlgQjKdZvrSoKF0Bmo8/24KZqBYPyph+7mcJSRi017qAVvEg5o+S29
tqsLG3IUXlUJ5iUX3DPWWl5bo10nRex1dCwC1e4sV1Jul1J+AuANGt/KkbZmS2S974EKQpEshLHP
8dr8D5ZRdPFVwBE5xzQ/dUjG61J3fuMIVP3kovc/dvMVR2g1sjhUoDr756jQKUhOIYji2wFMvXbK
Uk4FkZsDEA5a91xVRUHswts+j+0/Tny+0GoAypmwjttfu5xoSaO5aRA1EoPifCBrh/LBuzuBqIX2
Y5WQnII610IyZY2Buucqw/+WByDSlJqb4zTZUgfXDa6P0M4y4K3R5AG2s37hbjG+u1JpKHKo+jbP
FCbVVtwagqFAz2ThInoydqC87cnp3gYTUmBGWbJeTjFiFfHUDyYehMCFWWTu89reIp0sAKdgzGg1
RuumPgoQjGKcZAaYRjkb7PAx1VrSQgE5hjWb9smCnHtAdnQd+xu+LYHkMnMtKTpmqnVcvPUF7C9U
LT3Qr9rJsZW2bnCEhWh4rGB+vfwlf18bApO9fECP9vA6I3HOezFuvyVonD+Q9QF9ls+qPel51QWp
M48BzhVbS1NdixCnznRGXqVuHefUmR9mq9qtA5PZhJAvPxJ/93w492X54/jPtQQGdWc525+Bf4wp
RMhn22PvyZNvMhRx/NEQksYuKF/u6wGrJrPP32YmJ0Jss20Fw+dZvbeokI207Ie3VKnlS2lqtv6d
9lfhZykCR3psQb1RhCvPARHU7UvwPiNe1kguDSHxd/fEazfs22fQXTAY064ZnNInCL5R+Mx/MFnq
+aOVMbkv4nFeHX67sBN/NPUo6tHu2wHtaVc6BTrlgzz2beTwi8A4HBrZZ/sybIfAZc++Q7oaqIr1
Xf2BcCsqnHQx74CBtJ0pVdMVMe5efmf02uNLdLKbd+o+l8BxkLrjulI0osQp/uj+0fb12n5GMhem
WB45528RQoqae2bQFMk5cgbt2sSTzDq0VL+xtKTFf24PGS5f6Mqd8L0XZoPV2u41vVx761+mYYer
24YR7Lovb7bHsaasGJJItQX6Lz2EtCg7F9i5AN8r6lpNYuCcH+Gtn5hocYV/Y5/l4+kQrAWKuYCh
rQFOabwMfAd0TdmJO8AoLJHu4QaX86HRBh1pCPWI07Ni/wPskEMTAkvy5qz7LNcLZT3LNsWv/yDB
+xvz0pS+oZCQrLp1R8Ojsxp5MD6A2Jw1D1QbwjGBlP2pbo+2/hvzfhfARLLXOAaJc4vCUE8hj7gR
Y3/UpbIdOE9Hgfprqj5ndqBFs8+WA/fETt7KxDo3QexY7pdzOlpVjOW937q2u4seDXXJVT3FBRuC
xeWKW5SSwJbbG6aY+Bx8wYA9rXmfzcz7bm+Dk2JbNOhjReYeXz5Qw3/2rHfq55VxfrpVW0e6UyQH
N/QsBBm1piUmoYed8rvw5gVHhOzhfCA2FbtVemqOh8UvVYW9u43f/7rlzGLLNOdX/Os19lYXodVe
P4rLycH7O3jR5jyx3wyvXgXxtme+vw2R32J0CMeBYSN/9ZVYYAVr001b86XGz8ubuJA2qHYtu/WZ
HKakzPhGFJAw/Hl3dORzI47Zu5dAHFcSbBG7uvxUbFvjiHXSM1J7mWhZW4BIXveuxpoW06M/Ibpa
WGwHxGbee+HBHMrL0ETW/1qnjRx4zCP59K4anxreT3frGjO10gpPdEn+fJGM+I9r0C5ycN9viCjC
5L7cPjX3wMbGs6a0m/yRzVKoYr3GwQZ0Zr2vWaOu5y90KVK5Axs+M5sCOZilvSfVlkoOC+/LJIFN
OqKm5WFYTDJGSGXtlWkAjtH8QAu0bA+CRUbWRK00ptjil6k2Ph6Av/EESvZ4+t3y9RGMu/0V6zTZ
LbnWWQBkfTOCajGNKuYsjRhB32dvxYtPT80EQ4O3sXMIBWuWnDsnwmsYDGJ+8P6j1zdiKUjwNhbX
XCpCqSrbMxrSEsvutFkyoMgCQgq7V6XuQenzbyfKukWsPZe9we60079WGaM3TZ0XRqM/e9gFy8QS
okLR4VimhDV3BFcr9GokjKhJmsJNqL4f99Os80hVBOvPqWzJdTRNC2s03xyONo72MAusrkMTpEyq
lBoeqPyEP0S2mjBYxcwbm8xLnenKVlThZLSx95O3xbxvGlMwfsoB1VmLimfPhXQNgGPVNLOAYzmt
59JdeKnbgb8tMAbMAm+WiP3OnXqTr5eZ8164rITz4prs7kdr2lIF7Y1nMydYxij3r2tYH7oYOwZ3
dFyKJliy6gC8f4uDi62cRo7rmiX31NLh3YXuJcsXxnLIjfoQgeEXaS2sSFYYUTCb7fXXdp7Kl5uO
ajugvU+O9qwKxwLwLp7JJAw+YwqDkEFEw33Lf/VsItGMAjbzI4CpVWsx6esYVqIN9aJcljAXV/co
njqk25oNWeK7Dkdmv7GpDC6BI+rY8atwlKXMg+mt/dvnAN8pTGzUB+S5/9aWS68ai0yy5elcmk85
NqIHv+JVU5iPLbHLrWuBcB0BgFQc2ON+urCWPTx0PfBsHLG68hTKIvfhQMUu+NLkPGEnqB4kyBtp
H9y8mhA952rE9VEUxm/DRpsToHXjcCzsEliyZo2ScVJvlhshoynx447Tozgndr0+aTF6m37QlJ2a
qqV/RspSvzz7Zz8H3UQLPl1eiTmKLouGD9R4ibtkfU4vG92vOuYAfDgmcgo6cc5EWRySr/gkWEBh
LHg93cGL4zJPHxp+9Y+SHbAB/ISPV+Lq3Rz8SjaV9/gCMdGccNjHkLMcbvG4jeLPbyLMA/6Nptn+
6HXLUSL09Owm/6Oc287tMAjmqvHWlExQbb97xm47416Jn8Z3muGGi01Rr6Fj+GyWu+OxgBDt+Ymf
54Z4HCYvKCXYGBRhT1w2A5nlI3MtedNXSim8b1FHC9lNI2lXbG5jNoXGSAth2eep26adHfSspZDR
FcRWsghVY20pGHUTS/hmnVLn3ywTV8ZP4L82pPYGaPEnAeAICtJ5XM6dXsOEHAyvHpYHMjG0XAlF
ueJOG/hCcVDgV3APkw0i37vTggNDGZpLqcJEMo+G5A1+OcO2INLg+mbrA/xaEAiFNwjXyAElHYK1
AC5jsLhfZ74eHTvJlplmb2BboBxpesv1oiYI5S4rH1diaMDpQi8hpGyervL13ly0PPSciX3T5P5z
u8nUqQKfSGZ6xk09UAqXw6Klz4Eu0ffJMwKoCQCq9ydPFm1kKDDFlAG+Pm2Qdia8eWNfMOECE76H
/gj1cAOJd8z+7DO0Xu3BLb4uOubtP8KHYSmMhUwbHZrhbf3Ib9yE9UPMJAEb76ji64muCPiBOep3
xkyMBsYZ5xLmWG8u/BVR5gFnKczW+YxluncKy9TdCCpnlq4Hl8bDnLAdjbXTNKPQ7iEVg7hnOsWl
ToTkpHolIettpiDuIwQ7nr1YI9xCS7OaKP6eKL1eVLA8i8npabrvdRdfNLMIkX5pP4AND5Rkyyij
WvguB5iHwypwbJ1pQ5dn7f4vHwab37Ob0YJf3BsubB2XTmpBoeHlel316fexfNuqQzYPgSbINdlu
2zOfSeR81OmIi899EGpbkzmCTlpI/TEoMKDS6wrzI26MPzbih0t1DCYwV4E240txMICYE3l74LjT
BMr8cnytCRGMVLVK7Ggq+Nl6sJiA1qD7voJ8YRlr8zac0AJwhn9gF1WkLC+Cvg9QEjZ75ZddjgqT
QgU/UUNmcVr9rREzNLzn9jgznWc8UJNrr4iEhyqSY0COVZTQvNk8ExeIT1lAOk0htlzFWgmepSgZ
6Man0O4at3NZaJhA8tKnGpWS3AUivLCHQ8iBoudGQzfR4Wakdsg/qbS/7dRuy5Rmoa+yld6/Ivw0
/4tWV7geGsszmqedLlQk2t78kDtr+r9T8+x6+4EoLxkbnjrRytQffjVXrftAOwEDYiEUobApHkcS
8GQz4k54z5t/S0YjxHWba8+7qUZZYrMbfJUq0gx+YwZI/OTqaSOrPpYuBX2acIaiYG9k8RidkQQ7
K3Iw+dUQEy9UWr5lGFOZJfwmrSqZLQGreyfhemadIRZB7TurhQudCx1TMB+ox48ebkai8jYX/1VH
GoJDf8fOS0qgNRy7v69+rHyPRvkIStIy1lpRRQzGaNlVsAn7Bcxl488xzPuNcdBL7tP815LyLlsy
jAmeZ0tIF/TSiNEPix/xU532emVszV42MK+5uHI/LXoCeJmZaJZueI/A+BhOJ5+MvMNINMahR+aV
j5COuGoKXxhGX6nrYFqTqfuy0C7pTqyVDFdvJr334Lkb1mAHaKia44EwXH8FN3+BDI/qn0M7FpO/
IKsDPc4cAa36zKEvYryPHE32GEHncNVShB46Hd7uo+W7rQFX3hSnO2N3FsGmPoPMtEa4WO3vJkYB
9XxmFMON1Eiahm9bdYtN9dqKaDpeHGp5O3S1gh0qnGHGbpR2Kbi4wwGl1XaYgtXD6cpcCnr7agKA
io2cetSsxdQgCyU8nw2X2FyA3pFfc0Q8Yt+kX4+zGO1BJc2Qt3iv1Zq+9ig2Es3H0VmDklRX+N18
TYWQG/VmBDO1Kmxr9JL5dvA4wB23icG5tCQLEbcDMuPfCt9VniHflNJhr0xM8y9pM+dlX4RlHyqd
X4sfJauE5t883JsS2n0TJ8+s3NuzuPjneBulVbgU8PGl7LfH9uYpDSmPJzMx4REJzt7A+NefRKPN
olRca2FWjEJTxZE4XMf1XqZmgJVP/ijA5B+JUzw2tMC9n1zINNeYztbpT4DYmjPbPIFc4l1yvaYz
zAf3bqJ4I8qDyHcsKLLDsUf46WDf0si0MzPSZ97vSxvm4AD4aU18e16Ag+uV2RBV35AuSo1nKJtL
UpHOqH2Y3GnA6G2Nt3xYfO4/N1HMelvyRHKzvixNRFh2WxCvHDSUeCppdqfwt2LN1+EtpzdkZZYZ
j0lOf+qs4yq7nQ+eDqGgnrBdSfhbZMMXG8+e0vql3SLHRROzw/tRRg0E68tgdd4ZYNOHMg9AAz2r
ZkZXZo4tpbS+6apNFh9kzL4yWFnIBnid54dSlCB8TyXxnEDh5aQTOwaDceOos/D/MVtCms88srs4
vy2Cp1rdzesCe2kSDYw2XUwhh79BuzMa4qqAfP2iyMSJt29GPAV3CvqM4FOdxzY0RE3A73sVcSSx
OmXJGDMcnec/8UZDLxS5crAX+ff0SXuSvwLoItfwibI3LKbTEYdJHojtykEkzJbvXnVaOkkN5GXF
rMcpWjJrrMzJf/36fRCfWJ1lFWLPPHKxa/iJO2dhFN/3/3obHaMzBtOqFABYPcqb/dmPDTIUWjWZ
f0WOdJP99e6UkB5h8PfXN0rytGGyjYL2iDMC2ar+vMb0KUbjM59KR0RYLGSxF3NpUYm7JLJcqmpj
LZrc+zat4AA0tb53imPbWw2Cz1JhTIRMIM4tAQcb2G5w4/K4sElzT2LzOG7lS9eZU4eNYfSkqMNC
C+v1oa3u74cC7jyDmle9QQCaVueiW/hSIhxr3MZAQsGs+sSksxCL3N7bEEq8tggPWJI0chn10JEk
CcxQuj4D1AeN7tGgDNE5Gea4NLfPLfy75mt/dMmuWU2H3OyoyW4GUu9zfFiAjJBC5G5zKaHJYp/r
EgMLHRCy67KhEOjF1CGCgqobV3W9JZwelU270aOmF59H90m2DyuLojPiBLSByjiiPsmjsYvrTvWN
XhVe3qsobPVWzu/QaRHjpb8tHx3y/T/Dlv/hNxXzrWZYhgq0A9DPvSbfkP9i/xXeuUSf2158vFVZ
N0cwENTz5qJFwG3K30ngoIEw9BsFKSxp73Al1HFy/kA4uAXhCD6Gulab0E3kaRF7sdulX28Pk2kW
3FTgEl4YmHYHAP6SG+AZd21T8rZjL/8B1RCtQ5S12z+S5tB8MYYFx7kKnftF7IoQDYhc1EGo3Ncd
JVBrbyfvYrdH59LQEcy0AaOiZDG0iyNW1zSA3s2j/RyWnloB+ykyoZHmCeCj3MIAxdWBUoE3CZu1
dTZ0DtgGC+BycMJ6pVoFX6RYcHVDgSUx5OidV1QRYgSR7cGgcIRAMQQTb8ybsv53/8i7n679Laaf
Xp3+J9fsu3AZYyFfZ3bjC9Y4kDIzU+YXk5YqwcXbwCIw9DALVYuuZ3xdiNxssKQQLj25wlM7iTFo
CG93cvB92Xxc9j7TuMn9vN7ZlNqHWjSPktsQyjQzsTccMG0mDCbYxTighX7xdoVjSmICFJUYk1gY
FkEtYJrzVmJFtniGfusEuATlsOyVwyhLFQJh9meKHwvIqPpGofDejeAbUecfgq6Ugm8Kgu5lgiqf
tbRfDPY9LRXJDl4bdcz0bnBU5wRLhZI+2sTHn197r4PkvJ1ksBh5p2IYSUwagUvucSKg8dQCUlHz
0NrUnV1qXo9qvLSP/vCY/xPP/ZN4YhVqeoR9u9C6JkGGtgUGwvDf4cx3LINDMcinOhWcU3h+iL77
i23x/bQU7W+g9riL9uDrto6Ysx0rCgqjoKNPC4UijJuGgNf+4YAaKG8I3fcE6Er6P4zK4wFz8xg5
/h+9RLYwVNNz+ES2KeXizu3fVntdpo0JllD65OPKJFLLEm4nKKileGqYILS9kdgXRPedTrL02JjL
anE9avHpZYAYyevFnWMPpM8GndoXb+bqpKW/WfikeW58AbfH7Vi3zYhQh/jfw3SRNi02EM5iBFpU
7/FTc5zhxCHSZ2pg9nVdPiufSnJ8R9u4n4q7xkKjRHauq7sq6NwDfi6TQMn/9Zcv3tk8eE68e0Ik
DGc/7saToGOCXU1cdU760kDZeq69GNl7LPUFlRca3HTo8M1YpmA0JMA/aH/I+vFE83PFSyDWDm4r
Yqa7q5fOXNVDfR6sy/8L498sEx/NkjIfpklGF3ajy8MZIIudFjqP1KPMUJQ5UtqXVYvawcIlNJoL
5pQQvqzoacc9PBZKRFSfo8Snh1oW07ODYQN0rs+o471e5GMIi6DDflH7Ei8Oy5YAblo+WQY525pp
q/tpLWtpyt83WrN66+qB+Tlg7nk4VW7xhG9BqxQJ4iBMDaUPEMEeq1z9i0+r6nuwn1FMXRpJLBZ5
EPOmozJPzZJUfVgLMazRa2VCK4oQJl8lb7YZ7bZNblz4POz/0/qFWzMwShc4OgZTdVAYuQ3hT7kD
d1XW2/EjwXzEwOS8N9FfKMG2RhID54iXnHMXwsSGvNA5h+nry9glCAWIZuhsXn9lfgwpO4keVBRn
nDPf/YEnxE6s3XkfLaZXUmMuz10UWRQy9mMBGM/L6qaFezrU4Vu+FnYtmEUCWNut9rBQfKfg2oKv
7uXOjW1eqQo2gfg0X2JheaY5Enoj5AadUQbwBoUub5U6qqyFQ3E6/EJbbYRPBTr9zA1+6opwgIT2
6YtHsVxmncBpWgVB6TQMjhTj11s8xndpp6ktpvIcKBdouHFO3u+PAYGGDwcHsvIV/llh8YSuF2Vm
ODdNoQRiUzU6dY2lo+OBl584bGmRgitXG2X0R3DHRpblLCIJBtmslRlB8Y7yboI+nJz6mqp7sgss
se/E0blxocUTb7vqPCTCI7WLlYxmnTBfeRHOKqEbH/Y/k7QAX9CaxztE7w7G9pANFUlzLrQumUra
jEfmEg/sbiZ4pEJmbyhiwXtY4SKRcObOreVwcyh9u24kxke1shTWRrGxMLwJbJoCpEKMT26YRqWV
65yTVpcs4Q8+SjMQiXQLZKZI9TPU6mDdOvKR7NWW+HH0ZxqfzsyvYDRtafhy0OXcRj0L6LYayKOp
tfi+AjdkEclaitSP+B9wUOfGJwcRbtR7KMMdOt0Oz+s8CwWMOghshVG+W7m8ooAed4v01qUwhzqM
B9JdaQiBxPfbzN5fC40tUcZwg88jeESNVFfY5isWTxHbYCxkA0YhS+rVcaG79HwIAYzrhSknuCZM
3H70VqqihKj/eymZExZp/iKHYgowe2Q0M/fSP9w4k0OJdM2dW1Vsqk7FTRVtLdDDyqqtAhOixX9P
ROpkXA6rTMUJBvjum582ROy7NK8h5Tr8ESsJH2Qu83MkwG0qrafpXNCt0BfjdXJ6jk/W65k+/NxL
ZFJC5R5vEtDhDq/NWtY75pNKKPeQfUvKXBcIz1RGKBQtMmkT5OOZ7UEEOTvsKUdQsyCOeer2Nn9V
YIB1S7F7npAvqOy+wA==
`protect end_protected
