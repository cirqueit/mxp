XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b��&�;�.a�(O���M��՝a�a�G��5V75L�ݠY�Ʌ#��C��<���([`�fb��5ɗ���Ncَ��́w?�"b��K��<)��*�+�w���?!G��j�m�_��B�#O�?�O�)7Ec���	��^r_�X�#��[p�6_��0w?_Y�s������h�א�U��󄗩D����HA,�m�2]�^�v�"��mh�je�;4o"�+��g�GF��pW�`�P8��a\�:7�c	�6�sz�1k�-��2�-��>��}�Q�X��~2'���J�P�y�a���T1z-�츮�Q�\e��U�ꃪҎ-�x���sga��Y˻�*�-�9@�й2=�`���c~� }�7��+�'J���d�엇?������t\ɡ�d	�w����ɢ?y�t�V$#��هR�k��)�	�I�,Nr{�p�'�I���Բ�#q�#��m��*�<H�Ô�� �	�[�6��?6х.�%�T����z�H�tjC�܁1@�a�D���^p��� ��7z�����ژnM��-�RSs�ݍB^��Z�����0�-Mz·+���OڢM�3�1~�;n���T�^T~0w�W���U4��_�$c�k�JRz���d�i<�˷אm78�J��kj(�9�=+y�G<a��C��R���k���ͫ��s��G���S���X'����4��PJ� ����N�v�m�a�g�]�{�48ەط'�?�!%�y����҅��*�cȎj��7��&Eg $�"��XlxVHYEB     400     180���	�Q��&8;����O���5&0�ᨓ+�`w�ͳh@Ծ���	5�˩��8nd~Q����(�w���M$G"�'b�9]��������c�~�jTg�\�?)|gvb^9���Ś{=ѽ9��W{��i�����L�\��$������ 4��4�9��s������2�R�S�#�K��G.�Wgv����s��K�:KQ���Ƚ�[�Y'�rع��(��,���>P��ʦ{MfJ�By����`c���?���[[װ~{Ώ-��`Js(hoQx'���UvHqo���Y�FU�D�
@m�U4�լ�}�L�[fڒp�i�?��)~�9���MI*�C�)A�p�閹��Py����g ��Cs��w
��8h���N|oXlxVHYEB     400     180y����dPm�yWϻ�w����������f~�v�OǖU>�ǆ�L�p� &��%B5��4�uL kj��H���a����ş�r�����b�0�z�&�C{�.��*UyK� ,�m*�BE�̯���zF�Z�;�vTj��ы�]{m�8�����\�`�k(rӿ�R�W)i[���oE�*��#�oa�b]ٹx疐FekPe#�W�?:b��6�d�`�zn38�7*�QU'NFIV�{�@�B�4�E�u�����������Es��bk}�ކi�W�� ]��z?��-rpQF_��C~���_�T�m�/R"x�����q$T뙬�e��f�Z@��%t�24�Fj��o;���d��]��D�#	t�V�@�*m;XlxVHYEB     400     170�f����eeIdK!:��Q��~�g��li��^r#@��j��Q�Uf�$�D���@��y��8QV�K��\Ї���:ؔ� �Ӌ�U��e2����?��&�<��f����DD|�֦Ѧ��І�(ڻal��GU�n�X�a�8 ���4Q=��ūC7=P*gߺ��4ɓ[����t��g��K�|<~��P��T�B_QՖp�J�,} �����*�rn�@�J���S$��+����M����0��?�M�&)���h�\��al�@�4��N��Ѯ��pV��k^#�uqQ>m�ZAC���D�Y��=5�A���.7gF�S[��e
J�'���:��8ʧT�����,
�0G�Z)�XlxVHYEB     2e8     1203��2Q�Xn�z�cc�f�k��RY%�Q�� ���`��.���7M9�J	Ք��� R�n>@3�w@�͍j��{
h��"������ ���{mdk�6�:��ڨ�H��il:�{�m[J»h_�c�k��J��p�B�z���1�������?�7�@S��3���e���R�wL!C��p��\�Р�*3S4O۩U��ǁm.�_$��:&�Q/���GW��HAv��&�}��<���M#%�^�0)lt�D9W��m8�ݶ�w������0¨h��I��~yj