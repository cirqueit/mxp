��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����~~�_��><�
�l��'�P��3~l~E�3s�nj���1��������Ẩ�O����S����~��݅�����|�7�����q�-��p,e�V����D��L�2�*ݎ�VV`��.Bw�(OÛ�{���4�$S��nwR�6��: iw�~gbx�d�<�_G�`�O�y%f�M�*����
p��v�0��Ps�r?�8A��&b�"
C���	i2�*�h�� bEp�.�m������HG���JA�����C�ΦQ��!�φ�ɩ����K��ωZ��ɸ@f���7I.Dvک�
_���(:ro�~�R9ڇA���p�"��9<g��9�	�Lsl��G00�~t��Ԯr6\���;�6�����`����´�>=�'fi6s�֣��V
2��������%DؐG�r�{=�T��7�b�-��Y8Ga"��7�l����Y���^,1}�j�?��y�ŋ�K�4�]B�_-�N��&��aR�1[M�02YY "���3k�:U�_����.���F߳�@��{~*r�	���5�Ҧ?��p:d�0ȟ�Q�J�27Ue��<o�'��UZ��Ŗ\_�(������Q�m��e�z�:y��׺7�m����,ϐ��r��/���lə�G��з��l�\v܋0�g�B�Ǻ�s�K�=���o ��z�L`8MA��H  aC���9����L�ѕj��q䥎��ݥW��H�tN'����~@R����Dw�R(Oɪ��쌩�4�����դ��p$|_/7�aM��u4��7hӑ��=���o����41�ժ��8��S�+����#	N���yҋ�k��|01)������j��_�+��C�V��A�;<�@�>��l4�V�P��S_[X�'�}��C�$�۞��.�������ƨ��11��p�����H�m8V�0�Ք��7#����a�2�$�>��)�SgZ���5q��r�j�._%o�y=W_����: �c/Py!o�.�t@�5v@�v8E��bY��@a��P9�,`��j&)��dzl��PJbi��p�=��b@3�+/�~s_�b��C��I߬{��ֻ�����Ԍ��-�& j�UGr�8#��_�� �z��'�9xǷ�p��!���{��� 쏮�/����-�c�q@(�X��?����A�p����eoxP=��7��*����VA�TIF�f"B[9�FQ2�oU�����5���P�Zv������x72��`íQ�>X~��(O��x5p�����^e)=�ϋ�uo�-��+�J�i�/��Nh�2�	Z����uL{��U��%���2Z���`"%�5��(��@ɥƌt+t��y�P2L��J*�Zo�E9�OP�T�w�����3�A��S30 (��=�L3GW��� ;@�vJ����M�s `f������G���I�x�hR,fi�%/�I�A���\;NY���9���gI$^D�L�b �iu)�M����
��1�r�ҷ�b�6kY���^��_��� ���-՟��nѬ�l�
<��*��,��:����:��0�c3��K��a��;�%k~��ű��Fk���H]��_"����ض{c2����(g?9������b��n���*AZ���7e�:lc����=�.y�+6�!�d�~_4l�� �!�Uc�zdp7�R�r ��o��g�W_.رl���'P���+�s{�n�zV�8Vx�=$	���)��ޑ4�XII�Lr�U���/�ʹ��Ii��.d٨�����d%n>o:�+x�ΘڑL<Dž)v|�^�����^�
=��s�N�]30l^3�K���f��|��ϧ��Q�]�DX=��/��-�}1IK�l�=�ni�!���������^Ƹ��9��%��a��;m�*Sp>�tf��
҅~��!<������K�$.pt��g_���xA�̖&us�V���c�݊����,��\j]�0�]б��<��R�m����<I.����*��*e��`֪���߬�z5��46��c}ҼK�>���|��mY����6��/{��1�=���*V
�y���}�`�A�H���`uQ�*&|�S�V��;����a��=���`���)����/(~y�w;pu!?:�!��k��\�P���i�bI>�u#�d�+�5lM$�A������C{���E��i.������`I=կc&�೩I���И�.nn@�M�عc"u�#�Aؤ��] �]��࠾�f�zp�u�d�#q�H��=��_T�%�0O��3�y����[Ľ����A���"�JgɇUV�yq��Z��f}ڿ�ʰO����k��
�=�
GK-	|n��D�y4e�J!g{��#�T�w��W�u��/�P��7���݆_9n�Q�.��D����ޖHݲ�Y¬Hأ���)J�09��T7&�{��(�-���R�'��_���{�4��y֥'C�y���h��7�_�<tc�7'J��%-C�C��tg��P�$�ؕ��/M<��F��fΗw4�C��(-��5K6?�"��qU��j�J�$?०ǶK�,�S�ki�c�g4��nD�n4�z������D�.A��9Q���RI�O���|D�� �$��~�/�5��~I7�d{���lV�H0X�첗��nv�k3�]��i��}�����Ďҭ�ԠT�Ax�̶���f�9u� ��m�f:���!�13�O{��7=�� ]z ��� )��^cb��6�f�d���l9�9�>�u����X^	q��E�3����r$C �fT���(�g49h��u�ϊTʵK�n�$=�Ix!a�P�a�@�=g�8�#2�1p��@c1'a��u?��}#?I�n�/�֦���\�{O},�A,ɶD�Aui��ݛ�Jsh�f��m-�T���������ja��	ǜS����q#<�x�z���[��2dg�qp#�J�;�<�N(�L���[a�ZDq�K�������]��v������ʥ�Q.�D�ieX���e���|����������l𞷀�z�vkb�.��a��[��ZD}|Y�j�<Gڻp�x����"���e��\���4j�:wU��H��"���M�����0@Y�]��U��%�\����zy,$�m�'q�����Y���1�D7���.�&Eq�PU�<�����,};o�O(���@8\f#�Q�C�<���9~��'
�G�����)Lv��6^WD�_02������22��b5j;�&m�.3!'4PO%k����ID#��2������;��r>׌�\5����I
��j�;�����oy@�~���^Z��7���S��a
����Ȓ
#	��P �gV�z7[���os��{%��;��2���t�yu�Aځ��28�f����Ri="L���Jyo�}!�e2���G����;~��čҚb&�j�Zs��m�4�Qkgz4�ҭ���c��@�UH�@����M^U|�e˰΃�&l�.����8d�S�t���}e,:W�^���"�c&�7\���ɠ�ѽ:sx.(SX��{B'�VS�L�#�� �Q�u�Du6����%�h�meH��#���0K���E=�\�l�UD-H2��em��*���Ci��8e)4IJ�d�1��w5��7��X
X�T@O���׽@�k�"k�w^�A�v8�v�S�tY���Mq�z�.���H�W�5g�.��f����[>�"{�z�6�>x)ا�}���Jb$�.s�H�=8Ή,����xxn�o�M�`"	��VcȲ��̔a&��ǽ��l��l�AKBU'�R�0=������A:C�W�@��X��s5s�sa'��+��w^�L��H�
&׳#�M�{1ղ�(�1�Uy�F~���H���S^C��y|{�nq}LRQ��V��a��9�Ǯe��[�=wG~M�H>WTP��m��z����wf�P/�"ю0a��d�i����f�!/�v0���RV�A�7c)$O&�=�EN*�\g��F�4`�)�Gف\�C �v���>Yr��<t�_c����ۦU��J�	
�(I()�_1�WTdo8�~�JZ�9`[
Dj97Ɋ��?�(l�!�0-dC��L?��*��^���k��#x�+݈����(��Co�y�'Nx�uj�� �{'f������G+�sܻR����כ	�6��*g�s�i7vD��͕��a%�^۶�Ex�R��B&[	R�j�����W��<_���8���'�*�P���E�>�q3��TC� 3�$1 �?�0�2�0&Hb��U(��	�5�{/� k�SߔyXTZk�#b5�� 0��_�o�5t����󽙢�)v�3��XX,6=�x�b�]T�j.��(����\�]1/��ب��/�����	��^`��Ne��^�q��ц$ڌS��}`�s�%�3�����aP��QEF|���qL�Ր� ����Z�ܰ:#��
��&��k,�L�b	�)�!����g�Wٺ�|���[�V_X3DtN��|trP������,�� -2����)O�t]/1�5@�T�Y��0���nr�J��FS^�#����5�PU�Q^����������[���~b�_���@�L�UA�U�B�#V����bHeb����~�V�|Y0϶ �L��M���0pjq�O/c���d���H�lpK�B��拙ǭ��%��͉; {txr&����,�KTI���JH��w��B�ZjኋH�WvT�Q�DuL&Q��xI�=���6S9��*>z�B��x���}�������+[p����������Ϧ���nʊ�Qn��jƕVUf��G��ZR��!|���l��22�	�b����R:����6mē`����Rn��x��z�`j��q��y��m�Ԃ��� �)����b����t^��<۶a��8S~f6`y�� �����N����s�8Oߴ\��&�[�Z0�??c�O��O6kw���fr/����J��,�8�9th�H}&�V�cW�����e���"���Ik�qx�+�;�0o(��|� /B���n�����P�͒)`[����Dd�	��B:��Nw����<���=�����6�������_Y�7��G�����.+ǣ|,�Yҷ�o�RP�7�N�9�'}ǩU
�yI��Jٍ�)�/�06=�<Q�*6�͛\�������׋�c���RE���t���φt,�!B9ፚ{�C矃�r��b�9e��e�λ�g6q���D�|�5tVu�D�����d�1�:Ԯ�8y]z����,���5����!�K}��$d�+���a���&7��Ɛ�<38BJ�lo'�`�<��3`��b�j�^����N��x??C�F�y�9!�+��W�\�9?�7vr~�_�Ի��7h$R�m��y�$�ԏ��콧ɿ��r|����� �O:C�O���;	�����7ۦ�~fR�i~MT+{�0�tՙƬ^��`ޢ���c���0 ��D`k����xaQ�r��.~�t��6{�OP�{ŗ^K���Z晟�d|���*���Ϧ�B��2�a�A|j�2]ʅ�����q��|�ѩ��� o���5�$�Y$�@Ԃo��:��N�8�.�G/w�W���:�J�e�cM{��b���6��-��h �K�$�����j�@[�EY�QX��C:�pB���U$B>ݍncaf5�ǗIր�W[:+;���$ϩ�\1�zP>*G�5���´�f|�y�-;zHR�8���`i+ ��ƅW�
y���@<d�oO���|�h�G7�vc3}fѰ�9��OYAI��~�z�E�l����d$�rF�ΰ�*
��{��Y˛O���J��Si!~M���߾���rD$�Βz�.$��Vͪ6,e>k��l��.�sR?�LXҟ}�q/O�j#�k��l�>Y"��d\�>؆�v-�y����q�A��9U�H���KG�V��+b�?V��4�C �[��1�i�LA���b�^��,x��.c2����X��ʷ�2�(>��ژ�`�%�=o�Y��ȏN1�W�UwG;r6�^(���g~�}��x����9��ZK��t��W��{��T����DGޛ#bzhp�9r,�І�?�PX$�<6y,."�CmܶR�h���n�M�� >^Z]xJ��e@!ܓ��G��N��%��"�Z�G�ܶ$B��i�(�A�MM�����3Z����b� �9���NŠA��k?a#2a�F�A2��|�,���-s�p��b[�ñ�45�rE �9M�(��\հ�t��t��6P�"}�!��5��3����z���[��6�����yS�e��4���W'���Du�k�G�LI�cU�'Cd4vޑ=����͗X
�K%n#�R�;I)���|�i18�Æ�2��!ѦU��%�_�/�H�pv$������'�D�_f���#b];�1ff�1)����.˵����3�
QJ$+
�7nS�h��w� �����C��q|f��Uwv'Z߰fck��Җÿ�P�ofθ%ϋ�Rɠ'lu��������eZܫ���|��Oix�nc���*�����T|B���rD���oIN&A��z\��:��F�ťc������3zg��L���3A�@]����).G�2����b�M��b���[l��XG�J����L�7��Pv����(��gΞ:A=}}v��~2�+��MQ0��
q W7�s�nC?97T�ݽ_B��D�(�Q:�\ԯ.�{4��E�l�D`�ۣ����H12�SC?p­L*P4C����Ό`��g���Zv%ܛ�F|m�-�#���M�_�Y��f^�7���uZEΟ	X�t�j�pj�PU��(R2cb.�֛)$�Ob��1�mn86L��=-[�����0���.�f��K"@�����_�z_â���_�z������"�|M;�+����Y����!�'/���i��-��s:�e| ��&T5�ipI����o�I|T�4����fj��V�}�Q��D)Ɓ��j؇|'��-u�Vv���]����bI8�@U� �P�m���(�}��d�z�T�X����%�聲u��a�YnG��Ef�]��l}l�*��Eq�],�a��2�بv������`w�� �wAZ>�2��O��๥�dl�"�ީ�_��/N�L�I5��8�*�/�=,�x�4f��qi�y�G9IX<`�bٶ�R+>ep����*�\
V�^�ja��A�	������gJbp�T��-~���㋅TV�d��c�EWr�_g](�o:���R��̛�qG!�RV;ɈW���h��E�����4Ud�{=�w3�H��dfU+�{q }{�D"	��j���v����V��C����-�=γ��Aӷ ����K�W���")煓.s����9t�^��ܵ�.���E����sV5�'�X.z#ʞC��"-\'5�C���F�_�/u��շ�m�7�s�Wn��;f�R��%��͒��U"�.D�Ag$���֏������L�vz9}������.eK�eu Gl��[��Iy�b&ۓ=bŲZ�I"D;���Ƨ��Fny�;�����k�M�d-A0!��HĘF�dEXԞ*@i�d�*�vW�E�U��[/�æ��!@��d&6���bn�>rI3j��V������yYE=�0�sء���RD쓱��ֶ$}�)E�*� J�93�D61)��������������"�;�0ǮyՃ|�.���7���w�(;*fE����~_��bQ7�q-��Y�g5~*�[���9�zP���Pg����J�`c�O��
Ŀ�<��|E���3ο֨W?(�"s�\��\����r�� �ټ��'����pu���ʢ�b8(�O%���Nͻ����]&:R�6���9b3/�Q��Y�ax�/6�\�A1�ƣ.����4��7�cXʃ!CD��Z,����A�!��?�Hg��i�`=�H�S鴄*ok8��4�N����ꕆ�� �gNӶx{�;��'dǷ�۝����-Z*3�
� >�[���Y�od� hn��yq���q�*UaD,lB�Ȍ�ﭹ�++��6�Pk�)��3\$_�;�m�A�ܗ�=�Z���I����*�
y�*��Ը����������|dku�q�8��&a�"��LF�M;���Cފ�,������g�ey!�*Ϣ>��� ��� ��K�>����Jv���(�hb&�ֹ�)ܳ�����CʣE	b�1��~�w�{^2���Vy\$�����0L���;�>�Vi=���1��A�3�&��vx�:^��֎f�ӕJ�\��*-&��2M-����M��HOm�F0~�}�s��u�����/Y�Q���Ұ�,�|�6 0��Ӝ�\�*H�L��R��}m>D�3c����4s� ���J��2��f���qI�Pn-�逹��B$�N����^$4��BM�R���|�`p��Y]��S�	*������ fj=�:�ʁ�p�a��-���j0�lQ

���V�b��䮓$��z%0773�=�v�����)��Akf.�Bu���o�Oj&��u�2@�Ww�2�.2}�T���]
��7*W�ݪ�7�&u��jH�J�è=3���B��G|�yWᒔJ�x:q�����jk�����b9{������8>��2�yhv�3����V��D!rdc�)Q�W�ת�*�Z�Le���{T�FNJVvCAa�5���v{��Y5�;p��oE����p�臙�Y U8~���ۊ���!9�bB��0GME�x��<q6��lE;_�19��5��چ���}�A�l�jj��aLMJ�߿�z�tW\��X�n�����������0̹�S�Q?��8�#�X���E����yA|\ZFDЛ��=!��A�X �֨�X��Z� �r��j�*���sD����ɟ�Kܩm�B%�<�\��[�I��+���s��r��} �R�*���n���+��;�]�|>N��3Z��ȥ�l�`#��#9���^�@���&�Ũ�=�?ˏ{��DU9��l�.Rgՠ��7!@�X��>��ѥqhM�_��&���:~���INf6X���'�]�VƐ�on>MN{���	5곟z�Ӻ~k;�
��i�x,�,�(�O�i��3b����X9�P��1T>߿a��9�P���F���yT*�!�?��:v �~l�E�7���ݹ�wr=1%�o�J��a�B����Ϡ���,�kP�AJ�SwP�4UJp��HJ��
`m~T�7߭FlqX_b]���
�N�.�|Kg#e;ʎD<N-I:��x	����u���$���wf2����g�O�����)�{��([�����F�����#��*�ybEl0{��|on�0����^'K���`��:bgq�9�*4��z�+������ʜ`Y����j����T/ۋ�5$�U�FŌ�9Ř���)M�<b�o��Z�7�d�p|�+x8\@L�3�h���S�'u���<���kMo�^C��}0�'T����i��@�!�QBg6���i�9�-���*D&��)����q��~��m��M��Y���<Pq��׮sh�0mTӚV�������G�*��{��8}�Cs3ٛ���ll���dN6e������n%��A@&��D
�g#:+.�?�<I�R��2k����_�I�#��?�opB1'���,�� f�J,ugk��<ϛ{���zΡ5}���COwuu0���W(Eo�ot�ݚW�������m.w�f�>+�AO�}�<�X-��=˷����)fz@z�̝���jN��##l8�Z���Up'X6M��a�>y�vy�w����UER\�W
$�y�Ӎ������4���zE`�1 0C� 0B�N���si�Y�E}e��_V���n���`nA�ޛ�� �dh�d���!��ձ�?r�S0��k2C�Q��T�X�b,Βۂ�>�G���D�ă�R�e�U�)���~�gIYph�sˎ���� �M�p����A}��>����ڌh�c0��E�2d��IA�ѕ��Ȧ0��	"��u ��j�F�(u,s)�q� �_��k��<�+{X
��@H>�O�L�4b������s�|)|�Q�� �2����r0�LJ����8'��K�p��Cvi��9[�������ń��{���|�p#?3r���p)rǡ���?�~IR⻿����
ƃ�J�E,���X:V���SD�w�f��'��a'�t��ƬĴy]]d'x�u7�>b�z�X�W*Ҽʈ!��ؔ��{��B�˜�(r��Q�זBn`Kƶ|�lO]VԼ�&\u���P�?x�#=��4��%4�c\ �R���ryO�3��`�����5j�3�[�!J�w���G���������b�?��'���̲�������!�-~n`��'C�%�҇ܜ<q�1��@���䟐Ё̽;����uנy�;��0=���E�9S��F>�K���ۤ�îVb�y�+�Cz=,�W��A÷��]Ye��f�.���nnk#ܩ��c�ê�]�,)��>�Z�b�m�KވWU�CD�2k��hʚ��i�t��9G�&GЄ��u؀�j����-WG�ő���i�B\W��Ù�̱�wR������e�=���