`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
dBV11K7ogZtwAqpnbmi9RCV7PtdnHEqs6CkQCwRSXMH2wBn+QhKmc3DXgVyBQ1kejesogojEAomD
kkMJXs05q2PwImJCa5ibv2xmlLTk04IrU00Dq5I2Vi7xe2WeInzC/4sv9053oOFsBcgHw1z7qpAD
dHdfaI4mbFw/S7fHrd5L/3+w21OnecBZuRbO155KdMlHZx3yljIkZypDXLnsYOca1GeG75ghvT8s
9yCqmigueTWw6803/onuf6s5gPu+XAKqQE/cJrbarxx3RxmZEJWHRf8MDmdv46PkAHPJytxj4JfF
u/mzFeBqLgLtR5L0tBVrR3GeVKcWZC9sILmqJ0cZdjsR4qsuxpJl//uLC/QKpxVCnoiUMkWzgxDK
827bMwU+wCU1WvZN76PSnwQ2lXZawBqOk6WMpSz5YvmhvankalXBVREEy93VvsxJER3fy6lKeXxY
X1xZEWjaKKd5qkuVQGHI2zedNrlBb35apG3zSrvbNpoWJyg/chOwfiqSIx/4BUxDnZaaZBjZG2xS
qbkEkvdgSAaCcP4YQ2ZDtB2V5JwRKG7lp6FXy/Xz7YgstXNQSqjlnLGCpD0FFbkWPHdTAuTYtaNI
RHTshTiak6S0bhgxzEXW85UGp8cnIcuBioQXhHahHE09NVkANd4pulNIAY0PXM8X35PETjK3fdhg
zbfX2f69vg+U+65urn50P7lG+kNEiMQTW2Odyl4WUcwBl4KVjTEQLFaMQvCQ26L7Tav8PEvpUsHW
o20vu7aIoZZ3/nBoxl3aYK9YwlN+cvLyovm+DAwUUScXpGds43Sv1N0VhQJu0BS/b21Bw00pxMg/
gCGXyihSMk/nAzxO1E6awZ7KK4uycp6wPHB4sUzOsdISj7LpiPbTJlAnPGYyJx78o4qbPTnhr7zo
i+lJV86e77R9hyFJIney0h0IoaEM5osua7JadyjqBaxNLYKJZkvoCPDdR39+etTxPedS41MxobIT
TL3b5pN/4IOXlDioQKAHJOUZ20oJSmT35/9F8C2aRNIPqM1tfvmIDmvoYo1xoySOujBG6DmVNIAI
qlQa4/TBDUXUGTafmL41JQEL4t2Sb5YD83Y5CZoduGw3Al90H3i/lulSbHrmTc8RztyAiWaozsry
TRx5U2rsT8ZQEgRyajvhFj7Jhmb+3da56/9HneFCjLRus7V9bfdghYDqFE/2GCf/LHVlksrjJd+7
CjQd8varNGfL23FOj/M8RQxwU+cD+FEea8jYbwowkCi0efwtLA6Lh6yVUZGUxOczgq2gYJrq+DEg
7jjGMU8Q/Q6MQ+saubkqmmMY+UkGjrcE3tdx9lGu5n/GBw8ZjsewNmZkIn2mauzn9c5EdjyYCjbY
qz0rttYOSB157aHoKv5jEq1WjivNLgf2GsBowg04TmL6abhUVKS+M9dINhX2F6aTxJPPdNQK1ZQ2
Vr1xA7lRmhWMn4tA+Slat3LhNSgk0FTAbT1MwmBPwJxRoreCcP+dIUW8T+JqGnVKXyje0j4dgQlh
z7s3Lnekp+CXwvT3+4VpSqs6MD6Ud9tG82U3YrqSNqb5g1m91IcDBpiucK6h/npI6h5aH6aiXwPJ
q8+XCZyrFohAAxNwEm9xB9R8nCzIUSxNV+Cqq2ViHymEDOzXlgd8gPWaV8HC5i+DNsbtpeAN8YeJ
yPdxSR2dWsdW6hqnY8ootqJ6NBl9ELMyXzpzo1nwizZZX1TVooTsgbNjOhfRNe+iih7sE+Nejflg
7uIqRsK5uKM572H9cHvcxeRdpTMs18b+2/CCs5k7zk5M5ixG6B1IINe9PzfxfCInCwvpn7vogb3R
CfPKCtjsA4Cl934+VRVGrPh4ha7fgirOh0u/M+vImxwvg8XWl7u4JP4eYFsdCKXNja4n3srLzfo8
ng7uu0SOj09thXlPfqDAQYQY7sl5nWW19UQDFLfN4UcHqXnX0OGmw5HbfPb3fr5/tjvTpVCTxf6X
9/axGvBFofX5LQtbbWcphcirIswI4NkzTxy+fjBq/orME3vctI1OGqBvvEqte33dzel6xfh71l03
gMxeqWw/FscxDeR5UmUhrHYIlHgNvRptC09WdEK0NcSyl4vYyR7bRAI75qotScR4v4lWLjOxds5r
1VuG19xydDZxBcJWchhmKNCkd5QuXjGB8UpeMbDR3gjlBNr+WWK0vR0jUAd3zi+RadoRptId+L0r
Eu2IwCw8mN6JNsJu5lLUO/2bXQut75JJ13Hc/whdsrFZmVBQNWDePjjSMOJMx/LTHYUp/a06f7oq
gUtYjhswe89H3lZYkYZL1ZJjWU6c8iYXP9kqBpQ/3Z15Hl90LosFlplnSagqbtmuA2k/EIXvsA8U
LKKU16sdU8bBlnYnOLeXs+btZLM1cKgmRHntY2BCSJMSW2eFGL/zdgLPAtx7L4H2E/hFvrYa/W2M
ffHPHKPEhrbsWyPdu2fYyVRklgkvupkNeh7pRhZv1oi84KwBaD64SBvLhSmUyAqreRq5IEd4RZ6C
JEBsBRouqeagQfnh2KJ0sv7k3yALeIL/VAyX6UUFeWJTJnQS0IaVnNDdp8ocU8zJtjsF7WHS84S8
LnA97FHa4FlavBUnld++dHVn3jsmLBktEwuar9r3c048ke6ozluCjgyxRZr9uNMPrSnKL8fWZ2b5
44haeSeJb+eDvBipOPAj4fgeonzeliTJDq6gSxO5TT/JU+HcCgJvhxk0DNLgT2I/dPCAoFPrFjSc
3O4VDBnHf6MPe9UecPo4VQMQrimvTMDyUQoJkHjbu5wQPbwGZFmgg4kNNxrk4PxhpQZos1vX4rjS
GziBli90j/b7PStaSlv0UEvcAlumfNrBvMSG7k5IFMXIpPw2RR63QubZVh3u1CTyqb2xi3w87KvL
YBnBl+1YPAVFU4OsOvFtEfNZ0APS0i8beDYNY+r0Hbeij7rT/6y7JIBL/xc/WtQ08jI6LlvrQDjM
YRKySPe6519EBgZqKbjnXfYeSA/EWPpthadeWTKK1rkcqo9MhnhF4VQE939ziYXaKXUhzFfn2Pu/
nUQaou9fhIqjP1QnwWa30ClKEWbMlHfeu50jM8Vl7EXDoxPzyvLQHQp86LTl2e8vTxaazp+t2zMQ
RrD73Z2zQlDpAfs+SmefkhhXJy7ihWp3Ku26Wyr3Q1GaXp8l1WXBe/FwEAbiLHutE1PIF7p6FuoL
x0VP5B/t5c3A5DXCmTZYKXksVoJKjfKp2fTi04aQ8HX+xbW+74SydldMJ+J28GWkI2ikC4O+DC7A
fna0SSlLmRgjlhrMCpvftPIu8c+qh41utIu9BK++dpJcy7h4wbmrTchx2BSy4dMATQwta2KFA+Sn
9ZIWS4BvOkICFFBy4DGNHqlM5Am5Kp6JYzOuOjZO2iAZTjsVcQigzu6ZwzA6yd6WcCzISO1NpOi5
6iWsSP+1fhm/j9RvLSG2ODQHWdgQIZq1MqpF5LqhkVIrVQmGwaIzhxaQUnW/8LrVKNwKBSNylxUW
V4lsDLbSje5nkN2eeQtsYXllNiVpTSJ1sDAWjaridrWM2jLoEmhAQgFSjDP1vTuNwRzFJv8NWqyD
vG15/dwuRcIwj9c1y6pLxZ+cqOUUFpiTHv3SlNdX0vIlp523NLvTLJLG0IfC9d7UIaJBGfbAohz1
+J8BQGqMGSKO+VjlayZywJnnFkUlJ2qzZ8VprQdJ5R5atgXAdrlJt3CsvXHtFbrM6mddEkSSotTU
BHxDHLoyl3XRwghVQNoYBzHIycAdsH+NcDpeeAcswwfDj5k+hbVyROTW6P8Bm9k0f9VVldtmXYWK
3Hp7JA6ncHuRT1ijmuX1rjlPK5ACeiAphDg9Z/35fMyDbK8H7C9oMkvEz3XGjk5uwxTfIOmaScoE
m0MCkaOmFnSF+FOXs6+B7h3/3SA0N22TkDS/AVSSCthap7XL5KpuWmWauOT4kzEC/cc45spA1XG/
b9iOUkZXFRlm0mHfGvLQUV9WjHDt6anJsaSYfDH0sM6ajF+XfpupSK3GFQTwU6V8BH2ZiG5cUkDm
w1t8jVZoQAZQSA2fuuQ93dbIWr+qm3T4FS/FBLTc7bOB7k2m5jgGKROKlt0ibAN1XRyT7you6UCm
Lu55mr+SWZOwYC6+EbFfwtjYk7mJGIyE7hMCNOkNfwd07aw/bU7/vfgsON4zdEuyKtBz70NWtAfN
yO+hUUd9wht42fG0JvHHULFbS6pYIa2eo5Xk54O4I9//oHydaNXryPoSSX/ZH1Nt/nP6P06SoMPq
r42zqV66gf61OKO1uv8qgf33e/YZ+4VfThCAlkQpmz8JDGsW5qrXn1ROFGeNmN38gr12J8cNQZDw
qwSxrDahUoOaAeYfC2H1r5dsg9+vjg+LrI+CqQyGtFcbXo5RCz/hxE2vLuVHd7k2BiOQ32pW1ULu
/o2NsFtO0z6SN0cFbOnB64UOmWkxpXYM+Cn6C/xN6ac3Bk+43AQNqYFETU8ZjI5Mcz8i261QajG6
klvo0a+mnk1s/SCSGTw5g7APHdxK2Hih7UhA5CJpPgJLZ0crg0XlTidMtz9aJPolgG7i+/lA76w+
dCjbY8QQ2F5waPeGt26Jl0dTbAuFp0Frj7deEO97fWJSmZcOrkZcNe0TI51CHOzVvWkwR74bJe0Q
lFpzHoLok48zDaAhBlUERM4bp0u27dFmYvcT+7z4keQNNMWGm/x9N5g0+gTMKdJFslNjwJjHsN7T
dXp1zWvnMd7slExcFJAdn/36QysOytgqUw489dPKPKhJBIj5Z7Q+s6jUq7RdSqaeoFnUmLMBFahl
suo0C2NcfTQWGeRXJYFefnHtxDiXYhCNrn8Ug88mFZEji4VCmrPjk6K6tz20RILvX08fGgX/ajbb
5bSpaZ+fHzYLlylr+kvYQGLW3Jk8o0oZjwJ8H3l9B+WmUJNl0Wmi1PzoFNDudx+iaa+BEhUUllsz
ZknedEZnzLstkzfhKfATo/zKi4cOCe43fRbbw3+VTqgr4T29CmuMk63M3LpjsRu7zRLxP7xLzYFF
PKsnvp8TduHxOgBMtNCNeS4lENAk4EGFIt4NNgN244kksxvHrtC7G5s/98jav1oxVPH4x1rfs3Ph
6HI8c/RaRi3OenMEJPeJZMA6MK0BBJJodzp1IKYPBcHvVbcC7DzDtste8ZxWUv/sUG7foVNO4zo3
ruf0WAfXGXU1ZJHELsepcqk5ZGdIbXRobAbrt4f0K7fGwxR8cewCyVp+BsaLQqPXf6NcaJ0Ms5WO
bYtcMlWuXcE5nHICPwho9rlYpSEPYOE7KvLDk80LrQ2N6Z+B7Vvu0ldU8VrLEfxAixrqa3dGJBOp
XxnGY/WCK421DRFoSyQYH1MqQLUc5RB/XHp+f2MSlZbT5YQ/QL2l/7sutqkKlT24lbR9B7T/JXGb
IDLwXvcmomYwYlTEJjXcgr1NlgfmxhZPRkSDvfougywUvOanHEY53POXL8TDDNbWXL8K3euNikD2
B/T9gTYe9gpHoS9SbQ4BKiiAjBD9mkLgTL3bdLirj1ntrUG2ZO/UpoxtaIJwPesEDDbbZnBuU1XH
zxo1oW4v3cIs/yQUgyZcSJOMhJXorKxL7PEARgDN5mLkebyj6xKTcTYLRHharYvz4iJsmsr2bUXG
qrsoWVbHChp6Cfbc4GgVI1eLhQn7VJ2AJYp/Yu785Ru/JNdrqGq/pf9qazTqN3R2DKB9EyhKlrMx
7XrqemdkEdRwIPLgNTeU6A3fcGbXaMSohbWN0tRe5TT1mGDOvodC0yKwlCLw7CFuGAmjxOYOayAh
aAhYe0VIemf9/TqM09LuV4a34fVlq5WnzpSpHANXPO7NFSInYxrxMZa0oqC9SzNoY219keffLTmd
ehZbcjlhbtv5D8azdkykmDzqo/ytxgqWUNsDESzdMF06+wcAS3J9MkI211B6Qq70waSSzMzZ0vjA
bd58y447b4HC2ttR31e41n9ee1rl2OX+IqjCBW3HRsgsN1rY92wpoLePEUlRsCuE3qMGJvQQ3Eye
VwNOEqw3lg3MdBGVZhnezEGkLNqT/Gyod3g3cXKgjWVbUi6iIX7kankliByiPsir/pj2sA/1haXz
eXGEQa54rLBr/mG/qoPDtfUM5KXshA4SxWvQp6UlIhZ9nUVu4zLHLTUlK8aNK0Kr/h37az5E82Ip
/G0x3cNgucBNIa8w2SHTw4Ma8yrATOJvNMfK23Y3Sv2wk4CBFVqfWyDrk2KQDreNhTJvGdIDIoxT
xnYLuWZ7MAnXoxJ+b6NU/yN4JIUOFH4L/kXUPcYO4J5EByvK/sMfsKV6+ark49Li2aiK10Pgba0f
k1ka18TgmeCKlG0H3wDS+bmjnvKytLtjxcTU/ZBjM8rjzY2Qa5ykC/GMpu5/hh8cNHKujdGma2z1
K0CdjrkUCSqROKYoMfTyXYMxOfdc5YOYAcUaCREWnYYSiMpJwml1fwOEj4tTaByUfj4IlljYWsQE
PjmGeJbji2fTTz4fL0KYUBiCXuAby5kpnx7gMeJmky9m1LF0kPF04JjisEc8qsBIJMqZgJrcvXPZ
pizJ2sN8tMRTOsj+eWoczKrAwueciQBCq4KXNiCJPMw/EZdXHBvajtp3Dsh4uwOzNOCBtDVzapoN
sPOnAhfbHcg7uefafe2uTt06t4b9VSHbDWaCi9Yg2yv3jFsfv5mRl+HEtwJXW03KpKREMi0ggV3f
FcEthTbZiMjzbBvKM+OQXznQKji+lRtoBWMIXU6erWj5AruTJIGeNf0uDgmVHoXffLzTYiJsTIkA
G4TKc4LScIJWfm8fGKK8rRT7Z5BbxPQYdUTCi1AlyNdVF6zAMLbek+VgABZR76YohNan72qSssNi
3UfOxgGZIYbKhJ4FIlxEAMKqOG9A0wDvWjFlZSaRFb2UzExfDH/7TLhgKheGMDaGGToM4CbNtjpC
hMAZd0uJ7IbyjoFb+oIdOIM/ZMxgHhPiwtDvDYvHQmUZLg8JJsKPAoc3mEPu6Bv1dwNrSphq38WF
T2ccmubdcJaeH40tiYrHtptV4BRAAXpOJjFTckaThLd21XNkWPagR2k7KZPZFOe4AO27aQpFIr5K
W9J0xbBCdW6jC4PceshXCvYe8LrNMWWQ6fZE6q2Jf3ciREcZe5q2d2JkDMcSDmv0L7Gf1ECqDB4u
DbNCYGLrGg07lS2E08MG4r3BaP86+bed+2Cb/Fqbk5UOI5smYJLeeZF2vkV9fod0EZ5IjcDb2TH3
CWzCynetMjVlVvuTRa/t7U1oMWsLxml+uqhe1y2ZlIzv12DplzZ6htoMGLMld+YGtRRJyH/Jzzan
iLdm2HgwvHv7lftJB0cvp7MeRakJ8KTSJrTwV//FuSMi+LQr7ns7UDw01fSweSVxPHBuwZ11AYyV
kR3dEUoGOjROhldhhJ3F4XCQvRTAeU+5qbIPN1onnUYqr1UZLucP+zbA9RDfOgz2YPBdHumM6V2a
bS5A6HYkigbO4cHZ7xPjupgDR487NKs03YSXMb1YPq65x0Qw2eMiFDj/lBl10XUhmEaoOP2COb/r
c/fKgvJg7UL/iOPGt5F72/56rzYjhfspEROvZRYHS3m/mZsWg0sVEMb/GzzGFg3n2y5SibLcO3w+
WqaJ5gY5Y4lal1ISsTp5TdxOnUOtAIrjsFEEGWZJT/H3F8eCLz8SUsAVgaYIAa1nCVfMkMOJaLdp
YjAIr5vo4+S0/gA27FavcESrBoSYbDrTLn9mnnZc56QSQ5K2nYjRyZX8T9ps8moJhUHwMJ4vlr1q
b64kwmmMIlJrsJsVdIp27pS1AHL5WsFQskFZYDa0kMe35RzMJgdvo0BPsC+DCvxi+V4BbIapvJvC
pEC6yc09K+ERNRzdd9sCdUvMwsVekm/xQwLXF1reW1HYTW19Rw20UL2pm5mk4WnadnD2VkFCd9Ln
I2SqhEbGOOMpskKJFZocA9F7FHE80YQ9TQG2cJkEB07OuOeY3iPua2tMiiBMLbH1eiwRRTFu8Ij/
ajY0PyYkeXyzpCdDmypT3zAKQ1lFrVyKu0TCHW0phdfOxFE8erRSkXhgqRK0hjmjsqvQWP6qflvr
LMG52nntZOyi/6ovnEBqFDrmyQ6WdcKvO7bCyuJYccccHmlXcx7BjN7r8s3cbZJYBO0Fk1imAs+P
gTm+Ig+Zw9PMxVz4zQg0099bAvUeMIbg0kisXuoKldbL2Hgzmo+YRA7BUDEtVDii+hBS6Gs+BBtu
86KWrZB6Blnw/dOak7mwgyBu9NY0kowrg7GIwtRKB+BRdMA7gFkcaRuzcXomoj31w4iWeX6y18gG
tIt5jyx9Ds2EUKThjgOrw/WFckkUOOlMPz8XaXsBBFx5a0rfOXz3uzqI8sif9vZZVokL+bbKXPgq
ytxJClpl22UIRAxCMkl6IEW0eK6CDx44x2WKsx8DXbf5c+yfTvHqkvxf2gelU7mluvYUd9k0n6oi
i4mBoP+3gKtIF4C+XMxCNWLtrudOua1Blt+W0Y4ca2RaFDM4EX38ekjuEeSscCawnxF8eJtatqKE
OPZXb1tXtPqy4Ipmm2Eml0ERB5YLlbFm13PrNNUjoBrdWxRVxz7v/f3T7pLNKLrAC5Rdz1j4TWNU
FWCrXU2Jv+VaHhWxxb0pUeA/xYh010WyQaxTGC0VofazOiW4ms2bC0zU7v3dkhA45AN7ngGRMh/l
IGqUOQdzKDSEnesBo88aOGJrbNcNSahU6pnFFNiLSEB71eG01By7xuE9dyDefy255c3Y/gd27RSP
vtxHlnmaI6SXwBpyHyvqQYde8eyJidYaAeh98dQU2xfs6l7DbSD6Q4qK+vHb/7LKM8x7whkL22J5
ckOOThB92cQnTUvQYOYfUTIpD13/EgnJXdRA66Q/l3o6cfiozJBAxQTCMPLrTvRGtgmP2jVh4TB9
gsOASbYzWCr6tnSSlo8n/4StPpFZ3uxq7PI+bu5TCEr/MHTj4q1prtu6aRyaozF4EGDhwHmYfZVD
/3qqnUwHfLlojnASWqYjy61/8/GGzN10ccxJjq9qa78n52wcQE2P8HYqFTcLZIHOpDLrUVztxz8j
RrGrX7J8vNw8MtAGns5J9XmpgXysICskVHV14RZGyUlMaMuUM+xzwYKjB6SakmuqWIEFO43Rv3Hf
fo6T5hAnSKjHosLNW4BB6N7+uXRGj/+NaVC2sqRcwXFiR6mb2MuFU5A6exL5mVtfStu0wMH3khvZ
2XppMJKin4DMipM6LV9kO0HyC4QmqMovo/9XJxGABrMvfD0LeZ7mfI4d8B6McmWa76kioYYVHR9s
YmTdapdupTbuzlaxUtFlqPewDo0PK0vrIztz8qx0QCodYi2wvY2ROK1WjhP5EGsW8j0YR9WLUUhw
qavLnVJ0HGCRdkVOPiuOu9Ns++u/ucbU8HWHSb8q2SFuuOGv75qOiCE8gVRTo4vP5vWKBhZ5l5um
ew39vr91kO2kyrRK1swRMfZy/QZb8f1nj55HZmDklvWOjkxLxXVjUmaABLWEg8s7w0rAoVTWLHP/
fXdGbcLl0ssxgLx/M+QCdhTAAixp2ILxUtwOQF8PZNJ0yYK0G74AGoY7faAVEQ9p6kL+/TXAhXfl
LFp0lkjpW+s3a5dfZZEEIPabI6pgo7r1Iqxtxl24W3slMCXTPTIJ7+qGp6VrT+UJFOKIJceVjCc4
kMX2zvc8/iaxUW/RfT6QAJE9Aa9471xulCad1uGbwISmrcNfQOYOFVCpYE7qoLlkWL38HfyT8eMF
YlxipKaVYNBq9HhiXafkgLCct5LOj3yGL4muNFmeDgFVDfZA0mclc1Orw3QHbTNn4YISvkrMqj3M
BOs/0rcy2BLUHVTakO0wwsLi8K90a+BfI7I6Tonu+fxwnEUhyKLDCSTWw2yg+3SAiXJmQ4O4SoO/
WRj7baxd2HnfpnU/Wam3AhQtz7egirIhpk0u4J8c3zRQ3fpgTH1K+DMIkN7HVyns/gVuAiKqHLLw
jgye9mGKl+Znock/tCJrTsOM72WmpiBRCmr8gKAtfF015yXHUnpJhzGDHvvjfafKB6wLCM94axID
QyTa2Yn5YfLvAyA8vuyyjNIE2MjSdwmS8fjzElmTwhjqtWyYQclH2oaPM4jv3pFhp7uJCuNcT/Pd
TKvcj9FjBtQNhstKCCcN4yc4a53RG0dXXAlbu19oMGZItIYDjTvqEfGQbFDgh1iOiHhqpfeHoZfq
dy9LPLdQYE7XKKFL0ivkqn8ZvvDpLAVnIy/9R2xi6nC1ZYIlGSkVg/atf0SfC565586i/6vo4p6p
vzSK9q/8zsB8ZTNGK/MDdQJiN0h9l3w6cDDIAJ2V1FTahrd0gdCcJV4r8w3FDroRI8W/mhwDwhSa
bkvfGtYEuR8kL2ytDSUSvZoLBnkCNRYysBktrFVGHc5j3BnwNCgMQHY9uIhXdYGC1z9TM9GeDFcZ
IR8kes/+4bxIQ/3rq+AzZbF5pmgrQW/5DPbcfmM1neeo2OmY33fXhbXrzO5B68C1lr++GtgZ73WW
vpruWNP310Rn+DQN0YszgayzW0EuW5eGq6jyXbm1PBtc+QxRmWszdub0g8mnLpmMm3bpkSAANr3y
VAitYwRouhiUcbweaS5c4UTUWU96HQODSXSCR9Y+++oLKZdrxRU/1VPXWa9TwJI2ANueR9nbBz0u
tZkGlt9ThYkj/ZcZLV5NWA8170GKVWb2uP4PM5FiuAr7CuPhL8EQ3cc+fE+RCzKZAzVKk8b2P+ZC
L41nVRSLHMYLoOzY1OfyM9N/vzspKNja4EhKAFx8oC/RGKIqzXws1J8YMoEn5/cPOsi+AgJ2uILX
6a4biKfcJsoAckMcj7h8RfW43zKwesYl8da47HTydAxS+DJ31K4bBhJzmFwtDxmZuobIQcE9Y87r
YXSa7VjkknxuG+rdoQVmpQLY2OM3w7OoBSdZfhWZcKK+OUmIaq6rb/L0EcgMfsqR+DUxHkjJLhbP
l9EHHNj2SiMpX/jjlt/zuvq+l+uJoIqMU5Da9KoKDVm5RFLEeVENmEPA7KA1EfxrpczlHAlpehlG
OLRPF9jhPNkDlAUlncU5l0XVI42pSoKSmb24C6wJ17dx+f3BVeCiLQbOV8TP9I5THq9bgbzuYxjc
FkC23sTv2fj2RhmBO4G6cPiO7m/2iUKeayfU5nN4IrbZsINEKQ7K1EvUApWc41/I0hhQvt7nkkw4
LD9xmQnePVT2BZ7nLxYbHvY1a42IHx6ZLwe7rdV+TSCqkc6nY0ENdyeo5UwLT54ePAPfeKEzZyx6
W+y+lLkMSbP7VncYgmTijRW+SC9Cvk+FLdpGhOmlflgIZkRPkEqDVwkTRb0TpdSr6pH+o/E5unVM
womuV5hnetGH39Aon4Drfxej1vjq0Ty1dl88mERsDhlFRZBfcOzUamgSh+t64FTVCCLvad2DrBiv
50m2AYdhvXLASpIfiOwzFbKBamMefmoE0vauE8oxngsZdtFOL4dDcdl+Ege/ozZUIZ3To3m/N8kj
FehDR3H7L/W2S54GqN/Q+7elUztlyWabSDT+xKq3Nd+/0AslxzYemZPrUfYpvheNWkyUE9aItf1m
rMRaFhYFovlbDB0QV4lO+MPIdjC74TKsZDIVpAo+RIT4De87eWYZwdWsxYqYMVc4J/r/vVWLiqvt
jMWRGsLhiim0zDgB9+9bwdwXYDDcn/Fwnzuev3dZFVoyfBDYm7zKlH+GaP0jviAduy2gUL5dkS0I
NSSmf8ijJHfFY8UfxAwJVM39LNjXquUe9/1UeihlDM50gvXi3C5x8i8cHtvGVwIjVtuHBPFMtxvI
qkxzalsoejIXY5TRSHALmgfoH2wpGXghvcZ9979bGJTOR7767NG6S+DtG5+YbW8xa4ZybRlbxdGc
A7o1/4krEUc/YECilK+aDCcrbCx9EYWLcOdi89uMGrefPGPTUxg6J8m/z9Yc87b1VhrwVq/8Qcsb
08C3zbdvc35eOrIlmuLPK7FoNSxGzkZFoEWH8EsDwReuSFql2JWoSzuklUZ01g+ZBo45sXxuVuwb
Xv+z8IvD74CO8oScAhmyC674VfRSykSp7eQS0zMViT/cF4BHG1VLbqRkhRsIYFQZfA9BHs9lM+Sc
yX7yWVqtGoECH6cGcI5PPfp0LEuX1ZPOh9Z2xTb0z8qkYg2n74bn4bZhOZgOaUreA7wWI9ej/w2Q
BVK5EOIbLVvr6WE9w+92/8InGAXQsqCdJrMMAWbYEknMtNyqr10rkHUDEwcSXWKAZaumkTTZSEpz
LEpc0BREX5SFwRuGSCyhmhWWRFJexHORPfQHEMye16VPmKXNnykIFJs0keO0PWmLOU0ckOTsa0su
VZBamyoSwkE914dJbqebZvCLCeOyhmi79tdz9acKjp6DFS+4VK4hLm2XkXs2FePxvnk0R4N02jpM
NQaB/RbnJMxvW2vylD+zguHyyovuqDr+Lw+H/LbCc1/lwtuHHJ/b7rZ7U4mUx/7bmK3LkBQCJ/EW
qDruUQsJc0AUqHPIElp7WrML4LmzkuYAZx5jOjgtYLpiKsEzThGtmlPU4NClk6CHzq/KvGuEiq8t
9vmxfuTGJTPU1GZg5hVenP04sGn9/hA2wjKoQueUxODdEiQgjejf4fSKsLUF73CZs03Vc5OzigF4
1HH59uIoqRq1CW7Da7WQIBXzGgPwZX6QLid+CNVRyKY1Pcq56pwAUJTqDKr/SYB6hKtc/pVtZOF3
VS6behsK4RsnJNdGreUpbFsBeMK1WJqU5g8W0St50BM9MI+BvQ63ol4tSW8LD23ZJ96CsK1YLkwz
0YAM/cTNM6KZKU/uQKAB+VOr33f3vXIiimqRALruoaFuWoe74R9Xb7kB1QOdTTtSkd4oAd4PKrva
YgA/QN4cvKQAvMox9SN8ZjKDBJKkcv2p9thDZeNaWmzgVqoDlTuxJmHzd4nL4Z7te/utopQLGe3b
/5fKMs0L1oyazFj75WFro7225+ckVteUu+Pm8ld8tPT3v2I+BDxcd0+Kzv4wE3UFsdbj/vgBEB9c
OYKDndEpnjC9O8HD5MBb1wnuyEPa8X3rWy63qOvbOJRE2NinhEpUQKch5XCX4lAxTs/lgmyz+2lf
+neGKuiQB5dBrjOO2RtRhJF+X/TT3k4jIpIAOauWZ1XPLhHMdzEXk1czhALqXWSQmaGuJ8N/GHoF
jk69AKKDVfGSfW9q7sxgaUL4E71RYqD0K9Nn6rLZjoa69BwBTDggbb4yJ9oFzDbMF6bOE1qP2xit
/DhsXsn9Xezol6z66ie1w0mcLiY5iS+Omj/NsJiwDBg2uTkg4MhLEKXVmg7an4iBz25A7jobSqaI
I0zjuKvtU0WYBRngY2kaOwW9A7bLpia6qw==
`protect end_protected
