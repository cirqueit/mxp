`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
rRWrpd6hjYD3K3q6kM1NZ1ODiTCcuaWYTL+FSF5iUwTK3EUTvu2ycgpZAmAdkEyCFCMcu8Y5aMRN
IaAyjEIjp5yTnlVDr/qaEK2pn9HB4XoPc6x3+7NFpFP44dUrXj2HfDK5rx4HBxydBtHvmzCOcoYi
so2DxrqW1mFLstaMDyZ731CXJdDP2LnvOz9z7P7qihTzMq9oz8fJi1THNK8ch5pmIIVCRh7JB5mE
rYVjPdLwlnGqI+DRAduUdYKFee56sREVpVImJlCQi293eRdWq1/lcAnnimGWsynX9PmzL9vP9ANZ
IV+B7uPBQVYIxDh3CLz39mzVUO52nn/ZFUN18IZknnL//JQU7+j6yQkxKg+vkiR6cMUJoHkVkg75
mc2hMcryThoeK6yS3EUetFCWCGQDrhQiR+TD/X3lBCVZlgcwj/LfVLgnwDDJNaQztlYOiEZCPQMz
tv0grE66/2j4uroCUQGCNGXkNX9KguVIUCeEgelmhuTffwbVb1W8NRwQC9HjqRN14TZb4GJ0YLxN
E+RxW+ksPIUd8Gv8iORPtVwf0poqDUL537+CKdvkwgtj4ghaJLR30cOcwuZWi9rcrRrCwj4S/qQx
8g2nz+u0OEa8dG8iJagtlhpbqPAFYtzQaWst9U0mO0SHS/diIghzMgnzKbVLvPc2yFtxUWBhZ8zt
hxxIyiCKBTX0yn7dzIJ7JwTETqlC+uGiAZuUJlvdwHpWfBAgcCMOy/X+A4R9s06uWBm2Zh8hTh4M
UgXN8pfWBaDkxVytCB3jBStv3MY6osvTRskvYPvgy2lS/Zq185kPkUtDkybXW61tTCHau9jYqfL3
h2zCvQFq7S9llHnLYY2AbY604hZrktTKIPa1LoJkBE6cTQ5SDurAh9vn+QMflmRR0b2DnI6mdclr
dw8EJT3e39ua9tPMFsGMk1ke9+g/ocHWr5YeDujV1iPWUSuQHYIsTSVciTueTK78tjf2AbrfUEMw
beQWeUQoqeHLfLAIOMK8MB3R43+vRENSnLjYqs39zB9cXW3VnijoGr1eT9Y6WQeHixGSX17MaLMg
Q7PYZ/9+Risy0OJXc6Dt4dfecp7tOxD18XDIhLOLjuuftmxLU2CNpcWVaQezcP0hJHHl+i0cSZ64
JL5N9jJagoUQslydo5q9Pt9PxpfqmIyprQlNfuF/rIw+FSJIOaghntCaVGXX1gQ7T52lfs3bEB7x
ChMnyVjTNz8Lt82K5jJDi3BxZTnh0v9Wq+UWu4BJO8JeSSePkLwYWUqnJ4VIeS790UpFWJ2EuIrC
6xT75axbUuQQIU52QVi1pkmJMcqIargVxwwp8p9UG7eSl4V8YT5SYsIOeCuPYyLhMG1pun+iui35
+WiGNGZNhjHOKlzwhdDoUB1YYroNMI3CZ5y6WNnd0scQhB/R/xQfNMyIegtJdxlUcZPnh+bJN1Kn
rCNowkyjtq+mP1IjY5yDFuIAb5KWRO8CB3Rke/e5ntm5P84/cU3Z5VQTBa793e4W3h8GI5JWifyf
ZfAxWKtI/XD9B39QVmKanEi72oUXiPo0g/dPO8FcqpeRl6aY6GoNicErcnBCIUEC2uPK5080kYhc
v+Ph/VoXr7Cv9Bc4g/fFSbLJMAdETmQGdGQBq/D6hsgcaUm4Wn+AXeZRCJ/mxbEChdFVXyOGQURl
w39+iFkDg2KhdYU7OSV35mws949k1LEcQ00e3J0gC1Cy5wgadp1qkiI+NZeqCA3gQILV7Bct/CFv
iqhy321Aax7K8n0QS0pB4oM3MhjyWffsyTFU7JVGLIA/3+xC9xDgpMLETAtHAVyO/5OcxczkPdMj
fWAiP3gU20Awm+t5M5DEX7E9NkK/fMGRwYdQIT4H8LwW7eQaF6avlLlndrc09a9Ob3Ag3u31GNIw
fGSCpGxfHJhxqoLpiDIjduYqVd7WMdhtcsijO3bsULTg9rtevsgGi7z58HJI/HxM58vAA47wTIVY
9Vf4eiVF2ijxr1UAWxMyzPxFm6PpC+eaKboH4xaV9C+2aq2B2zizwbnv4bZOB3gXPlVe6OObDOhA
SqN6rQ3O0BPH/av0FZaZApGHwuACdJsxyVUJt2i+OMgtnd34bFvC2Jokzd4N
`protect end_protected
