XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ۊ���V��2�#�ց��_4�@������i &��i0�8�v���qe�ڛAI�������&�s����v꫗�5�MQ��C�X>��Z.����a3~�#�s�(�ڴbH�C���g��ȊT:nqOb^�c�U�+�a��p�@�Q��ՠo9m�=�(/�zp��6�u��~�ED��{@�.��Z-��a���mԻ� G/ĥ�;��G���Qw�A�Y�� �B/�A���N� :[F��O���&��,�����5��}���)���� �bq��#�#k}��s��#�ʡ�/9�̶��؇�<8��bb�_?Td�����+��x�K�Ĕx��^�Y����v�?��r��/&Ü�|f:�;u8�U\"��$_p���(�)�!��$q(��l]ܶ�W���/y��)������J��*��U�XcU@x��UmD[$���Y`1�P*
��Q_�FHXb+���kp\�:RO�I��V��e/2�J ���@�������lus6H?�Y���^�/~�1�1��ȡ�=Ӻ�E��rK� ��Lv�'մPr���o�8��?(�+��&FIwoi��6+�!���������ҡ]{� Y��v����*�J���׾���Ȥ���A�b$6G��|��I�~��=�ĵ�ưe�O�Hp��)�4�
���Oi�A\���u Peؘ=Q?�o5���_�������r��e; ���ĺFX~E�N��N�ґ��H��b6l�`#r9��/r�N�hDAXlxVHYEB     400     1e0�e�dj0q�[Â��F�ɮ%bu�o�3��&������Ciq�9��gD�ڿ����<�v�"�=����w#�ҀD-�${^7��X���`[�0%�\��ߍ���Z�t�A)d��V��}@����b�2��Cȸ�CС��{���J-�cQi�)�
m����Mj�͐J�&iC�-� 3�Ԕ�R� �ꣴ>�Ȑ,ʶo{�, �@ :�:�S�P4Ow�۫x+Xh�����)��b5/�w6uS�A����O�Ɏ"�|��>��@��e^�r�Vø]I�P[��ݱ�����X����C8��;���IQ�u�Z:P�@Q2}�*ܡ�m�ӯ�;��Q5C��
�d[�E�;Q�~aض��:�#��E{���S�&�~���$l�mQ������G�%Z)��l�~������7��F�hH��b�������D]�E�\�l�{�F�����n̐�/�XlxVHYEB     400     130�����߯D:>*�O���R��K��c2�3�:�۩��6��U~�G��l�D������ˆ㑼ˁ���(�X�Y���e�XeōC:����Sx��Sl�5�;�����cL�_l*��խ�/�y�idA�&�\��%x�h*��菩�b2�K�����.�oJ�� ��&C��J�Bk�%�)�.E'����9��⬷Oih��F��R�g�4o	�0uw������]���� \���q��+%�ޭ}o&(K:XU�}�G��M
���X`ʐ�-ͭQG���W��| ��5&�O��9ѩ�XlxVHYEB     400      e0&��{'}6�3ظ��w
#�nۮIe��M1˟^�8�		�*8@�RS���N"M]R�/"�j���{����ٽ8��x1�˔F�"-�����0��5w�3���{^?2B��#JZ�K��e��02��{��	3�&I���(���w�/��i���'Cb�z 
\jB>9������-�����ҝ���zj��i�]�-�P�}��f{�f��ݽ��DM�XlxVHYEB     400      e0�.K����`k�H���9��n�X���2&�F�ǉ����Υ벳�S4��i��o&^ӈx�X?H��:�X����zZe���s�4->h�=�cx�CmS@��<�zX�Jg�T~凝�kCq;���I�ocm��ȁ/�.�Q����7��n�oJ S��q����Nk�7��/���/��.L�� �79�?�i���v��eD����=W�@L�����>��pXlxVHYEB     400      e0XW�b@��Bj���jD���<xZ!UJ4ӣ2`ޣ�C�����k�4���^|k��?�N��OB����r�x��	�ՋiJ�l�MY
p���ϥo��2���7����P�9���j�o��{Ç�Ҡ:bF�1�^�iN
���7�Eo(�b�J.���}N��Am�=����(:Z�I���,D��\S�mp5I�1/I*J����?����n��5�XlxVHYEB     400      e0I]kIU�ٟ]!2BJv^�ǟIA5��H��{e����T-�
<$OP?_3P��_*5�w�L^�`*��Z�⼽�^��t`qt01O�A�B1��)
W�s��ޕ�0�QW����nA(�Xk�3��cLgF�)�f�cV:����������R����j"�6J�ܰ�����.'�[w�ʚpL�gdn*>�>��*���-��NƳc�Y��agL_�]]
���*�XlxVHYEB     400      e0�w��=��.��%����<K���X�N�ʒ���k$�?#q�� �h�n)Jje ]�Y�>4kf�Z�ԃ�TL}�_kط��,A������� p[�kIq�Z�y&:�VΩp��g(	r�Q?;���|)Jt]�K4��F���)i�)n���';�~&�ҞT�c�jjk��4�g�i[�Q�l*�3Ԣ�h��P�!�ϲ�_�3��ݧ��KY��iˢ��,�y�|��XlxVHYEB     400      e0���o���J���QG9�5��H[ض�L?'����g��k�WBi��?�_��?E����hK���"��R�)$�M�̓_.������!>��H���i��]���e�Ԅ-Ƭ������[�_X�Vb�`e�m$C�{戫��G��{{X%�w���F[JH�[*���4�'L���⯘0��f�A���]��nQ�x��%���q<���z��=���XlxVHYEB     400     1a0�m
4�%$��Q�o�/��5�������oXYKg�(d�u�M�X3��
�KW�}��!<|�͋��Ǟ�1\�}��8��&���a���YMY�,A�y.]����n�q��l\%2O��yi�gۯ��d�L���2cP}�����K}�]�鷟;V��-o��%��Kc��j��B����Rz��	 	���0�^���J�����T?��G{Yؤ_{��=6���ʮ�,��(N�?'�/�Z�_��MMW�/#	>c�'���V^��L�Mńr�F*��0�E�>8��r'f�����x�Vg�J�i��sTІð2@��rBK�Bej�����/���'�����tXҮ�Jm�>�A%lhI3�����8��;���G��R�;m�rJ����,�=m�.��A�
���XlxVHYEB     400     110KW�5�P�e&�BȲf:�t����/��y�����0E���������R"�=h�#��ʗ	�߫�c?46a�_'�4�!5&�@A����HQ��P���@F��M7P��g���ʤHI^�sC�!��W���dq��u4AK<?�g�&�P[�7��ٲ��i�����߷�_�6�Oz$kԌ�������e��xj���}>\�yY=\�ZA�4K�Jx��uݔy`GABfA*PS��8��6>GEW�zDgj�a�H�ߞ�C��Z}���XlxVHYEB     400     1809�R��+��%��%,�/�ǫ���D�y�TQh��|`Jh�J����(�[�H����uވ��/���N�g�(NE�!�f>�S��'�d��ܸp:F�<l��Hk[p`?�C�Ne��a�8֑V�g��V��)l��d^#6���W*o�شA���<�9���Bj�z(kz�Y�~O;}s��"����Pk$YB����q����+�W)�R�R����uԟ�ͯ�z�Jɀ]G]lQV�y{J
�m-��-9Գtf��b����]�t�`/19�{�;���#W�c�d�gH@�0�_�܀ϋ����������F��7l艵8m�)��,���$U����pӥ�+�=����_O�XM��z��� 9���W�XlxVHYEB     400     120�WvI70�{�eE�������$G!}Nu��aˮ29�0��3��XOb�8����Դ�Sl���W�y����p�Q^�x�D����%�k1��o
Rr��$5����6��=+�Y3�=ջ���P�����;�����<��V���ߖ
�M�k����5��W��$����8)h��� �qIʮ �H��=���r\?�at�r���E��h6�ˬ���:���������{�CP��8-���qzK�դ�W��@���k�m���Z-[��XlxVHYEB     400     130�5<|�PALIDQZ��90ᢧn\!�ǣ#��گ'L�'���� +�?�pO�\������q�᱅Q������������A�ݭq���hR@4��T���^켲��4�x2<ޮ���z��5{sp���4�ڱzӵ����[9�Ļ�t=Hj�0{B�+���Ti'���b�l�k�MY�S�w�z�A��������?Wv�'�9X��#<�@��d ����!��#��^f�� ���Dժ�{�����sf�?�1����͋l+�;�Sd$������Q92����J1���C�Y�:I�fXlxVHYEB     400     120p�A7KJ�1(>A#8(�u֗����^�O����Џ�$���	��~ ���FtB���.%xy� �t�@;ے��ǁd3f�=�i�� È�׺$���s��B�*+jpǲa��p�{<����=|��c:ascDQ27e�.o�����P�8 )�s:��/�c���h��w�]�>�iWJ"�G��3M ��<������[��:Wѩ��\�y�e}~��p}�&pYX�O�CS�(�o{!�b��/���*�ڝ�*F�?Ҟ ~�Ǘ�^l�pq��~�XlxVHYEB     400     140������
�i�=y���洫w �@"���X�K��5��w5ϣf�I�h��CXC0Xj]�����lG�JO���T�ބ�^����ՀNu\�5�s��������c�>�.ǟ �!]����;�[�� 5u��[�"�2��r�B!N�|̮������4�t�<{X�����1���b۞Bs�l�쬜�FNϧ�r�k�mvcjz���@��(��Jo8-��d�uN�;��iJH����VkX���+��V<�L��;�������7~i�>wW�ȭ���6Ѳ�a��~��7������_��<x'����L�#��'?�\��@��=^XlxVHYEB     400     1403՜��� bc��* U�Z6��ˌ���#�[�]�xS�ʋ+h�D��?���I�U8�[p��C��;T�8�a�0�8��t���qɉ���B�KI�<<� o%O_c�����q:b�qn*�B����K������;�d�a2,������p!
{k�z�!w~ ����Y�Zt~oy��&�ˏ��?qQpb��r$�������2o"��8�=�$��ݳ	�g3��Q�v3�,��"����w�fB����\�Lti_�ɨ�Т��1�QhE�����Q�F��$?++�G��}��{O8�㘣j�	�)����!@C�XlxVHYEB     400     120��i�Î,���_{��n�uTa:�P�y�4|c�K�٠�H+k2��}o����'^�0�OL� x�.��C�ɡ	����;)0�8��sM�I*:t�| u�3�l���ւ�8�`j�bU�Ք��xDC��Tu��嫵F$�>ƥ�|�EE�E+���k��A�j��2�, c	aO���(�SJ^�ya�<�8��B�m�o����i9�E�	1���J,.���n�#��v �F�g�\�3o�J��{�DG�7��g�;�4��׍�a񘼥�9C�s�/�ʌXlxVHYEB     400     140��i��Wp���`nG���'�K=:bI+Cd�rs���)]�>�BT�e��d��f�Md5���}��҈�u�%�3��]
�&��,�75�|��z���j��$�+�F����rf�m�6��6~&N�p)͆��\�����ed���S�f�;1+.��^ۑ�n}3��wK��#�h-o��<Y��%]{�)��Y�+������0�k��������.��=�w<_!�D���u�C��\3́s��=���p�yx��Ɏd�G����vfg?��*�˿|%��,E.��E�o ��U[Fn~������昡�j}�ћr@��_����sXlxVHYEB     400     120�����v���,�wB�~A2܃ݠ�>�#��y�H��$G�K���EV��]8c����iWaѯ9q"�k��5u-�8K ��*�׉��2 L��!7��D�ۄ��½�s<jz����B8�C������x�T;s	���4�,���w|��7=��Կ�������YY���*�\kh��Q��x���w�_u=��?3 ˣ��g��5�X瑟}��W�� b�V����T�6��*��qg%�%��N�HM}���J��#���Z��>���j��ŤoN��ŕ0�X�	.wBXlxVHYEB     400     1308�R�����_4�ˀk���!�ķn�=ԫ�����a�ԋ,2x���EP�ѣ��}e
HCN B�^��ɴb��(|�6���.�X�y�qx���kB��*��5>��n�k���N>���Þg���Z���8�P�	�KJ�OT�O0�R�>�����d��K�3|J��ꔌ�
�b��x��6+�< ��t��>S�ӳy�a=d�,��c����ײ:6`���4Q�S��Eץ�G�g�E$�h��#���S3ML��ܧҗ|!�ega*�n5�7D��aC��ĕ��H!i_@b*�~=X��ۢ��+�i�� w��XlxVHYEB     400     120�B3 F蝕�F(Ԯv7��,S]�tk���,Vy5*�s&ƭ<�@xEy��W!��b6�:�x�7�E���R��ۼ��r���`�U�)��'1ցt������Al���#��E&����+�IgTOrF�0�8��� �ә�͚��e�ʑ-um%��D�]z��ǉ�~xl���Y��|����<h6�l�P.�j�&j>�pc�X O?B�3�RP'��BZe�-5��rR�D	 ��X��&�_%��S�q�"�U����W$��>L����������8���0XlxVHYEB     400     140���H�\���X������P�l����|y��.WNɰ ̋���`��RW�����gv�Q���N���L���n�@�����[1S�x%�]
O��`��n�O\�	�b���f����N)G8]<缛�e��8�]u	@�J��`�Tۓ�#[s���y��k��%b���dŢF�	�7K	����R��c��Y�ꯅf~d����ԋ�gp�h]�h�,�c���ڙ$�F%�1}�D�KDL�S"�
����Z|Ȍu�2�}tș֊8ݜ�:4��v�h9̨E'����Dj�����=�TP���82��5H�:�^XlxVHYEB     400     1403՜��� bc��* %#Z-�=Fq�ټ�k6��|Զ�%�2��N�C��aRA	�D��l�>ah9]Q>�pQQ�ʎ8�~����nL�l�v�gřdL�=�A��8z������|[.�)��W�F���b��o.�ʹT��ڐ�z�/�5:d�8�J@��6g���(������+�7)�_�VԴ� ���#����s*f��𣤺����ѓ{�P��~��Y�\�,�x��X�la�E�#$��u_8Z����#o�d����ow���8 �1��_�"�U�!1���Qh5w٠2��M�H���Ϯ�_pXlxVHYEB     400     120>��|x� �H��]�Yɗ��{?�f�թ��+S�B-���ܺ���z�`��xu����Ű��x�"(7/�b<���������%�Ҟ<���X�^(O�C�fc�-Gh�S��^��5d�oMʊ��l�N.���<]��X�'H��j��n#�z���e�=t:�����"� ��[;,Y�$�IV_q��}�NN����Q[g��`_�1����i��:N�&�J��x�.�t]��@�1�~�U���̐�� na��|�N�NY�ٵ�O�,52ΚvY�j�(����XlxVHYEB     400     140�ͭ��J�< 15^��sN8!���WW#6�,v6N�`2�}17N{F����u�CGUcn_�3'�@�Y�ƉA^�=�C3/�:�X��2�RK�ҕ�N'�M�w��;�x���ݾ��
�I�9:܃��ru�m�Ky<b�,��T,K[�����4E����f� �)2�`�_�FUY�"���-yq�p�6��`�2l1b����6jp�����@�[p~hD��(�a �{���)$>e�G�G�)��Ĺ<V{��C+xL��@T��\�1HU��]�JS�[φC����`� *��5.R��z}3gWG)�l��U��GD�XlxVHYEB     400     120�����v���,�wB�~�I��x���!��u&�[ �f+l��[������E���t�h�W1+8��-��&�J9lϗy� 2s�od�vS����W�g�o@x"5�� �������J9�B�X�w<������&��>ni��0zg�)�����+q<�&b�0c�4I�'�n+�n�Z����ࣼ��-;Ć�K� �\N���Z�8��$��GW��'?P�Ʒ��b�M|z����Xs��������N��S	z]���!tؚD�����E��njsgh;��9�XlxVHYEB     400     130�ܔ����ʽ��n�0�x��jqw���B�gyV���Qt슍�.��m�Ec̓Ś)�K/]��+���b�B�������륒ԗlb@@;��.�<g��k]|&	�=�����1�6�=��ft�r�w~xJV�i�'�BJ��!Sǖ�1g�!taoL��c﷢�&cĲE��[��3C,��ps�;&%>d:�܄K�|����_[�h�H9&��IC��H5���y5��S����A���<��B冀>�tM� �q~��tۮ�DN���%Y�}�)�+�FnGĕ�b����U/r��XlxVHYEB     400     130�;u�y��)9�K|0�o9��Ū;�.�,�1���E\�>��XBl+��i$C̻Ra��%x�"�����6��1C��@g1l޹���`�����^q�V�.�TB�?6?MC�p 2z4����Nn9���#�`���e��������^�"�P�9�C�k�*�n+��^	��J��]�<[�W�r��\��ڧ��y�U�/_<|��C���[�B��w�dБٖ��G9e�&O�;:~���)1[���H���i4��[��96@P��8�qp�:c�{��S�q�@Q�S�]�0�l w���y�XlxVHYEB     400     140n�����*j���N��؃Ŝ=����G�9(�h�^�в��$��S�%0?�a����m�;OP���6I	��FLkY:Q��IWR։�����%��!j̘����w�n���I-���m&g�evU�C"��:Jg5���8��n�>�1��\$5v�z�]�x=G�s�NP��.͡�����BٿQ)��vt�z4�{?k����瓞���MY� c����M��|E�]l���Q!�H�]S,;K#w�VǄN�`��N�z B�8�I��{���q�Y��4�';�-+�$��XlxVHYEB     400     1503՜��� bc��* ����"�d�zt_�q�7 ���ќ�A;� ��AfL;I��#�z���c�S�(�1�˧����5��U��f"Ѿ�޹P����3x�Szk
>�|H�(,D�s��&i���Wj���H�+���n�K��h��+0�o��S�F¿�-z{�<=��l��N��4G�����l��?����#-���Ec��㨼�����S)��>��9�0����=pΠ7h�#i�I�� �N�{���x�jYj���<�VJ�E������r��<�g?�D2Ly��#34�ڠg�3���0�Û­�e)�Wyl�@��9����A�XlxVHYEB     400     120P,G1/�Y
3-G̳��d�C 5GO�!�o�����j�XG�d�5Z˄h��	����5x��7<+�����-V� �˨�k�$�l}��e�t�5Įh��I�����ƀ����xu�`,]�%w ��˳�g��2p�����Ei���8�[x��%��C��+8��ƣ
����P!o���L�5�w��/m�R���{�����	䖪ȷ��j���QQ����<�W,�G^�r]��Nr��+Z�hR,�Ǣ��u8���O��1�N��8jzP�2�U��7 �%Fk�yXlxVHYEB     400     140Iʺ�o+\'B�l�@.\P���q���.�8;��V��>�<���RU�K|�|�0��Z[3w:} �+�����W9�j#��ӟ�HiKH��+��[ܡG�X���VXgj#��i82�5o�BB��������yt�F�EcPz����ǫMp�Ȍ�{IN.���*3B��2�Qz-؉�-�X��+kzE�����b8�^Ŭ-�eC�<.{z3;��8fA�y��6��҈=#>�	���3���F(����pսS�!
1�"v��rn g^yS�0p��+�6���e/�gJP���h�9�c�z)m4,XlxVHYEB     400     120�I�Ǝ�ӛ��9n9+&��D�IT������`֑7�`�����P���G�$χ�b�I��wӉc�2掵�R˲�\M��??�.���q��ߓ,��tO����1�Dt�������F�)�P����f��VCQR6�@�[����	{CG��C���x��!g���L���$�*�,���q;��-T�ۻz	HK���V���QK��`�%mGW�o��[��I�N�t�\��� �L�26�4/�Q���3�C�+1��i7Q�_�a�jR!r��hT�\��Az-XlxVHYEB     400     1308�R�����_4�ˀk�ĥL5W@��MΗn!�<"	�ST~�kk	�h���������	��]K�����n�3�5����[�7r�yytO���3���z�9�Ss��TC�~�ױ�{�B�
�$d�݆��&[��-�w�#Y3��W�� K[H�����;{�	�8d�PG���}(4̛��)0s�aQ_᫔�bs[=�C����R��ε��#��Q�H����vYO�x�j�0L���A=^��b�~����n��ׁ7Y�P���a�"X#(����_��y6�5:K��A����0��XlxVHYEB     400     130�;u�y��)9�K|0�6���&��U=+���0;�߯B�K.�uAI~1���R^��ڄ������ғg-�F�$�	?�ĕz=��I�Z�41���q��f\�]��	oi~#�KA���?��C�ᔺ5#������|�#k`Gq�m�nəF���oj��//z��q�
m͉���������5�C�U���b*~ �!��0�mT�A/t�
-sS����\΅���:	�<:�߼�?��A��vyIN��h}��-�n!��{1�B/{�zza�v�,iW;���ӌ�XlxVHYEB     400     140ëX6�^�>^�8���:`ޭ�/t��+m��	�6��/::t������$0�"�)tiHX�y�9@f���4f9susD��E��W=/�7�q��t~�R�8�w�&�����E{�#Ծ���c�+�(�X`���O`X&���k�#Z���Re/YZ1B_z��*��H?EM��:�&>IaL��f�4B l�O7K�p���F��T�G�ċ"�����S�}��Yր�c�i�yrG~m��X�n&���u�zT.zQE�+�������"�Y��kt#���re}��Lf������΢5�� y�`�OuC�)�$�=XlxVHYEB     400     1503՜��� bc��* �~�{��X@��Yi���m��K��
�Ɂc��~�c��N�1���5S_6�ys�	�L ���W��j@���³	�@���8}t��À���o��l+���-�~+=0�P�n;���>�P�: ��0 ����G.}�ܥ2�[��#���o���9Rn�88=㢩�=�8�U�:�bY�0Nʨ��9��*�Ϙ�g�ks5Q���d��!� �3D�CL˲�/�;?l�6C����&aU�s�~��&�{.&�,��
S��f�5�+u�/T~�� /����9���+�� Y:^2�ܿ/��#d���d9"̉ӵN��|Y��XlxVHYEB     400     110�Rax�h/�4VZ�D��Cî�9S}o�e�k��x��r��!<��g�M��p]A�U���|m�$o`�
0��sO�֬5q��t,5\�7		���։|��q�۸������_�O�Ffs��2L�F��
ߘ��S��mm���24�T�����_L=�އa��U1��wUz���'B���N���ӽJc�)�Z�d�*L��9l��߁(�}S����+�L�L���?��]`�A��J`�T�ځ�s��r��FkHe��t�
��;��s�_XlxVHYEB     400     140[)�8"Ip�B���C���&*?�C��2��� �A�G9�I��80�	 �!�2���n�~��:�����K��I?�	����Z	B�����5�C˗HsR��3l�� f��+t8dOa�+��Bsϰ��˝4�[~�~�h���t����;��c�5�XgB���`��䳦�4��p�$%��׼oׄȰ���GzB�Y�f��/��x�	P��M��4��e��3�|,�
�+UL������ �հhbDQ���"�zq��v�m�)�G:���(F1��6���̟�?z�����q��[�=�XlxVHYEB     400     120�����v���,�wB�~���C4	a�W"��/��JU���'}1��-��/6y�V�ahO	Uz�&"�>Z9x�V�`;8&��z�������OT�\��:������t�%I~��9�{y1|���>�
��K��9����aX�+#on����,���H�o���Sa��L4�B�0�>��5i)j *���y�,�W諒P��C�=�y"jq+�wH�+SH���/Dq��\ܯR䇠=�T�M|���Y�V:$�ӷ@HEi���/�G�IӇ�Y\L�&Q$XlxVHYEB     400     130VO	Sr�HN�����Q�d,7�8,N�EF���j�� �6�GX�����\x�WX�i6����Y[�R��v2�Ơ�x���~�ifm��x�3K�6En���l6��u��k�#�1��
,��*�<+�a�wm�����$_d|���P��'C�Akh#�H���w�;k��٩��^S�Y��A윎6%�J[�C߾ZVy��5/�JH��4�Dl�[A��
A��G��e^d��?C\Ƃ�q}�_3�S%������ʓNU�F��`��Z�P��_�Xk�\�(��71I%gS=���XlxVHYEB     400     130)d�<��S�|���>�*Gk��.x*<��u'���4��l	�P�1޿���l/��7�>mѨ!�a�h2��5�\�Ú�[f ɨEs@�75���cԺ�{M��@�������i����i��K�hXS#8�^�:f�!��
%��$c5�̫"���kJUά��B2�Di�y,�n��u;j����}�H>�<#f���f�r��4�*�-��,Miχ�jgI�4F�w��&'������6���ǩ�����fLȢ��`�>9��zĨ9�F
:���摊��oI-z�=	,"$�$��D]j^�=XlxVHYEB     400     140ɏ�� >�;))����đ[��w6�5w��#J{���J�	@M�ٜ�,��y���9B�M�"��GD�?_=�B������u���~�Iey�
,e�����4�Y� T��I�t�j�"I�E���}Z㻉8
��u�"��F�����x8�m'��nn7in�6�(����U�ߜ����P>�2J4�~�� /�H�Y�����:Q+��o�p\��O���e�7/���$��i��m�#�'X�h�R��)����+��78;��M��#�����w�b�Q~���Z�;�<��%�R�p�mA�e����W����U"��XlxVHYEB     400     160kYH��������U�#K�@՟�����f�ܞ�=r@��p��\�n2v�Դu��k��ު�iOͫ��%>��)t=6����N'�-
�<%��`aQ�MT �U��l;�58[�L�63HG���t��B�ֽ�_�A^�n�ώ�����&� �Ap���[��~�%�"�wZ`�2�ɣ�z��+D����8��QH2�3�ȿ��>i�Z:�����zJ%b�6ސ���y��}��i�ɤ	��/&�o���"+�i��Y>akZټ�;�f�}����u0Ф�8���Hg��ꗠ�۬*���&�OF�D�H]�u�[�hF�#�&)�M�1tѕ���Tl�~���k[XlxVHYEB     400     100).P�\�x�^�ʣ�<(_��Z!����@C�����O�2N�;n��E�4�&�7f5W�ޟ�D#Y(ӛ�v�5U��D�%��8X� ��N�<���0]|W���@�i<_(p�[ ���Y���y�9U��%�pC=��TJ'|{��.r"E�,����t� �<C�����=� �B-G����U��P��Y�_
�33u�� ����%1/�7�@آ��ä �t�ӝ�A`��聥4v���U�R�?K".%��}ݢcc��~XlxVHYEB     400     150G�mf�v�Z|��A)���<xI�����q�W��=�XKu`�g�5�-GP�m�<�iU��V%������UG�K�l7@b����N��Ɉ��0|�i��*�V#kG:��]�źF#���\2���l����_�u7�t�щj�~���}��@#��� Y�s-!9��>O�V�w%�w�//�{�����-��
�S�d�+�/.��jn}�K-�[��38҅��Õ򜩀b:X}����7�{_Luu�vSu�+`�N���ho+D��"HCT����٪(�z@�@�ޡ+v����F��]ȷ4vз�z3�B/ٍ�R��EØ�N���=$�XlxVHYEB     400     120rJ�}0��ì����%�x�D�֐���:�𪒟&�����A��ܔ��f�&�~�:D/E���6B����<���Q�v��kCQLr���ݮ>8[�������w�
9� Z��;=�:=�v[dbb5��v�\p%���+}s�C(�뻊Ǡ���A����hp��;�}w��+��A54�,!��Ոj�;���'��'���
^j-��3��E_�*�Y�9�Jԥ�iP�q�r�X�$�k�E
[�����
t�,.'`��B�Ѓ}�Y8�&@�S�I,;$bQXlxVHYEB     400     130ٕR��<ű�_T�F�o ?��ӵE{�b/�ʴ�^���kF�4B�Dʲ(�5��m���\e��h>�0� j��:���We��Ed6�^���cQuQNq�,�����G��^�ߙ�͜t���U��,:O���=�7��s��E�F!�T�O��U��OѠN�;�e�.>Mn�:�I�p�g/�S;&����Cr4mi���R���Y*?ڞD��ɳ�+<p��۫(�~]�&� u�2%�΋�����%��cTI���5kκ���	���`��Q� T@aNm�-VyG!�$XlxVHYEB     400     120�����.zR&�.vf{�7�	�1��T�23�@z�#}(���T��p�,6'�0Ht#6����=�Vt��Ȉ�΀�i�\�k�P-.{��8�
�' ���G�n�� �tc3Ǥ�� � ����#��������}��c�w�H���w�G$)����~��$��yUNlBgG�i��0����!jl�|zkԳP��9
��W��l)��E�we?�#㚘�'����{�:V�{M��N�":��w��{j�A��<=`����6C)<Y����GNI�R�'ЙXlxVHYEB     400     140�`��#w\9�����:�W�� H�[^.;���y�z.G��{���U��VŌ+��;޵A�ˁ��A�S������~�u����[��):1Jz�+�M̇������?��Ce����Q�R��/�_^Ԝ,��ifq嶑�1�c�S@�����3��/�e����#���L�o�X��eQ@ ��+����9E�Ԃ�(MRik�`�"�n0(}����|�1��Ւyk�Hv�f����\oT�����h���:�޶ �4F& џ׫-+M������?r�!�RN�=��g$;yd��rq�r��θ�
�2\l��j�XlxVHYEB     400     140�0�'4~x��6,�dxR����l��g�����G��}�k()Ԉ�k����`�z�6ڡ`M�3��Ş�V�,єN��Y����u����U�0�w�`��I�K�����ݑ�{��j��O$>�H�G1��C���Tκe��f��]Ȏ�o'Z)�G�&w=-=kFچ��|�v��Y�w��3d�z��)@օ�2�P��u:9~��>'u�:2$���!K_��e��)șS|��V�l��_�R���՟8l� �J?���Fj�T�Iq���Ɯ* ��~Ų�����s�7��#~�e�pBve�Xb���+�C��R-XlxVHYEB     400     120���`���W�Rݦf��#$o�~$٘/dr�[�Y�d���s�e��8�
�~H��9f@�h��@���qb�8�̌���K{�w���3mӸ�!��]��t' >��;ɱ~"�)��E.r�7� .t��L�.��ﴐ��T�#AJ�o@d k��xFf<�����J��)�&5�E"d�Q�Q�Io�~����tz�p����	<֧7�\8��G�֙�F�	��H�V�#��$�!o�[�(7�dB��i�^�_S0�$�r��!a��.9�,r���Ք8����~�z�=�$}��XlxVHYEB     400     140�V��o Mhh ���ߧ�v��|?�x�D��������ׯ��
��< ��S��L�J��,����#6)w���P ��e��*q����#�o���0=.���M&֍+�QW:��"�*B[
 ��Rm�zl����ȈN����\��0UaM	��Tt�{qܸ�Ws��MR\�h ���|kE��v��)X�G���CA��o��d��:'D\x��/�Θ���,Cv>,.1)>�1�ژ|���,C��@�uṈu"�����Ӌ����SUi�m��V]��8J�s}�����*�n�~s���oo���XlxVHYEB     400     130��Q?R
6���M�$WZ��A���'f�����9���hBQm�	�!I��4M(k5���F���z���m_q���4�6"���-XyQG[�S��z`��h?���i������n+D"���t�R����ꖚ��K�9�� _[(�ftMWv���
ރ��"<�3 ��K�-�1|�����W?�@��ƇU��wuL��G�G\���܆�g�]��P�sO�]��l�i�\.J�7��OT� �K����*�r���hDn��k`��&�mt�tC���4X?b�z����3Z��XlxVHYEB     400     160�~�.=B]��P�x�ft>�ośz�9�ב�:IA(z1aj��5V���W���k�W��Ry���q��gf0�� ���h3*o�HJ�D74�Pz���Y]�t#��ؼ�HT�i�X��X0�)�M掬+�w�����C��cm.T��W<Ou���B�	�ώ �e'$e�OlN�:$�<��=��.D�s2m��,��຋𡥐��	�_w�W2��c��d��xޑ)է2��mj�A�y�4��0-ܢ�W���㳎��"����'r��?ܧ7���8uv^�fI�T��_�Ɏٍ'Z����R6�ʪ@Ě���!H��n��˗���*8\��n�XlxVHYEB     400      e05C����ƄG$�"��G�ط�[K�V�Ni���ޛ��f'����
|��C��v��e1����iP�D@!We��O?0E�q�%��i%��"�'~3��_F��?�ֈ�:��C%�yk��F�h��(���dy3��'O4�[�AR�!�����'|�Ȯ�a��4��RPl���J�+����Kw'���W�iHI{\=쫐�-�y�M#��+I����G��XlxVHYEB     400     150�.״;�z�3<#�e�.>h���s��\���<$ �=2�Q�J<�ر�@d�V��/�`�A����9��P��?K@C F�@�,Q���)� f��,�@��V�~1��a�t�{ˋ�L�]�j�u�ҵ)��gY����"Ϯ�	<�i�([��Q���M�Y��I��v�;dNQ�
��R&�8���O��A���>-�@N��k��RM;0��.�۶?ƕq� ����~���7�>��lox�Z�X�/�ϭ�$\�\Cb���$ϑ����e�=�AEo�����;d���'_��?�m�<��`�H#�S!���QXlxVHYEB     400     160'��0d�He~Z�ozfe��ώ��!��0�m��p���y�l���x��/����"B��g@!q,��z����!<�����W�;�!MґKlި�ݷ�4Z �r��`����IEʇzwʳa=�40���hsŹ%�#+�up�4��ڴ�9���ʹˊ�v�H"=�UT�@8��B	��� K��v�9�@'Y�����䳣P����mӸK�^���[_�����t>|ߑ�kC���R\��^0��]X��}V��2�/�������G#��v�E��!!�?^�x�%�*8�/SNu.a�m�D/���$�m�f�+���|�a;.����D���ow�ڷXlxVHYEB     400     120���`���W�Rݦf��6�X�NT[΃��̲.�?��W�N�ä����S5_���h5����i�XK��׌Y��j-�j/��|dZ�D���<"$y�$a����6[���`=�U1����Q�yQ� y�g�����:�Ή5����&�C���E�Y���3�c�\=�x�P&;=3���}c�2���i�5�k�8b������%���sŦ�(���^���G������X��d��x�=Ą\��KT�&D0���hfR�n��6sXlxVHYEB     400     130�`	��i�(j??I�pF\׊�+ w�z:~j�|�ޢ���R��He�����B�ɥ����[ϓ�SP�+U�jV\9��G���AX�^`�;KUa5�q2�q���xQ^�p��2]]��r�|잫H��Sy�b�<�S�$��U E�x.�.O*�2{�(/��P��{ժu��P�� p��r�f��N���@�� ��Ƚ:*�P�Dܡ����/��6{ؠT�<�&9�"���O}Q�X�Q���ኵp1�yU�:��wqx�>P�+�̵�Tg�N���c�5�O Z�i']XlxVHYEB     400     140��(Ҡ����eh��?YI1���Ta�[B�zzh�����	���T�:�R��%�Ȅ�f��t�S��o���+X*tK��u&둶8���*,�4���d�����*8�"����8����K�|kO�Hpk�ȑ�C��ZZ ��>����|͠���_���	_�0aOʜ��L�
=]������)���|��� >_��1K�����d�(���I����'i�`uB�q��n�5��E�>U���Q�5}[�#"ON�;}��y�o�pm�6��F�M�D�V�$jCq���,�-�见�1Ꮧ=XlxVHYEB     400     160	y�*�3m���y��8"�;u�^K{��i�t�R�n�s�S����m��^��v��6ݱ�g	p��	�p�'ZO�Q���˶3�F��SzGxV���#���-�i�s�X���b���m
��jE>����LM��a���%�6B.ڀc��t���O)���3Ӆ��:�7�Q��$�U+.'S|�f��>�5��M���1�w���c���kH7b���5}�M�y���V=���-�k�9���-�O&��)�ȡ��bh\�)ա�L)׆��� ����O�Ϙ9�����S?[JF���&���k�Q6u� ͙��T�,9k��se��V��_b��Ac~<d��XlxVHYEB     400      e0rMhR�vX��l�ǁ�<^yφ
���l�@yL����Ʉ���'�V�~��0Day�O*化��1޿�������j>/&F��D�mR���ۙ�m�FYsG�f;����:���+����UXq�V���;��o6�|;��^>��S�v�?ӈת!~$}Y[tԓ��� �n����>8�		�ߨ|��9nU��?�ED�{[漯�mĂ��B}�3%[�OXlxVHYEB     400     170�����>֟�i�XM9�~k��Z c�^��,3����'_4��7a1�lW��~�,�O����3�x�2C����g�EVb��M�u|���kDE�����zxv�r��i���u��u�n����π�-"�c��3`���bGW����!���z��r��^7!@�I)�v n	���̋e���[�Wץ2�y�gN�EW��H���e�z�~�闘��M��/����H�:7������jQ��j��y��˾?��?9wnTMv�|n6��Ì�n�Zx�pNfb/P�.6���5���ނ��H�2uX�lVv�:\ ��z�?������bbc�B=�9��-�C�$����XlxVHYEB     400     150`��]e �iH'ۺ��Lǵ�u!;���þBX`�٦��X-3���B�.�@�}1Ȍ�To��`o	w�>:+�Lx�kֱ��6A_��6?#��}Z���7�U��E�/[7l*k�~���F΋�i����ǲE:x���c�f�.������,�7�P�kM������kb+=ge�=����l�Ǎ ��STMu�>A���mx8��nD�_��6t����p,,�8��`
�9PШ1{`��}���<3$�گۏ`]�T��N�M��K0=#�v�A ��帓��>�����$�+Nntk�4uy|��|,V�y�XlxVHYEB     400     130�wc'�0 ;O�d�{;M=��vw�@�Br�),Q�!Pnʫ�k�~[���BLnmfT*����I2��׭�Ӳ�b5���10�|t�]k&W0�Hxp�R֢R�ϺF0[�����p��#M.���9���23��9'��ɠ��|R��b��5�6�֮�z���T��Hz�M�M���$�_��R�Ed�<�:;�r8C/�Vvg[�g�)\�����TZ�ן��#�Ofo@)�Q>p���H%�M�-iJm�r��{7�3�4�ѭ\�����VC��]W@��bUGV�P���v�zXlxVHYEB     400     130�����j���	O�1ŚG�d����Z^ȡ�-�)��X�x9�W��� )�kk}4F�x���H��y~s�`���6�R�3(	T�%l!�aaV���y�Bd��	�3�
�����i���a�?��>�I�g�4+5(��?�O���Qױ�\�*	���ڤ/pwoO�t}��l^����9��#�1Q �O�,�}���N��9#J�����[	s�j���B��#n��F�"���y��8r5�ؿ�J���O gr� g�'Ȥ(�V� �b ؛n�
������^�ǋ�$�َf*
��uXlxVHYEB     1b3      e0�~�r�"�xN1�)Ȋ�P��
B����5���5ȼoup�PC������9+;��l�ط�}	^P,��YOk[�o6֬l�
�O����q� �`w�c-� 4g�P��
�;��RQ�),�Ț�Y[I��7�{�[Ca�i�H��s���%Mʿ��O��DŽ���ru�tp0&p�
�t?��@�o�~j�+��Bi��\�s�W�N������<'�#�0�a$��p�`�