��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���o�*��]�1qe&���K�f`h�~|�X�Rf�hj]o�̦@qG�f�eg�2���Q|~h��@�ɘ��*1ϊ�\[6�q�$�N,i�&�Ez1uX*��~��yGH�]�JW	�S�V��e6�<�v3��ߚm�2-��&���D��맓6��q�w>��Qtdl,u;���ڥV��`2�~����j�A��7�y�/^_{}�7�ܣ�Z���~Bp�/��R�tm�F�6g�Q9���W+!�R�Ak@@ ��CK�0k E�؍�Z�un��I�cr�89�_���ulR��^����g�V��iڨM�a�T7
.�'�n,ǽ_�ѕ9A,ə:7+�H�F�L}�؇�����|�k�R���U~��Z�I��)8P�#��I��c�+�]q�6V�2�ħc�S똨�d��D?�)���/�gC6wX�񸵚�mE�͗_#D�`Q���l�NQ��K��ג�*.�ڎg"�#V�(ܴg�M�����QI�t��{I�͒�Jk�O�x��4������6��������ON��^$��,٪� ����6�|ϻ��*�~N�N�d<!�i,D+�Uf�!E��\�ƛ���b��N��y��h�A��u���Q��b9�Ū��k�0��<&���������#g+="A�Y����r1�rU�,�C�1�^���y
]�uTG_�23r���������FK��X��M:�����L���Dí��AR��>o�s��1'J�m��8c2k��"ӷ\�t7�c�4��e�o[��j6J�6#�5�����:�\����������'M�����|�I��ҭ=�H�G-�'�W�I��ވ�|�������H�nF�G$��z���@�Po;��ƥa KŒ���UGiJU\^��tuQfȜt���!r�;`82Ҟ�>�0������d\澢`��I�,�8Y)�x�U�_0X�n5����"ܬl��1�� ��ݽ>HM�m73eI��Wo� ����*"�ӗ���j����Q3��C�����Q����5�����.��Y�kj� A2o,; ��;s��OT�(����Je��/J�r?�����/q�"	�j/#��m��\�)?�\�m�f�,�Q� H�؁�k�v�0n����~��?T�[W���Yl�>L�-��{�K(y�=o[9��׉J4[$"���s�J�� c�.P7�D�j�7�� ����<�솙�V����W�y�Ւ8��٠��yz�h�dw3&�8���� �]�\͂0���=� 1�[ĜMg������z ����4^U�B��c-�YrqE$A���Û&��-y�U��dV��mi�ZQ���p�? ��,A�2@PN͌�,��#�F���t$��' $�m�.%�[�;�>do�Ȍx������&0®�P=knw�?�e��n��]tI͖Ƞ��@��d�e�y�I�PG�82�#E�~KW.x���+����x?����m_h�o�
C�� �����YC#��DA�  �V.5�Q�C>���39!�kд��~��D~�&}?�:T�z0c��o�`��Cx��؅�J���6,�"��%x�I� ��:�ſ�TC)sP�������w6xw�lI~��*�׮p�����D�^Gm�����`Q�
:��q��F��n��4�Ȕ�Ķ���z��m�o�tcF��߃v��n������;�4�	#_{s�Rؖdu̒F��X���[��j�T�}4x=惉�6o�b�jq5��+���Cj�z���	@�y��� ې�)u�П����b)��ք�!p��V}��=w}�Z��0x������.ȃi��I�������X[���4�]�X {�F�,��B��҂�i	����}�)v����#MWd�:�K�Z�[M:�K���4��IV������&�i��z3�͉���b!��<,Z|
���/
�!4_(��oF�Y"v���v�$Tj��ft�����[���6"˽Ϊ�/h|b��Gc�Q����e��Y���U2�c#<�� ,d��s�5�J���@�q8�,�z����1.��=5+7<#��ͦ&2:�; ���՟��$��蚪 4�����;���'��� ���"�S��J,�#�I4Uv����&>��_l�[�isMM�d�������Y�g6���8�� �g�Ywp�㖎�|0t�7~Y&����к�K��^ͻ���C�i��@�}^`G�G[�f��"x	v����l�폒b�xI+�#ɚ�}x�R,T�7�lU_v��\/��B|W�>�sn+^d��>t��)�^������bY�J-�4
!"�����i���w���$T_�	����|��L���'_���J>��C�gkW6r��n�&�m�P���]"�B��LU�J ��p�#�d���S���J�ۓ:MCM��?D��R��x�g��XП9�������Q� rC���jh��S��S�@w5�B ��)������ˊ
�bUAv/'b�B-B&��i��:�C�tY�Ο57��Z�����2~��ޭ�wҾ�勛�|�x�ہE	��;���&��ӑ;[EFyi�[Zs�ɬnSl��ђ{ԛr�!]�XqH3��X�K�$��`{�C�l��7Z��������jw�N�+ߘ:�+*��vZ���A��q�Sa��Bń�� f�޼���üd t!�G�V�=��x� -�OJ6m�?�G%��'|��Y�a�X�@��!�tf�k[;J?��C�±K���e�W��^��:=pz��L�`\�H����	"�7�'_.{�+�#�T�̐/
�G4�F���X����IZ�Uȱ�"	̱���Z��"�xy�r�L���	����~�3�Za�U!���3*gߒ!� 곛
rp~��/����A�G?�0~'��!��Z^��������|�a�=J���j�(��8r� ��Y��d�d��$)ٻ�[߬��4��p���58�Utꀤ�\h�ם��i<�e6E�K��X��p��P�����xZ$�K��m�w)�}�=�1� da�����C�m�d�t�re�1Л�H7`���2�9�A�Gg�q�p.��(`)���)��Z�C���*f]�"V�>ە�V��O���+�]ڰ'��������_<��t�"�w�Y��V"��cg����b�(6J��nQ�g�������f�Øs�8x���]A���L:�upޚzSX��pe��%�8(����ԉ}CF"��Z7�:Lu��O�B0��>o=������Y�����C1��}��w��p��'P�*Fy�}� .
�Ϫ>&��9�-2�����D�!�m����>���(��S�.U�M�єLd�M�������Z�t���Qn~9�n�3,�\CQ8�h��
�P[s:�J�|�' �t��!_�eoաwD_�������>�0Cs�^����Oa��0�r/��<��6�IG��⎪ n�\;J�i�aB����|�fX���_c]-��!JO�}6|,�H�:�#U-���L�I�"������q�N��Q@pR+����%���&zM�z����NԼ	�`����:��ec�x
g1v����hkU$��kF�n�;���g�-����\}eZ�I�9�i�`b>w~�~2�.Z���h3���Ur�_���6m�qW��)�VY�_?i�RwZ�u��	!b�eq�,��͡�']ٙ�u���z:�W�mê�g���0qC>3͇O��[e��P]~����⠓c�m͙�>�~2)�)�^o��������[�ʆ�QdL�J��H�jw@4���N�_�@`�	����D�6� �F>� �4���tx����N�x�����4K+��3�U�.�?>lI0�1΅'`�%������L�K.q��W�a0^�6�2���m���Z�K����'>I�gW�O#ڍ��y�oh�Dm�K����/%7��� ��ԘF ��/�X����T�3�@��0�tcW
�VrC&��pE��LJ�]�K"zS����V��^��������xg_���,
�t�W�ڮ)fNE�#����f�+S�@@R�[38��sSz`"�"kԎ�D�2g
�ʢ����r�v4q|6�Ab��Y[�{��ֱ�� d��
p޻�#�N{�졙6eg@�D=� �h]�!�hq�]\YJnJ�Il�n����,��S��x$y*ДԶj�҃b���Zg�b��S{�%���s.�I�6��������� ��d��,(;$��}�M�,�#hx��6���s����QF���2S��5����);V�0�LŮ9W���>1�n���n��l��S�Dn�$�| � 0�K��`�����n�V�D��a�/k�V2bٝ��Gj�>��E|����o�,�;hib��f�0�k�����w|�c1$x��_����f�΁]Ɇ���?�\̓�*�U���/Q*W��AN��*P��,�q2�Γ��$T��,@�����ճ	���K~�,(ԏ��(��OA�*����-w����w���������n���,���#�O��B��I�:��-�ʇl�X3s^��OZ����%;��egËU�V�"(2pwU�hR�6aM�f�x�ϡ�5�c��	3YC-�ΐ?�>�9Ϧ����=�j4c^���U�_>H�硛kS�M�}QH��������FE��&�v6�F4�j�1�r�}Y(1�Ց�q �8��a�ޛ�^��V쩩�U��8g��X����T��"��j|����0���L��#̒;�P%�L�Տ�g��t`��]YA������na4�Ի�=���|��ŧy�FY���I�:hk����q��^&�*����`H_a�O���N:�Ў�Tk�R1.���e�&�xIj���l���by�K0�"�=�N�!�_G��kѱ^Cr �C���bg�N�Y��d�fW���Ti�	:Y}-i;��Tm!�~��
Sf�
��;��&�Ghh�Z�m�IX�핰h_C�0�Ny����&N��6-��ʖ�_;/���;�LP�b'�Q��	Z��ޜ�rcr�9S�T�i�r�j�)�����N���b]�3Ȫ�Ia�{�@cD|$�����q�T0��
�$���R�@�r{Ak���OǑD������!�U�N+��-�]
������=����&��3tnK���]�S, e(�} �Qz�D"w��a�e8�-��ʙ���#ۨ<��9�z;�hz�a ��Gb����SX�Z������iŢ���'�Y�)e��ȉ�Os��~��P͂O��ވĉ0��ۋ�\.ns�����L6�ɑ�2s�L6?^�nr��ù�]B)�6�|�x ��_'Lh��E`�No�t���Z��c�{V�pX��Ur�2$��h2ǒ>���w4>�s�Ab"�TFTI+��T��'��4P�D:��Ђ>�b1�굴͛�s;���>Ҵ�p�"FJ�?o��*c��1�ǜq���sy�{L�#��f_�$��>��Ew�F�H&NZ)�o����8:��I�5e���r��A߃�6),�΂|!	����vj>�V|)�Ij�m�){W�c�o"dB"�!o��֤@�ޗ����'~?>IV#`�[ |�����eC���4�K��g�������Gǝ��g�m� {^Q�a��)�e	�����M�F����R��4�u q�;t�E�W�s�pc/`$�N�VW:&Q�ۊ1�p;�n����pښX�~�����@��v	m��jr����t�_�~3EL���[-�U��1=[����8W�D��oǸ/���b�6�U�=k����zD~\:��B�Z�h��a,yc��h�q�XG4��ai`Z�ol�J����4��4K-�B~F-~��M�	:��b{ߥ˺�F
!�%EF!���]�i��Y*� 	t0)�R�x��:���խ����4T�S�͕�J؉/Ne!�y_��0���R�Z۞c���дfN���'�é��Y���*�l]i�wI�Eǣ8U
7�j�D"��g�N���0fsʍ�ԉ���AI�!�'��z���r­׽ǔӍ��=��Q�ל�O ����>�Ϸ��ܚ^����a��j�I��ke�3��vM��Y_ܟ��\a�����q^�0e��N�hI����/��̵����ɛ�Y�K(��SՒ�AY�LF��F��̔���aY����]ʀb�x���Hp͕��
��W՞��!���`�/(�ـ��t�x�>7>�����_�	�H6p�'9�4��Ȅ� OQ���I��Ri�r����QE�����jʧλ����r�M*x�Xk2�[�<¼fr]r=�^�:i<�{��gW��H)(؁�č6�0�g�ϯg�6bB�4���g�r�p*/	2`����b�~� Z���ve��6�?,�
G�m���qPjhh���$5����}���TY^ߥ�DI�g ��M�)��Jj���C�n�a����O�"����������C�^=91T���L�g���L����Zy�e���bS��&���7�DD������l�{��"�C�Ҡp2aQt�N�� 6戹k!�y�!�:��~ɀc��\��������E�-�R�I