XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��M�w�s��S��*h��)�V����f��D��h%>Y$6�YW��u�c�k���ӾD��	\GT�TU	b�A�����b�6%���-��`�K^�o*�E£���*v����o^���U}�$'�Y/^���f�n�����	}���Z�A�9�5�<�0d���	!�Q.�78/8���쓹�,
�bK�>�|���$�7�2�q����#�����R�b��N�/����R4J_�r�{��Zӕ�ԃ���ݴv�w�s�*>��oG3���G��!�%����i#>�aM��c49��>0��\�u�v�O�V�q4Go��
Z����{���{�����bF>��:�%qᙖ�b��"�����e�bt+<+3j���@���J�L�(��*�'f����M,q��o&+w��Ր�2vFo	���F� {�z�K�tq�^�7�U<�^VL3��ܙ���t93N��|@8ƱO��iБ�����wo�]:yB���U�|��>�V���។W��>��d�E��B>�ҷ����ajC��t���4N����.s ��ux�/2%;Q�"�JB~�s��w�n~��Ƀ���w J%�����Q��Z�{��]���H��wj�����g�E2�Cl�l�։�d�J�u��0�`�3��
���yr��^�볜Y��!`����NR���p���❁�1'��������f��Z��7����'�%MQ�]a-3#����j�9s���N����`���H�B��XlxVHYEB     400     1d0}����˽(�%���xK�+�Z��X u yu%�k�����ȐGJ���ήLD�|n딀s���=������[��f���Lk��ת^'�V�0|���"_�h$mV�CQ�y;���B���_bR����4#�u7�aH-�#�1��aa��ܭ�F#^�?�߀�T��/i�BO�9v����t�吤aFȩ,��u>c�r����UiÛ�?j���'��3^\��v��N,�+Cz�%�E<]2хQ�{��]�vH*�q���$.ǵ�j�W��n��S����p�W�ۅB6p�1��L�R�(����ew�p(摥�+��l�C#�cS(�w�@5���Ϙ�Y�l�< ��z�c<w�=P=@u/[��w]�7<��ֲsT���u�>��R�&�ib��w~`�VŅ"ٕ�%m�OI�LӅGt�)�!z}\9��S~����C��Rk|XlxVHYEB     400     180�X�ل���W�S�(8���<.��G�6�o�$�0�O+��܉e���d�ŗL�9YF>���/U�xI �)ǹB�� )�
��F%
�VR#Roe�
�^�^F
r��<W�o̬Ʃ��e?����c�c�
��N���@tK
<����yAo�à����1�^/7��ի"�I{k���p���;�仡�K )}��dsB��å�3�*�ofbKfr#Я�e.#���]S�r<A}��)H*������{7?��r{�r����Uo���E�W�rb (��
^���� ~:/�4J/����1�0,�����׭��*��깛3����jo�J)@$�j;atua���s�cE�r�#�޶�Me���%ϳ9XlxVHYEB     400     140�9bAZ �4�$��k�G�����r���]�����ǩ��˕��X��E���Z \����q1h[ۗ�����o=�Il����F��>��s�(ۊs��@��ɛc((�X`y�![Vh�_��MUr�'���Dt�lM���A@W*���.=~�Cyޢ��軣;�j����� Pbȴ�n?,',ڱJ\��u�y��r3��\����Rb)c��5$�&u#i��p��$�ȓ��[�m�6�O�
��L�F�|���H)ꡂކ�wg/vɟ����y�w�:\v���ͥ�����:�A�gza��2�XlxVHYEB     400     110�0:I �%����hJ�Cg��҉��9��Z���J��52G9�Fzw���:����6�ڏ���؁�x��	�cs���1�4v��H��T�yuj�mD��L���ｨ�"RJb d�&K�'�����zh��l����S�?)1E1�+S*�9�s	G:] W&F�=(��u��w�㦩�k<2�Om����(�����4����@�*%��8@Bh�RLv2�∀�� �/E�#8ߑw)L��	��;1�6膶!��&lZ��������\�7�XlxVHYEB     400     130'���}*�0�j��,��x�r����"&���)aWAk$u2Z�g�2��ƌ�,�h-��QX=��ۍ�� �C�5���K����a�bv�Eg��Z�,z�z���i��ܞ 0�R�������'���L��,s8���o�X_JFG��-�.ٺ�1����l(�����@�G�)+V��M�w�adk�bL��8!��DHW6�^��J0�ג���΍�"˓�����_��D����W"��P�XO������T���؃f�l�
�d�#��S��^�eb�[�2/m;Sa_# ����'�V��-��XlxVHYEB     400     150H᫨�OZ69a�[^`Yv���r������`t�p���4��Q����B)�' g�\�43gZ xY�Cjm�eT�$�Z7�?Q�{%Y�fix1�b\j+�u��xiR&�I�[/�1����=��-̪1�DG��o��RZ�
OyN�+'��g�嶳�n�6x�2P�k��ÛЄ��?�q�,����l�K��+�Ҡ�-��fXJ������G/����Zg\S�zW/��0gsQi`t��d���M��6���f�d!�q�j��c	��o�#� �� qQ�k��Թ:i������KE=�0n��T$ =t��g
�dn)�a�-���AI�x�"XlxVHYEB     400     110�����.����u}����P�)�,5�����Z�x �����Ԃ�'0ݝ��K]������jnqcH��%��R�=��Y��ݳP'ʌ�[���)�=�R��Sn���O^�ك��p��7�Lf*����R�+�٦y@�j��AJ�͊4���������ö:ڴ�u1�vKV�d{� �#�����5�0���8m��+H�����e1|J�����T�z�����6ڒ�df�*��`�8g�$�z��L���aY�����q��s�XlxVHYEB     400     1c0�hHN�	�(����^���/�~��c���${7�#80\B�)
� cg}�ȧ��Z���T��*�$�}ѷ�3ށH�>���젘�Jw����$�ϊs�׽�D!wV��O�q�R�7X֒Ǿ��smQ��x��	��w��0F1���{ue�����iL��o�H��CY�U#0��Mn"��X��J�)�R��ʬ�� �2���zE��T>y��e��z埏���v(���;Ʀ���AJ|��;O 3	�O�ڌHͱo\�?6��vq�y�w��6�@�t�&s��gR/�'�� ���p � rq���R�4���t���z��6�`���m�W��Ww1	kF�m�[��u��?�vƏ_1 ��=4�t���:L�����(��eKF�$]�oQ���[��48�/�CÐEJ`��q�i]X��FHr�9����QղXlxVHYEB     400     150��w�nK<GS�[�Cs���?fgi���N�u�C�VNA��W��a`F��DB�Q��(��>A���.?b��u,�N�/����
X��zc���$,i��Ƴ��9��6�MR?�YD�����8J�~t;(���fE�i�����b�:�J���λ�Î9K�_ /0�su���&E/�����`��܉\��[��d^L�"���H�[(����n۾��H��r���On0М0�m�%s�H�(|�Gzvǣg�oʝ�f�+��m�����A��:�6�C��İ�O��*��\
f%_q�7}�Α�FX*�^�C#�OH���s8�XlxVHYEB     400     170�0ԁ\��%B�W5�+�M�*��t&7W�q���_�ZD�"��Nӱ��%���[]� Dl�S�N[��b�7C
@�=gw%��jU�/Y��~f� ��\Ь��R 6J=�9J���z�O��C�Be����\�t�W'���[��5��M�� �zD�	�?0!��:yFo��A��YCs�����X�����5�.N߯������=�j��++l	p)ɶ�ʽ�����d)��HC�%���2*�FS-�֋.���MH�S�Ŗ�j�J��P��&���;�˻1v1a��1@��A�nG�!R�Iצ�G^+�A|�N�F�Db�V\���2��;��k=�/ҝ襉� �hb������XlxVHYEB     400     170h�rԇ���"�}�[��-8jM*��T,ɹ	+gʃ�to��riU�v�uJ��r�i�"|Q0t�PD��⍁�A���hVu�a����\υ^��9,1|�PZ�;�
�aS�m_����t�y~ʪ����]e�rIUA����=���'y!.��z �IkI�_�"ikҮ��|]b_~��=���F����>2�dP%rrW����#[�1��n�IP48&�����}�̙�m��k��׫%p[�_������*����P�Gw\�F�נ��R��v�!�+���ۣc�������
O8�@�r�_���eR��b�2��A�X6� ���Y�u
3������)D.Б�vn�d�̑��XlxVHYEB     400     1f0�i�>@hB�TE���(��������~�0�XYw��}r������0�DBm�\1��x��J>�M+��{�+{~� ^����݄�2�t��uI�*��h�	&a6V��c������Wg����(8�x�BC�\�|a0������"���
kK���"�E<�i��}+5Ta��[i�ߟ��6 b���eĹ\�@�斳g\��Ӣe_yZ���I��ool�E�	̇����2�	�3,�0b�GW�sM�ZK���6�>����+�d��!�sd�=�����K�����=�Y��0����'#��^f�"7i4D����8���y!t������=�D��E��W�6���M��Ho��	G�Kv��34� �2)���,kZ�x��*��e��$h�VC��ϳ� n�g��^�&h��������M���;? `h��Q�r�󝱌<�?�9��6���oxo�����c����,XlxVHYEB     400     170-{a,�\Kp��<ӯkr��F0ڙ�ZGFHY�Dcn���NZ�PGS\iRˤ��v}�S^�Jt@@iL�=Ob�,��y�h)��������6�5|&��}l&���͙|o-���*��ؤ%I
w1^���Y5>^� KZHM#�� �������d�)�~��;O�w���m�;밦?M�($T����HR�J�
�g���I�N�V�u�+��8]�Vw��"'� Ⱥ��ЛB\Y�2󨥏���1��y�!����К(B���Px�`tZi4�;ۨΪ�/"�?�j��c����@���rQ]�
S+(gH�i���'m��������/�6�x�������������`�?��b�H��XlxVHYEB     400     190j����OD1#9���N��#X�g j�cĭ��l�ܖR�zU<��9�R	��jl��9��6�pSa	z9z�\5Ƣ���.�=�%Λ���T��|�	��Z�0U��![���&�|�b�ݝ��@@fc�8��AQ�3��v`���b	n{y�( ���ګJ���u?wSak'�2�������w췉һ+»>�S�]@6�D!�sd�L���/��U���J޲��)��PQtp�jD����/�Vmi���Ga?m�Q��Xĸ=G�yט�m���5 ꑃ:~p��X�f�@i��F���;8\*�9�H*`�m� o����^�_P�-u&�3ȁ.$Ư��G&/FQ�7Y�L����S�7�Wp̮1z9 �`��W/���B�^�M(F�`ݎ6�l��ΰXlxVHYEB     21f      e0�'��%���F�Z�{1���M�p�X�{##�{D�%�ߖ/����t��
�hA�X�娪D���u3S����������!#4�� H��3�j�~{� �֌�h��,p+��r�vtbG�M_�{1M�l��{��x.���@g��yrry�&7%�w0�Z�J��3�J}sX�d��Ra#���%��M��*4(�����)��t�{�4�aOh��6r���~ĺ�ݦ�