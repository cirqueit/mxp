XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��h�&<�u$���#�V���7���-Վ@ر�~,�����a���%A,۳�'LW�i�Rq^�ҟh��u3�$�L�<��g��!���L��ț*�Kӓ�ՙn��O�S��F̘� [Fo(	����	J�ȫU�䣇�{�a�K-��@b/��Ł+Tc���:�����`��"e?�$ǅK#[��?E��׸ܕ���:3�]o��]yN&�`�Ǥ���e58h,S3|�P�����8�Ҧ�`�Iә���;<������<U��3~sx=ރn�N�<���^M��.���VV��\�y ��X�i�/с��$�k8cFAV���m}G��!����b�{CAm�7߁�\ �x�ou�xј/�Q}�8�Ԭ��ĪÀѴ(#��F�������Ybԟ+�ݩ������2���4��0ٷ���k!M��P�5lz�@ ƃ�so�]LIA\�p?H�H\`��s�$K(Xy��a�y\�,�LT�]k��A�
�cj�+�y�1�ԸFAjl�f�H�X�u�}��֝�e�o��%ljH�"C����A�v	���I�:r�'����0n&�!J��k�hb"?���&
Íc��{j���->k;OI���.�����N��G@��ѓ\	��ȦkԤX�+���F��|泓�3>yfuy�/��hR`���������+�sLuۺe�b�� a�����n�`���
K��kTt���,
����(0#]�JF�q:����:3��@R'���m��T��XlxVHYEB     400     1e0��0�H㥥����؞�yղZ�If���X���=f�P�Z��)A���˕F^L�#~��OCo�+�&����_�P�H�<�T�ș��9�) p&�eJ�#�f���7�B�~��e-��*�����*iL\�����"��^R�r�\V����v%۩�8��.N�=��dU�ۓ��ì�o�(�N8���RNl�+?"��X����4H7&�f�`�A�&t�5�3{J��n~����M@O�q�R��}�gq�>������Z�~D���^GV䫧���9��m��5G��G*�?C�|��%�/����c�m9�xM�S��LQ�� g�a�����~��a��, iwc+X7	�?�t��z�G��Ta�á��T�⊠�
Y@��^I���Xߧ9W4�����j���n(���O5w�hW\;�柆6{�ߋ�[Z�w���[UJƄ�������j(ַ^��Ĕ���}ЯJiXlxVHYEB     400     1f0��3H�3�<g�ָ�L��V׿�>L	:��E�$��q�Y�vB{D�����^�U��J��SkDv�3V��MB�7�E�>m�2�b� Nyfe�O��9�<00�zn�h��K����O2��z���W�m*k�7
_=?�EN^0�=�,Z�W?� 9��ȉ�f4Q�/��/��E��)r��#�MO�����p�!T�X������X�
�-f`���488���n%��/Aᩌ.z��RϨX>p�;���|�XSQXT������C'���#ކ�I$xz4	�������x�n���/��֛�J�	M�v�W����r�jѰ��*>Y垫��S�	K��s0�#��kُ<�-ߌ
e�Ofئ�i�S�0�A���@J�n�a���E$�pK�O B�D�#����p2У�G�ē��ȚpwK�HD�x����<�wI�Ҷ��}ED��x���ǖ�,�n"�8�/1��$����T*l�Q7�>=�jXlxVHYEB     400     1c0�j�n�%�Й+;�#�14%�A��������n����j(?�6��TH�#�xu[�	z�-�ӑe��-xL�n��O&��;�J��1���|7�-X|�^�@�:K(�t7G�mFQ��1kvy���3;�2LLg.#��œ�����n������ CwTQO,�;}:��vl��� �[���!mlG�8)��a��^E�W����)����E�^�N�����-V�K[�#{�b����V7).-�f
���	ˮ���V�
�!�fH����i	���W8)}3JoӔR#�0߄&� ��*x42P���TÏl��O�ֿ��f�;K�y����z�-'�fm��Sf��=���Z��PuLa�$c��u_n�W��	j|`i⍫�	��D��i�=	kٷ��磙��ƺ�O�"�d��8�t<����uw�7_��q=zOB,n��7�'�%�LXlxVHYEB     400     1d0u�/��]{��D�"��_+�a�8�o���t�YWF"��0���Ի�ɸ�N��|��!Ձ�Y.}��Gj���N)�\����b*�Ql�Y��՜�ٞ���E�D�zXNo13D��d��GB��6�3/�&� ���)�,w�,�=�X�3��ݩ���F`��L.�A�xL�De]j�_�Pw��Բ��J�ͪYT��(E�3����E.Q�K�i������ߛ���x��,��RL+m�;�8���pYT:�͖�c�h���\ �o��f�u�ۚuF<yQԪ^����^f��2O0Gd,���_�������rU$Rd�L���N���fq�$�W9�Ql��$�*�xW0?=��n�����	7#=�j>I|J��ت��}�˧
�?�d��^p���4V�H�h�!��i�q��H��V� g7:�9����nF�:g,�WYn�J��E�2�L+�mXlxVHYEB     400     200������3�E|S�$�f�����N��CN�7���/+P��P��m�F���^ɚ��5t;sl�2�jEc��w�����/����
Zt�X:�ke�>����Vj���5�V#	�dPj�\�َ��7��>�_�j��&tD�1<�'h��P)1���K=��)�r�-9	x�u�R5��1@\�'�-GоR���^�$�D�4�;�[*t&�*V/�����8���SG��ywv�~��;2�q�O�Z������k|�6?.�F���ޛ��[V�K�c2�NJ��k��v�r\jר��'��Wa���9zT��"�;���#�${��h"�'�UDYT�x�{Ҟ�G��fo���N ����Z<X|��-�~�{"U���nNq����4h:}��O��S=���k �:Ḯs��εS"��"��r@*��Peݠ��Z�זuu�l,kvi�|@��dac���N-���-FC.o�=�)����R����L����̠�2���ݠXlxVHYEB     400     150��`����tX�~k:}�%(˦|=E1�ƣ,��-S�§��4��8>��|��`"�k8=�⮲��h)4�ɓ��J����_�0�z2�ak�����a��4�\۞m�^pF'�dY�ʧإi^�B�5:7�U�+X��&���1t�����;���*���=�0�ފ���pS�r�7�y�P=��~g��s���w�ok%K��y����k�C��sx�~*H��l��S��S�p���|.���.�C� ��F#�ح�Mʢ��g�f�X���,j��V�fgkf�+�(
�H�x����	��bݙɀP>S��l�K俓�b�lzA|8� �����IXlxVHYEB     400     170v���rS�(A�2��HH�T`�D/����U��k�&tZ�0��J.3��b^JNM�N��D�3��V��F#+pƽ�Ք�����)�.v� ��j�6��T|�lQz�h	���Bg��{��ܸ^2}�Ώ���#��r��RR�ʞ�3�#��8,1:.ނ�/�Kr�)9�4���-if���Py�� �f[�|+��EDg��-�&?��]E��h	�=n\MM�?p���H.�\�X����Þ������{�,bAp����^ɉ}w(")wu4M�z5�ۦ@2C�'�D����
�Ǳ�¨<ݡ`)B���i�(�������y}��_^Ŏ[�>��c��⭐H�(�1*����r�菑���m�T�x�^F�XlxVHYEB     400     1d0��L��m���L��(V���y4<PW�e�3��L��a إ>��V��bw�� ^v�ۼ�$0�0>��Z �W��g1��+_��y��-GևV�R�}UV��+@ʝ��o���-h����E��c���1_�.Ի�W��zx8�-��iFl �-)����������ʠy���+�'�u��k��=<2���ܱ�W�YԹ�"|Plm?F"&&l�@߰O'���5���r��mh�,N����e��zi����K���G�������6��S�z̚�/`��{'��:'._����e��._�U�Q>Z��@w��>4��#s�������H�u�Eb��H�yM&��a��{��7���pM�_m{�	�p���!��.���Pr��-�6]��k	jݤ�o�Y-���#��ݍ65����F#f���� ��7������7фΦ�Bt#�(é�&5֊�֝XlxVHYEB     400     190��gє���7 ��I��?�W.%����{�|�`Q�!r_�g�����P۴�ch���PtdU/mm�����[�9pZ`�̳&��8v�\����sʀ��ѯ���n	'\p�n�Wm�)�fUt�1K	&���)S���|�;�b�n�)�K[���N(6��5�t tQS%z�c;�s�o��ѭQf��Ad|�H�W�SQz ���.'58v���<S����[Lh� �KbkŲu���w�q�Rr�
h��ʗtIڈeV���A�'l����;��dQN�!��4*��5���{�`|s�f���N��Y&9N#^���,��extunzǣ���+�VUٶ��pKye\���\]s`�w����j~���}L�w룾h�q��\)B��^2*XlxVHYEB     400     190��ﴞ��I�dcc��%b�s���'��>�sI?��u�l�2$|�0C�N�.j�ֲ�����X�o�˦�],�~�4�J��SW�7�����UD��N�b-p�Ox�_t=%�3��|ໃC��g��:���JJ����,㔭nK~( �O�r��"�aL��~�/B�!������V2�����Z!�T�;�M ������-�H1D���P
�rc'���hH(K�0@6󯈄΅+�$u��e��7�	�E��x�����|�_���y
/˵6,��i��gP#gO��m$�M�U�Q���)O���=�`���NGtIK][+�����=���'�s���ݭe�	 �*�k��6c��������s5R
��~6ر&
>�� 噣���t3+ܲs[DD�XlxVHYEB     400     150h6f�1>E��3��bq� "A��8"]ٓUIp'2ζ~K]ױ;�r
��Ȓ��;���!P�FQQ��ߕ�RR���V���r,y�Ҿ��(��k���<{cr�o�sԢ�e�D���������b�j�\��&E�*i	g�kx��B��M5H�\�ѷ3 &@\CHR	�I69�90��׎�j�b�<���������<~�[��������@�h�Ja��nQ����V�V��`�޾*���F0��{�*P�]ԅ�eLn��̚n{��H]��wM�sQV��~�P@������/��L�H�����|uk��y���Qx�FH����:6XlxVHYEB     400     150�y do���NU���p��h2u3xq|�Y��Rr[ �'���I-C!�zl�pϾ�x��"?��S���{��A�/��w*{�.2��m5�)Up��������	pIv��dK����}��Z�ό��Wr�0���4s��V��Wh��Vtӹ�c��v)pZq�!4xK�����(OFt��6i��4��f v0��]�-�-�H��IЕ�Nl��P/����`y���t[ש�rtnKs�]3��h�D/l�ϞL��hJs���u�}&_��UY����7�E�3�N��Y�I��s��� )�_Dl5�Q�y�,�t�!�I:�r�_A5�xXlxVHYEB     400     1c0�7�-��a�3��6Lj�p�c�X�o�/" W1���S �
s���)Η������~N�U�~rf]��R������$q��m���%�
y�EO��
-e�S�4��k��qZ�d"1�^�.+��a~Q|MA��b2������7�o����봪�v�U�6�2�g!\��;���0'H�s���f*��7<A���,�V��ȈC��.�����A8D��M@<�cd�Q�c�)��(%��Ҵ�5���T%�����~�%����J� nI���}�ajd��xo�\�C%����F�i�$[NPA�m�;^��}�J��<:UW�.�o	�k`�Ԉ�LG��uY?���/�Kb��w��~��� D�eM�M�\��-X�a ST��G���iKN[�����Y`p��X'�?��tj�C*�9��XX��22!�D�|�m��]YXlxVHYEB     400     1c0���+y�aΈQ(�a���	V�S�k�,K�SH�	��)�xke�T0��\��[7H�!/���g�J^��c���Q��;bf��)3zF�3�n�z-DϜ\��5d��4�ڄz�����ؑ����"XkPQ�58Y�wp�ͪ��V�$%h��'�ۘc�8��SonZ{��s�U7aV��0�(���{��s�U�6��O�T���(�S2�O�>��u�E�A��"Q���䬓�S�l����s����MVZGe�߁�X�Ħ>;�?��|m
���Bl�MY+���C0b�Z$�H�����&u2�/f�so��f�q�Eɓ�`�z�4�|���uk��J��ɼ�5}d@Tr��eT�#=\�ܠ��Ŀ&�cB��
�֎����B*�z���@��"�G�7�$�4;�$f�2��_��	.
����&�T��;9���"�����M�B#��P�T�XlxVHYEB     400     170T5�%���]u��r�H�`����#�"W���g-������:�D[ӧ�.����Ti(� ��l�����H!��1�}�Xko�.>������Le��15V�Lt_�l\�+gmR��*��hq�s�w�S�~�kI���|�Ӈ�)Q�?�\���)!ΰ�'v�ɵؔ���?YBfRU�\�}�:T�(5���v<xʜ���L���ia�Kmg��7WV׀���q<�7�7.M3a����qD��K>�H]p����g�.#D^���E���S��"2j:�'R�1��C�I��B��3���Q-}��"j�r���N���=�,P���(m[����h�i��iy��u�XlxVHYEB     400     200+�
�Z�^����an%(}p��8�%�����V�YN*�����XHLg�����#�W.��~�݃G�R� �ˡ��JX�HV̈́��Jh�����ոh�v_Μ>>�C�Βt�iD�RxO"2ܐ$k���Z��?w���:������ޥi~ް��&xo���j��vc9B�:n��N������v��'~`����V�C�2�[�s��'����^ "�%8��=��ukoS��>���ɗ�b��R�t,������F����eW��	\y<��+���pXb�]zP����uhSK�*�k���4H�'��� ��^��sN"�(���wĈ�9&��V��"6����"��fcx~�Tjj���z|���X���oŴ~}n��:�������UDO��o��O؟y���q"�I�O��o�Nn3�ƥ���e)�Hw��z��[��Ib�v�rd��@��ܬJ���-�;xAOw�s�p�E-� vJ�:8�T����<�o�����~5*�&XlxVHYEB     400     210�z
���1�&f�t&�l$�)d���w�i�+���D��܈Kl��>MXK)��n���m/�g.�4�x��*��&��\����#��,��[͆Śy�O镍��ǲQH��<�^���7	��i�ߋ$&�lr��7��i
U�����$����6�B�nn�g�K;Me���m�s2B�%�'����mp��?��'�*��*�]�γ�:t���^�+]�/��@j��@$�#7�U�K�$Z�V�t�wd7;^`�?�L�F�U|���}�<��2i�vvyz���qа��Q����p�M	���S�⚗ Q����gL0a�ML���_SD��}���|8��OUt@�,8�Ž��z���k��5�LjEL��v5%Fq=�X-ߦr����,��S鴓rR7�
��\��J+���'�����5����QV�O�_քM�94�Cw5��xM�����a���,��9��
���?��Ks�aN��U�{�ak*�fM��5��u��guL<���^����bU1v8�CXlxVHYEB     400     1c0{��P,m�����Q҄�n��h
��K��B�.�ntu��8����7<�m�����H�:��iA�d��C�ɤ��~�j��Z�u�폏��#_�|� �����Q�U�Q�=|}����?�^�b�kp9i��a�U��]����>E:�][u�	���q�4�{�ź]�����f�)9��v��mλ�q����X��1\�aO>�p)Q�Ă�}!GQyv!���(��:L�j���0`28��YW2J ��/e�Lk�0�8��Q� !�*��}�C�ݏ֒s�
�T�杭����f#���y�o(��p��=*.o�[���;NX�Ld�ezqAϖp�Iw5�`�d)y�����f	\��]�s�HS1���6ûi����vQ<��ʇ)'2n?�
!���.�g;�bW�֗�P�}��")#��XlxVHYEB     400     160~�'�)%��b�pp�����B���b�4e}B2�q_���#_����EA���,�pHg�Հw�;e�o�˙̙�2q�z!�Q��ܟz|]!�0��ˣD�Dϙ�O�l���O_m_��6�Q��ֺ���JÅ���;=�e����}R��"ܿ�0�U�+)�&�����,����,v��a��y?��ɧ��ᝄ�3��2�ۊ��]�U:x*�!ly4�:o���F��+�K!3I3!�5���ݼlY	�lK��ם��Ѭp^Sl��qT�T���������Ld�(Ə)z(V�^*��;Y�o���%���m34p����-��c΁�.a�5{���B;\w��C�+�HV��XlxVHYEB     400     120�͡}ku,u.e�44vd�|�g�����W$I����m���/�$�Ue��q�.�(�������<ƒ&{i��dkh��*�k�+v
���%A04'23���8�J��O���_�5luc�X��}�-q<��F��V]�Suy�T�9��3�|Τ�>uA.�kP3��p�y�{V�7N�.Уk?$d�/����T~��W-`�M�-�n"� 	��U� G�g���n\�l_�X ��I��T��q*-��ߐ�?e&�i�t�B1���g�|IZwF�'�����p/bXlxVHYEB     400     1600ڪ��oNxG�\�wR�ze�Loj�#�\��ӓAֻ�g�)z���l1�'N{���6YK�f���\�Fo����	T`���l���:���}��φ��O����`F[ �O�8C=�?Z�:s�� 7�$�����kJӪb+���W��~C�0A��o������dM��v��A_҃BW0�\������Y�l�t���q���3�	�����8��T�!���K3�\	�%�Ĕ\����WT*!��<2,��p,:���~�|Yԟ`�?���a��q�	�"/���ǻ�*�
��F�|�E ��n�Y�M9����*��!鐣�0���2a�[�(v�'��`+S�XlxVHYEB     400     160@)V�I8�~��D�C"%M��������:)l7?������}+�\���p;�a�o���x�9���[�,>�g=��nCk�#�}�v�75Ȧ� ��K���?}�U����c���9}�>�v42��_���6��z�4���	FS��E��c��J-�R����8�Rv͞d������P�������^e��1���<Y�T�I[������54�ļ�rI�v�S���W�Ea�a�-����P�B�o��U��������rčr��A9������hG.=��2�P�R���S���V�f̴&�i9ZĖ�
Q+���m�ũ E���% =���S�ɷ��XlxVHYEB     400     200�8+�P��N�<0J�+�q3c�l���y�]$����F�I���ȇ��#g܍�TM��V�Vp2�^�a�qS��G���k�q/G������p���6����`)��T�����r,��[l�gK�}v���=��[i)��U���VB�2�lv�l�պ�G�4twa��eǌN�"�:�6B��p��o��~
��BO1�]�?ǪuO<$	�n��~�)�4rޖ����MF=��9�x
liO��Y����o��K�S��T��	Ф5�P|5���"C0��ΣXϚg���,��F;Ħ��D�L�43e����ZM��^S���¨Ѻ�$>�ߡ�%���Z����OF<eTQ�k����u]c����8�7]3�x4xZ���l��x��l �`�A-0��yb�.������0Y�*��qu{�M�r��ði�� }v<�A0�0_JY��	�#[b[��1�Tb�?	h�HQ��>���4��?��咩�*�{]XlxVHYEB     400     1d0���s�Ua���g?�YjI}a'QX�X�|�,�]��g���i�Ge��㪈��;Ø렪=Ix^�����S�OC`�'?Y0��r����mSC"��Bfl��)�����X,���Zܵ�Y�t �V ����5Y,���
M�����q�K��D�D��JXBF���{EQ�Lk�����5kuB����3\ΙbǊ�ݹ= �Ҋ{�:��h��yݦR3�� �E�ԓBzI���tRl�Lx�O\�� %Y�	���s��v!ʗ!��U��k'���MdZ�� �bkòSkb��!�	�4�)��b3T�G{]?(c��_�ЌR��0���ߓP��a"
Fp�6�O5�&~���_x�l�9��.��
j�r#ޓh
V�|������������`>� �t����iY��|J�%��Rg;��sp� �1��JMA|$��C9�U�:��|m��mXlxVHYEB     400     1c0�}��M����l#q�H�������A�g�b��~f���*s�K&-����0�I�0${b�n�7"̳��޳�#�%�<��]�́ҕ�8ɠ��a|KS�(�t�7�,צ2�'�f&�y���೮���i��,���f.��#���!��$:ǔH�N���!�:�M�n�G�+fLJ����?�H��O���޹mp]p/5��G}��͖i<,n;�~��Pa���`-T�QVH������L*�T��LYv��B�`Z����z�`�g�׊��Ӿ�c��l����fiN��Ly�b��>? �;<���W�:}��xJ���p�!sdC㓉�����==���J�x*��&��>[�;Z�_դ��=Z�Ym+�P�ZHiY2��%_�%��
�&n����M���0���f���:��)�[{[��&�*!�-'�g��;�XlxVHYEB      42      50u�w����wb`���O��<U�!�|��J̈́+�BT�����V��RX3M5�4��pg���u��=#Ac:�D�y�W�G��*