`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7472)
`protect data_block
5Rwm27jrNWuZQk9YWD8WcTA1JdEzdtqyckTfdy9cU9qNRULoap7+oLSrXrKqyFi2wau/QnKhGrQ4
vYjSKpj0RIEEpBLGN5BEmMck9XS5NClmn4V4pT6A6oLkXAVwxy4aChTZXhBrPBKqHFomOYam5CD+
FETnbSIdS3Sotn5u/d2J6vXIQ2wb/I+4625EpiFmpYurq0z01nPJYjuWUwwQApJskeQvQig4zVbR
ubUgECEnptS9MCLAPmhzHkvC/gcRuf34eczmv3mHrI1fedKNdrufyyOsyY7jR//6APjhxzzmozl8
EbyIA9Y7EWAQzKqUHAGEFkh6WRTGD1wzfzurGY7/1eR8XRE4UIuxvwFWr58KPxgYN3/lQGLI9EhX
1POConKNDyXFWEPjojKgz5zYNDAnesPIgTCEtxDKaAn0ccgiaA2uCxhgk1JQANAD17NFzSPB4xkF
ibIT8GrPdUa4sqbgAE7CCSRL45d+IukHAzrKC5ALxMIWFdQHvDE/68sadqk8Wm4LR+FABvlMAcbt
BTYrol3T/wbvwy/39xZ96jPQ8LruUCXKA7YbjEFfuFIfUHATXdasvguJw8Rb25FuUe8pAGs4yZHC
QHG4m+GPUkb7YTL2E8f5scPz0GkTnI+TM7LPOd3mq77uBtPrnuuSbehdb2G7MZ2IZbJAEyrYqOu8
Q/pgFtY+B5ouPdfEYQKqxcDioWz4OSitVlRMRVqqjDtauW434OLnO4vlU+srx1fVqTK5W78NHmTz
Mt8p8qEGqKN4bDPP0fdVdOrAEgSZ5KLFc8htziHUgdfhL+N9MJ2m9icWnU6PSKfUwK83eoRwNpek
B52U4IkL4G5SMbkjqA9TxiC9yHlmSMVYGHi5TFmqmuDFi2fPjcntmQ5u5pE6tC/RYqnmGZhl70JU
9C/9feW5ohmwHmWUZcnAC8kRHNiAvgsh5AaXkkP4UVETmBYt/85GLyL2WdSSdv/N/rx1oo4vJuk1
MpOcpz7Lh0j6tigVVKdpj+odADb9k4QHfQPIUM7XTuYSbrIST4UN88muIarG9yx+i6fXrHuTgkXO
J6pBO8wx/HgGJt6LTOmWFu+aMtW7PYxsQZ1iiFaoJs9XeH2e/G9611HbzkNSOKOIQ2iNnEXx38Nw
l3zrmrRcS3R/YatkXWRz8iMCpar//by7cCvmAY40brw0Tul+SSki2VaHh8GlBPfw0nKLevcgmXjy
l/2OHXKxbY9jfVIrEv+dPV3p8lpdJCfUR0rmuW5GrhNKbWSqiPG8ZaqV+ALixXhhMaLPJVP6DIcO
ysSSujQIaRlSO4dN3xKHWOgub8wvTIqjehpDvbJmh9OGVuFArCFTQdC9bIfgx2J+oMTH2V+eNpI7
pG4yazG9hEiM2n4JIoIMwZfCbXFVivtUmhkkkr8Y3/MYe/hUeWmpc/AxhpJlCgLWm9smw5KEF2Ek
za4gSq2b98xy4ow7IUaT0U3EN0GdRgEuKkdXx8DHBxzaBlUd+J/GhzkldwpkfcNtiPj0TKda8F8a
bdA9+KvdyPwDUBS/JabSOt34D5QdEVFIyFL89WTlPIvZzJuIoTYLtChBaO21pfwXoxItj8uHIYPp
wwpwBpGZpi+NjuVSYRmuKsNo8tQvwm0GoOuW+4se9oRGqehdCJuiOvXoSNXW96fDWPLOt+xrI1iQ
e0KvTim0GkEu3u10uWF0Z5AjvPpqPPfyfYolBfiE4jg1ukXxTPEovTX6DPMKccQ2+YranjppsVMD
7afWsuxLOu+AIByFplV8MFu596gBoZzz04Y2Iszs2JmfyuPEd3AThdZBHecdM6AvplFkIecB4Cs5
L76C9tA7AX2Oi4aoGw2491/kHaTFGe2lOYSVweI3939Z39nzz/0/nN20C7ctKngASI3ZrW2Gu027
NPK46QdXk953/WhNynbW5/hpin/Vss9TtJh6m36RV3I2uMDPbUyWkQbLs4gTg6HotE/jf/51Phsa
HfKPctRxJKVeuEE59pJc3uExiLnPmY8vgAfmlkD+UQIJcn30/0nvwu98zYa3Vks1ofORxqej/y/Z
3672nTX7DOjczaMymnDM0gA/MABZz6eHgnhRviFZkA06PZ0GBwkHrOWh3K2Ko2O8BsTAtk3M1TEl
YrqHvayVkiOQujLYycaieGgxIqVdt/LXWA///JGiF3+l6nxFGlxMTaR0tMT2piQ6tbaUB8+4ychr
tmfU38NUj1WLO3AYvJhlAGm2rtfzGgf3ggKf/Kkn2xlTTGLoKEeWIbqcUUvZsBRdkdrIW7GZDA6G
hjR1v4yuUXTZEDD2bqqgHh+SlsrMvRLQ0+4hs2V0z5EdPi4zflGGCwL+9ylzPSvTVvW0Dob7xb0B
CedM5mFw/868hEOvVaDkVHq6f7E2Ew/LKhUxwZH9J9gBP4CoC7HP/uKJhinYUyIEo2wU4ptYOiPR
flls2RXRXH0VVT5m/rDIQ6gsfuOgZZF6oQInwq4HHGVQzfRxkYeI4v7BWkZOtD0b/4smO9Vj0X+b
c5JljGNiBsmcARvwMF/PCHxs+Xdl1jXow5jS21S4og8JP1OREfXoDKkOjgXHUbZ68WYoIBLVbWQH
oFioNVG5RmSia2qO+O12BUExs8n22iWRUHd+Nt4ONw8wihpDk+mOe3FjEbOB6NgNJSlWJ3zHHyRg
x7XSy325I8mxraDhQK3KlEYmlRAjyqz3BIjRtXr5xXcA90SJITs1W5z+7asXlj4tEhZXtsToS0OA
uXFYnolNCbZPTSQ835+fo5HCgCX+fWcVHo80kDoXan06DNp4IhQQlvoK5EMz/I4DQ/gqsmiOgQbT
Gg+xytwiPLwsACCKXwvPwvA0tm4UjNnwTwRmY7yDgQIprrRvTpeUkdBfpd2z1N1c/V23g3710woA
9PBNdHyTb/rrxM+e/Hr2uvFTXYHExrfeA59ulslYF++t1jmjMWBhQXW+u7MNkWsIEOXYo/oaIuyN
OOJWj/9BmY9pd0WjX3+wefvj6GHs4kofenoZUF48HGBG2f1YyKsIgixBm4nhcntxgGD/ev6rMh/v
LVwIv4Jo6pe5nBMwjBVPrYkI9AVKqqrrY1Sb+YEUaDED8gLVFKz8HOo3Iw6bWQu7OX4km9B/6eas
bzEeyrLxhGG9L1ub9uVlzvzQzZxo4DpwWr62JRgCKCyzEfdRbHSnDkULktj+qUF7igaNFoqY78cw
4PgWiXHB7U/iVofGscksOaL92+nl0z2qTfbM76nSJdIxLatepwJT5lzEt/FYNbI/a43iHWMNkrCw
4MNrARkDWduvoYx5w1x8ezpK6SJBlR7PqZgf89izdQQ1SZWsxPutksZpIBlePynxL6buHsu0cmJs
J0bvhdcsURRrErv31vIagUJELNszSw09bx3PxF4B1bowIolW1OgvuE3LQj3eUBUtLwQgkbTyMtd+
WJqS7wOzJtuPdC8CY/wi6PLGdlqfFCjON2XzlprUq2/fZwAyN/WdxO2ND9PHDr/shgMhzPl1HpjL
K3x4IcCkaBSqOhDAXl6BjVgOqj9yhBv7eVEU7qgS4m1BAfiLLxvO9qzB0bxdvAFob1fqjlCeBtRH
mWuUyqUn7bHQpbDP/Yfy2JwE3S4gUWTgWT629ODhEXREZqDbmgARCw6HG3b+n5lH0hgKyyzK0Buu
TdQ5lpiR4Fl+z0n2IGMBGprLfOuEPfV4/SgVPixIVtpAIxwAqF+Hc7kSUueOvEVZ+cSdKzWNSIIu
qyjostMK/2McvMFWLQipz2es7Mrs3AG/eqBllJIrdVlxMmSZosC1FqZgG9awxe4ZkZLOoofmEZDj
10ogo6rKnJGBRATkFh+ZpkPfY2UofUR3gdkQKpl+Pejj+M6Yh6ObomVR11RcoDE54tMT2PWl6rUE
orVMWIv+7hm1E7uxedCMq14Rb3tKiHPFKz9dhFRsitsCnX8MLJt9+qT4ydpJM4bmzpDKxmo78A49
98qY7lBZij6kFOLsskPykrWHezlLrXfe4VWuxzEasBGzNxeuE5KQD6lOFpIzfoC+ssmL4QDUjTWW
gDbDybVDTyG7/gf2zexCa5Qk8KPw/PJO09K8X2HgIUb844I1HwkbRAa4ou9pAWWWv6JF+LH3ME6t
dq9lJTaSHXovqAh2kczXcsgVuwK8overK0adn91E99bs0EO94UjjlKTFSfzx4vmLFJ9F3Q/Zj/t9
CwBCPMPK5AdIfyYXm4a8T58KUQ6fW+c7u+6Et7Rwrwkj0e5g79A3O5sjIpDkDUsqoOd/2p9vDmxn
2WXBhBNgdJLeyh1z1KpKRw96s5sXqo+mCdF3wl+MzVbnArQ51+IFSPgzl8fl17zWPJT80sTDnx/O
Te2ONseuZ2F/Fe6w/q6sCgv7RBlcpvoF63zXVt3JVySHU9d41ETZacdcc5d5+GPLsAX9i6ZR+C7J
S9aQ/6KFSRFfmhPIjAomm0eYZ5yJ0Zlb6uvJRoYN0GIxiukNo14olSAkj8Uy6FHsS37DWB6x78Mb
+qDyAzAqvOYCPTipeC33md44CMGzovOSIcQgDZ7+ImE2GmwUKERPS9ZrSZgrH+SGaSu/YabBdmUA
4dzpIbMLIpsw7nmsF+A2rf80VMaV+/CPCGliB6BVdU1ZL6LQ3eb+vlpbeiy1R/qBfIW0BUjOQjXy
76SGvKvo/HN+RghvLSlekA6uctoD7SAU9TRhFKOYB5wdu6qOado61EMaqk2Pmj269Vaq3aHnKMLn
A6aBYXjfyk1+MRKQaGwhehADMpnPZUCZNlgFZbC7cWiAve9VyRz3FQtC20To79hA+X1/ob86Rwv/
VovQedfJCcUoN21ez++w7nUUfc7Iez9kcvAsznm6+M4P96qC1nrPE6nNRKncxwGvmx1+EM0g/0CQ
SwPYnHiv1Nc4fm8MW0Fjy9dV0Ew4WBbMC1W3phLb9KxVWKmBqYBOZQNwX2A5qaxHfrYzeOQTNxEZ
5s9RgHnFrqRNHgUo6olhxgersoB8/HOhYgXoGEBQVolQnfRvpfH/Qm9v8nr8LMHuK0BOS836eA/+
Tm+M5T4rhopCuKBFvdT/qLy7XK1fDiSaFZCjg28tlELrLmEAqI3/HyeT0UpPmL1rsM8tV5cx8Km5
Cw8MGRmLYZMO0hVJinFZrOgOl49C5nPnR0UUD0wLmI8kYqvtmAv7eJMPNvRJN97AmDrnP/JJ8maj
3Jd8CNRoIQXMshqPg7bRGm3tOFWXO5V3+3BAIB9qAOB87wFQvLXQ8b1AhQa0NK4tDEnstL9MuLEK
OH4q3r5fgODqgESFxej3pIdGe99D6e71z/SJUhN4dbgDpod2CP7oJm58UrvziZ9pcjNa5h/kdmIs
is61PkTAP+ZAKb1EaWFwYIWJdG2yFo6RA1VQcLF6MFUSCG5eqsqUr1ZsDYAnPLom+UT+ZxfMB2/N
oOZSbQKUrmDZI0uOJ2gzZhbVpsZJas0pgsitYuDZ0nwBviD9rMr8IDZ/R1sgSeLRi2iyioVbjXbN
fM2uSVUcyPUgO5OmFxdFE6yWBBkpk6eP6GBZp4DeKF5HrihQk63GWpcMbT6VllexmfnmUPuVq4Gb
nfe0/yXwgB3YQCPbMvVNkrXLyr1VKF8sMyvGlKmEHh9+I3PY6USBIYQemjxeC0ss1S7H7Rp1X5Gz
YXMNo/InJaZn8Whm0I8OwMGSzBwc7ggpzA0SE2aJewLC8wjWT9xOQic1YS/jSyMgG/jMD9cpH4n9
LmLO3Pt4DE31QMgBI09uM35+MDFJuqjpuEBWXHISw3cLwl8Yh31cZzbulBOG091ADzz9Ztoh9/Kv
32yD8+jw6SLaqm3BykPxGBj11iRYZccz+liuxtnpdEUu6OCHQmUq2lyK1e5+ZzI1kGyA0hywtHwE
OQqSABP3BV2FY5UcBzsiAQQsl/AGjQY+hgXGrZD0j+CX5uN2xsBrbwPj4Y9PFGiNMtOWKD6tyrc2
KH5wcbGwrfaErvPvQgkeV07qSZLeMrio9sbrOXlX6R2pAT4HoD6PYyfmhjM/h7CcDJh66mLggpf1
gdax9f5uZKeicIBwSb2coD+q6Pxr4lB9s1LpS37c51M3b8OJDScqw1KsuWX2Ss0l+9OFDu0GZsUR
mOVs/xl0yXwSfUppRPPNUOphn320O9kOrqQrtSF5Ldfbcp/FdM2VaSqx+JjQO3Vtyaie7hI3z3zt
5mKbw7BhPlQ0u0TrDa+9fF+AevLvOMeBw3sKjT1IzDrGWWCqH44/op4xBJOB3DScpjbLuwPIQNK2
RVLraTdWAAhEv6+jVdPFdiE8tbYdH2g9qGuW/En66UBlUmQg329b+cGUUehGmGTbetm5DeOgiQT0
RQEayYSodt7K8AjlKvRwsFbU2wUIvKZYbSTFZTXiiPzQMmqRh1gqqP/n/IZbYQ7e57yxd1G1utai
TYcva42IKktrwfhL2YJgC+9VA2SUlWCp3DsCn4zVjOT9h+gukXxU0ZBTc2usvnLWms5a+BPNZ3LX
0bwf6m6zFm+JaLDgAE3ns0tI71Kl4ilYB5UiU3QpWTKfHuGYMNwdQMmO3qLNGzcUHmy12+cWV7A+
rBDp83nhv4eceCm7oQKojMlMls5kT9pU6yoTOzI1pGIj1Pe4AByRExjH1mnSqVLocnxl+nSkOLUU
hHblvKFm3AVu6c4VOOG4Ye59/eeW6Mlcs0eeSBAORyOPXfznrtRBrppPkNb9lcyv+W2/vwA0IQJq
GRdP1x0S5K3A8uMAJNeebeem3dTS063gPaKCO9oRul5aenzJR9VehO2jDDeMCSdyQsNrjA8D5bP1
a+XVeppsgJ/L0ALNopocbl0/tDx0shPxch1JBT8cy1Yrf4jgdtRZUzzjqGJ4oP6NtflAS2vcon/R
udv+U3qV+m7dOIZUWpKwTcxHTAEAm1ZW7Y9lBRNx8GzLSOHECn9eB4zv4nYx2GbayYgdX1OHeJWN
5UYfY86VSBmZAiQezQOBRgFydtrj3KNHcvrbNvkvrZTWRAxkYy5L9RM/5uR0gZInXayslFX4gIdd
K1tZEBOteMD4X845iBsRoike+JaMejLBu5iRPv6f6uPcEokMHGCwaIeZE+79F33P4I2L/rTg4A5z
q1eSgLMp75SXJbignVObDbKp8fsNW2h7yVt3OY3P0zmCnBYtIJwBvqedB1KkEaly1intNaxd0ovA
GX/XZOOekxrSzl8UxVRot0BemnZpLuZ0RV88ES5R/8U0gCbD1Ug6+mQm1jgt8UFiTXYVHVO5szDn
d5X5T/FUIqQgfN/EjLyAEFV0UEk1iV7cSZF+G3PySmQ/XD4VKY6plndglhcb0iz7C6nbPa3A+qsp
JF2wR+OOFJhwFmNpsRUJ4BaquTMcnJmrCGjyYgAgFl+UqgiVqXqgBb92WTa58V/CvOMaIHKpzMMq
/BF6ygHUVZcFGpHq5U6ouOT9X26d2bckOMtdF5tCjGrJLGb6dJHTdynQ+4aqAQp2h1k7Qg+WsUmk
dj+tg3C1mEoDQ3om4/OCdjqFeVpnGARknsIFvxsQebuMAbEQ7iVodL0b6XJwje1Pkqn2keLE85Ao
faSVaNyYU16NmHSaFduiFxlgHSBTtyTcDjhZLI4cgayAoyLpS60JvQ5BB+fDHQr2/PaK1Gk0sdfh
A//A031Le/aQDr3+B5nkEzzi1e3jnPW2gZTqaeXDrzfS2eO/vRSfnlq+o2yAv7hQLnFif0tPyN/8
es4t/NRlAKvlVdRCksrlB0bayWOZGoyyAfV2Q9fYjwiXOm0845VB41q26zTlpUzzfFWBw+ZpJohB
gRxvLz/nVwGQhRx1qU6kvHS3fC3ygyGMtBQJHCYKK1n9Jy+Iji4O5rgqITJ+AkaGLtlAzmCZYwSv
N+85j/Wt1HKd4dR5rs+v5EFJ+L4jHQKJ+P05Q8KuvwTkC7wZvAS9GcNrkrr6/lA9MxzNCa2LRHEa
0kfdMp3voI3vZfTr8KzERW/HolhmzqTuQK0j1d7/JFIysWEXcQ9EsuibqqxQe/AE98EHxTBdNQez
8smyfGWaJ1T9s9CuBXoD6FG1OPtUShE67E6a0WGdmqsAaUP1tVkQrFiB1anbnGTNeu5Ij4kiCWuj
PH+pLt7LzmziWijD4gXT9hqjt6/hV38LP61bKQ16rG5tQiuagy598ZO2TEhTeP65X6jDQ5wjoeG2
QUt7dUtaS1NkgdtQTBnN0Ml9Jk4ENEk6wVQrLPD7rWFZNu1G232FuZjm2rlMdUIKio+lCR9Ie/+r
qwvy106OJMekg92yJuUa2b9uNEMU2RRYZdriDfdLSFjo1JQF+XfXPynSqkopWKzYP6tCC2wpYNTh
HNpxYIkpOBI8BMHQ8NsCjWB9wjbEO0lpyNjaLTH4V1Z3cnD9Cf6B3HlWj3ckXrXRe+K85op5Pqek
RjgiZVMHVAb/XzMVJJC/mBqOZO+MZY1zpHdgqOxCHOZz6Hh+AAj4v7Iq+3llLCchiFmN/DnzXl1J
VyZ4IA/RWIt0QOpZ7eLrO1qaGWbEgL9TzCt/m7VmX+CustQ8m0nmpOfUzNbPAFUTTvJh+fb+AgiX
PQAjSyfUsbvVytJJfZjKC024oPH0edltZ0DwAkFpBXUVo24oyBat4crk76sCRtxSYb4UZrvXfmu3
w4NKNf6YMfQb5NlEzw9zEjf+F6Wuq+fOHGwR854hGaSm1F7gXCd8r8UG6pF8H8Q9rXkI8FyZr1Pi
AAvt7bGJrWrnqjllTfhk7cLTxmdzjJXunzFzj0ISgxNSG81NlSLcVfbJPGih1TySAYFUJpsqn9YX
vinpy1DfliggE7swD95yArdDO8L0ruNQxT+WDtigmxj/1lbaTLIcNWb4xtCAMiaB7Fq/Z3JvHj9/
7jXDPWMFDYITsXl8ifizwoAPV8nzrsPh8jm8QNv/P56yQ9api8lPiceItjp6szJ0eY/J9/NLV9td
+y4VgBfW6heEwyCml923IhiQBeD7gvhPAQDLp9fDXcA2n5k5bmqXJn6Rg+EiXWqi4SFA0QJtBWP/
WoUO7mzeDu27cTNGzBUtU09ysj1Q61TPUuZqnXV0UNkcJMapCL4hCVH7nxpyeIeeAJnqM2nUXTyf
kYC4ZFM/q8yPKol4s4X8TlOPOQh5QuDRunDXKD+H8UGL/sYfGAX9/KEPsqglKEJL4SyhapQlO2dc
jScpu/KEuTesU5WKSaIjOs7sUcSMZrAxT0CNBBmniH+clk/WLxFYFJV8ucVRUd5Y6O1CnkWK/Y/U
RNoVTqDZ8bX4wauQaoK0nN+phg7Mxq5beE3Pb1+IfwCfiGGhLg3vrbWgfMwpFXDQF3U3q21pfFoa
pI5nbo5CbRlj3E35yiD9an6RMQkReTwO+SKaf1nTyrD1CHpWrx3OkTiTcuHt0ljOZKEJ1tjZa4sY
Rp44ZWk+YdnneAk7tUhQTTgfPs9YGBWVnFOIQyEmw3TbVuAcd5OtBQtAo4gWwbYC8CV+7NIsdxTQ
3rKKEjVTBl6o8Yzr7Uad+Gg93F+twJfw6Q7dTI2Q3InKYBGL1oMsI7qTvN4jQvqgpkANhpnwbrRv
l76Skm+2yeT2pO49itPl9QMFIv+iobOxYMqCBf8H/a/Vq/cYG4enkdps3xrh2GYXvOSPvm8exW8q
38OBiCv9ZsN4xlm3rWZcbnlmaQMxzfKErbGPBt5USaZQmaQA//8aRaaTyY8dsHwALvGBqafN68d3
uo6J/6BHy/uDmnOgSKO3H2e+Fy9byqSUhRmruLzDOdIC/mjwhruHsOFJCjn4r3cHTGf0TtZFl+qk
YWjdEggAr6HemoUuHc3sf1sObfxEc1v1ZAPy+JPLj0cLG0vTZPyaCbhngA2JdcwWBdgcO0i2bihs
42RUSv1ZuyKziDHnYsjLn947aEZb7we463xFIGQNPN9tQgZIvO39nyiOCBdYNLxX6mOPcgjHN62Y
LNbUVf6nEnvlaJTa0AIOBVhi5lYNzCyv5v0Kby8ZezGBzHWxq4MbXk6kuqYdF1ISB5E96KFkSQQl
EkkMU+s=
`protect end_protected
