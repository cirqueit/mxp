`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
MoRrf2TWV2LvNPWuWxP8uzLqans/adqhK6EZCOzNMQP732uy2NEbSPXXYOhRq5US8laGRpMb9SW6
BzaGq9XtB7WI1uGSmA9fdn8pIgQPrG9TkXTg1K2wlSTwfJM3u7+R2RpZ7N+DRiRuP2DszQrA78aQ
+PJJRfMK9iOc9qUv15kxgECy0gA07s5aiUiJ+nH8dIsq/mgdiHhRK327b227b5iLpl0E1GCd8v/8
qBPrEXC+b/3d6H9epi9uSV7iHG/50d14YSt+bcPh7t87NUSy1fqU6YoJUADDxcnTIOJWZr7IKmjS
vFsNAcOyUhu4evuIBOLh+U4CMA4XtU63PvhCvP8AZPtV1y9qaqPCW2h5nPVJ9dyWYZHkQRBSJIN5
RyhBGdlIVshBBadsIToTzmNw7pKdutrE9z9BZdmQlAsRnOGPgZlHihdbMV2KKb4nS4KFgM3d7jM5
hN6/SnYBbuDGiteztsom2JislYdp+oWY7qYBolw0NnMS/w6oQRzjmQM2OsPfDEBmW/2Cwp0bE/IK
Rz4t3dTj9eFvvrUjOjY0dC16Alqs87sPaNbLKHX5iw9Y4oSDxkQiCQlhj/wQC7VF9qndoKHmElh3
vZtKr2eFMvDBsyv5z1I6gPUJtDfmuonfCPv32sLN1SwJIrjSk4ZLegEJrnwq/6oT5jP+HIqZig41
HgYZ8FrILopOpiXDUA/820BDwKxCtD4rD1IfuPUkbswnU+4Aq1/jFrDrPV1+3V8q2/ShcB5bXWfe
fnMSeqWLzHUR9dmyaQRfWxU2zgs+K8mx4mb9/yqpfQ9zpYp3bjtSIwczxdt6mb2X3vW6LD9zSoOs
/JZ3PFd+9I991vkyCyKnzJGrbm5mJeATEq1dYCr6VJ8aUEMqe8b1aTetKr/p6lgXlPOfkk9n9qVK
3lsyZTAf1u3Q3xRuDupi9R/YlpnV4kskKh7hpeM029jiiy5Ifasj/P8uMtL77alZc6i+5p6xSqZB
fi1ZfGX+KPnR+sWCr/icOQEcchVBIT+AUsOAmzVv62Py+gdylH2Y475Qr4vSOEqRsIzmj2IWMrIt
dFPMWp7u779dojh5ww3eUu69DX1rhWZnw0dNA/la7pCrVprBA6HvarY8yUR3tikXc+n32t6ke7j5
GjN2ETIv7okrqxOHgkvVpizfCrQjNn7AL5qCLABShtiSscuWnA+H6+V6F+VZB99+P8jWqwDjouzp
JyZfhM40XyWZRxB/itAnZ/C9N3n8Ol/oCF6J9+p4tbL5y07mddkeyt3CC7mdpr+HBJ0eHfuUdjUl
VIEuchMkJpLu1dO81KW6Ur2/92xjv2r2hqywtOZ+OA9WWE7pKRcoo8q8lUqvayJi9qNz928lajEg
STlEdT993azXwuD6eEoeQW/PyvtidxYG/xsKbho/yD18gfhLb0lJfh2hqG8YwWNPfYMaFhrY5YKs
ordTAoqq2t8qeY3VJgKeDbqq4IDTgMQjxREqU7S/nMRt/ww+frxJC6RP0lP/jyRyJD8OuaHx7Fcb
SqreZygMfE2DDLQX7RSK/CuacvsJQ5NGvEHK+JZiuVQti0OB7jBhH0OS8s7aXm+S21zBR44xJeR8
16QmJtP5JI/0wR4/3nmeHbhu5pisqmdhPSAwgF1/qaTHSX4ZmWOcW7h6vPA77+dEXwT/uIiraBDv
Q75myTfgvRe375ayxcFXRx17w7Z3fMs5RzAvLztpyWaKepJOblXyYMEelhdi2oh0ILwK3LHPufXm
BEKb9EtVtE5jBhaaVSLWq8JXZneI3Mf8zLpQocF9pcGToyakHBIXuzMFzVnO8KgZSbw9cKYifs6e
UDjmicVsB1iToF25hYV+dyUPQPg3p6Z8w04FIYqGoFvXoFEtzx6ipA+s7EgPDDp2DPISC7coamDn
1+zZ9oKIJ+E+q74mQSYWZUsyAzFoH2/9AgFPdy6/OTgj/y6we5BtmWIpK3GZWOWHh/UDLMIcKsSj
6qq2mblKQSwI8l8LA4kXKOtJC5+pXXHjjWJqa/fjvDFLGt2cji/4vS2mO0lM8VvMA4iRb2y2Diev
G+QEn572vPchoDsukfi8nHB8AFyeH5RQBX3aNnlIY2b6vlbsAjYNRIK9BZcrvwSVqK73+wnMTOTp
VBx8LxVJlEIjK30zkrDN5qnYRDt3PqNLa8L4KHQ1OHtkYyvidXW4r8HeZwkyjrQrWgdbOQ5u7eIl
ALR3Yfe5qoxPJmcmGpJRwoU3rMUr26KiTXh3XDq//eXQuhEI1w7IOCV3X3NPY5zpbqnjF+W/MXDa
rAthOP+9RFNrFe4pYAvBG3kHFNtN2YB0O75dy6l/m6mM+kY0muq+o2oq/42W5Z3/mCN4DSS44WnI
skFWjcGhu25JW6AzrpUUL2P7ZdOSR9NwbuVTVjcyA58oaeMUVxHgFA7HYs4QWg0O5jzrUAxx2TwA
jieWNSbJZ9/VTb/mpaZLZoYxcGD31dnyXdzCq2ksljSYi7Z4y1jK+mvNl7XbXMRc8G5LQjUomWjo
ZkVDyczKdgoenE+neKIz+pJYY/TdY9zrwA8F0s7FUIZdsr+l3Zf6vb1xbMus+u81iJBHqlT5L2hZ
5YC9wEHRvH/PVtayzNWG8cGgAMTjDz0FEHU/zMK47jpKJaX4+olz9IV1NCYKqKzSHOSQlEM2rIPl
8CB7XvAe69Udk4p58id1zQt5LwjGeFxaCMSBVGQINE8ViBXr4m7qmEa7tAS0uG3En3Z11JMG2C0l
iwDYs2PmBPRUTemkvh3hWvDCWbpO9n6Epw8r/dNG03WfDgRmuamwf/FooemzmL3UrpVKsImLHEYY
iSaUmsPGM/9gT838lVktZeuuUddtoz8fen/LWFOMub/bRIXtvNJunxUr/1UFRPceVJXCRGpiEYuv
eiVxAs7jCUtvQmQwBod0ErfTN3SgoeZK8T3guC4XotpmwMRkv9uia58/CnrApl2GsdbEJk6qEmc6
21lfb+w+LGyn9uAVZH5IplsSm7ErhszB851CrfpTO1kRlr8SrX9EuBRwGVSr45qcY1cu+W7dreg2
jvrb88pDvt517Jz51mfVYvkSP/mKF/uUnQUVLSl7505KPgFEEySbY2ImkN9odMt6duRKgU+yaSKg
JxlDdagTevS8x2z5f+zYFmOxwqAILQW0g611ANawr5+nwGBRauC+2BTRCwYjGJcMQmnSLiCC8f7W
1uEv+0SbI2WYPSOVJHYuo7c94MrVJSCQ6od1/1fuPZCaUEibmVFKjXyfOFk4mTjb0t629aJyDVPo
ducjq0bHwpDf6BnkW6oVIGsq7fDW5zzPD3xdwyVB0UTYlj5c+0UbQRgXkqlmge0sUrF9NVtQI7Fj
mLbMcvS7EpBlHnSNW+vtofjCHQ5EGac+nEsOupYq9xG2hUm2SlgqMiOlGA7jLk2ccpExZ6rRTGCJ
hdmT7HAvnXMYoGy2YdgQSkrc39XmMZubZWmrGeMeEQNKPWTrq4E2hZ21BwjsPZIvELpldf7OvEa0
SVmRri/bDfHo46NGfbbnRIoUjEqDSmAviIFddaPT7g8rJp6xjS8kAKqbLeqlmjWWwgIrKLZop19v
hExxLrS6Zk4TtgzyFXK62ZmF+ri+f3uJrIqzgugBeSr0AD3bxCLSz0pd/78V04YEy2ZU8rmEgRTw
m8n/ATt4sCr+MjfRBh4RdliGAC4QlBRHYq0aU1inVkLUht1ktbb4/ig+eji6OiUFbb31AzhEOVzz
2jQA6gGxyQGNwq6QPeqTIOfGd8gCSeXO0fk9ISVl11ImTgiy1mpgbyEdO+0cmiVZiIGIUig/59tX
27JOK0GQRM1/cDzGW7wEGqlxzgWcx5HJ26RmAul3tHQmM3KpAeUPZ44ie23cGgJmAz2uT0VdVdoA
UuM2eENGVhdtpHK+KF1QBB+9sPJiegAq8eqC4CjlTUg2fGQZp22kXlw4ZHXkZSVGT/axW2hlzMAS
0PmnraQvpCE0D8Oz/LGFYjfXiEGCTbW8fd2ORr9TeRmRsTSQ0Q544r0ElXSTJ2bbvm+n3ZREGSvX
w00+JVGZPdkqE0RGKB2SAZYfHRJM9sxohCkYkQ3wTOUhVU7LFJ66d81mM/5ZCfPdHX75WTpKWhXX
HLgWgqierb3N1Mequq6FZqxfRU9KDicK5ISnHNMTx33wAuR9rGWaGQsMebFzfhKsU0yhvLmk+9MU
MMRXcABtc+grWprvcQMm6zZGLTboN3bv+TZpoAp7Ahs79tSaTNaJZuqA0EXOc1LIHf8JF4Ld+boh
bh3t2ONdbkO5YKDOlMkejzVFoxLFTztMsKiZhgY49fSKEG1GE7qPCf1tlj7/hXc4wHvsPhIuDdz+
SWimH8yYI5y4Hlgxr+K+FjKfK2jzUpDkVHR9OIC9t9nASruv11IjGZdacE2QObP5RdHu/V0OYOy7
RelhWg7v4aCzzMZX78YD+Kb809fE8KBT+zeCqjnhOxf3+gWSZ+mo3UQHGTcd0fF7ZzRYZDlDETBK
fGawaN4DTN7Z9HyVYqCE7oDstgHsOtlvi/j26yLTH0QdSjztNr6k9CIxpuS/MNhLGDAcrgAlb6PP
4Oo4RHmzkHHsy+KgUiaQAvaHN8lqPWQxqt4agh3Md6xKn8p/3MKKUt2zPKteQh5zNuDA1AZzR7+X
yR0zZqC6dgBFkcLpq6gnNHVogJ6Wy4DWb4ekK9/ruacGGLLEdLtK2IY7o5KidKzRFBUumAzKH0Z8
ovxQGQbGm6FZgRTPJQrbQDgsaPOFVWZo8xhEmrjEJ9NjFAAZqnyG4BkzMfN8EKyOwkFt1Q6bSzks
Xp6iFYs8fdpWl7zWS5fxmILHPcX9nYIXmokzLLv3QBR9ASYxz71uhFfAi1Gbq5eHrwPHK4reDud+
Ntl25iPgHTQIg1PFgZDURQ==
`protect end_protected
