XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����n���'�CC}���c������Z~O�vsW��M�K�Ôx�6Zt������i��QٸL�'͓B�P�L��:L�*{��MN��_��pB�"�EQ�<o-�<���k%�����ܿ������&<�����{H�~�l��� ���U�'�q�w?�ݫ����#N�0�,�Yx%������"z8(%�|�6	���ҐW����|�1���j�����&��]���L%q�.�L��/
P��ѽ��tpDKm�����,_n�A�GAQ�؀C�|-�����>I��?*��[����r��{ ��%���ID���@ MZ�w�N���<�g�Ƃ�6�T��H��Tن������;B�0����#ϕr�؇���E��f�VyK0B�Z7�~Mm�
	�m��*���:�ͅ�n��}��4�w��C��z[y>A���J�n�$��7#%����547��{|s&n�����ʻ��x����Lxg<�(W��u��u�zC(kt�H�r"��a]��R�/��ή���܇�r|^���N�&�z���%��vu�������iLN�+P,WW<!�I�<��AE�����_{��ۯDJ8����U�#�Qkؼ|@3Vן&�;"w�~�E%Ln���VΧ}.膈�~��ZI��(Z/�'�*���`as���)�ޥ
�H�/O�B���HM���e��ʔ)�{l��g��MN��}�a#@5���iw5Qٮ�>:b��|�P%� �dԀ+Ӯ�XlxVHYEB     400     1e0�`�4N8�تY�k��<�(;3v쓗���\��]�.:�F"	S�HX���>Ej�$v��������
�f����KHS�1��_j{ ������&瘳�{�kn����w֕��L�ξ�4�����]Ǩ��G���R}D�5U;{K)���v�Y}�ca�)�z��ҧ*D}`��C�X�;�9t�綣�=��9���p����x��5���?�?�=t��mhnb˨�T�
~�����v�k�4�j�`L ҍ~�\� �K�v��u]�PO�J���n�������C]���ev**޷�֑]�t~��R��������8x�����l�$�ݼ%�0�KI��I�q|G�8�{�����ռr q�rR�N��}��C�(8�ZW��d�"#�d����K�VҞ�����!p��Y����D�zNBe�q�z�;��:%��}��;�6�� �탪D �p\��XlxVHYEB     400     160aAGpU����b�1�����z���b�@���^�zBj��'���x�N�x|��2g�m����T2���^m1����H)��?|:�nK��W�+F�eYx�|�p��#_df�l�V{���-���a�l�\�t� <js%m����[���Xo��V�?/2*��N���M�Mt��1i������v�wF�\b��1�wa�	�C%����1�RTL��A���U���|��|H)
��Y2bÃn8x�=��K�6�$��O[�_��6�B�����9Q&�?S��;����h������B��U� M�59�w���~3Q"]��w ri �����[�����Y�\��ܔXlxVHYEB      50      50H�1_Ǽq�BI�
�ļ'ɂ{~���#c�|Z��Yl����r�w�w��B(�Yvz���k@�����T���