��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���ɋ�q����DI�"܃ �&�"�r��qO���e�%P�j<��g]6k*�x�H�.��`jd�ƆP�6}��*���]�"�Tq�L�A�5�G�"��R�5��`��p]�/���}!:����ȥ`�"9%&�����1]��RZ�ɔ7T~>�;(�M[ �	��f�.BB�$�cz������@OP�^?�.~�ЧAF4W�"�q��Fy%���[.��C¹�)���F�wC��,�Z\�0�a5�]8��Μ�V:/a<l����	��`�i�,�h�6�nJ�Zv�:Ӵ����ꂜ��oe�����s�}>��3Fn�ސ��YO���>�W�L�8��!�/��jX�"��4�S`R�dËML�!�w����NK%��Gn3���-�Ah�%��o��b���m�3�Z�H���4Z>Du���V-�D/o����\o��D]1��\n0�"c«fs�
ͬ��%T��뿸I��F�O�ӄ$��?�^�,=Y&pB��}�=Q���*d�}^0b�/�[�
&%�;���&�P|0i�o����V'�^��@�
�	��dG;ǉ.�;��U#/^`'�tv�5i�Y��=����4�}�*-��?J���SU��^���$q�<V!DH؅�p[����:��!i��"����N�P�9�f���|�i�Εr&�P�&��͙�K0A�� ��@W_m8��x��'�_xa��A�ŧ���$o�+�6��+K]�q]C���s�I���$5Ed�r�)��Z���7�j�F)��w��ی��#�A]�x��L��l���7���r=v���*����n.����g_�g� �Gl��A�D7��7��`��]$�Jr�ש�z�@*����:\9��P	��L������.%��i���֯�xc.?���J�"W�����I%
c��R�L���PH�?�lU<�ZU"�Yي֯�Y��z)p7�&cj�UͲǗ�Ɛa� �4�,b_����8_�+L"EJ���0TT5�;CS�Լl*�d}[���,�1O+6J� ���	vq&B贉p��M� ��0����h.�k|�K	�T�"�Ph�Gmܔ3)�x�+F|P�C���+ϳ�+��hq�&���d�w�)i��V��T5��Tz�V���8�;D�'��Ii�N�s�$+}�`|��n�)�X�{��h��q����RR	V���$�2#I��`��f��h���[�D�3���۲�kQ]�-%�w���(����6B��JFx��)��ag��d�"��<�NE��ש���ND�tl�N��Ľ@t"��a�`Z(�d���d[�����z��+:�i�����E>�>�A�c_,a�!����?:�ќ��(2ʪ�~׻*'��B�!dQBP�N����
��I�<���[�C�����tӔ���E��ֱ_�[J���τ;��r���ce�MQ/fO�뢳ʎK����Ϧ2���.�R���e�k�Ԧ��D(zS�]�m����E??�������g�����P؞�v-��@|�Ѐ��r4��sB�d���b��J�f.� I��҃�}R���y�=��\��<�qE��o�Gí��1�"�q�\�+�c��ޑr��[�o�j��`a�j�s��Y ۥ\�,U���$L���*���x��YT����`S��y��{p�Z�ו7#�v�5>J����&����B����h�z �d1�d~{���.��5:qk�ݹ8[�/�U����y���-��0�֙���2l�r����?�Ж����#�G8Ѣ_�@��S_6���m���l]`���+�s�uPJg�*����0z�)i*�^w ��Plw�\�*{��9/��ۺ{�"xkv�������u���=EO���C�	+�t�Tq�E���6���9Y�n�A����=���1��Rv���B.���b,��l�Ĳu4��zV���[�oDx0d_Eg�WT
�_�0B]����q~炝����Y�tÚ;/�.��8�M��-���Y�`����|)"��5�IFŀN�ݑh�U�NK�MtHk12)cV ͦn�Ґ�5lDL]�oB� ��#��q�iB�;��.�����o4o�_&��L��
��˙}��	���L*(~S�3�Q��Q<��aLubS�����#o|�b����D��ζv4�4	��J���D������a�6��U''�.R/7�+����`�6S&����79�{kUp�� z�q�9B�inl��[Qi�pw�XM���>���� ���و��{�8��7��es6��]2��Q��~4�ЋI�q�{fa�x�S22�<�Du��ޡ�Gp�G�E���@"�,�Ʀ@�f��Q/�/s	k%��D5ga��h�n���~M��[2��ȧxs��0�J�e��-z�AreCB,�I��}<m�k2�;�|0�ȓ�u� �i0�%nt2�G9PxB9 �j�W�rQ����� @�8H6���>A�N�}�9�=��1%E���?5jK*�kK��ȑ.�%��\��ER��A���/���������=����~�HT�q5e�f��B���ԣ�=n=��xS�w7J���w�#����ے�9I�8�y�U��e��WRk�ݿ��%e�`��7��5v����8�䂣�J&�O��w&4C�=4:��lƭ� �l�Q��XS��FG@[�x�3�k���A��\Z^�-�o�Ɓ�Um|���E��V�!�i���k�$��e�q�p��m���A|i��Ḗ�ٴ`�\�Źx�^��,2ҵU�k�A�J+��\��ˀs^���]��6���#:��OBʳ�E�5����[�!UC�ˏ���{�LO���?�/TV2�ٸϫLx�� ��8��	7�Q	ql�[��VrڝCvP�,���w�1���D^�;R!���Gq=�jV���g�.�0��Z��ˁY�
5(��R�3pj�X$��DJ������P��T�x�{��R���>w�+T�WR�8�y�@D��)kQ֬w���`�-������P�[4v31��o-��:��JZx[�]������4�I�]-S}�.�]�yl�2��-W��@�wi�h�FC������z��nB�Xv@g�`Y}�hC�.����ƶ鑍>X�x��_b��iC
3��gݪ!ػ�ԥD���	�6�Dv��JqM���f�t����(_��Ի�Q#-�5@o7�J�����l�X�|�<t#�w�H�9��O�&Qt����|�j#WL��(ni��e����pKo�IĆ�4Qb��7:$���n��V;��1W����co�f~Z:�o2�6R>�n,'CD�W�i�Da&�z[������ �a��x�@C4����mWU�y�ϓ˼�ܗy_5��ה,�
v�p���ǑH�/�<v�:6�ȩ�����[�"��=�f�@[?�_�*K��-Ґ��/J���-7	��4�"�	���W;`�8.��s��]�=kKF1�I�5{�T�*����ZTF33�哫��h{�U;��9M�:� �W)D�Z�E�}�6��yJ�`	bܮ���ϴ�!�j��{#B����{Y�&e����g���^,%IB@����u�;�AghN�+����jp��������J�*��NW�ed����GU����3�r��Hu� �a�m����m_H	�`����0��q�����m'�/#U��Ѝ��B)Ob�	(�D��j�U��ʕ�� ������(��!V�*�*��Me��H�R������Ey��#1O>K�Ǳ���w�Ç<�߽Z��N���i�@H!��f�<S���pw��!���H����Z��j^ӓ�S�H�Su�;2�W�&�/�VH-�n��� pF�=��b�0�o g�9�^ S�4ؘ�X��dC︴����)�[�.p�e�03LIY��Ű��h�Fo�(cB�oE~�m�C�#&�f�(��^H�w����f�u:,D��R�6��h Ž�A�/�LX ��( 8���m���g �ČF6����A���7a$�soI}�8	ɨ9m��J�	�iʐ
�����7et���6ד�Q��߇��J;\��0�	Gs+��z��D:$ ��,�֐^�t'���A�ƒ��{G���X�,A˛���0���rN�Ċ%^_��\����p_���%SS��b�"e��5>�_F�u�#r6�lE���qL�םL�����9lx���� ����� `�=UV�w�k��c�^Yـ�-���������z��CͦZ ����C��K��_	�~��/ �����~>�⋫HK3n�M�ؑ{�-d����sh}e�`f���XJ����z4Q���]#��]~����Úk�V�M���tz�����[�K.�3=�>T�@N�K�9��vYD9	�&[<��k��ŗ��R&��U���,M>���Y�VT{�%g�ߤm��åuHO��vј�jbݢ�E�y�h�M4��J/s�	�L\W����ǣ��Эуr�+�ɹǿ�ʩ�G�f=�:�`�&�kʔw~�l��6T�1r���=R���ѵ�Z_7�ȕ8z��9��p����ȇ��O� ]��ѣ��O9}0�b`F�Wo���M�O��WYlމO-�dQw����F�������&:�:�l�f?�Z?T̏&=A& �����i,�/D�k�n������7�y�$���JJ)nHDxC�d�ʍ��A���5P�9i��Ob	� �ӽy�?��h�[Ʋfߦ6�Y��6qA�.,]J$V:6aoYv�z"���t��Ȉ�
_p�׋����s
���R�a��g��[xN�t:
�0��� ����0��\$���_u������e�!"=s�əI|�N��j�ӹ,��b�ˡ�ͻ��>���lg��4�i��g^CQl?!�-�Q��,��}�7<�i�����p�:6'��!zHE2��[�#�V���,����@�������F��o��λ�Ѵ�C:���f�f��U��Ė(�pAv�ֽB/���=�dmX�#i�.��	������%���%�ð��3��Հ�&5��9�S��`��v�J��}���+X���a$zb�����Z�0��Y 4�D�q��W(�<00� �Y��
^w����I��J2r��IZ@�%p��Zt�#u$^
H�8�`���s'd(���N_��������%d� r+@�Ms�����V��ف(�Z�?�Ar��"�qkO�e,�ML�7uF���E����'��z��H}%���{^�:�1�p@�[�z����
d���Gnw���<�&/��<{6е�Wx:`]��~�<u<�Lvsΰy҄ J�~��񺦵���mxl���A�R&Slb1tVU��]q#�Ad��*z���������>��U��)��I�.sEE�s���.E$&�>����wH�x�%6�j>�W٥�P�=WWH�?�Ak�C|�s$�Ԡy� ���\~���Z�,��ڢz��;�.�@�e�|�H�ԛ	}dӳK�����[N)K�}��6F�hw�KPfX����¸D�5Q�E��qQM2\b�v�w�2u|n�,�C��ng��I���cZ�V�S�3W&�!ϊ]�!�u�l���A�o`>�2�F-o���2+��gcS�:��H���9"`�r��/�`ەҽ��~5O��lG
9h�}���q®'��*}C�9W��f� �9��}��6�5<����9�pT#+r, j����z)hL"^��Eݼ׮���n�g��
,  �.��v��w5�cM_��n�E�o�U:��fƣ�G�a�"�t��3AX�i�y���ru����{����8$�k7v�2q�D����a�s�c%�mN��â�''��;�QP�=���N��]�rck&����nk�����!���W�Z9x�����?-��>4k�����o\Է���' ��ϢUQ(@RPK�����LnO�x��	i@�G��Q:����M�3�O��%c�<����Ez��HS��ΫS����m�z*���Ld�$TB�C�&�Ҧ-�ke�������MH�EZ����!b���j����@�n7HT��'�������\df�ĕ9q��yc���:\� ���r�&h��ܓ�"A���_4����o��P[=�E���6�>	��e������ n���[�h�������J[
�QG�i�~AR��ӴT����S�C��]�gvRdr_�17|�����e�]ѽ�%JAb�M
�M�T�z�Bn1:���� Z���(�V�_�2�T1oW2���9����M���<`���%x����ܡ��|��Q �6LmN�8�4�tc�wQEz�2��@8��y`���t�mTh��Z������_�/�RO��2-g�������h�oԫ�`�z����4�x���Q6
x��j������b��FD����3[��Y��$LfR��s��,[[�uiF}�6���lmo���͒Z���I�Wa�x���k�����'�ɺ8�,#�.!s�� �fnΪ^ѐ@5�6L��w;�XS.�=\�K1��ׇ-
�tj闛�>�	�Ң���5?�:yW��ut��G]�Gʨ�?v��a��f`-�U��@�
(@�$�LL���@C� 0�Pd�ӷ�]�E�U1��Z,��	�P�o���EE�G0�ʷ}����O���8�^��ٿT�T��kϒ䮺����g@�2	х��EcX���'��ƨ`�P�9�9�T�L���jVxm��xjy�	�d�Ɉ^���$�+�y�:	���\QԂ� $@.�綧g|�{{V��xi�]]��7+ čt�oޮ�t@"%��F�R:��k����j;ۗ��������h�;H;G�s���ۢ+���1��%wʾ5mm�?�Hy�@EJ�Mʇ fHBB��$�@�����i28�Xw3q��ة�N�����.�و�lb�4O��X	����y�i-'�'X>�\c�B@�-���.��TǕArb���c�]�U��ꚺ� ;S��������Ha!U_�P�T�G����;�H����jf�zZՉ����,A��{*���AlZ�v����ˉ��n�l�k ���-��{"�M�v�����Ջ�a�uC#�?��_A��@�/�>Su�ZPi�,��l��&�9��s~d{���<Q��Q��p<�27�+e����\�{�&ʦ��g�D�a�� ���)U��q��ń�w�xۆ�BY�3�T� ���M�	E)=��f5w���mKC�{�4����aF}�9s���a�ú̍h�p;� 6)�-H�XJ`˅�]5o���ޅ��n�"s�&�$ay��0�ވ;No}�V��@KH̺�3fZ��r<�/6�c0�w�Y��8�W����S,w?T���7��q��!�;Y���G]�ʍ�Љ�T�`|>q����]��P�4�phl��	6;�D�$�ClWWI�I��@F�IE�@�O�ZW�ȡ��ΰ��E��Iλ�P@��b�N�M������u]l����[z��:�)]$f�{��&�~�'I���M�I�����vz�����d�i�I9<��ɨdD��5��Tpn���_^���/�s��^����3W��t.�k$��!�6y�����k��i�U�t�,=$����À  �m� =�x�����g �������>0��+l��$�Yh�b����J�$���S�f`��ҪS��8�p^����.�(�[05�im�\�QJh�͢x/�����]�sx&�C50�-G��i��5m����C%�*��.�v���T�I~j��r����)�/"(����m����t�1lOdM�Um�6l�g9Lą�?-6B7hh��zJ�3M��f&s�b�@��G�� ��izңI�Q�z�����7J_S�v���7���]��6&�
��%�E`x(zG�w-�3���)Mv���A�����c�(��Jʐ,@�s�A!��Opˎw��߀�)<�{ �y��L�P��U���Ɩ��|�d��9�ϿZ#�NR����H�x���mm���E쇗j�9�A��
9 I�CC/bpz�h#�����D��U�=ĭgUZ10�E��VJGv��FV!3��S��Wv1�}�,?�ub���3��RB��$�w{+o�D��9G(��ܶh�c�$�%����ER�U(\�I:���j�Y��mPM�bNs��'>�`��h��˭ɉ�HKŐw ��c_*�E�!ݏ�~��^�P:VN�wLnT|8��8!OW1]6>�B�@|�<���p�Q�I�^�C����T�i^�=/����Pw0���:��T
�B '����cF����������Z(�}i=�y�mЈ}��ڭ�m�ؙ�:A�����:��FS��:
��Nd��*X�$*�i�XO���z�B'����)�
P�c�MF�7P��(Bp�헪�U?p߫��ib��MZ2�5H;��Q�If�L>�[��ch�گ�-wu��+���*�Ȅ�5C������N]	��g@6�!1�!հ-Z/R^��^�a�yp��_�-j��cs�>*��{~)kk��hK��8�E�?��_�!~G}T_�`�DB1ؤ	X�Oi� {�� �?֪��p�C���*8��-�%t�CM��G,�������a�d���CLܗ�1��-�W}�T��%omq��t�p�Y����ls\� �����S;ɮ1�����Ќ����k_�f�'�̈́����������i��k�ȁ�_�d<&W�6�vj3Â�)R3� �2M���J��5��=͖��cy���#12\�O�ܜ��z2�F�v�Iu|�k�K$]�X�ujn���E��-`����]��tz_֫�E��w���x�5|k�х��k,)w#�w��R2���e�h�$��p*�����d�+�11/�o�91@C�$�rG�'�ڨn m=��r.��d�}Y�!�x~���ت�/��InJ���6��H��L�R	��7s��	�q���G�&@*���|S],+k-�"�a������,0t�R�V�?_K{�j�>%xd?���d~���+ܜz&6!�߈�a��^�ݔs��tJkG��M+hp�͖Q�}*��Yr�\!� ?���amУ(^o~�O������'[@Kz>�N��H��DZ��E�%�3���(!A�9�ۨ��W����sN5�����ǉ^c4)����Sm�����m����R�M���V�6�ة�U$߉�*T�����"�$7q�r2[���ɖ�K������g�;u�S��H�sy7���F���r�AKrF�����N�B(K&m��Ժ{:cf`�QA=e� JJ}�d ���p�މ>�nʃc-�h���v���2`&H.��n�J[kE�h�ŋ��@JS��&�x\x�I��#{�_�j-Ū���@3"%�z&A��^��,} �>謵��ْ��3B&�]'�iYh)�r���p�E��yVw�w�T�tٌ��H��[�ES^�����nC�%�j����a�<&�'���������ג��&�5�S'$��L��p����E��j������k���,O�7�+Fb�,ŝ�����Ք���~��]A��N�*��="3�|
;��8����؞�jӛ�y��V���0-���*��)�y�}.=;�_�6S*�!���A%jV�c )���ۃ��d���ey2F�\�G�3]�ljVKR��V��B"�#�}�S��fC抛)��I�e�'\> ��Ot��F����]���{�2�@��X��XN>ߞNm3������"��6�Ԍ�5�κ�
>m2�$eͶ21j����Bvs���v1�����f�-WR�9ٶ.�9�*X��'`6��6��A/s�4�!M!��[a
�����[�˩���Z�����U�w:���tY�ً�SL������w(�*+��.�L��ݧ;3/A�����Q�6���:��e�����0���n~(3��$Фq�n�ڤ���.� ���;�_�HW�cP�j���7��;�����e�T$&�i�tz�e���S�%x!��u�4���SZg�R�2��K���4F�݃P�{C�+F��t��(� 
�lW�@�;�����i��ᰉi�nz��R�ܻ7I�������P[�&hwp���#%c|�qf{��]�fߡޏ7
�1]�������+i���@T�z�g��gG�M�^�����0͡�7�I�b��㚶�5-j��e�������?S�O�7\�dĉ9�@g��<S�lU�n�c�H�eۈ�3k���h�jSr�w�>3H�(U�]�JN��㊵�T0'�;��O�B���L�;�_��=>��t�� tӳ�=Ƶw\�8���Li��E�{��by�᪕Ѳiy�d�y{5�AlAunbp<I~&��c���T��S�$�)��7i�ë̊p;��?�E���~g�*Q)L��v�6Z���8�*dK��KԔ�1� BGDh��*�Id���ߎ�H�L&� ��(na΍���`9��e~4�SÿDTUw�j4�+�J���B�2z��f�L�y�`���̡j��7����wA�j�U�]��;�;վ~ڞ/����S��>��(����y#x�]������3s�9�xɹ�I�,��`�Ƌ���K�?*��ǥ���1x&�R�ڛ4��h�#̙ʦڛ��T��	-!��@W_#��q,ė� ͷS�Dѵ_b7�$�2�ձ�6���&0�h�1�]����T�۹�2�_`��|a"f��v'��_)�#���C���m�3G��,�yw��6����'u�[���2
Um����9g#�浺�+��%�m��9��d��ƥs�I܈�!���1(az��ٱ%~���@�^F����}RV�~��0�/Eԋ�\��P�d`��Oϫ��_ڟ�Y�F7�'_Y�im��W��Ļ���M���<���7ʑu��M��-!�8N��2��h��T����g�'Dn2��%^K_������Af�k��:M:���Ά�R� �Ȕ�T�兆B���x2�"�!h0�?���I�#�&������K��Ӫ[|S�Bʸ�8�����`O�5�P��%{��&aG�w��H)|;
.�^�{�ka�2���ʬb8�椔�P�,�I2�(00~� �p��3�i�u�M��Q�f�6|`�	�%lT�J�ްh7���Fފ� QUE��0I:QlB�m���H]�'H�uʵ����:���[�nH
2���O2k.����ǎ�p=�|רj�a���ZԘR"c�ӐR�-������#x�7`�X~��ұX%�w�9$2F�2\�9�!R����:�_�[H>-	ҧ�Z�߹�ϭ�gs�Ր��rn*��~��pF>&�Uǚ�Dh=�C敊�����S�2ݯp��cڗ!�h�.���1�I��>�3�"����.��N�Ri��LvY�+v^���2J#D*�Lr]�C�y� N����($#���:��9��;c�����	��[jʤ��0p�w��3$p2�ᔏ��������1��t/�xBE��\���	"�$�C���ހ���N��I��-+�FXx�3Y����x������������_V���L�Ј���acYܑTb΅9��cI��-��p��6�U�/���Dm5|��+���2F���s(S��^�ґ��(\QܶT䇝!�TWz�%yZ��l!ň���m����ͻE���$��OsT�HlA�/M/Э�j��n�TU�n
�FJH愝�Od��䖈:�I�d�`F ]9>�	�=��Z�d�	���op%�ލ�+�de|���[i҃������b��QL�6�[=���Hi/����o��}��Ѱ&�k{�c�kx���[�{���D����g�͍���	��$]�\����Q�~�A}��!�Bԉ9����y�lX�O��z��6Ӟ���b�;+T��ȓ��5�d�(�7�Gżg����<I�Re���W�)��h.��>L*�$����|���)XngxV�j���W �ݜ�hl��{N�ρ���L6����������='�bU���	AJ��l`"��y>;4呟rsP�6C)�ݎ�C��s���6��m��x|��)����e3L��t̚5�׫��BD���ay𶟗?���Z�sp�KˮK�nLe@��D�	+ct���Mi\*�Ǧ�����i��K٨��$w��&_I{�"�amoB%(�GM	�_/ev�n��j�A�<ҬJ��<�3�} j"��|I�
�F��P$��Jy[B����;p�_BGz�9���Q������N�6���%׬�$��f�H>/x;dt��{Ki#P+Gw�����n��	%����	\ '4�Y��D�'���ING�29Jf'��x�w��)$�)�T$.�yC	G��eb_��=r�q�i�������w"��O�CݩP�<��9"�\@� 5���<e��8�?�e,��e{p��Л��BGq�e�]O]ߦ�_0�"��O?>.��?�����$B�k�M#���*x;��ŘOV�-W�k��ʰ(�~�M�Xݡ���s/�רXؕ���>CTJ����SI.�I� W��`��Hh�x��Nf^<'�1��BX����q7��Z�����8�؃n�w2��C�C~S� 3 %g����	�:J	X~��r����5�;��cGJ��;י�"���4A޺�e�&�&CD}���ggz.@-#� �f\W���ڎFk[�_0| �t ��&^xל��2!��ڛ{m�&"��
��^�R�]?� �9F��g�؜T�t��*��>S{J_.|Hc	dc�H�#�CU��9��raV�sl<f�'����pQ��8j�k��s]��-]K8J�7����*��%��C�V�'�-��]|��p�Ɍ�h_��aU�wҗ��fD�pq��T#Y-T]�ק�����~���>r�'N3���
�ĮU�p{���7Yq�Q���4�W��$����j�/�)s����Y�(G��=_�8�JMj��GM���:TXX1�o�'����S:,� �m�� �Z����,S��M���{�π�_�
a��yh��R���e�li�?�t��gˢɿ^4v�Չ9�]L0�>ϧ'��T=�Q_?������0=;�sï�鳔W� ѷ�����{Z��A����޼�t�����O����+���Ao5������'�)ع�0/}���B�D���/�@�P�<ٳj��!4jk��,.�+�&�����h��T�\�b���Vn'��A��0�nu�C��E��`�����T�T�x�>��n_@��u��o_���LJ�ʇ/�q���Q��ֺ To�q���G�ן�R��Q!��9S���n.�=T�m6g�Hì+�Z[�2����3��+��G�\
�2��C罩�G��ra�9�掤�O��R�R:J���?9�����S�cQY]�����0�B��N1����1�7oe"l�c���H��%�7��zC���dNPYA��@�D�s:�D�u���f�3a�!���=�������3#uI�\��w$t⣮~��ߔ� 0a�IDs���0;AH��=U�J/�9��Ԯ������=���7VB]�fn�^�A��Xq���:J�%��VY����XA�N