XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����AG�6mRƠ��y����"%�U���'��p/�!G8Ǖ�a�'�-ƒ�֚�Y��Ɯx��� �s4��U9���\��K�rÂ�G2K.�h����!��$i�Y$�eN}M��b�H�?R��Ya��'�����Ee��䮓��ϙ�]���;��^���>�^F�X��r>L޸��L'�y��U2Wnu/u�����ِ˺�	bn{ҹ�8I��d����r6�,�pUۯ�z���O���7�`��Eئ��d��Fg��yc���}cb�]����Z*d	���&�U�#��&���m��>u|����/ҲIL�x'3��0�����0]4�$��ҍ��=�!�M�a�{Χ�=
��S�-|�B>�s��Ce��Y�(u2�\�Lm%���eP���jPPl��m�w�=��5�Al�P����,%�`a��8���`?h#'�i�Zq�0:ѐ���h �`�r$�r'����ւmba���<���!�C�Qe;d �3vR���|���BEv>�)un�=�̼j�t-Y�8S=��c4^%�b��Hiڽ�l-����V\�UG����~|��~75�հ���Oa�c �JԖgyL�2_n�����뎢�{$\<�؍ٷf�~��[E
ի����*,�$��JW6�>u0�`���׉<7` �\��>�i��f[-;0���K���N py��2�6p�B��G2���s�uV�(�՛��>x�7Q6��F|8�M>ҁO�&k:� =���ՆZ�	��XlxVHYEB     400     190�,3��Jj��Wc�7 �fO����ּ]Cs�3���{�p�
�L��䴺[�}aJ�с-<����?�K\�����A�ʌ��*+%�Yzр'����8 L�d;����X��?D���i绎�Ϸ�D̓	��_7w�s{��q�<����dz�zJ�I�o�ѻSĕ�sA�-t�� 2���~����Q��7�RHQ\O<�W�����H��"<t�
1)e`�����yFޝ��!�<��<,�&r��Ē
�T���^J��T{d<����A�v�mdz��b��F�]�^h���w�^ � �������5n�Vm�,j�jI�X��h2�u�Ԩ���Z.벛0��/�FɃhC�)t.0=�g��lO�˥�$�9�b�-��O����F�@&XlxVHYEB     400     180s8�^��2�%{�-t�*n�'�����y�9��G;��=�VF�,og�����A��O��d��@[�h�/���-�-����[/
�%��18#3�%*���G�oU��B��Nq�f�(��D�}'�ݳK��z��r��t�k]c�c�p�P���gX�2��s����E%�~�n�a����H��{�An[5��bM��*�+���F���}~�����aO��$��!(}�H��8�ls��c�m�]�Ri"�sQ��A��q�؝6���SQ�\�ԌP���r� \������2�L���*�#F�ڇ�&P���p, �p/D޺����c�4s�O�v�����Dy�$�b���R�/Ib9f龉�_��Q��VXlxVHYEB     400      b0� ��@bRI��+�a�����О0��	��E�"7B�bs-�D߮������8���̳]$2G�����HH3J�ĎEd8T����'bh�[ �1����rdbvߓ ̌���[�r�d������K�WbA�r��;D(_/���e{�6�OΏ2𧄚�%>����'XlxVHYEB     400     170r:4�c�0RK4Pn{�l��P��k~ckb�Ү���pg����S������u�CG����U���+ă�T�R%�q���|ku�����P �8{��� V��/C�~Z�[م�bsr�S�����f#��J�S��Lc���+�Ap�4�`m�7^.~R��Y�e��}O���
�^_g���s�X]�����&c�y�l�a[j`ZI'襺[-���:}Hy�����9��ۅ�>ct�/+��՛q���Ӿ��"̆�ׇ��Vv�zӼ�T��t������ev�OB�6������AL�����!7	���bs����ߖ�M�W�=��t3��J��G�k�I)oPŪ_H:Z0�4�}�QYXlxVHYEB     400      90�*�X�x����q� s�6���M��vyg?�"��#e@��R�~V0��3$ݟ���zF���X��ԛE���?e���F�c�b�N�o%[9k��
U����]7*�J}F�@Y�"��\�A�����*�a�lXlxVHYEB     400      90�[L"M<\��U��3��ͨ.3_������A\?��Q����O�bź�r�������1D*�:����R	�����$��XJ���� �����
�UuL��
���w��"�]xQ�B�Z�Aܶ�AgM�}A��^HZXlxVHYEB     400      90�n��%>��G��y�ϋ:�T<�r���Om%?F��[��J�����?�Q����	�5�1���PT>JP��G:�i;�U��M��1g��XGj��fw������Nu�O��7>F�{��պ�Z�3�5�|4��Nq�5K�AXlxVHYEB     11d      50�?G�nɔ�M���4�F|�������Kԇ���<Z$H�����Q[�f��R��:5�vW��Ǹ�s�/���?8�'BՁ�a