XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���LpU�d�7��,X_��^D�ۭ��tUlŔ�"�p�ޙV����[䟗u���w��^�����Ȣ�U�*�Gh~�&�=�t�@�i��c#���*42ps	� �\٩�����R����-�SUh _B"]�M{�ol����(�����CYI�#7}�8�"�i$�X&Wq� *$������+�}�JwȜ�{���vǁ�E��(>Xe([���h���܁#[\ʄʾ�1���P�s�7�����x�3�k�/N '6/��vZK�Pk�W��y7ڹs~�-9A6���U��/}�p5�c���e� XN �X�sO���V]}��'&�n%���ޡ@��a:�7����4>N��$-��t=������`���ڟ�S�f�+�MG�Uh_?3fW7qJ�lYk�Ɉ�kC�2]>�Y��PjLnkL������dR���)����{9���ZXk"	~�%|��.�mvm�p���ϟ�3�蕡��nՕ�Mu
CĲ��
��ͬ;잹#K�=���<���N��N�,cT)��<�Ò�xkz���^�+��ۣ4ꖠµP��Q*���^74�#��V�8`!����,h�WL[����S���u��d��k��d�dPN��ALU�f�e-F�$�e�@�2<�]������_�fQs?�	�ݷ��Ð�jew'8=��&[�[X#qr�l/I���Dm�%m����&�Ӄ�g��O53;'�m��a�qո��� _*��f�`�ݴ����&�аL����XlxVHYEB     400     1c0@X~��3��$M#��a\��t[)���sw������DIrT͜ek�2�̆��VR:����^����l����Q���i�ęi���I���o
�Pq�+�b ���o��,﫨I��4��>���0bX�mz�(��)�����1/��օF.�� /���рX�kۥ���ۈLS��\A���pa��Rawg�]Bu�	y�e�)Fzo:d��m�s~�V�5��z��̦�g3']�'�㈕��C=tB�P���Mr��Iĳ�V�++6�3yʉE$I�=��n�F8i�웨�*)۷
d���t��?r����p�k�R���w8��np �q�`�4�#���X�R�h�+�w�b7�(X�N�R����MB��zh�\��l I ��f��� ��
#�H�ӒWDC������Y���t��е�7������l9����e4��XlxVHYEB     212      d02��^ψ|:�m��?p �D�n\0P�ϥ��� �	_���_j]S�]���V�C�0��{�FH7ڊ�S~�J����j?���&]mm��^N���3#��vD�b{��3�Oʤ�7�6H��O4��6D{ojyw��w;�DI�|���0���[��Th���!w�V�G��ㇾ�ؕ*g,B�-�5���c���5�G%,�55/��_����