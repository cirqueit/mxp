XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\��yv�(�qi��A���ú3k�8��@�L��{�N��\�7��W�k�BR�1	����s�D�U� !A�i2�O$�c���N�R8��==&�����G�NXb��e.�uz�	������n�?'���� �'M~/�f�����'�[��޳�đ���Ȳ:y���mb)@��]#-wA���"�I���j3=ogI��p�B�ଳ�������}����V�k2T�{���H�V�6]�,�:m��qH)��U�4z��N�p1R�^l��9�@er�8VZcU����
ھ_���"l8��N%�i�3>h����A�G3~|4!=�ͅ�	dWB����1D-*/U���rjg߈9-������Ǭ��$�h��s�9�.��x�?�`���A�)������Ȭv<зP�q��0dTٞ�E�l3)��5��XIUEs����#��m�\���ʲ�D�MpokD
9�tÀF]`�ၧ�=ݱ&{+�,�?0��m),69�\�ͪ����ҵ�U��e��N+U^�_�Q���&I� n5��4���P�
�K�7�����b���' �.Zjx��+��L{ke���;�f<����XD�+�q���d9�|���^��yUP�Z�]�9L�ʏ�����W��.�����d����Y���}�}�v���㿢<\��t�*��٥FT�H��0�X���҂�0jW'UP�/�ZL�p�z��}�vL�+��M�V���[ٯ�b/���z!�$X�w�����s�o���n��\~XlxVHYEB     400     1c0S���@����j8�]�;7�`F,z�	V-츩�:����CU��-�)>���_x䉙�5a��٬N[�_r� �͢��]N�a)�j̄4fLcN9���ȳZMN&��A���i�-���r!\�U ��j��W4���N˷S�=uޫ���$�zʆ�B�ɯ�w,x�='�Y�b�d�,�}0�f[2|^�E�!��gE̋�y��(_WN�*����Moe����i�YԦ����g�'��U��0Ŭ��x �;�`^ H�$=����B
���m�i��P��?[�&���`׷*�]��:=i%�����[7	�>��ͭy��b��{E��>��8~O��|��5��0����<gBù�5j@������JA�=�ʛe�摅y����=��>�������H#�B����&�Ϛ����Kr�K�E'�x�m:ҙy���XlxVHYEB     400     160�cJ�%S1� `��>β��/��0�[݋���C�{$,��fw�v�6O��� ��Q���,�Yt��3�L@ѧ���UY��3��/d�`��K%� V���B% ����YV���W�N���BS�-�T_j\tӱ�6u��!�oMH��L�_}�3�]��TcZ��gF7{V�n\/�
-NA��L*�!��|�-;�I���I�e�Z[��ZN���g��6,ɖC�-��;�"�x�e>f+ڙ�H@�X�z�B�"�Sb8;18b4����ei���r{�6��e�x��o�C]��	PK�ϐz���$��Z�~}ISV2�^W�@�2�)<"����U���� �MWwRbrrXlxVHYEB     400     160s���b��	��_*R?��8����FM���u���ݓN��A+�c�c��u�?6�4����5� ʁ���C�,�C�����
������6�I
�����t��A2�W��l�z�9��m�� �s�6���v�+xL�	_.^Fn��b`��[�Q�m�"ŷ��i_��������䋆�q�~{i�����䔰D��p�y2�8��SOo��NhQ $x������P�\JAØNV?p�v�IܼB9�$,tLڮnn�RUua�u�,��.�hy����`�8�����9�O�G(y�H�d�r���6�܂�#$������\��
T���fFߝXlxVHYEB     400     100(�8��H��)C� ����ˌ��RY���A�cQ(�k�����_p�*a��5���S4^������:��PyY�!xHO���r�P[9�#!��*$&��".���϶�h�!��m���b����l��ꅺ8�xs���pFߺ�H!�d�ܑ��~C3NV��=��	c��3�n��G�3�B)��x��+&@/%f���'�p�4aZȩ$Mّu���L��f_��5�m�����;[�[,%C:��k�R�N�����fSXlxVHYEB     400     1a0��Tý�!2�m���%��U�J��k v�To�It�v
9�D:�Dw������N*�%2,t�"�d&�������2L�_B�SK��w��bJA&�,JS*���~��^&���"	�Ri��瘳@OA˚��	#��\)׭Ѱ�]I���uT��:y���L�\�2���e2!T!�qꤏ�L4h7��x�'[\_�F�H��w>���x��cn��R?��)cҭ�J�cQ��E���6�&�qU;w�'%d X,3ք�mx*�m�nہa�C��X�)fVp]~�
Χ_�^.�5: C�?����˼	��r�4Kp�(�����jpv�I�vd`@}(��J�ܼ	6g8}]�ۣw���V���,�vA!��rZQ���NGI�|O<�ۄJ4�~�WI�w,��{בֿX\|XlxVHYEB     400     14083[��e����M\��C,��f-%
�igZ ���G?#q��fVZۖ�W����@���[
��D�"��v�4͊��V�,--��@;h�D���\ ����S+�Z*uD��V�Q�V����F�+Y�k��n���b�I"�vX;	8�c����zzkt�lY�xU��(Q�):� ,�g<�xJtqᲰ5�P6�J-] c'���4Y�L`�y"�:m��m�"���`�z4��I{"�m�R�5��gƞ��S&j6=�ؗ��������F�����G|�t�좧('y��H�� �#����MǇ�V���
�_��XlxVHYEB     400     120���1<1LE�Y�۳�t����U9�mP+}�n��<�k��0f��������f�}��ᬾ��F5�+��� �>@y�C<��Ei�[�L)�UD�?/�l��P��9@��F�&E&�䶰��J���%��N�"����Qt@h���l/�l9ǚ���K?:J�M(����+q/�n�o��j_�F�:-�ej��hn����	�1�-��G�1�[��@�!I�9����.$��0T�����uV�����`$�S7"�V��]�Q�����;-��	�E6�XlxVHYEB     400     130;[+w��|D����a�C�ן��K�<��
%�A�$P6�s�w{���ڈ�&Q�&���3��4�DQ=<��aO�}p����a��> �����,����g,
��^�0�3���\S+o��4�qC$����\�2͚��N`-s�豈�<g��B_�A��]�Վфɬ�����q��G�CZ�J^���f\V�ee�K��H1z�j[)���?}	��"v���.��Y[a{�C̝�� ��cO2�=N]��P���{��3����d�8�����j���]t|�XlxVHYEB     400     1c0� vr��ɢ�|�$�+h���T�L�Rm���,�(o

�)^�ӎ�� ��n�5��e�
S�*�����q�L��J9�\�=��k�"'BX�6��^ĺ�p�y-чv���7/�Ú�=tC�5��%Y�-�FH!a��(�f���+�Ӏ��(�Q���Qs ҆�i�l.�|o����j�#���_ī>&/��;$�3/��C�ZL�j�B��-�%��O��8?�>�e]\� ��e�2+�a�/J�o�]�KS��(+�$�o��O'$B�|��d�O�O�({gX�RlL��3�F�|�ё�^I�'��_��z�|0�8��$��`	a��7}���;�=[˕��K1�I�����Q?
0P��� ��s�9�j
�U��!#ݵ������������Z���
g���&E�݂����+۵ʓr�M�XlxVHYEB     400     1a0��p������ĭ��d͘���2A�o��a(y[0]��]�$��찄���y��`���_��7������W2�����=i@np�)Χ!4|f�$ec^0�� о��@�j�[a���`,�;������
����F\�MB����׍�~���w��ϋ��wu�TW���ǖC:s��������;^�AM�����o<B8�qvB՗�%������ZKXz�e�ԴE�x��W��Q����s���j�"��f�L0��8b���IX����0��>��XB����+��U��.G�]���7~�e-�b6�! ���,r<0�W&��@=�-���'V�(�I̕���(Yk%��o]I@M
W�'w`ׁ��x^���܆�b$��k��|h�t�-`
��~Z��XlxVHYEB     400     1a0�T_<)8-��`.�{��N2��uwOV�A(_����8% +�	��%q9O��<�⻻$�\O�CU�"=�t8o�{�1j��9"y�(/+��A�lك"���B0z%�b��XϚɬT�h5��{.��V���٥X��7(�X����&`�����
�Cp������ن(a��D�߅����Hx��!��WEN�i�G�ی��+�x>u{\�"�a��4w�Y�r���[o
���)8�㤪�4��T�5H2�qB���y����1uR&�@�?,�^����ώ}z����0�-��ә������QV�g8�=z�UA[����m}��'�8�)�:5+��4裹���k��Q�!w�n�3H$s�:sr;���/k'�_ aE�ʫ�X�Ck��XlxVHYEB     2d9      e06�qV�rl��ȷU(Y
���k��	��P���x{��� �L%�|���CAq�KƏߏ+-�Q�5ҭ�ve׼M��ƍW�@9��{J�؏^;�wnn��[m�f+�-TdlU��f3�ȸ�M�(�].sY� �$;�g^t��	r�v+�p���+]��tqH�8�����%��D(��a�O�"���j�i:qI?.-v���� G47k�����