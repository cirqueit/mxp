XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=�/'1��MF���P���#��CAp�W<�ixřQ�ݿCU�k��utJ,�F�G	�&���8)�{��]�6�2��mS `��գ$�f����l��F*��g���z.��vT��>�����l�Q�,w:C
�@"��P����Fnգ�JM=F�w�*9��8#�����/�&.$��.@]%A����(�v|�r�kE�W��%a,FǓ��\Z��n1��6zՉ�9���#�9QO���!�n��J��d"0�������#��A�Cqp���``f���gaV,��&��2�I��~��}k=�e���A	a �	��!/�K�Ʀ�,M)��QI��Uay[����?/��o��,�Z�N�Il���Ā,n�y��uVCP܉�KK��ƿ���Āj�˱}�%�M���C!�0�J��5�,�����;�W��r�E��ymA)5ܘ�w�� ����-�ыcs7����Q$�[%"�|yT/�Y�q�JY��#ښW����8&
ǹi�C����!�l�E+��z(����2@�C��-��о}�/qᰓ�o�v�9��ҩ���z���q��N(����w�
��͡�⡛(�??\ɰ?��ͽ]�e�h�1|wr���$�� F�6?"���������z[΄�Z(8���F���o
S�#\2�>�P����#=�q$vH]]��<P
@�LJG���55�u�X'���=;'!�!E[�s�@j����r8߰��i�K�1���XlxVHYEB     400     1b0������j���L� ��������!ǥe"�˃_/�1��Lpt���T�^��@�E|�g�!���nA�ߨ`�)t�vkr��=�à�k$ε-a�t%^<5wz�sJ��w���۪�^9b��$�+��k�x*ʝfp�e�3�E�~�o޾��s9Z��>6C��R�{���{���W��I�be�w��`�Þ�XA%��I�E�W��&�$0�~e��.��m��X&ۻ��2���o�ݜ)��bf�2�9P��:u�t�y%:�n����+-�: �~��Q��[�� h[gO�����m���.yY��k<��v�����`�����Ą#=�3Y��wc"5Vd������E+�i)�tIHI���p�Sof�7Ÿe�:�ר8�w�[g)�m�1���R�aC��G�ܪXlxVHYEB     400     160K~W�.D=e���+5t���"k��3�K���y�vm�	t�6R/Y~dX�$�0����������K�=�p��s-+���,,s��֚��)���ψ��QB!���>:����a�M��������S�$R�p;�:���Z¬d��W}߈�a/j¿~���z�H���CVj�ᆌ:��^GP�Y	�[L]��k��M���G��G������ơ��C�8y��?���FL�Ղ�n���D�U�FT����^� 0�NE:}y��`��,��� jd[˭p��î2�����w�B�(ja���͊*���Y5����7$�� �X�j�`�0��
�,WĚ�2�V7�H&���<XlxVHYEB     400     110�~`5aPn$��7b��e��re�H��>˃�=��W��ʀ}���22|I�5��3����W:J�M+�&=d�H�����I��F�M�n_�){=�ނ��})��Ͼ����lBH�ulf��9�y�֟���~$?OFD]�~����H4�u)]>�儊t/�
,�<�������|�9����Ӹ�O�C=�+�����	pZԛ�3c�Ope�,����PL5=���}ZY�&�'Gc4��Aa[C�LvG�)��"B?�p�)�eO�9�AXlxVHYEB      42      50��e1-}h5�6�+K}^����UW-J	m����ϥ��cE���8���'�)�:��}.��5�l����no�U=��؋�s