`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25184)
`protect data_block
uUUIXe+iO5MTqTFMmz0UygAIDoRKPBfW/435yDntA80NeKTJ+QYheCQXFx4XcyToQTLptYTsg8yc
Ijdm95f0oeuIiPEtUMURwKcHFqp37+nzcRq6xm9ScHNn/IK1ALCiG43lDUN191u06LSBd++N7glM
/MoWLlU8yVTmPxJKhAM74A/l4i38H3bW68KTOwVbl0gjb7dPIqUeuf6ctr3ZqFx9I61yCdSi2U3k
0bxq0gVvb2jhNCe3iW/C1SwEp46/jaAZwRuJvt4z3vd/IKmVtJ7sRrnkE0C0MAugjyWw2Dg8YPiC
PD1OO84HLcu/XRte9jwHTSQVdlD58y/RR2VDiljzQA3p0qWEaNczM4noqgIxneFMCWy3eIDxsHGj
2Ij5VcURz5ZwZ0Zd1xr4mQC17ymRnDLyj2CnBBvcJSB/L7gFkv6hZLLyoEzg91zVe7iCdYrfLaYk
CAE1JJ1AW7KF6MPadmoniF7z6MUwU4s/+Smt8zyJfj0ectgHCfOuzR30qRZKKtmv6VLvugDk4OuS
OYdriakcjxZ1XEzpy5qcBZgI+6x/r3H/ASHtxQPJzeyKImqpwhjUcx3QEyXn3D5zYtc5FBghe5aw
MZXjg/zMcD51wjxupHDFQaEGkJQlKfQkmx/modRFIESanR+iS2sBZF/pAvgQT54XQudXa/u+fTFf
Hams13DjR4tAHtZPi+gvkio/KlJ0MPq8vSvn/b67xX499znAVwApRSfnOVpTsai4+6MzgXHzpYOj
OWnlq/Zkki7nHB2HRy5jUQGGLkDx+6VD7o9vx4fDTx41AIW1mQB/lMGmBPl+ZYiQyH84xEkJYDDx
HcLhnVCS/7Q39/PCa83CQu9Y0k4P/V3qNSJOx63N6GnKr6nFI25oFXKTYcnwjS7fjW0QDIEzJ5SW
h7qzBCNyegUoLmXs4k+2DsoFjINEh11g9Rcr1gGFaC55N79jyxcdDXbR1BOSQz4y3pB6yUkEQxqS
dfrRWqKLA4elredD+TVWRsREzdH1+P/0Z1j5yxXLpSeejkg3ttLUAJ8VmoiU43Ep71DmWbwZlboW
r951OmRu4TJ2L+vzNs8ZWJkz2BM57q6YVyV/Np7e1t6wKQn2qv7E3OjY+mcEGAEbYhmXdNZmSjqb
hISFUv+Ag/xiQEC0P+YpsfO1dB58Yivn8fY8XugM9Rv8WYPeaJXBQnASYRBlggqDIhaphOQEgx2P
huzwblptuH1dSe9OLuRdz0SG0xZDyLxH4RO+wD+nuIwPN/zc6PGwxXO3xYJbTPvGhtipsqpgjBQx
BpnJXKdqVJYeB8+E0znf2NdZrsBGzHeAytpSxwn+gx8N4Are5TaKAjKgowBzEcEN2rqkxr1jKh11
H+rQcsIP4iNT3XI/UWvqyIBd1aRux1ShCYNHKqGrZjBgBAPERm9oPc2B1f1sFavHtARJGCVZUXWC
DzOHozamRPX04HdHwO9EISCco1A5vsiGG5tmcgtKMB1+sOVZY4zid6u8/FD1TMr01HoiVGm//Yql
ZxIZodKCHAiHaeeWlq50mFZQbvHm+/YJJiyW38DVHNXKR/aE5z6XeenY/ZEPsVRg5OBxWv1b/BAc
NPe1PTewlIo0JZLXmdUOjAmt617Ve4L7J/tx8YSD6c2bNm59YWTSi0hwqskkN0MYd5KPFAiQ9evt
kgXT0u7z+3Z/qfXiEBNfKWLXs6NsytejNuetdj1Q23VhvJwFZPZtC1IZat8XNfwp17cLumB8Ktwl
QxhtkU2xqrohlo8CPwTaOck58qaVDghomAPQ8N3BWfBTP1Wjgxud1vKGo/il6tP1G1GTbdokqwX3
I7p96ucB7k8mUagK1ab5j9Q7Ev5bz1KVqLyzi/OX9/HLaSQehwnXH6Rkh1kHuEnRU5F6VVcArAT4
AYVI3SWpWI5JqFJrHttuWVJJrQ12v5o3081jKPG099vlcnohPKCCUUegH9UwRNmfy7gbjO0EDySp
2IqCQdhdeSI/AEFHMVGhRAzm4LX7FaA00gusrr6lSJWYZbii5Xt8s/I7pw+cqDTrAt+M815gaxqf
wU89wWVaHlUr4ciwQ42ywpOGuOS+GiQQZ48YlkKO4WiCH/gAznqQV7bxYGY1ZJeCd/UOPmGbs7px
tXkOFU+0+CaG7s6ewl3iAWxUE7MVLzQl6EXee3QDpNgABwinxsIRn4keLTaAcJRYAUV/CPFByUeU
1MBaIIbAA6ykeuyKuNDAZDtcuoe34o3Cn+9raVAvuCO4JSYc2O2/vG96Hb9uxny2Eo7NEOtRQ4kH
Cq7hRoxAukxmIFbVLHF//cTmkR6tkep06LukEn759cTQV6kgdXSUlLvrG5QXqN2qjOLfd6WqWvhD
JDh3Lrv+voUYBiLXlZTV1sCvaTv1BYOi8pAPsJJRxbrdMkvqk6sjf85RxHPBsgMi6K4BBuBWPnfC
63O57+kxVVNnQ2LiA5OW3Whpc8kx09atDS5vBesGdCwg1RaSuqSoww5ipqELAs865gBg6HxteFbB
19bqFaZOthRE8L7S3qqjry7S1tPOzILtP/RY9lK10bJrxAnzB/u2Dl80olttwb0G4dFiWnx7G+3u
pVqvRvmLUlEMBm7uwjz8BVOQWxYT+EYA+VKCnU9qh9T+uX0MxMk/dlIbtg9N7vbn/71sxtUreO9M
8o5xFTHCYl8SjQWSCQRwiLx1t/r1Io2ZnQrGZsA+9FQAVL7gjnGeok+sd1Si/SS7FnCJRZYy/iZS
Kp84wTvMv0RdwwZQQIGZCf3AUc6w1uKU6vWmGyP67YBNTlymrDsllgV+fnH4ksV4/3vnKFerKEdF
LsznM+J7QS8AkEZxWUetiDpIF6e5SnmkmkFwof2zN7djNE8Im6cxlpshExE7PW9C/RHkuKXfq9Gz
IWRpNRINuYsVUoka6LZJViWK9zj0Ee+odaogn13sammM15hbH7mF6l4TNp2OA6PtihfX08vijIJ5
P4HnhWgS0TOjvrqGCYefR2ur7j2ho6ZyJC7MxEL2pe7jb6ztOelGuCthk8AyFhGycP5Rrb2eiQFj
os8VQm6sLWhGcoCkUK7kt7NneHKc/n/KCxEPSUQis/OrRW6YnNPG/H927c3WFYhNuAAgYmCyuas5
y1lyZ8X2lThaVmpIbZfuMTRfgHb4T8rdBMasof41s6AVLgsTDHT+X0jHriMsDSMec3CBXYc4K395
X0qD05v4+EiR7tzyj0dHF6T5AWGb5ZlcizsukEht6Ope1uRUq0FDs2ZywpPBBo5IYmrd5z+g9OHm
+5YV5F/PG5MAYtd+Wo3OkLZFlzR8bArZi7xelM4bKGXfIkxK854nwGDbdMn8kgFE147x/kPL/rtY
hoTg7hwkMnF1d5zZaphbxJu1MGP1G82d3jymHF5UKOy3lh0Pc44cuDbo19Q62je18zPedgzzUeMa
/Mk++rUR0MELIZ4RWUKaxpugyuDyGeskolI8Dc5PgABm5+QtHjEqJ5/Yn/U64TW3opYumn6UIcXj
wYbVwIF3AWdYSYfkK2802owxkRPpA19X7J0FSgXs/CRoEcNpNcehe66Q4RCvKUy+QZFL0wdQ3Exm
OSxQLpVTbZVhw0JXQe+csM1jPs5ionbuy5Wwk29MmrCyMzz4njhxh7f8xenjg0hfigVAV1zz1UgM
hUV6BWH84RNX82dfqkxRRf7e55G7INiY+oSHZM3c31CM8MRVWCrPp2Es9mai8h9ttlAYNW7xU4IU
HFbsBk2VDvZOFLZO4xYVyJa50ULtmqq+k/v3ngIjaINjU59Cd2Z9fxcSUZE+PtG58HKM2ROUfXOp
i/hr5WJbDO4gWvavfw0DQe4zNGhaVsgOpSEY8bOcS0pr764yLyyN3brjR/QsTQ7b9UY0IB6/nHPQ
PEEKdDxpXc4aivW5HW3hCS5+bPkXcUZg69DWPzHmUDNSp6HOvqKlXbj4cbB6yN5UEPctoUxEq99f
In/Wk6SjJh5hC3AIKYAWisLpP9fdaLloR85ZqR9g61FP0NVx39Im9n9f6hdZpQktAHm8j8EF5R7r
XjpnuPMT0zJPhVY1GBUXeFuylFUo93O9ci1yam9J4B2djpyZHtk3U1uJa8WaGUwbmeDLRoEhQyf0
ZitZ0fqOLFaev3rUsOAwJ6y8KMVFTZOMS6HmIWY6Y9+hRQRj0OquevmWoZsedjMpHsvLZLBPjiRF
o5b5X+wGNOWsJfBqM2AMms7agafOduBe+cg2tZ3XSiSwnRIf9bkKEVD0dqb1g0HOG/o6b1+I9G1U
XmYd1G5trTnxSTh7ZS5D5BKPhxjZl3HNrJQmSwjontuRKMl/kFRampyY9OXU58TKUClB6btS/6bE
C4Vupb2GlyAykmHpmrFxlmnaBDvWuck5ExPk79izFp/QHZWzOAvN3u7yARJUhIL+sjbt9nBhdjvM
AfEO8N4rDgGWfT2H4yImyUGSOVi0HGkFejtfM9dCLBVh6jvmG4CShNDFcrM3TRttG9kLvtH2TH9V
JrRsHOPFqQO6F7PoY3pUdFY8k+GwtRV98YHyQszRhlVCRc7nWmCqmEns+TOco3XZjNZH6yUK446f
OpwkLMABqxFNdpKM6wXpsnCBB5oWzTuUXLxwnsMXNd/E+6sYZLo7w/OyIBmR8LeyWNlY+K0x4y+D
vqEvIvqEiauuYkYnkgIfjaWIzVZs5yxHpgEdqzYm6oPp4oB3ISVBfbVAaUK1jShNFI67qHn+N5qn
1hQod+nxY0ef1Cmcekwl04txgruD8ZTUCJr1DvkXFPtVpoKWiUon0+Jd3j1MVsrkw6QuZGTyVHkQ
Bgexs5+byQksSz8sAPErHA77dFZxv5jQT1PWVJjhf1j8vD7fvBU9nwl3xfHrxZSUVIzSW9aVbOQG
PbLQ3mZw21SsCvm0Hr9DiuGgjo2ZNU4Qq3erYwzGtOafaYocQCmHve1jgaYZX6Tph1cDQlMr4tQU
TS1bz1xBqdCIKfAllyjfBEKBI3GH7OZI5P70X5vxw2rE0mtNiA6I0TBJ5wKCx6SVVVMJgvieunk1
YV3KzW6jJzHm50I+A5gPsC1MRcj/ljGv8gDBggZxrHaPRBZgjfxRGe4UF85UJPhbtRU/fs6iWx5K
SWH3UpgKcn9Ylv7f6q3Y7OyphP/INKXAwUiwjvSmfX+xz5XXriET3ObiXohmiwEMGesEa7WKlC2Q
3wMzSBbv1EpBi6gjcwN1YB9XIo8lrLjgwk2mF4IXNyLhX7QW3lKGJUcIvA1VLHqLHUPzXtwPEcTz
2EhkrfHo2f49jduaBUnxQp/hea3F55FUGm7Mwk9iQF/l3+utAZAFFpv2T7g2lPsJRK7D0CdbCaea
A8du/2AAqx8FaZFCAEF0cuz9GEZO0LEXW09UDQz842v0iaWKPZZJu5lhnEPAPnKqi20f2/0Ik1lY
4n9ltrZLSDQZTiToizP2JKZBpqQNvfXP+ryxmgQf7Pqmsec1jEkIov8+e75Lf3BpORPkbVhvw+AE
5IRplENEnvMu+l5Oxg5pIk3EffWRbyRNMPjgY06KFLTyGHoDYWfRDNa8Xcr7XV+bZDvn+s8B/lep
jiWUQhbf4/sYvBLoV4xHLLSYly5IQYOc+HWiJzW1XxQbkXEnML6H0VqOximg7Q/sU8gx0MmPXqBd
ucVO/bwP6IRTbrOMTcvr2c6FHOxURZPzQpdiqXsiLe0VDfn1xfSkH4AVLXr2jjK97HDKWs6g/f3Z
0N6+LZz2AWPrjbf0voaSJvc7NzDxvW5hh9DZAqUGJrOuSCyV+ghxztsp46OGi20PKpsoLw9n7SQQ
Ak3qPXM9taOrrRcTcHuszsvDUc+W8URbFWvcoER5/tlTtakSrYu1pX9U8GekpTYFDz5qMOo8hKaS
srd+0BCLO8FT/OQsF8Gc7yKkhENFk/csPKFG+vi7rCL6FNQJfRZ18PBFf0fU1wx/M20Rvr0bn2n4
c4+zh6T1BxKA7HSCcjW88T8nnA04KVDUbf4cFilBu0h9taPsPh/ukOSGgGGpitYyDMY6DftRVMts
RzQzWNWibwdUaeb4pP3Px+IDNWTtwrYjuenoZ6DvAgc7M49RvHxW6eNfbJOZ2d/5o1oajSf+zQE1
xHxaxvcr0DbxZ6ZJgfllE9V7DdCCSJ7uwdkkLUbtd/vV0JN1BnD8QbN+c2STPgp/VLq14tjJRT3Z
ljInx4qJeoc8dCm8C4rR8k+iJx+lJ/791scVCC7h6NGCBWQLkSxfTTR3jLjjj3ZfbDArBN0fjHfP
eHLl705LxpwwBfpZmRuj3hGxZefbCgmTdr5I9d3DqbwqmQZxKdURV3ew+09sFRjtmdu/9odFDS47
v1hbIGCplypWHrxS/mqjzr4HGWJF4bSQBZCp3uhQB5R7tIsMUZqFVIIpubqenqy61rT8PeqRYtMG
6yJ4A4yErTyFjGhsqScqXHVvOcgP96ElHtGR8WOSOHC1aYruv1cX2dSP2XoE1aavRfbG/rgsoyRn
FLvD5XyReCKqiP/YGL+6M1jkTpExAkVffgXOnhKunAfIabJTjnB1kkeVjNACC9vcvNm2qF6P6JUV
ktc2DqWKyAt83dEx6u0VFXhVqgpVvRaCsRwBMkiVZ2Ndeg+B7ei1LTR8qzdzO30VFRcAfJiThed+
OqacVQ5WBIP6IxabddFoSPVGcbFPjQyen7pQnvE6QOrMk8iPJ+zj6JZlopKifz7eQEvAs5CgNs2/
sMtJu1du3ZP8TVwVCatb4qtslztIIBW2w3AjPm5Ps9rzQ8TxuRcAXaZ46Gf7cKfKMnOkFl9FKoI0
Sgqkd1fBI4UIOBw+Pu+AmM8/FdF/0ivFOshuB50NrcfTNoDG3dLALKEQwgTgkATi7sFOtu2MvfPg
LsNTFw9IvHkBzGm/DNwO0kHgdYD/qsVV5u4cu11kKpJZQDMDzEZU9sv/VUKZ/BulQ26zkERYIMUz
WPXtfKKlmuOJLGvADehDuUhkdBSqrMJe0XoTfVGrCyXK4GPIOSgLnFAcER/TAbYRNSyAzAv13t+I
7kA5AAGmfqXX/rPVCNVckxb3DRhqHv3v39cf35LBncMEuqZnEdolYFSsyvokO2HcPSy6uHII/WnW
T/f4L3E9uFXmoRp6+b4j8/GCUKMd2wIykO7Bki00pZUhQHxWyfvVaKDNEfbnFI4VMOciyhGTw4y2
sWa4Wzk5/9a7z2LQm8wEKeNtMb5tbi4jf/AGzpCwt5N4D1qWC4LJHiSA7paD45qPEyy2YTnwumoI
+7QjhAPiNWWKcNLbRUXU42EX7g7Zth9XtSArTdiwVcsCQUpN+0MkHM5Dj3Z3Yw68z3JPMCVeMUF9
clPd4OiLmJ4L3fTNL/JeM8CCvW9I5p9Rsveh8l28YQa0mYvGM62T+0zsTj4yzCj9mAhFAOYkLlN5
Kj/AS0IMLTTAlQGPaBpAop9Dnqi8435mB/3ol+QyRCDeugTvLOCw04c7UCmJd2gm5BzGMuvAIKqI
TDbndwwBuxoJQ4FspdEamiAndBAe1XBt2H7tWxu0NYqtqDoBcNRNolO0PUXdn1ZHLwOtYj+4O8NC
cbjmioWaGa/nH3ImuP4McUMdGvDkz/oivGIsyPKnqVFXy8GwqS+GMKkeRYu9rUNtQTqkD63qFsw0
3EPrug46OjGvOHcKxCibop4hhngNRlgukm3DUfKNBbRV7ir4h10F9X+8zmFfkCqnxMnWo3bUpnfh
ycXVO9vB4HM8QA0wCLTSsptdyhSel8rcWl0aTovUKH9poRhpbvNH15loNoV0RMkzOibY1KLlpmAH
2i6O0RwVayYT3fQs97IuM+DvCc5p/e7IlejOzBPvSR8JQzg0NcD8ck8FHhdmKjwCjOyj7HIRI/mC
aUVP094AJKBuC9tAGwrhipw/8VekveyKtn1+ANbLBiSbowMsLA8EkexqLrlQEpRx0I4jtpTOsXeA
ftv1mgPts8F+OuW4sgjxk7RQsOK95I5iTRppg17WsTToopbuTkUs/hrdQkHzjFhcOplsHoR+8JqB
O5GQOkYdSLmH8r/5lx3hK08X5wk20GIqmNStah5o3q3p/s/XxgPQlvERBS2hiNVyotOeHzZ/tyMd
cY7y4YrlRqYdWdKLy4lv2cl1HTOpl5w9dhGh01n5xIzbIzaUSniyfUnqFc829bNy+3N+OzoXoXCd
5Yq4IzzQPQeAUQPKROYltI12l/Iej8D1pkd8W0hl32UsRhI6RmbySCIPrVAAvz5OyyY/htdRLeyp
ez9jASHpCWgtQr62tPQe8fvBZQvD2yxyTfc9g6qc4oIG6MVFwUBat0kKpGnxq/8LTOBZiqdhQX3t
RPI/RRpzdhMY40V8utEK4v1LVKW1qBWUj/OnSnGhlzuq68dWc87nMkImlEzzAhhK+caxXXQtiM6J
DvJYdx6UzJHyCGEch9owocAMVf0RinV2crBj/P2Dg2VY5AteWK+Dfc/2CYp4UUiEFZFIjuoxhK64
sbi128NleMZEpYcwbKUq65RwbqbKnqtPUuWeBQHUrg1cUdAaQ3C9ksStDr9dtq+JUQbP+/OtnNC7
HPsWZDQvks7HGtYkpO3cUa6Ennl1LbUedF3VPTUWiU66cPe771CfAFLGR4xQiPkPndDrokQ+BJeI
gEDmt5Wy0ymGBKV0Z/LL1qzlmbW8CI+Lv2uObO7134G9KO4jzUCIA99ljJkBGd2hQfIaNt20wBRe
Yl7M3I6FvK7cCrFZPD1EYA6yzzBM9dSZc+J8RMO3K2mRh2+gUxwb/EiGc4QLiIwhjf8OrRqzLLZF
eDOFTwCsCA5Oe9P0xOMgxWiLG4aShloow6yRahyOj6so9HmfA6yRsfgaAyxWdQ72KxyDcIXf6E1t
wo7CsJXxSmvvbeVb4aKFvaVAvYjkTZOCdxpMEFTXiFMeRhwvEbOVs2iZyj3hcKbgQ26SW9INqIo5
yzTGov6uM2+2VjNZ/+3iZEFE2PTOLNVbXzz+RtcCz0ZflYBA1NdcBenjUCsqKeYukZrxg2dNu8MH
qtTo+UT+WrLwEqxYXHDTMHLMhO2btJQgfsNF+9MJSr/Lw6UiuKmFrREgpqy6lSi5irRg/fRUmruI
mQ1buEyxNa+tEc3QVAFEjSI6v62znZjg5g02Z2a/eER7EBaWuEt4O0te4bDkoC407+3LmtUp+QDC
grAteTT/EupQ7LturJN/EWGGXIMfJ+p9gUaEvzRyAQUIqvb6bRmiPCkst8tZv/s2EQ5pa+ruOpKc
E//jzBoZbYC3oFRm+GNXl8RyMGmw/pDC+FZCcOvvKQrbngYk3JZK5yIvM/xNcZkWBp1rHD1VMM0P
x2ZfbwXuvo4KQ2zwvaI3LgiUh5bm9MRelGIOmIWTSuqsS7IG95dXvJ+bU9gx4rxriMS4bllKNQFi
QqlXKrD3QBhqvlCbNckrBcULCAC43a9eZnvrukI3SK/mMFvowRMvShxErzmQugt6/ZrF+Mc9cdXB
rrZkwcVBylXQ4X5GOWGCqvWKO3xxLuvC6ja1+hbfhcfzcpSf0x620MG7xB4yqa+77hJgMVibzg+f
LcCuSpGm8wM3cMNlKIcbOQwScn436DxrkMoxejulKyHtooJk/vQm0gwGFO/5toUkTP+RfAog/SlG
EoNyIkRwbSuCDPYyc6S/LV3SVvrPJXv4xluNT/e4MWy7IPZgQW+TnPg2cAOwcTaERZZtK8VBXAHy
pyP9CgpexgCveOARjtCvZ4JyfACfoZ8OjcgiP7KOYQQt9tPneEQxT44VzKjbZz18FANexF5c7U91
d6waVIu7nGNOXJMvrjXug3qbsu7YRjqDkMpV28elEXpl63OErgiLSWPAf4Gr7gwLkxUMkgwyVKT7
7XqSNrT8ehGPKEXZZDh1pPHaXUCzXcYdyJAjhvv0VLPxsVfQiXZhVaErQHUJTwLMtolq9H78eVB7
q5mgbjm74k8XocK9QWyXCOYeXBPTgk8N3i23t4s4VOH5HUUDxuHvsECU3Ft+xYG9VFyTi9CcJ9TN
fckzl1LWE/V1GTbg/aN7PRv7kcnnRQbE4MWmRuPaHqCDvT4pg2m4dUySCXIuZXFf6nOSr69WdOeT
p/EswmV9GRxA4BCeMoOcZpqIn9cII1pmR95QoXnd7WVynArzXMutWwH5Nl0YEYB8b7w/27WaicdR
C4+Cz08to83QH0vQjRLDImQdCa6RY1ybLNpfjA4d3u/lBAGKPaGIshGvYPDG+f1i+OKtk6Ewv7hG
tYnF+ysy7YwBmthEAPBdsO/jiiziQ/Xg4dbaymuihWFHY4I0wYXOxK4mNVcHekD8d8lnKlYRxszu
/aR11sL1lJ0IlY3YFZhIhSfIL9pEYrd+KhG1rl/6QvfEXZtHPrE2YRf1rh9ca+gx1jwuTlHfiGuA
IjVW9zcaQI/GIYyD3yEcsuZVT40sG41Zj5cHeg4eJFQZQjDcu72zC1hSgBGSQffTkd5kQznT3bjb
RLYtRo7/dcz8TiO1qxvpu3gKlrwQ5dJccKxhS2menBn0RyvQD22Tn6ANwYLuld8dX3wfwSGuP0E/
GCI+Jq1oXVPBZwBbnRtNEpCGZVia8n/qA9HN0Sa0PBOipIZLGoK60gx2wS6jRjCcx9isNytTpYWY
b3w2RcPx7wd5/tHqyGhH84D6f2f0DH0Y5nxh74eHNKk/ZC6zdEMbTQbEiO6+CPbHWc9ZN5mNeit8
fb6uAD7lern64HnnT2ObwakFCBxsLOKE7yEP+Ijfejc1D+7Mpx9JmhlNz3irQlI9Lp0KQpx8arKR
xjvI/IQBapeUj4UgIEyk5QfRr9aTMIs5/hFb3UwZPdvg/SLz2Arn0ozvX17xpSxeQKyN1JL4NIK2
itzxRF4pzCJhRysngbYwB3AKSvyCEkftDCSR0Fifc/3oran4KyDwBmtjsaJc8FBz50X1qP5J0kEL
WlEaMKF1gK5gdj160tl32mhlIVUHWUDRi4GqTjKPlB3mmMstz0LHDZNPZF2FkuxH+s+C1Fxn7TS/
rMHNSzS9ifWp5QjKvAVSEsNj/SCcEeaV4EXIDW6ZEqvrs5o0TyurekTyh1Tf9JpI7VsUdUVEC8c7
zx3ZZtCAeI3o+dpk0lpXXarcIJJhssWacc3PnfXB4DhKuqLcLw887w0ojFjXG8zyubGvBPFfvF0c
lr0QUrWh5lrFidiMsfYNYIMocf9lnVePPxO9ehhk1POi90g57Nht2tioB4Uds+6DtrHoMvRkpq7t
nu4BA1+HVgNgLItc1PBys8d6aVlX3OLtPSjcXcFrgkklVwXfRGipwqQeYyitYO5rb8TmeTcvX8vC
OWNO+bUSq6CnzXr5CqvZMDlWMuIEZbWV5BrBFmaZNzyG4rbV2av/KldbNu3ssI/15b/iM/xgxcwC
A4OdIej52s4BXjrfli945V3xLUgXMaPr3ym0UdyvBGtld6UMU0wlAn5NPFgF9TU8rehzcZrU1Oe1
+KFCeYUerdOLD428UWs0ruAdemjS5JmRpZnlI+BX7H/9EnBCHFSOKxf/XjLjIJRHatjdhfTzGjlT
dMKgb8iSpXV7ndp49G73+QshaErb4z46vp0dYDc3NJgIgvOBjmC7sBby1/yA3msbQrO9ca7wcL/B
mQSc0xLXtWxBLREYvFYWR3dcEYDrp8YUwHTaWstvqLyao+Q7OCB2+YywpcispShXIkO4WjkMaGsP
BDasWcYHFz7gSqrQCeprBGbaWC76rWaEKCMihMhtlG9eur6cPEc8QFMmz0HKfyO+ce/VTNQTp/wp
7bVrsWohBqHTWJRLwhv4JkxVqwXEcRmIIULpEQh9mw7wukVKv9J30kjN5AOdY5u69Dej8/n8+SG1
moxg+JDSzEmZ313pqKUzw9wv4AlKScoeK3ZFDp4oYpa9n4iX7BWgu/BZGvdS/TI1IbP8Kf+GHjgt
zNz4U1DhIPzj6HPvqDIg7JwZhEh5lyiq7BOn14FJ5RkvaeGlVgYQnVBsii123aRBYkoOEMgQX+EA
HmdSVwMgSgzLI6g5udYSB/uG2U6gyPaij19SjnVUYJvFJFr618TvD2twTDuCuKmVBNCAxvRSJW58
JzuWE5iHyH6fGqbKy7fIdxA/GyCWjrw9Mow2oPmsGEW+5nH0Myx7kf8CaqxlFEe1QPT/s+E137i9
cf+Rtvq+csYK+oJcTMZYU6ZfriF9s+grPamg0ecO/KSA18LD1aUMPd2wY2cF7nszMvtGkdTBYezo
JmDjui6fievxKDDQSKD9tXt140JywE/kvWc2rw4FPSorjbEYu4+DaiRMcRh+q1k3tFTC34HSrB5h
B/7jOTsfFbq3y7swrhvF/i0l5ZFtrPz7mHXMBE2Nq9lUu6Bz+VC5IdgYKmuKM2OxaPdzGoNtvGH8
P9F0ZW6tjqhOFtLcYAwKaYQJXTKbguo7lDNdP72NWFLxLOH2LGlyXUZjzDSwJb95yCygBbXeT8FN
CKUdisvNVgt4/uuurVVWbsmZ9W1DdnwzgrvlYBB9DGUi/+NvQUSfsWgAIzL4lFO4MX07hXJx2lNj
aMMC6dqdHtcyvzkTyfRHA/lrZkSVLfT1gvAeh3Y3MSJ5g4AQ9gFcEep1OuN/HD1Wc90VvRH58awb
3sBT6Uu9+zUl616Jg3IIs6FScxNFdMVYv9P35bTzyG3g5tVN46cNVdOrypgUgvmrXo79HdFHWX7D
sSj8YvXiTpxaxQSdK5FNI0q6lk4Xc+Fge7K/2F1LgjWLpcwC4JYbGsrQCnbJu9qXBySHdwpXalGW
J/mNXOGBbquLlxZcaFmjxapXfv5aXPVrOst7aztdJDjJ5Aw0U6ATWn/HbBSiIStJVMZxNCn+wkvY
EvOkj/+hrw6yOH9MtWg0dfmZZvgUMqpefRQHzj7/bBqAlvOLlUztrNKR86pVGR8wucJFi+ekbIk8
GaWuMrufEfrdisvVhBkvUDfhfhXHXT8ptkO5HXBPlxYu1eG0ceZ+yBWOrX/bEjzqS4MLt4NAJBXK
KLznDZ5UWbvt4flaw/Xm6lwgHalJ+M0d8OR97vi2WoUgqbMxBqDmbgEvGz40eGi0pZs6HgzdJolV
Q/97srePGuT4F4J04sXTGzTdiCF7oInpJkUULK7NJRXMXpiVjYxs3R2h7RcgDNhOhpPo9BZl7VwU
T274fmVxNA/LwmCZ0fWfY+sn+3ddzqhD1S7kktC+c1N8m402Mp4jsJYcnOfuuq2Y5SpUAU7kIkHj
1MdD86hI8j41gywpXWOQxCPRzvNSfDYpwYe8GZ0zpg6BpR3yUFN8Vat4JnehnAb32d99DuBCcZgU
Y029f6h1hUffXLL9AkDzFKf+utMyzZQdc/C8xCcfnhqJ9FWS+07g0JgwAvVc+OGWb86UHSPHAX54
pntGUMd8QR+tixB3ea55k3hmq8+ifnHyo9uaTryiVMd2wg5g8ayjWdouUbbuTh8YpHq+SJJZtTjH
yJedMmB4TWaYe4WYOARMk0ncZjnOueBnWOPoLtwR21Paz4ycHcyoHyXGF6zwmZAEnreNM2GN2Y9U
xDToiYQBCSD1ykTrN2LhUt0BkXqapdGwcOiKf6hecGkuag84ateHXlMB7bpYHVbOME9J5GMNaaxk
gT3D6+GkS8S0auZ8Nowe7oHMWiQlZpz+zgWfi7Xas/Uq9MhhL4dpUfxQ9WMJ+j2gHNnKLd0KmShm
Lwbw97gPc+u+V8X3MK4S5hpZgrvqONiIEeY+eznh0y0GL6mwxohKT/PBN5EvDcMpCNX7MvexBCdb
rJ28erM8KxBVHcIv96Hd9uOhi6KDMoUkel3hyn0BE+nD4w5Z7bWhGoZZftu5+FQFeD115mmN2L1h
2bARorlLyVp9HONqbh0dD8AVnVdOXdIghrBNa8BvC8TIPJjYWzoAvb8sPJQhFF37nISEEvg3781b
JN7mcUcPqMA0+gDmtM8RnWGqXJxHKuTwtu92VouY3oHT3Tj2B0diGB9aS+VJM0P7VoqVcDmOYtxB
U5p2D61gSUchHiWSOJ4ZKtCO9VDw/xgdWA8rjC9l0+Mw/fcbt1PSLJkF7rjPiI6P+DOOmM5dRZP0
dDBAjV2b03SjhSFJaXbcmJcm4ydovgOumHR2f3QiDQqjVTp0TOzp7Aipi0p5WS4cKTft5+3UF+qh
yxpEHwXt0hcLAVXdG5/XfumB9CXQldX5jLsYsgsnyLJufTuBLWkIqWZLT9MRRXfA3qCuEBsdli36
210qtYcd/nrEryLdeWOPE0TrwFP7w2cqaST3vuKB2aJYASXn6nNGQu9X9sJ8Rc0nxpGcELVxpp5D
ME431iCB1m/wnUD87fDWI67rR3VCdJTRCb9WlEFa7Dy7tAESlUgTGMnpUkuYNrVkySsZzoVumZ51
SbOzbsRgt29dKwRdDnRdaUuarAxkC6/qqBZznH7RMSbt6TR4eQNSLKMi9KubVyr/4hGzW6AWKQ71
3J2MeMQUmHAtNeQ0PbAv7ghDlUFTzSdO35c6FkoD/wkLdP4MFJdU/dh2oqsAxqaQuMTxQNAQuOiA
b3mFfU89ZEGzv/P2nEfPj9w/S1I8NtXQjQjLw0ti61k2a2oyi5f/l32SAKwjoxgGSzcblXjUU1gx
Hy8tIcHYmzPptfQgFWq2zSQfX/k0yRmpBx7TThcv9OXsTO4d+Xue3EejZZ4IRulgNl094lqGiJKJ
A32dd5l2mo4Sh9j57dW1MebEz5Eph6J5eR/61wAgG3V8bk1MjbyQlusQLqw83HyiS37HmZcbP1x1
leY+T6nBrjWeeXck/ZIzeD4e0pyoSnKZH4RkiZnK9EcZAqWeq6pDZVidZ7+TOEp3S3WxrkLm1tGy
IMw0dswwMET6k9vpCmEf8Gv3JOVSHHDIJ4ngNwQWwgJBtxl3TMn+sivcuGK0QFWZUkbLkA2ZWydq
n21pztvtJMQZyTolN+Nl9drE2xGJ8x7GMMhENmkIYEWqEr7OkPrLeLQ0qdWnypqCoxE2wKlIHb/m
2vQ8G9mWpp1ZKPmbNbQ7q7Phf5wg/kZcjsphNZWZ0LWnoGWYA3ovy7GC+Z6t9T9zzhispG9yWZWr
4HL+2qu2o3pMe9BsVow6JzPgi52l0ifZQ3lnEObQ1DyJInHAYDgbpFZSXCjpPWJj+JvJ8qV+jcJz
ltEKIbGcbwvofZdeco5vMZjkTr8BuXVUZJM7Usi0ZAgNsWgjSOsuZYQ8FEx5aj3ZoNQ7jBB0g1Tm
nclAkS2HpSFzcg3VXAn/bBzctfHbr+HM3KV+NxWGkRe4EYpMJ4aAyyWQEjolZ2JtZXw26VtNIzi2
imjMW9Nvs65UlTiczupbPtk1ZEq6HSdwEPDdfelklIA/QNWudcF23j0EXCZkoEFdBo2EZI0PEwcr
6C0Na2GBFPeid1YD7f3+VaiZ54Q3LAUIqFJnBg9d5HNfD8pITwxVa6qwojDH4iGKKNdnDvPRm+p5
NI+tJTZxtrFNFfDnoUabo/jJ2x7+8fFFgOCPwjH3M+yLt2Y0R173FNkdGMmRopbqe8qHzDKj/Teu
u+uMe02bEsN8X617iajHbdPGRchZix857Gf65Ro4BRlp4xd92sTvWTVaILQVOywir27heKcm3F23
4OKkPGeV9uzgSm+870DpgDaj2m0g1f/gWjz6OAlAMN788OFIafelSLDq3wh5JvlCSz69iJ9MKWbV
to1s7vxH5k4WvkADPuFKNfH++woUA7N36N9CKXYKmwlBRPWLDuAyPynV3nl2Y2XaAMoXCsmGlIC9
2GB99MMa/gNQczsq9bE/sWTiwNcea5OufW3XFfSIJHPI2Ova01p6a9yuISzRcZJbXoAyV6WwJAZC
GCqr8F0rT5yyJQn+pW+ibA7zxSEp/8buQ85saemrMd5N3Z/8qEA2qg4bQ1TW3zTefp55f4ojMWyQ
qdkSSF1RUssFhuTvBzY+USq4+CYgYHMKs4ytdF6UrK583IVsfGGvhc1E4d1aQ7oCiKoD8/gH0Jag
mqku/nwU7M0Ovuj2D3ry3e1h7F+2aCNjgNfkCVeqk7IBTDDLmZ90Jk2mCvwWa2JArq5pEtagf7uH
RIG+GOpsooshNAHz0zK/9WWWeGIiTg5Rh37S8Bk8auXhuPsW8KdDsofIR9YO9350aNCO0mFzs85x
efrEXODLlcB1RkVVVqNpjQje6gJGEnSw9hDbGJLL04wGS8upvJJu5McGEWnh8TRqfo0byMuoZ41v
ETYIEdDO0D87qfQZWhV/u9KfwQtCYjV3vC8uiMW4NOnH1a77P8TFGso5OVHyq7K0Gd+OvaOQl2rw
Vh/rpJKMCDJ0HBU0TNCsHZ360fs3oOhHhPKLvdTWvGy7kT2lXH70ut1oPesq9Z/2dJB7vJ5y7T8s
7EJ8H28T8FKqwAnHPPeQjrWkp2cx/VBY/emmWVrLH83XLxBBbB4Apcyb8Tmrm0ERnKOuQHXD8s+1
Hv3D3nygn902kL6Aw1Wd1860ys+P4gY2ntAWQhE9BNMTrX2X4C8MeICM2WKKckuiyatnPfcdULWK
fZk9z1NIw/EfWNm4sRfZXxODdc/Fx/p10JPSWW+VgoAhSeSqzWh+KwvvG3oU+ZFbO4I7dp0rhVF5
BT765KnP9Y1BkEsdQ3xQVZMglEGC9Ver4DaQc65KYcVPjW02Nq9xzlkPUVi2uEWVhoF+tEooQedp
JOX3E7PDBowtBTBFNG6ZGPJ7enAXtRe2EY6OwDiLQPKq1rtstaGW70Lma+hSfEJu/YLcTpLZUOvN
RfC1KNHSpPD5pwls81wTjpFvU8/KlxPeL8fremLc3BDDNG2+NoAWU7yvG6y1/ZU27npdDzEzgMn/
UvhtYbmFPTC79nmhVSebCUhHRIS9Xhvml9oBvNxrBDfd6Yfz2LJzrPeqy985AE5z5bajrd+YBM7Y
buSCGDlwvtU4+bdePRHCM6kSOLOMKqADJsidyC9o5Z46dNritSk8RprChS5OOC+Db/wVPa53VfOU
TtTIAyGafvnPLz3oDtd+WxDIHY9ISOoF3LgyEW6PhgnS6eUyjCo8yrDO3SbCTC9+IG/MQV/e+S8Y
s7/hkH5UMZcRWvICEL2W2qg+KFxM6WblMcGaNFyH5AVA6CIA8PjTnN5gDvsAVRVYCeREVdnAvMGG
IUsLjWVBIoSBOJAORcmJgc6Wq6w7IOUZvWT7YxPAilRTEzp7siiSC4B/rVrKQqIenz4/19FH6HwQ
m+kjtRs5HBBWTWW/v+b8tUdSRQ7/K/pq1rWVlLLk9GjZ77llJbRUK3FaVQYx39uIgFNj8HoYTRzE
t3VRX0Rbbvs+EWz9uBNu0JlCt+thCk82xXPlNuXY6IkGoPfhQcyQ/YsGyl1LPqZp3r/szZ74KV1K
amlRebG2G4vC+yaJtmEWGkEuHlhAA7yhgUQhtxwLDDtYmKkak0zzKQDozYfKRBlilS3oRllSbQfV
iE1Jgbe77YBYtLqUxzZxTXcswgiUNba5G803NfhJUeEe40RTrMN/Qamxt523AUX2VYK+EhA3q1wI
uGIFDYZTUPIQkn76JfuO4jVbzgQTPbR9bZB8kxrY4zQIhEFsxN2+WYXSpOw9D1ssdqLHuYBkmXnX
6wK/j8imSO1p/0Y5Wru41sbHZShwYWp02ZyOB/h5DAobGwylZK0Zux1h6Y8fy2njl/tqzK3jLkkK
9V+xhEccx61e553wiI3Dr1KTVB8V2rqdcs2/Qt7Jgl5eDrECtul3Odf3etkI0/AjVrM4HbsNNER4
8k2xnMB/cODYrLlO5NbhVycJpBELQqv9KClncadGfGN8PM9jmK8gJNJ6wzRev/wdDGCaEIJUTLBS
3CwtxQdo3mKXP/3hFkAAHgAIX+0hO2qItWDsis9dYsfW075HJKku14FC4kPy+qN/+vYeeFipQlIe
DaY1/rdf78NqYec6EYCC7BMrjqLPeqUBbrybIC4GmAjcm0cOCpKffwvqHP4942+tFOC1ApjYGP/K
6aixXEV2pyPSJFby+TTwpDG+69MNe6GFZMnH9m/j+LPVo707tQN75wVA5NsvzdSwQbZpedS+P+07
gQtkPL8tesqukSJFaO3yE3ld3vEyMx/dvtOVDvKiH1/7/FCrFpmyWBlfYCAU/fe1hxDhNinJRwoi
EbHhnufyu2gcvyFCVMXSGDsKvp2y9NEVkoWrmw49r85FLOWYo+2bTp7ea5E7HMuIZ8kvUF+Zzv/w
V4wQaUuxfJTrJEp/JQDTuuMSN+C04LkjV2NoaELoVS9SkE8Nwyxz6wWazkb6K3JNeJln6lpFmG63
OZvJhkYII9S+i4HvP/1B1ZtD7q0RvJGoQ6cBVlPWMqYblykUfbhuQMci0enPkKEBc2t0cYLt4IwV
j4TCesh7SRljLAGCNO8GJyPJfJB+yGu3wb4QckEwC3QP/1f6+Uzgjr2IDibsJ46QGMDo/OXGZmy5
FtEyW/6b6rhATxZvaJ4Oggu3vw7YU+Y9taJXdxpwF3mlmp0IPCEII72VqC5xlLA17bCsfHS3NmNA
ATPSPBAN8f26pAIE0B5w//vKwZr0dijoFl5BynzmSPYVHgFdy6mKErVT/oFMXOcY6RJuWSjbDvqd
KsqAuq2YJUfEKw8U1Xx9R6gVuNMcH+YZbbwXlzGYqxdNJdVqujeOdbY2J/fnasGrjde73RhbC9Za
ssTs4abs+CWcfQF69llgMazDGyKXDrBsHgKSQqzK+4whQkG1Lm87JHDqS3g+Zhbfl2cWT12Erekp
XvTdMbE0d6RWnpkEGnb0S6d2slwLLM2dJYTx2k3oP3VqHGfOowLSIUXbGIt/B3duASUKjAJk0PuQ
HerdN8FvlSnB55tg6u6IiofTvhNVpinBBblbJp+5Q7X3q3hq/0EIvM2+KBkjSu1Je+U2Wex1MvbV
LVC/lraCaUc5oU4/6oCIMYJu64BhoSIOYcKxr2DDTY0E8ZkmAY6CjeayqyNn52n47rbouQWh+tL0
7qibMknkW7OeSaNm+RfYCps2epUn891UhibW44s+LtZOOvnyhbv5kmGnfj8fI2NXJtXThkZfclGs
8DT3WpRmHAciwPLM9A1lHp2fdFDTRKZZY8wfIcd4JwqvpPgrlGRQoeAbWigyLE2j/UfRE9Mvpquo
G3TAkijGaPiVqcVMayh6aOSgasOiJirpPCjee3lvJr6AfGMh2RoqQGvMG7UNNjauwtRCPlARDeXK
1BIaVsAiZ3mgqixk/ZADRNbBvHDdzh20JyE3GqsgJcWZnOJGaxcn3yFj6Hwq22dujB+VpMTjx8Y9
Nxd+fxniz0mm7olinLqUPh+LftAuk8x1EiTzFPx1nGi1G53phkmAdOUlw2zB2E6GzPCdSH9PETmH
y8p3PxUWUatiOmaVlUy90x3fZ05OvGn3raXUq2nw/it3mqQDACJV/Wua+6M7bbMljOn3FrnTe6xN
w5y384l75zR/VxXyvoAvCN0GHZSEdraBUxKGaBcA4Vyv3ZK4iUD1Aj3EIB/ia4zzD1FkQjzwU7yn
Ps8XC5FkKjn8Yxej96tx6XxnYlrNxDs0R/bXvajC8EJQ+QKIMjfGm0NPFjaYtnYhGHcVFRpGn2zR
MSRuojRkie8IXAjlkB2C228aASo3bzzDT1nOGugK7cJyp75lQi4nGVKRzQt3T9e8GUh+t6ecIl7b
LbPMhCOwYYNajgW66zlB093UMoQ+da6xmh/qum5uDOBu56kcE2We88oL38KscHMN0VyZxS/HBu+k
aZcSya+WQZM84pdiSbzlAbhV8OxSwS67YzhFo7z0cbIDUp35rP/jKazGubVuMKFuxxhb9HO+URKM
+5Atqs+DJiOwIDTKnytxArfr8qhDoZf+1aSdHhrIvUZlHUCItcFbd7ahQWAtuYP+eooOwYvoSc4b
CtKKFvO/cLxAMkIjvADDnaeaXSeKU3QGZt5HOI92bpTYKJpDhg2oZIa5PlxJ9zBLlzC/H5mw7ek9
4EjyCYP2fK7wFUMYaumbFCyABu9BCzPN8HO8t3uxltaEeT2x1udbia20UWtsE33g6ABFXLMOJZnC
45s49v2F2fzd+mfNsxmr6aoI3Fyb7i4xGm8Mm83A7Iu4jbvKJ/ZAlMhrkWCA1hwWPW4OvLjeoIMX
OFTTf2Nb4Kuv6c0LbGe5poLHtECRwZUSSWEuZoAj0A4gSARK8n95+gBOYQngFmdZHepXRt1yo1QF
iUxlMruM98w3ND9FsA9RQ8NCBnx+7BdZGOg/4bwhF6kBIQRIPgJhnN4NR9N6ko5hKD3ITTkSRmpt
qrnhyZlVIc0+m4lw6cxOHVBI6wAZVQhgqycTn7pQvomd8Dpvxlbd4jILBQ7QYrdoFXvx6oaxGiiY
RrVOtT+WXTsMH2c5PkQK5HuuwYxB26uPocP5Taf/Vl4OQhJoMyb0Cwy5YYrY03mgrpPlhBu5oESC
PVqEmTzggElqxRCNnqTeEBoyC80/CV6AXISr8HEjH9KeTwgPNfREqpOjzZw6mdEH5c79q0sSbvSz
vEFwAJWkgr3FTgFtYBlPmBlCsoFY8lHx4s+Vsm011pGJ9qAHCfpYFP1RuP/tqjKn3s/IV9kKRbDi
xFwAKHgLS6r/m1/Y2B8Vp8GblglheC0RFtnVajzm2EIfbfJkEtrluroph09NTMs3LBY+NfLjY06G
Qm2OKt49ylrN9lN94qu7yh/hYy8D33JNZljsmawkmAPC+Rszvr73dqP5Sv1ZS1FYhDQ97R5ek9+V
EXW1LQlnOCF4d5YVPbfr3WjGXUz3gWej3uvx+hom45WcZISmiulRieTSPo9YxT3xwSAoiiYTIDfM
yDs+Wv00IVS12HX8lo0NP/JuUz8e/jpLBz7M/xsPRsMdgoq7SZf8C338hZ5eEVumNWNo6ck7tZS5
Tngujgv/vbQoyVk4M8hrtjjveA/fAD+z8Gk2z5G06nhUOFfvH0dY7bhsEEc2Uftj9fLQW7xVDOy2
KwIKemk4MdGVK6CN01JVSIHeRbHm0JQrXPwHvXya504axw2lA0m0/79du7e7my7B3b9tQZ8Pgf7y
n3UsN29Wn+VE9uWw3j6mWw1LKh4DTNEnxMDwiRajFJ3H0wOe243Wyi0gNCzqW4Emitwrz7m06wEA
UE9RSN5zWZBg8boz9UykhQKdsIhxQKEpFwcHLI287Wqn731f5q2XtcwIQJdSoxfnZCQTR+LcD8+J
oDESbAJ2lu3omWgUcEdjEsMsa/nLXJMXx+gTpUEr6qYbqeJPhTgAZmFAJimFHid42h8pu6jmpiSb
MkLeSUMBZOSTF6QHb9fv9bqARXsBdjlNuV+C6S7S4r1d/idadusIALcpnKFdOw7xS1G4RfU3Y98/
UwDmsISxI8QZNrwsGXSlUQMEF3ZUynfxaXN3M+WPXqrerzWCGtJCIPgJnTzvy9C5Sy6FUFYqJKHZ
mZzLC6qAC3a00xIQlkg//T1uW2QZWcVcaBUcfHGjiQX4ZZxKf0LACJFlclUAiV1nGaSJblmkXOXF
Mbiy2Qj/ikzqyvIUt+N0vn0gkJimo8I035jCwuf9RC3liBBSLZwn4lW98LcNGwKnAC4zefeiHrXo
GEVeySe5J1Q9J4poKmeAcrpRd7EqhRiOpAOCdqww6gHnEXM1gXQTEuOqdqKki6fPvSWl0vMJn+cB
Xn9cG94H74wMmPmxJ+jK8KGfzim+RFSrchpFSODSjSTrkcDObSxcKbE3PeNC9mc/G7WLYWhIBGOn
+kdXiiYYHPcZpX7EqBydwn+XXO8FV05Y6GFMufB0MZgqqUEq7tF282oNiTsXUdw76lmPkl4OQqkF
qAvNyYr5HlmHrqkeGpfZ+pTJSuSMglngwB8cnal31bdhlPAnDHTYW/7aSLb/d0fFB0JWDjaAjOfL
NeYb50OekPhvxvVdkw6J/4bljtPJQVsLyhcaNI6wXHiTxCXdQ2+vEaVpf1l7IsvGH9rneiVtq5V0
HgXV0LYExkayFUYzsvsTWajORA2ApI2Pge8Gvvv0XKpTyiT5hH6qzSVq7C5jo7sEuX93u/Av/NIo
azH58vFjVyyt5ZSikx+Wogm7DYWue9boVIIuVQcqRuqAPR3noANZ/x+gOpAyTfl6H9PsAClm8m2V
zmpr5uDtmaQUClIgHpl8J1DEjf2eEpm7X6DWflUS1G6a3g1buH/SFhNP76sdZdG3dVYlQGh7jCr/
p3SL+OougWEJ/lkzR4ezgXIwSnOqBPYrBsvKiR/zTg/PXZDGJQQlI94ssC3+1kbAFRf1qO31+fep
kU04ioHy/vbn0ixf9oTbJRsKeWoHkugqeItt3OlfcNpbrtjpahrpVPPjZRYPfraezUpnmfHiuHJ2
xHJXCFdcbK0xYs4GoxPm2fbxuJjaFwzd1Czsm4GNMNK+9VXlnnkaCgwrHfb9sUA5rsZTOaQBKcah
XKOBlZegRMsHITEvXlijMIM2BflrZTD9fp3OWZ/DqATQ1Uxv6OcR+TCAliJLRyS4MYbYvgbHVc95
v1ZIjsVDiSi6IQbalOxufNFahIJ9HcgNCVmKc3UIjvrXV2xXygoCvj3Ooh667zqE4gIEiLkCpFin
EpG+rpgRSa76SO4ZiUlA52fqvAI/ogZb8Y4OmL0HMq/n18jnABeZk3X8PPP7a8cIr7TwWOpvYpUn
jJG38Uwj0/TcxDMnZMFuhXO/5qj6v5qgU6P+m2mcQUJsXFrrA/mc1KDWnu9CAJNTDuwEc7XkdRJ/
AusQDxr/9SFl5JXvsZtpz6xbpkVrMU9naMo3IqQCpbvoPipOzwQ1+eu2Qjw6dDZHMfBXyG7es2S6
rp2b8IGsnvZd3KSlMClDZ+wcpFMm942jTxIlYNEKP6zxzQGhRL3gxF+Mmyb6qXobLzspKMC8MJ83
CeYuOmNRKDRL2NhC1zKjLlye4fjs/AyrElHMrlDO8K+F56ddObYSC7etGDskXvmlmplHHecQ5LHl
6ILBBjAqzZOALLXWxm5JVvDmqm13gsUsrA9OsjAZLSEgGp+uCeiJuL106MBflz12jvA4uVbGFiPx
8oNeiKOuqu+xV7L+Cra2uX7kdRZJjKo5LukguWtNaufRjrBje9WgAnzorXAzkJzl63HWI63nz9cw
qIsEScEU25LbKJ/2nY1S9BOB/o/GwWWZRj1XkxPzjaQfl/0IqJHT30k7vxxqCvO8rez/BrYO+UcK
N0ECSszil1qlI0Pcdifd2oQ2DL5F8LWwECcXoos4yMGe4ACa/yA4G1e+l5dT/aLrvNio1BwdJ8DA
0zi+lCiL2IxJAmWakNiNhplyH9CHWMZ3k4Ns1YQMCGcS9Z2s0JWl3J4xBZp/Gta4SkNe1iBhArgH
JOkhNItOOQ4NlIWBJy7GypCq7Wg8JV4a12UmdwofJKsuNObmef722V2+ya52t3X59yaARE3FcLzB
6Ar+1SwHavmLq96QM78Laqe+Z/QQpZuqwsW7wyRfAIbGcvFHYv9Et3TG8QwAkUlJMHAQ/MsyUMQv
wyDdrzK5xdTkKwkanPVcyGDKcVkcziybvEbzdg0zJTsO7xzxY0Fu/m2glBs88zagLvZ+POuTkAR5
un48TYgn2UlNP4iop6VX68AlDaE/8fR0yZ2mG86t0oFDz/iC4vSI7QBw3xDw9A3SWmXjSxgp8CWZ
bqIi6ETEsNgerBIr/TfrlZVzR3g50JlZaFygCUvHcqC9RvTvYi8ZVw00ZJF4hPjps+Trt0rg7Rwx
QnhdNySpgt+jgk3e6m9te2HDbbIrgNhhWOBrl/iGdvvCblfpMCVbeDRMkZh7Qoee9eVkLd5rjMEA
5OdYGfKb73MRDQTdnw8a+GlM0pDD4IDkO4w5ymZ4XM6Ioy/qWr0/LSfWcxoKQDHuXQzMW22fUdF4
bi6sIqU2NIOgqKqatQ3qdXv5SautpGwcs+lwZ1laLrSCqUzr6RfXFCSsLyyjwsCikRtjCFlY7tC4
3GFNG7H3tSLIrJ7F96TV6wn7wVilD/BsVr9zrnmP8lifZzZq/Iq/yelL2QyvZXJvPhtGaZ5bbNn2
7Z0ew3zaeBUMR0d4EN1AZdkcEhNC02cnuMZY9e0yniCjNtV4ZbWD/4DBrEKpU7Msl8wJG2I+mFKV
tSHaOZ+Yq0PaemZ2cw0xiGiU6+olyHMC61PhMIwEHEDEWSEmYI1+sHOXaSKAHnr51Ev/Js/9s6dn
IIH2Z9w1a/eTb+JZZniLGGw22X9aK59Q/4oUa1FVf/BuYMYKf3Oa+d3M/8ORIlzy5V4m1h4mENAo
m8CyMBMkiX8KvtSBeDT7ImDrmdAeOcZidEvDTYdz/5rhUz4bJ+10DD5tALetmhjaaKjV6tbHOhG4
eYpOpwDL37yUBjJ/6tsHxa1MLapOBXXL0l1yFfJP1qIxXVlh7TCUAGv4feQ5tBcNQHsys24xxG8+
eXhiYUTgM7NHPuYAq+O4UY10lhCleCHhavTAbsqJ9LatHiZlrQkwUORZlDcPzdgYm9eabO7KpHOq
Kt62zEQB0t6k9NMTzgC5OUmnCrYSyb5nW2ggEpCvOkJqybqDS+JgpiTSGogzD6W0hxvNATAVjZnF
kr++KsNcxHboBRlKjBMDRIvJd9JWVIdyn2ydMHmAi81/Sp0mCI/R90jBb1+JaYm2EoZn6k8wvRLA
sAuWugO9r+mSkiLn3yeQFpB/Suvi8w1O5RGVkBVnjVmQDt0SEZiurORw9eWow5fFC23m43VBeN5M
ndPlmvH/H8pCiD9y6Oq+dre5gdlkNfiMNJhVHvIaxyn3mGmddYXlPZtv4r1+rDTHOG64GOZoQsN+
fz9BkXkKLQP9rYYFUhey8dotoaE7zyRbQ4D82PAOKR6z/KuZGgu1JKOUyUeqoefJEj+04fTz5gjD
WRsIxCRAMd4Gd5p7LBWF0AYUTPbCCb/MXfxXYsNR7hrJmYDcm5zNBbTxG5icYEkolxIC8H4MMwGV
+w1ipTEsdoJ7OxtAjZPlOnpsk6V/lQ+BNKxcdSFhKEpfSlyLJ0nPJOcXAcp8qkmGyo8mrPT6oWaK
frEZ796qM/9cub9i+9EcKnvZid03O0estCiqtjfK1RJ3+yHUrRRGByYkH0WXodhQ5/vTwZ7/FYwd
7ngsS6RULBBpMsLZfPAa4CwFF2DsirD8Syos3eqPYYYmCDehv7Fl9GMLjq+khBtZjUxywQDi6qQ4
e7iAF5vZc12NYn9GQyV4769F6DYxJJMqYNJxFnpeJD3A0QE9o8MRn7DLTIuNb97zsKMjkyGx8Zbh
tcia2dzjqrPfaJaU/ZFg9RfRI4RmOCBQxQ+wNzT3biGrO8K3F+Gu4NSablMGcgJQHr855VpeSNsH
xs+Wfojr1SWt4aqcX5MikFBfzXwjdaVN9TB+EL9qzcynvTNbP5kbtLlk4bs787GTkUexZGLHA8jp
qFXnD1Gk9X8i2ecmSMK10UTBaBuYtzOmAsV56ByMzzk0OG+lhWCVNU6KHv8GIQrl7hxKHP1B3t7m
ugUxb2Z6jfvWi0BYzRfQ4wk3JfdrhZpmCAkuajcG4p6wh5+XuSrieVcuf2Io4/FUd60EqfqWr+rf
c1k/Cf3y3maxx5icAgfPE+ddq71GQsngrV/wXJQa3vL847agVPxPN+fzRuZcaYGi9h2kIHfM3l6M
+9lUqxX9MmMwQxTpSLdIaLHzw/xEGd8AhTFECEPRYGL71inlpypZZ5xWp3NhAvIl6ozwaly3uX16
gaBo0HymR5H7y0YmDsTbzGYWpV9vs0hQSLEZRckBjgVncHm8SvgZ5O+tvUj0DQks/g3NZvqh5nKj
17zJOd11tuIgGo4DYUDy7/o7rFeLqHgLT2oS1l6pJsr0SaELQiG/zkJVh5NjAgi+pogUeeSbJvCk
XrvrIxezMZ5JAtU0/rxooAbksLRqCedQyjqU5NCSAqs6y0thk82XlKMjy4ZyqR/B9ZeQj1f7UXxc
Iiu99DOreTGzKzjGvExib8WydWxWZtFYlGScaV/a6MjUgiEWyQerC5nhkj8ky5oGHIfxtq2+vaHL
lWxvuhya0M6BGjeOKttBdozqPckMPNJIZmSioeU1w5r3gIbz5eIW1UA66nP5zYIYoyAXzVh7hdXn
EiSQQaXEziEdp5X3TNvwZbg2Ngb7NgOTqZRYnewCqwC6ccwzYPbayaSuE+9zYTBPK3rDgF4dplkC
7HGctDRg8SC9Q6DGWp3/DaJoAz0IpEAyfprIQ9Qq/za0fiDobtVt0RKMOGB+//ubQwe/Vvi4z1Z/
pySXqslkaufhLyuikPp/icyhsZhiMdosEGfh0reUUYH0/R+62pQjt6ME7oTwm1fgvkfZmaQAa6G6
jBKEOxmylbmiGfnx/UCVzqZrkczneSv5SNan3YBCnUw4tLshUyzIr7c5qkGmGTvJ3dH6v17Q5JE0
v14T89/6LtQw5SrtBlP+0FWsl79F+Nalvvqf77jRkePD3ON85/KGTyM/Q0gnCAHQtWskmTmCvwQE
fLLIoi+H6Vc6xlKqJje4kq/+ohyM0kEOXJDyPsDwX6RXQC71ZeO782SGvC9Ydsi+ph93tgZ9rU9J
t+97XDCrNvobbK3RXjap+2dGtRvFgSW3mcpG+I+amA3IJeHFJvWI74zjsnp2ZcBy/7me4pRInCGU
5zDQjo889a5U1sQwrhzq/ufPP3ZHiO++g+B0xrHHSU6hS7feHIeMUfTJxIzSmQbfLvUE2c8j4UlJ
DrV2vMdoeS3d9/unvnjHiqhQ2jfNPiVTgKzlx2fzvjafB1HHwhsdAsWnw+rUgewmNkIzW8IBh1IL
2Y3ffO5+lC2Wi36YAP63huBBESG0qhVJsX3j9cC7EuwE7fmmkEESMyauaZiFI861+AbuLlZuJdLA
eBfJ0pjUSTm2fRSP9C2QbGxb53tWVgMeqcu0rJ3bkLLYw5dIb1XP8TEHcoJP/Icb6VP6vOycr3m5
Ca7Rxg1m7cygr8h8tpr26k+NGM3ANd0CubW8TrO+tunNv828F98l5W11B6Rpn3GUI7nDEN2aWv4N
AVEptRBhn5NX5YvB+vkP2JDvY0eAcDVQMMy4K4AztUi9zQc49T8wvmDgTyByBZSp+RVf4tIyb3yi
XFUamIC6HmGvIDv7JMW/UAzP5ivsxuhCf3NLUhWdf4in0awlPkmhgOJnKrj0Y0081Vr1ZBBVaL6T
r9Najt7OiP2tKQdoPbZ7KoHZpNf0nS05+9XnvaQuDtw6AiE2q1Q78c4EfHA7WQEHqSry05Bt6/r5
h/SVcn+n+J3RMJpw8mZayBEqGzuTBwpOerRS+u0q/UiiA5ms2qqFfNeHJQM53K3Bn81hHCtfuRA4
777QqwdYnUt/Q0wYzdc0NyN6wOyBuypl5/qoef/Tu4B/KL+JPKi5NjCBHVnbTSeTHBRYHFXuvwKh
d60/LiEOeZqX1O4S5N1PG6wSFTYUz+c2a6wFu2emumTOGdAZN8OpABqABQngcHyn57qgxuNDmeOh
b7+QP77K/ueh52zivFMxYBR86XlZhZnPRf9NozTgTHaEpRTD8cx7BmfEshF1CGULfq5NFcOVEicL
i+LXOBJGqo4d5BsZM71EnIhYCbFYeTwMm6cqX4s3DxZgf0n+ikrFm70WhCqJJ1gVdq942KRdXY4R
0c/W+fSJJ/FFJkSYRikVlLKcu7l8aCeq8Dy8fGxeeGjoV3wVtxWUxCxedfY8iQ8YuOZ7zwqB30Vp
sRmRQqRs2asMX5T1SjQ0ttHez9jfY8p8rGvmJhmTOk3xQ35VTXCrdwCEC9+f1+3BoouPsOEotZj6
xXDSxZ7JPkTQcjig97FwxGrdC6o44LPGJKHtGjRlEMtAYDb92d/j+W3Vj/WfEmgXSBl1YC3IgsBw
fuM7ylYVfo7gvdgoBnjRARSZzbnPAQkhinhIvFYq3pjlyMWrWTo9zy6ldZkX36NRj+Mte5wbXrOC
5JodRxJRiovnKyhXiQnCWmmBf2DoflZJupEAfM3VIrOdIbP84oxOmRyM5K4CH+qIl7B46StR0tS+
6+2BJ+tW/t7jA8JlH/UI9vT2k6DhorvQt2jJIuE4AP7BlRpF4nYaXnVP7FljOephYqR2LS3cl5by
3/1BWfE3PLJcezmz9PCPZc1SC07NoR2jA2rrvoNPUyhcPfgw4/DPmw9W/ANVsWyuO739GIepq6n5
jAwHAg+/IFCA2BJnGyKFkUJMV2i8ds9J6Lxf9oSo4jTtXret7TX/x4Nuc2q00+/nlU58OjDJW+Mj
jhmhBha8Y5sgO7cLeceaFL8W2iDY1D23TNYsuvto7cnrbPGCrxkCxSn2C+CAYqfF2yfgsbDeF1ne
4RVpcTDZHC1MlDRzZng1jKqzYB+mOEPDLDD0yCljK4uE2K8X6cnbmmr7a9eRPgyVja932yv6cb7F
HO66ziiPkaEjbYpgCd2vB3jCoG4CAFGst+huBQWk7NHaOIp+zxAhifCIZgreuC09aujw9L6vIGxP
8GzEy48I9walwD2HidpXyJhrFJkMeCbnB+NPdJIXT5shDASZBli1RvFN1VQ/JfyRdB7BiFCrPS+C
ksFzUoIsWiI0vX0V6/geP+cz9ItnRvyRBXkhUoHkq4iXtcHV6pI8GFQ1gCJWZVARF1HNi+jqrdtH
mU023cjhnrR3/pOtIDqO0SvFf0hPtFSHWImTO/9L7qEjAzfJIDkgA8GqePnRO7DRHp26NK8UVA6R
wVdkVHOuWWAQU4fwy5neJECLETblMiIDhCaqC4tJD1Yk0qEsWAsbXADyuUpSPVWcEqy5LXRkA0xa
ea4O+gj+hwamE0piWGsoYS56wf9AcBUXrka4oMpmLNVU5zSsJsP+L2vpuD4phmaIH9AfRZwhvruf
GWjs76Ix7E7SXyiXka8E6bhrVPCBWaUomnivyiog87KXZvlFTOVgph63ebeGxmYDiEmBUA0p7DEl
/NJvCIIKBihnYUMW2ar31RB1M3cVdy7IHine3oV3WClWKvB/ZUXIt4bxcyxVN1h91NLFsscDl2F8
yMARUS5/X4ODn0wwWS71/8s0q0GMvJHC9in8Kzok+PiCwIFX2tcK2VjZJRsgqxfPs4SxvqyaYH+b
H+BrPf19UXXzxweYIUiQVinz+bXRq4MfTPkOKpkwGlJ1LlCSmOPjQMCujlqct18UItBWYzAznNSz
RrmSt37E6XxbMPXQIEh0gpV99ul/cSj76urTHZ8o2Mq6QQpfZJE/q3De3p86+Z+bsqS1b4SlfM7f
5vAtJr+Zd0YawayCwMVB+sbQX2f9QdwX7hocVPh2LtnEG7rxUqfAqEWe7iImWoIGcXAM0UJu9nc6
OuC9heVahpeff+r58HEZjkfkZ1+iR6uBQqS3kWfeEdmoTZmZO+pjNqaFZOJ7iQDeer2ucT2JXoFn
paG2DeU75HFB5afI/d7P8HSi+/56MdbubypO2P7GBCFj1uCSpEQbTOQZvtc/PPP1erKCPswp4BbO
63HP1cKORzXhbbgqXsjjmWW1qGEiVUY24nzrJy/2qWWMMDKwK1NPPmgoVrrrjB7YkjvBwu5xFI1G
gEON1GB64/A+PsC25dzjWZEGVz0zOV6tyvqxhFKry7Tr+w/DbzCegOikjC/NdTCGMZBpwf0xKEpn
RV8nd9D7/EyGsRPszLbMy558qOpxpr5kZmAN8Bi0sGwZRjw1qGiiiBVyLVHsMl70SIH9GlSiufwz
HxIORJGnoOm5MW+/jpjmCuwKYUSh2jg+f0NT28N7ryC6nCI31TfnDL2wQ6hDH78vP7UWmzWzf82p
XSWx+WnS0ErijRSwQKN4RRJs+BQjllARsa0ve+ND4DtV6C1SZWl1rj7ZD1QSf0pee4/2sd+9BR1w
1pBovBav/9wHPJAFwqI7wTjzUDyGveo4uUffllSvQrwMRSY5yd0vaoWUhZEghI5FSNIDuorut+k6
cE4aPud5FRMfcqlKIpMJkEd/ySirdWzz7IyD5k6s/DZAZDS1UMZvmEfzUvANsNI7CMsEvTNgwf32
gUVybR7Oo2J1SqKHWKDJO+VQQHpmFN6eLrgAZWG3aXg+x1PHWs0UYhXoHYeVeWJLE9qWIUN9panM
aeSPccFKoUE5/aKiF5cgaXJZzdMVsAxbBfgczTrvHAReqrZO72Ltvwamiv4VuGT9ndUfGvpUV9tT
2Hwpp/6T1mOm1l0z3Dx+Ifi+WXsSdvQiXaR4Zte4GjnMfpnwsZp/2GWVxnlyA0NwPC5U4+1TbKHO
edBfXc+BR8D3d81TPoF3+Hz+rw1jt2aQWszPneQT2exTDnsV+5KusHpU5m54V0A7LyYRUHTc6wcT
CYBZrlr/TU/gQqKnlhDIVWW6l/JUdMs9Nbuu3CWBgI9Pc4KRgQh8w97/okj9s642qOzE5tVMy2NH
3xsrpM/lfjLkrIizE7EJ1lKop5ONQsRumuOAN53jd9uZJTxWJgtNWg2sHynNiNbK/ECWApABvd4E
J8q992/sMZfydxwCCXqlUhsAhgWBPjskqcYaNJoE9J/8GIq+DtW0k/5kpPZrf5iCRTgw5g4u1033
2EFvyYqBjpT9f3aMoPE7nhXfbooy1+Nug7cSrBdgYUuICTtAR79Q7DVpH9fQJSfCv7//XxcIviO1
oGMbj3N0PxbbmsjwbNR2cQ4ZalxQ+j0P03KQU9Ibmzz87XeIIdd58ElPt/9xbim27C3panPJ18wx
0ZDdGbbkstSESSEEI9iQ2C2nZyrTnLt0jkMc0mFZrMEGIVQ3PAI9cOdik0qMC3CDSbbjmPRER5ca
ixZeJlgqVR8oayH3GaZXA1CGfr2dvRbV+ET22UhLnx3ZOHh+dKyH3PXQgQU8AiuNz/lXG/A9TMIW
JRTHmcfJ0gs7/Su1hVu8LMa/eagsUEn5q+OpMopVWi9BFvvEzI6FVBgepPMaVck7oHcz0y++MXkn
nsjmcqBW7jXCvNAgNtaqgY9wqw5OBCRa6LuJ2UXcgjC4AfLoiertbRmNtiMOvTJKxEMWKrb2iNWq
IDe1a9nhSipCxvxjbAAqg+XYhV3xIoCkh7j5wKMg7twUsZKD+/aS2T5cgyRox8uMcrr392VgwixE
/WznE3RNg2LNHdQQcz666hJ+P/Sz3MJk1uuT5I8cD88HOOuRLYhvZY3qjBhX42DiTWPE6EFacZQr
oCOUqR9+yKuLbwqmbXASk7csesNwhJtobQOyC6dk51zBjt08Cc5F5gISMmoWGSjNP4PrAbvLnARe
QzEfL4U9CMrVC62KpusyIMTg4AStlQo/0PGMWSM0CECZ6rKhIWJ46dctEb6PgjnLWLi+PaBo4/Ra
+eFpQt2OwRCKURXkRpiwbCstPqhY9hThrcoTSFhgeBckro9L/kXo3DKpSkYc0IW0iOUdRt/gK5VA
OqByZlHha8RmR78JgmKqj3SLug/sYjkC5YyaQmAOrDGrnMjCdW22UvJYKwAGK4dVIO9c0a/9TrrP
BlgOlD/fiYaku3CJIm++PckZpMk681x/KZoWwj6+HMmolLEusnBgN28nnsSuqVLuf1KxE2exPPS+
q2tAPU+Wb36MiBLZLXBqoa7h9oJW8jwxq+XGYUuuCiH8Pzmtm7GoMeJ3z5zuKHwzhra5sg902319
yy3MKwIt9ALic0Esp/PWFVZ69oDubx9A8cxUqtOi6I1Mw9alt/DBLEvpnSfRDrVpEv3axYVrtkgx
+I74DdpPIrDwWqtRJoBjkPpogWWHJ2pxPlt30PCKNwyCVEERmsqZC2BzAE8tjBcqcvgXU33UwpEA
Hrvzn6yt7U2z15L6F0/9MOMHPJ9/kL6NgGNDXuV/BVbQUww451RY2VlZajL6Fj5pETO6Vmm3ZR5i
N5FTLN7KP1soLy/Ph4DXPFt7Rk3zeo6aHFuonOUyN4n5220uketlpr/5ycH/j2T+uKOxbCpB5/Gk
RKbAhZOHnP+XhhnWHb8JtTxOZCVmTKZV1zV6ibW3GL8EoUVLuVJX5qe/hVmk4b0pXWtz5OXMEPsk
AdV2LE/F5tP/M8RhM3J+TNb6h+nxGovhs231C1LD0O0PK45hBR3ufmWaOSGvUgcsxI4gP2iqRjSr
HkmsKdUgNKAS7nMC7PvKfaeyq4RAbQYH8nm4gNWFbXtxGQKcJYpBPFlofd5UMNHyuiVdS6kJrTQ4
5ghpnSpY2sJrVm54guGY0+lbc/ezLw3RyLD03zBdt1mpWbLcROAY74s/tIaYESUXYS19QO8c+R4j
VK7THYgWYBAb4qNKvE7izBd4NoKWZdlho7Cr1JlnyDo/Pd++g0GSy5285E3yIgzgRNV3XCqlUxk5
MM67NjR9f1kAgKlLUikQsIE9d8eCMYj63H58ahxOp8F6OPvi4NG+oovaeCThu4+D24odMphBvB+I
EA0Uz/zmV3LV5jvCVR4mdFLhYVQ7yg73qapixV7Uk9i5n8PBSTC52z4xPbf67nz0KDthH0FBENvo
9hnpKafHkQZXMiouqcIzt3fPX/BCzcq3DICzyb9U+EyQklU4Eip5TjorwXlKmKtI81j8pVu3gQTJ
2r5npvDty01yZV9I7MU6QJrUxf1Lq89ZEI9WvPlE71vWHmRAwUTGyy5N7K4nHGLOEMF5PrP/u4dQ
YT11YnTzquWIy/IH96Vuex1D2g7EDc7uUxFmXe8VE/oQLaWJEAJZgFYnLnBMZ00FtgiGjbjW4B1H
Jcnz+7Bg/+YuYux0j1kMZIo/4tR1LKMLXEkiEHQdBQMTSeUFH9AgmkMy5w5D20w61qQqe4ZO7e9R
6o5bMGnnJsEANU4VPleRmRSlU9Rgahu3GW1ywhfqDO494DtSSXdP+Qjlya2vxgUHZnGoNS05muNH
IfzXJMbzRdQhc0kWE7TwhLC3hRAAUjXkTYQhyAZrh2bBA4i8jotC4f2foySlttghXaTUl36dFJFg
A1hxVjbZ0mj94Mvbe08/XPL7gpgIpygqwpXJzydpD/FLFunfLT+MNxz5xgZKH0q8syzzQM+jIjCE
6tThpi9rw2fggmL7T2aUnUPEB24TKknlRrtR56sMG5W+MOAU7G+VOMKy3aWu7gLl4JURR4x/xZad
mk7akmUbpVeKxQ/bITWBkKF5uWvEF57a/jwEGcCqthVKxkr9UYVMOJ6pDZpaYojQJ/fy6UGKaktd
Mx889E1tAAk/nK+IHZjcMh4SDaeyZBael7YANfZH16rFfIirCR65weS9OHHWvHOa7Vvl88sMwNxA
zexCpIvEmuGD++xJnb3bFhRqZREDj9JHX7r9BZFstfDtOm/FjPpFENXqrWA7jm6iMSUFs1ziKB7m
C308f2J8JjJCYvydM8xWQQMEn7xnf5zpWsCTs8Iha9NDsn4sNojovx1wtZqKlVwbrEkVdvgm5yTd
ve4lqPmT4SaWi4Ol2vWrc/5bqf0VDLKbozUADavJXThYi6+LCTWe6plocHGh1h3SuVYI+OxRsP5y
kR/fdNKB7pCtRbEbWhac4P8o/+yHqSFW3iSOSWhuSV0iCCRk4Cz3Zdrw+OhggJEsapO4mS0MyZa1
oNpiYuJPcRgiUI0PSmsXTnkCIbSydFMyabN3QRa440/R2MEavbaBdfQCMeuXB/U45BJj7GPhrFQF
2Tyi0Q0iifhegBld2RPku+BHhmKzAfYpU8AMshWqbuPV6w+A8XNj12ymm6GFTRFqXbcOdwucozbj
+cmQk+SVO7cIdmARy+JMFAKJi9PnUaD9asoVVBYx8GI8RJVAfoHY96Z9wLooFxrH0x0rvG+t62D4
3iHeCT1NGnmaR1eBOdqrnue+IVhAC0aqNrZrmPP2EzjYlTj8fYGo0bnbH/HjCgI=
`protect end_protected
