`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
Igu8oUvzB6WRll4O6LEbRV5y2/yFbln8yOgEAgldp0eCxbuQkiZzgWwEXvdj+HFX4ZM+uK+O137I
xQ5hR7GeJmSbxicDXkhPMUgnHeYPVRQEUqhWmved2BHtPcfBJJNYx1OrWYBJEkfIp1fC70EcLcvR
6UK3XezFBMQCrqCNpzwlSghTxQATYKqcHqjuIFMvu+9Fz6gCPNAPb7JpjuiBIaJqupa/hLLorJCq
btnzHrsnVmvdPfecyz5GMu2m1h1e6BrkBd3gaJuGLVFhNWTIyWglqvaMd7zk2mmVQKRvqqTkyGDW
TKwo+8NciKfkAeATAMhCex80HqLbtoI3ZW3LUkvkdjlb856uNFr+mj2KT1bPp0VEx0Tf22fA2Q1n
bNPRzjvYuB+4UkMY/6sEiuwBfwkd/IY0xs/5ZLQMu3ttIQ5PSvMY8weFG8BVNBE/JT3MJCHyi/DW
WPssyX2kPl9alFpY0IL0j8yyjdxpVU+7NbJIqHjMVLg4vgAsefbzkZwR+Y9XtGbvMiwGG7KvcrY4
ODy5M63IQJEx+VX7NLopKnvYblwz7fjPnlttTFTzDvs/RZ9eJfraESa5dQE3HzmFIm4TFxkxDQQZ
2wu146E1I1xlVHDGCDm1xC/Aedod9GNUXRGQWPW8spsuFeosngUUqv254/nNziKIEHNBPuOlieeN
id49enM4VAv8Pi3Vx6nwfzbd0MC0omwQRjCG+AHGU8AhmnONQ+eyhomAm4TKMWePtXHQdYdQs7TR
TrH/KNrS5wbZCS5uqgJaQdwvpssBj2v1uM13crZQBlqAO9EV2jN7Ml2VpZxjit+x57NZqabg0qcI
9ppMXpfIQ4/uMoG1XfmokpbqZqjaqJThUFqMQFjCxk9oCat55MBnHRssBq9LTQkqlyFHrl4tG9WI
Kw3eIMo4i7kXRibLWVGGKrVYA7o4Zx4xOab6w1lAEDcP5G8N8LHCrln32zGsWtnwJUmEGg8mxLz/
Suvoa3sLHPVz4zfhUOmpaMZBt/VxJfuT2Ot2tJSE6LIx7+gPOoDp63jMo3T55EO+bJfvGuTuYIfj
O/zYVrnELng4rPYv5XQKz4zwd8QeX6brppWGVXwrPwAQyVT0XXbd0/t1obFkZtX/zx+gXgkHpzT3
8FZFEmw7W+Q5KVIxE2CZGlIwB/Yn7WHbdmci6WWQT5MoXR94kam+PQfJDcboQlEQXGWOoXmBUE7D
6KLTmPfwVN64oxZNwxH6ax6hbcW6HmKU+ic1yEzILZ+hfdN6urVEhHTL1+GiF9lVO+i6rxGeRH4g
ks/ECpN8nQv6iS5RAnf1mzj4TJGwq0H6DS6Jc40bkPH6hsdgwvWSD3gxVkv90vyTFtsNhOMCf1+8
1uan3HQ9mcvRkQKCnraCPq2Ypv0t0g450n6Xf//IzT3gScDlXWyW6VvZ3Nt8aV5Dff0YsyxKQPQ3
emQb7A8B9midcvHrt4glFoXWp5chJK6G0glwsATANL3oUh1QZdGeMVSokp5n7U8aOLbZMpG0Zg16
Gu0g3Q+hUUEq907btOQwsxpurz5O/bBg8zXOPKhU5HR0+d32QHvuFWirArQQdw7UzApiDryV47TW
OiczW7F2RGK7srBX5KGB66BxQje7Utc/DYfz7fR9oeBaE8Ep27P3+l64JMHip8/vNbRwXrduXiM5
QnhOHB9azsc6wiy3vIgMdx+L5DNSQdfcSitwvk77E9mUb1KwZVjkQ+V5nyvBEzRw1zEVqrpBpZfh
X1A1FXWNJAQxevL/iUO7U/WGuGgsE858JanoVFwEen8VQD//DLfV/LEQBFzCS3TlD58K5SOCicMC
vpvd3I3/yXEaeMMQ0WrRskB9XGARMyKmQYsTJIa84psk7tRgH9UAggd6xcQWN91jpOCbFzoKoY6C
8rlgLx8GRzdkZm4te2jW8Sw3pNsw7Q6sj7qQNE2yV1YbNZJWVa3ZZuV+emQsYmQcTTKjKxqSQ9GS
bOpKBbbWZP11tgxj1mFiSFwxuUeYFrzelPqhEah3jl9bjA/X1phhXzm90oIU0DZng+1EeL/D9a2e
X3jJdf/uUfS8zse26uUw4KLhgMYyLUE4y8wTVkY/utelAz/yMui6gGYGWQEqV++DYu3XgSRyYe5k
+EXcHngo2jauC2m52DMaDPLnp89XuigCEHMwzXaxTvL+0ZlwG+vPILk15EvKH0gFxbf6IApJW4j5
PPHAaZ03Svwiuny1yD9o6SoenkKPszCwxeOmtbkIjyiHSoblzwuAhIuZIasVphdlV1PkH3KcU2Xf
guTsJKmgJQABbZove8gYG0xOqH1lzH+MOXlR6I4KU1TrV80/uCbMVyrfNP/wnJnE5nB2kBV4i8Gk
LubasleF2EkB3gHXKM1w29tlO6qT/QiEwJf8ioxecCu7AGmRDy+KuVb3Xajdmpsts1fnJRjqo/Ix
f5ILYhDdTiX8tvrmyro3LLZgzZ4zppn4q1BrjOhmqYGU0JVK2qgG4z/mbbheQ3sOl8w/eFWU6TO/
htrBzeQWjj3MG0cbAsZIf9CwJDii+iHSHufJeEfDtx3IkCXwIW9ASkf/bZuOUKs78Tqsbqubkvjc
OVniuFzbCedcmpIKlF2wczQHBt6aC2SU+NBx1KZDfLF+P6Gx8drQmfTRu3Axf+63oSsEZzHyhQp4
AszaGO4MckYz72GlaENsdkQ74ckielkUQt+16qTJiTi2mx6BtquwhygNsMR8bYjQojvgYDGALHJ0
3QlJTnKzA0WzUtxpcNQEjq/gc6aNcsbNarcu9TF+wZBM/LOBLc/M7dMUSvMkdudhnyCpfe33qmPe
HrWnT3oAm95hZnQb7AmA+TQOPRWdzRFzHMjvTCBu6qbQ58gW/LhI5gvG9dVq7vNr3rqPmUx3BFIb
/nBwlK6ZkjBfmxCyVFN6S+JH298IVS8w+TRv4oA6MiT3FCwKQLA0SiJtbKZ61pmAt/g2x3o9bhCc
FCM8+G9ir1O1qNztLJXp1/WdaHT902WBb32U0q3EqtCikGTzOkOH9DAWzkGqjRhfJWn2EqWdQfi4
kGt9tSe/TH4fwOPHn/Ku2o9YwcIFQLNm8455KMf2qeyb0NeAWVPIbMHMN6Q/8hnU/fzE6cmGq82g
HSEIK7Go86OtRviIT+VFUG6HAQFyrWSBhzNYKkq0RT5AO0D3lXc+8IfBeCutVdIHrGvGfSUa/NQz
8MgqgnMf0PFyI/fUdeHAJCjRY0iV1++/HfOyDa2aRiEfu9UC2T2QVxUSTzuN1Aay2h4I7jQyNC/M
knm/OytCaRMXow5U96p0FRVINFiZzp4orqx1bvltEeRNaFHsS0fmEuMKV/Sn5n+KdF7mlSMQ4DHC
sNe4/bNScom07WG4tmzlmuN2UN6sTsz9AGX7pa23WhJZl0Y2V7D+y90n6dq5MdOh7XG8qu5bWqKe
MDCbNDePmNXyIJlJuozEobTmwSc8fLQdTe0JUB9t1ChArMzfImtb9HbYDWg20HUP8XBPy22/ioF9
wDJHwAR2MGmV6jhCNJxlirilkiJhkVtHpg74gt+tEB+Wok1004rIqtTTO9raLplcYutQAyA/A1Rp
wqTRZywuyYk2ccrfTLsZmBN5Hcex9nyXRm24VhWZpPfw/ohEI4i3nswnbU4mDjjl1uDidyCMLf6p
KgiDH3IR7FPwm/U2tLDOBISdIosVonulwTKFZGaPc0GPUrCWSzXyshbZAoKJbeoZ+GWASt+UzBzf
qYENNWZmMrAo6+wq04L+N1ZxkmkGdM+dpdlK3lb1LGAX55GeHFS/3zTQLeAeeNDgmGKsCBtrdiaW
cfQ9P8SVeMqSRZe35KwmLGHaCPBOTgYwrPZNycS4RuPK6bxsoLTOaD1ol1XLCm+2r+vHxqh+EQQb
bu5Wo387cCQAYw1nC+W+5yjxoUbhGpZ78kwI2E742CSyOnsrNG9hVJgkRL2+H3Aiax4JoDl140yp
hNCozXZ9Le7/XXEmeQMMcY2lEJUDhcGXmDZWAXoak3rIJs36hQOjihP5ZL2QEGbogrL3bVja3rnW
OSQrWSGQg2igAjikAqNshH79ZiZBjtVMHuKn/TQDr7XoXPx5itvkVylV5Oonhe/mjIAvSBfjSoWs
uAxeAPLgLL2/qymWxBzml+0j5bBsvdA0I0kiqEe6iCGED+jWIWyLtbGiSa6P2Q8WX3ICpFUdEQeJ
SIe5yF6MjxiCakeZnQKcnGETBLL3z7Vsz3TE6ZiF1RHebzgoHVxk63SeAk8O5zcO/aEyst9MovJV
aJan5ILrkty5lPkeXwTfkaMKMb0aS7tWME4YVhslk2zsTLA2/6rhUJ6wHnkC3YOm32DImErH4ITc
7teqBPt3BpAPpACXsJm/TjEK4T2el3++u2Md5e19Hd5uGu3Q7h3LiLgp0wrBzBGaaLUFWoIZ9pkx
U+lwEZX3qCqeiD/U9UDDCRTTRFWZv2us8DOoEYfkjEG4FOt464ve93qpLvHE6NdBPF4M5dplSuK8
czgpJf8QdsXjhCtU1DVPQZE22oIsDHGQINN14FO0Lk6po/HsJDsNo2VCdC1wcFSWPCtWVPJPSs3I
Wl23C9JxK++NQotij0nZpZQv3DYMWxDCmc9sJNjHXItit0KHCxWXyXevSnxWE/MCpr66Gen/7x2/
HEcP+hzNm12adqnO5mZsIjOB+jJjdkPQZZBeB+uyAd5cDA6/RUtxwFe2L4anWh8pfkmiFCSBA3W5
3eFaeA25+MLg50lBucx4Mob4aRNW+MEBLG9y5YRv1zaZxPXenv1X+47sDFkM9ZVJRf7fF+MaPPeG
4A+q2G9+7gxZ5l6kzRZXlYeCKiqHaY0twnY+UH/FV3OHG5cmBeMwGilODBbbt7QzdXZyW4QuBzvu
VDdT+IdfvPonV9yvJ9H8v8IN+0GugYj/sqpZ4tj0vAva+nz7LX2/aqNR9jMNAYWSzqyGmrZxPPlw
9nDltQllIGV4l2JweI4NjOhqC6lmZqf6oT5aruN0HI0YvOziQyP2y2o9s2eSelZYDVEiqNJFMsqP
zW1Zgg9mvL7Rhty9df8xAMDdlZKNrYsqPqKUoEuLyG/2xj//qKxcPXUu2DvQGFy/7cuyUbe889rE
egwswUpKo+Nj+RHeKWdo4GhCsBvQuVoWGjyhkHNbguiKMhUUDr/nvqyjSTwZVoN6aDzhUX6JHK5w
kHWi9oKENiyj8OnjZxqxn+lUp8X/JysWoZDGUI3xoVeazVf8ONJWhYh/BN2VzakKuQF9Mcn1R6T6
wRmbd5TJhpkpM1JfdYqQBxaj4DwP6Zy1OQ9g30ooNc034obpZjH9tLC/3QWfQMZ3W1x7OK/Onnv7
eBJtLhvDP7oGXI16iDTxDbdy/AlvKBiM/PxydYaTPDAq57z6qKbMXGQMBUNKCK3ciHApONEMIcjy
Q0xoJPzYBJ8c4EqToTlhMjsDlrC5WtoFVoTT3+mjaoeW0rHx7+8EosozTlUZSds5cOx3SJIFVfOD
HxqY6XO2w3KXuDxA8fEtRHt3U7+OymrAodB/w4pp8Rk3EeQD9PRzTTGWyHpB6Ww9EamT6AGhnvNN
+c2xNvCZTeOstxLnjoTlyyJWqRs/9jVRZn7WhyiofXweWgQil3YRIJRlJdKHciyd7kJYbcbgVziH
jEYZqUNVk3IfgW+NtMYqCBLyAZsFRms/ENi1Pk+HH9oeBSAH9zxbLdarhtAra0fRG3L6uzPX3FuA
U28wmarrpNC48sg5zaKOX+z2oHy8/gQnD5nRxer87f+h1lvsPM7Jc3lwdaLHuvmGudgQ1Nor2qiE
Fkd8gRqJkG2ZAfbtM1+Gn23nyv75ZhIW6+3Guei1eRAI5r0h+0DNEKcFAlAiXXkBROZXHOioLlUw
m0Z2ToExtspp20z+IR2zNw2N23vN14tBCMCvEtwYZ/jGcgL2CtGSkQ166JEUaU44i8gvV6m0k+04
WJOPNz3n+LyWKCQcxo76J0aBX2WtOw5CKV3Pl7mlWO7MuBUVhdAlrGRxeaR71seIE19Q2HmB/6MN
sj4GNT1epRuSsExw+05Cl1BepAAPUOz0aKh0T+V7W1S+xDWPCqENNXyUN8geFchHE53NP+gz1dj0
3VfYvpN+jbLNyuL/v4fewJKnFVpySpS2j6kCA7qGuBJUhDYQZwyBm+o5LdmSqIhn32sSS8VgjDrk
k3Kw9Dx07sUEHSYokIS9tSqHPZsU9GO2LtZO2oUpXZDTaRgxXEbzv2FnCPbPLv/3eu7Af9ttYCNs
6gGH2SoZegC+Ul71GRSfYO/07JXWygjDuXxzyN4VRHm/BMBl9Ql9cTyZ4oTPhfJHmFfqwDXUxRxn
o5ixpyOou7/KVfECmpU0WSw3oWYL5KaQZafx3jLNA6fmrZJ9QCcP1m6iYxAXE419QhSTn+TSl4xX
TIfcg8p+oEXshstgS9mTqZ3Xf5JX3SMb8NZ12wGknw0J1LdsJTTStVm3fakZomHLCkhGMpXArjnx
Zy7LXttiYOLvRjTqQOBmlt/iPrOAoQyZb/bGtpPA8GMoW0AtreYrGpBEZD91jVM0RsRWrP6ibWSs
C0DFg+4pjG8AYRUON+XY7JPF+bB0/6+qpGP1dNWMCR4A1TOdgEX2ubDNg/1LIyV0ri8tNoTz69HC
dmUU2K4pKwNSE5QEDocFwMEKKVXCISagrQ2c7I6PosXl+CmUvG+R6eM+/nL1TSTKCOx+9q/Frdn/
F4JpIcwVuRBcnvaZoduKnUfmJT6t2txrycSK2W18vM4/yio1VtQjyuxFXMyLoddFMNqwMGBzOk2B
ISx7f1djHkbAH+D69clmtkracdni9Fu4y6ApnTrXmDc4wtt4MdoJAVrgLG9Bc6eGr61pNNTU5p5q
DWYSGo4pvdveLABDGh+52M4aDcg7f/M+xtCImrzh222ZlTrlxVd/hpd3IwIkanOseTjF5ZkgZgM/
uoXNQiW51/z/a2SsAVJK005j96kqVjEjYloXkAJKZ5UontYvjTIsQWlQIb9WPYi2yG7y/JZCrAtD
Z7fLw4ndNpFF3JlQtKx3kFVT/t5UOo99pb1I0VbwukIoNdnTvSFV5nWaVJ4/laDJxXOgHbf3Kv5g
fzas/zd9KaJ4+Wy8DV825QL2/IxXBLUbAxmRdiHtoscxqNBgTQ7lZsUAZ1jRaLYv4AJP1kOat+Bq
x5D/K/vfYQ+Ev6bxaNtn/Kqxk4Vh0QIXwCsKLkZqoB8UYWdtp66B1eOlEbQ/UDlGx3XVlUZO9jxP
wwI4dGAs/Was1cU9gwzTMbZNzc3dIxrK01wWzKTZuUAKX9U4ogGLMxvYgOGviyuA12sjcXzdU12f
tGX5FM+1hkmWVtdqGPPSurFYysd0pqijpAIeToQFbEw7pAXNExdxUuizJK0t8DHTJq/lHDoAlqWj
XGPvc/UnPe91ELC/K0TRpvnqu4q3btXVMPFXiyWT0U7SnzRM1dnJLcBke+dldnDABhVeHcELKbcu
FiBxlmJN7F1BIls0W5idYkdCfrP3G1MfK8523jhF1jlG8bl7svmwJaATxVVbOrb2as1QIkvm8p4U
GTYj0NtR0dhvbJqzAPXV3tVED7JxzAiI8MMPM6ohvYxIoadt2fVgWAlX0rmas7DyQW3qs0H3YFe3
elHaPsfIPFAKAeALNL6NUaC4yrA7jkKnfTL/xTBuQ70lWcFEbt+kdJSJyAlv/Bt0rOSsbp8pRTn+
ALsP+reLpDsykFujcDnMbnaTDaUrYK5OgydB0nCL9eNeqjspspQ6Jbh4ElqJtUrzAE/EQRgah0Rz
m6Fv3Nc8AM28NP+iCIBhPZRoBNwsad2CcmrMoRC9HG3b37ldGoGbUAdgwpffA0cWAOom/k8xcIpM
N4E8Mz6/rxrhXJTVElAQT4b8F6olezwx6q3REemgd/qHJFuRcCpjtpiczRNKE0AtOzDSP60U1zCX
5515VKy5Pm7nmCCLPAWgT2Wsijdb/NwBIt56IhEyYcn5YhBLoGSPtih90Pe4bVJujBKbmAZ6LL0R
GCTxoR73HHI82xzR2YXhIJ47CEdLkR3gIgj3cEiESauSMIiMjkqw9yI2IHQ3jR+dMhSX1Jz56Ayc
hq4C/FRO1Rm8LwhMyyEl09w+qX69YYoJVCrhOcQJbCDytch0ftH5F9befh/B7KFe2lODRYt8tP9+
bIsc+hjywASRqHKcdiWHSFHsSvuz0jR4EJLzcYpuqfOU6Mjza6oTZxh1IhS/meNaRDJ8tYmM8Psj
P7ganO+Rav3+fdCFwBC5CfBE9JqLPyZxAkGf+3WHz4gXd2yCfFf2NxxXyJSfBNdGolnCx6gFJhtr
qVIiUPsS0KL5rHaqHqJ69YSrcix4nXFiACdPlBtaKQLO88XkqTLFIYeiFfNHaSBLtQ96LwSXodIa
17t3J8aPee3QYvawCXMi16ut4gXh3DJmGP/dstNT8bx4asRRFogxPiVrSBNOi1Nd+rYZVOzDPZ/U
ARPOcLEGu7Cad6NCw/QOFVpUbZn1JA2AY3ReJkHjCXxY6tnY/XmrTZD536RcHEMi94gMcLQf3Xh6
6q0ZTKB5kB8Ulw8CY/YpqQ==
`protect end_protected
