`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11824)
`protect data_block
O5fFysBSvOxiWla6lBMnWSZ11kRcEfq6fBwWIxlbbP8JhTCqMWGxrlcEB5kBg+/bBio9iDJcnDEP
fZZQLEo/qYaYg4EeKfm0I4dwEZd5SP8BTX4OPHqs1++943H0NBCnawtekW2CMP8be/2vSYJ8xE3w
xi52RnrEgjRIqu2PJ+qhU1XDdELmab/g/x2uzluUZX4yhySGa4DAOaB1qiM/fS2MdW3+e7KLCM86
D2Ln0Gdsa2SxIXSPNTGdqMdiR/HsfehlW0Oxpw4o2BRcQl4DIIyxlZt07aXB7lCHV00Mbx3L3XWt
NINGEItarIX4Woa6l3pXMpvXY/cpeL8Y4+tXTURGtCBd4ZhSIIiTX3N38q03v8NJDdS+7TP22aM6
79nzNJzURI9EDkorCN8m0UU9w8FiU8WEpoihKDLmSjQitiTpPAEwfon9fHLzWmhLPBcnLMdSic5Y
/rex6DZqaRJzCVdty0k03HZSN+JhX/LiDJg6WnCRy/1kpeiRYW8pdYstUxs7AWK4kW8MfUZume2k
Yiw3KJSb1IkyMcAEKDP6PCZEdHb7khJnrNGgctxcTQg8ek509yMaHctWvsLmuHmZ//zzISZwJHmr
RqJGOs8EW4L0k6IBF6biUZkmpowoFsaN0lA82i4lXtA1G+xxAzdGa3EsrZ/P5qIluc5eBN7ZWBoe
EAn+4Mu765rA083f+p+TSlIogCQ6uSix4LYxNwxu9C5I20DTiKZO8ljQLcjLN3J0Xt+JK2R5r5kQ
hE8MH4AmTDZKz6vB0I+m5INdJtZA9j4nnfU6v6MViCc92CJryh46PaOOQEyk1aPQK9uV+O2zPbP+
K6b+s/EAjeRMlpTRkx2KH+ORgZhPLEgXDLBLPxziO4vr0kMmTUZlS193Y2NDy9MNC1Gz8yUQP5x6
M4MlukIP/FQCG5seexO72EFKbMbPyY+BjoCpXoJyZDmd/jS0EC6PlYE8NVb2LKRmos/88wR86T+Z
yz3e6SRh/L64fbh6SWMPOGPImnQD9KhkYc5jh8Q6CuW20RmwqkISTgz8lG8diFg7w/TfbUYlzRpd
slAkczUgQTRcS92H4xy8NAFmfUKXT0D7aWgiW8VDHDQx2J8PCQPdxA/+G2M1djPQnATuVIKpeBiN
cVxgRUQI9vDqKNGbYXOvS3FU52lmRKPk//qptzG8X9TQDW28DuPDAYes/ZINAHUBKRhe0gOgS7V7
vCkok7/7be1Ko+WnC/zVOOsWMuVkczM4a5ss8YOkSiAbeWFpCWYGT02H+4ecY0dLjWUMpLubAjCQ
s2gyv512K5+loRsVpJpCYfwf0Aa/KYx1P295MnTsXVuSy47XfEkD7g0c03LxfK9Ua/kxCE7RNDbP
COFIDBsqi6XbdtEbDXIWwQEMzDXIFkxwQXmLM82xItPDEg8UchP+bYW03g4Vz8O3ErKwWYh6Ahkf
I6+9yjkrP/eQ/OjXe10XwwrP9GXdB8E0CnoVuEchhcb/sHgEAWcCipwTFBwawUjUtsvYt+rMy6PW
7rHdG8TRCrk4Kyi9UknrMP7tKDN9VRITpLjDgM1EOvPBhy1i5hk2TG1pVPODehxbNI6kre6zN10v
s1ve7Cu2P1V2vmnsqoNQ/kB2HlK3GNiUk1J4xJUJ1LSyTHQQy7i4d46OoimLAMBOEbPL+8uqPtG+
GNDg3wFJui5VESoVIXf/b6PxAHlA8J1nHscgn8qCzGALDIcGZ6tIMe/6RTpeJdO256PG4+ZQSLPj
lYpOyJy9cx0HwaQznaxTNVqPL9JogWDckmNygL0uxdUJP5KSy6+N3SQszzxbxaQf25nVQ2UwZQsE
XW5hDp60gWT5FBohtAj6CkZUYOq0KYduzKAlpTsM+1iyzFf4/eJSok39KxzvOuKmlaVXfuruvkgx
w0HrLtD1e9zN6BJwwdoUtejoiKo7UI3F5veJs1MTr3G4A/j+PsZz5ZU3jFttRvmzxYqW4jl5Zpk2
FVZlZr5J57Q8TPCVp0ZFVM46VbA+GVYP4V791ZWnS8x9H0ApePOJC7NEG8YFxuziePoQfr4zgR2u
O53zpLrbHW8iS4lstjMu+AOuxW90dydFgGl519bnQz8343EqmG3GkBwnn5+7+mwKbukPYzciNfpC
tEcyy5++O8ZmPyP2p//RSCtyoA9OvlNohCsf9UrtcZnsO4BSrhhZjzu+UpNAHzT19BzAAnEmq0Qp
gGCCETaz021apz0jqpKYr2ejpwxaRiWggPEGHWjon2Jg35Beh+1GLnLJxP29gi2cumM1jXsK4feG
D5IdlIVatCBCkwCSjtcVVlm9y2px4MSSRNY//mmWVpZ8pd1BHmeVApO0vsXJBOilidJRjHny5S+u
LYCZEHUC7v3o2+SVsUOXm9a8iaS5J1eKXsfAzKRCBTNZ3kedIQ31fgaL20bfSy88o4WgozwXMPds
n32JcPo+awOaiRXrwiYIgOZxDz+pjVzPH5oB966qBWFJD2AygBRHlK1pyFFxYmBz65fS58o2lK1F
hPsZi6SneJU8QjbpBC792lJcYtUhlOCRuNz6+1ZqXodFXWezdWEDNjyx8xkbuQFQGuMhSMv89mjD
cuhCVCmJ4PdjdpC8wp4QmleMdo2SFGaTxFXaZ0clHYatAN+l9Zb88XJN4zIy+b6sA3L2tTDMWN/F
4Fjf+iXNYFitE1PQnS1Ynjs8qn0qsnF1T2nlGybFIij8ROVJpNSQbRHVsUjC8PpoMj1WMeCrIHQk
bGisqZilrKS6bQZoeia1KT0gNPZwRVJ/CWj8jZmyLSUqM0LSoxRMW/f38PdnNVpe+DP4tYtujaat
vDVt4JqBwma1U1CvKz+ZeRci6ffX30ak2fGCD9sUpo1dQmulq5O0yPv2/IvQYujJs46kgDs059j2
9Cm/1QGiG7rqe0yz6raMvHuX5SbD74IRigmBHag+VP57f5/o+V+BsImU8njjXgb0YIUn5PjAOj06
89G+eMo3aipVjTvZkh3PjAcFHxd7hnBRL9AGFyiK8DSX0RJ1sFEhIRQsdqUb7VAVOlqOqIYsJDL1
M4+zFMEzLHVYX5dbkiowl7+1IG+Tavkow4I4Qu6ESmXNpmfQwxcWZgaJIaO+qWB5bJ0pxJdmuIwr
MApECVJaCcptFLuOH+BxjAfh7A51NFfRlaQOXApxsrbKKYCTyU15MPEdxhdKvfghYrphQnJ1Ylpa
jggXMZg0Lzenyi8dq60vCXiJMytTqgWJYHRv5ghgNLIiPsMFujaK/zrBEkYVKJKHkDKXuMxlxj1W
NKoRW2fLpyiYD5FTThJH9v3gtKOg1sUQ96y90BoCDyXp54TkwT8KlOwtdMEnLahA1HzRX0FtNs+J
61DjMh9xHEsYzCpaHyyfaacmiHNcs9FPu9fPTv4f6V0IGvOcid2oPw1b5zUXQaHZjRmYfnvBbzKc
g3NLyhWrPsqbTRvKFpl1Uyfklasd+CEa3uomuPA2DhIa9c4P4u8MPoyAs4DFhbj6DHI+dngHwd5Q
hvHBjfAi2fI4HhVCdaBMh3pazZyNyrLT1Jm7iyT4mZeuVkIw9v9XAwJiv4x2caRCORjzaAPtbCjy
+v933bLGpng/FLOKiL26ZRFgEttYAcrHJvFWdgQ3HGfRtYDKVrFAc2FqPSduFDJnAinCbBKlIG4j
o9k3sE5mRdZQ6NPQfUi4wdiklZQSvnjpgESe03QtMELsFjGG/N+lW7H8qSoVLAKF9EAoqY9M482u
LdWxYBaJUowhretiifUFY7GUePWDYAk5HPsLc51eRx/dlRyqcbU14GMZr0p67LFOB+9cwxJzs8EG
iCd0U4y3+6n0VxvAOxhCoTXxw6Ag9Ki/wtB2CGgPD8jhyJI04b1pPPQda+NqaQfC6AOb8103Jupz
hfhbe8SJk6MSzNKi3DKRAoTKR1hZQRK2dDRujH+nHgtZJM/4Z10sDHQ+Zd6ciDuCYCUG4YwWRWbP
rdbTHKfYbVgts6JGmFLVCYQUhxp/H2r5aVWzW4MrWw6QiVrDNpPG5SWN+HoWTaoN1N21Ps7W4NK7
qBgUprnN4/XF1wzrbIbi1z7iTdRjoBtKYY7ZYVUrEpUNVGx1yXI8TIwT+VuyRjzSR6YezqPeoPvF
P8RpGJI2BSGLUWh2Q6cGfRAWHYMs8LbYb6VkWKhp6qIa4Fxuqh47BusA2A6oVbtu0o7GEB/HBu8e
d3dalOX06xZQfpZwd94v3vFcWE/UjNXWgST1Os11Zrl1OHHt0k/EIJOyNKx9ntpgvh0vmcGW/rZh
SiedpP8Lwqhts7JzjUKmqRUaji0wg/6kqdJjwajFkN3dEkIGQb/ArYZyGGBpVvj9SV7iT5rcfuOO
Q3cuurtAIgU3e1OHZrfalLitXAuP+83VFjZXHCG3VEEwHtVi7jfWG20Inetz/GNueQkaebghoQ3C
1yhj9ETmyqBXe4qOrvpNerqrOxawqa8Uw9oo0XEu49LQj3DPQqb5ZQjojxqoR9Ibh9nJIrCwbrMs
cX9tc6+ATHc5uq8a28J1l34GU4u2og2JwdwjLuC9BZYBTaRJhRZSnGt8HQoUh2BZJ4PVfVgcik2s
C4FMhex8eYXRQowkDOH+VZhyz7/6Su+ygTAk1/T50bBgJUEAX899n/UNk1VppbS/YGNBEuMkYCjf
/QJPecL2fNGTkq38tkVRayAZgABLhgvpqETHLn+8B7SqoVIcEDyeDno80Z9fAZbHHM0oOfP+jr58
cRwQjYgOsvQ00l3QqCPEIbnGQDCJ+LXuC/lmHOopgwprjweARooe85tR7mGLwsSvASgRm/4lRES8
kRjkSJ8IjUfSz8WkSGuq8y2Gs5jSXlGppqU7Q4UWwEScruBpvzrZar3nwJaAlQF9pqa1ihwzU+n9
l5dfX9e57BD3ZSkT236pPFjkqecsbQ/LiUWv9VAhdlaKWx/p2aG9D4cfRW8bJpOPTocFb4kk++MR
Q19w4QXx+qIeStGrtjPAZevmC/sIOimMn9rMXQxNFtJ7Isj7ae9iYu2d866JDbfygQldIIfOtcPq
VAXjI++LtwaRsvs4BWktC2CgU/r3/lReNiCBUKem5/tsSvr9YzTU3qxlVaU8YS0Uq7b0rl1HMfKA
T6Qam0YgQsaGFolR4TEwLl9BooVzql8dgopQrwPCwpKiPaFULxMuAp5I85lOFn1aJoRwq7IK0o0x
phXJRsZacs1zgWjuE6kb1StKEgd1H0gHdcO1FTKWVnamxHkBiBbTlbpBFKeP0G+get72UL2Qtd4V
pfAd0yAhtKln7qCKmpf35x6pdDSIo4RjbA1Ok4UcJf8GQ4E3O5xL8K/1U1Z6dGosb22ZbQ2au8PN
kv0LfIRKOJjGv+1qwtV9AQwCQTZQ2NClv6pMPxOLbvLehV+A9ym1zNC4pNbdnR2AIOE+RgtHCc6i
AFaAuKc/tAC1RJ/03rf+uoot87/ZS2ejJmv6HHFXMrgRgOtTltQbLNzJaGPJgkdLAyiGTwPDLkMb
d90X3A2/QCwCkvAVKu1IqzpezEqSQdYqpnLzMaWNSo22kSll2RqGEbKqE8oRi4SMkE7t2wmI5GBs
K5WwL/4K7odMnKszDtj6vzI9K/fA5RTqXh1ow/O3z7LU6s+Qv6yLHdEfK35ZNxGWXpnaPY+Jrq6n
kYdMi/gwMDsv3lN0fBDcforEPLuSHY/0Y6p4df96VmyjgTb7TnsnvDIyP/aCBKO23JRZME06wicg
weDZKUd0Cz4C4OBPwwukjTHEfQFwICdEi4TGNjjUNeUrgez8RIaiMM5LYzwa5k+7w+5wPZTmvtul
dT9EOi+fRhF/DDMXfVVHeXg5g3uCLm7dm9UmR5j5AGxjCT7xXlDi6l4lR7EMBdcXMmmiaB3WyexV
yGOklyjXcibr1DpXk0VCoyqfO3SIO9wwbAR3Yh4jn1SHpM3VvRlXe5jz+/muMWFOwdH7n/6a/EA1
dYy0BjdNwcKTpqSp2IHfotTMPUJlibh2lFumHrw5MfxFprI4b/qKHmvwJUAnsJfZ6N40Bi8JGicb
jTCru4X5YHecUgQtXdwUCxFBjrt0DRpsLpkQKSpBCQ2iBe+177w4J/ADUcQasH0BkTc519ftXZLs
diq8hYD0/d6BSTNIMgk6JVYkklCzbT/yaW0i8ZDc+21Btqk7YfoJXNh0BAGqzTMlk/GqXa51lX8b
Zl5wHVOA3KPqK45tgcuPz4tBiXaYHBSVavoDzWJFrigErRXKLmEUsBSzxMPAUXHAno2Gg8PcQrgP
VfHVWn141uxRfdwme9FusmGfp6gly04yTldHyxSralRRb25pyXzpUdFUA4knljzQlkGi6I06TaxB
3RcmFXlJEgqtElIy/hNyon786z4QC/3CkfyKcpaosKZy6YGMawNCUTx1D+OIcIyRVoSMor2I2bG1
kCDuGzM9XecEnYzQwOzbqDJNEmObU0a2Tguw3nBCr8KYkzDIM+cIchKFYTY7GWd9s6Fa8lC70EHM
7btGFQjDbraf2p0lQsyLJSw/v+rTatbx0tBLHOt2gewRQJ1o04Nwu7x+H/bYOIrPNwvqahGnGllK
dk5c9/5fBxm4hpw9suB8Nbdy+XTQDs8X2LIsw3FiWIaxAMTamokh1hOMEKwsnxH7CCPCfeyOpNRW
Z7Z6IBuAUneopFcfU7uTrsEKIl7ujco42x1gVgAA4zPplu0RD5JkocQC1S096yUJF/uw4RaeQz2D
HbrjKd7+EAvG+lwP4qanWgCY3MymaLltBSys23B1/+WLaOH6zhgCVnnoBYy2K8cSaYYmsNBMtSZe
tS6qGEH5cUk36hJMajiZARlE4zc5NTlYX/5voN7+eaaBkdvhjBpyHuCA53SNSzsT4MQa6zAmFeq8
4myJH8Eb7OjeXiubk3pY+5ODUvB/JNe89JcDH1/d7P0U8inTyuWstbiP0arGDHx96DB5iCu+MM7X
Ox4iD3EiEwxaPeqaUCRYsGdzyopQ3OJ85uBPgvDPs+JiLI6Hd/OaWvcZl6XyqMCpY6ot8I8u5FRU
zGdAZghj+EgCbPGgHyK1ShwG7o2HoCuKpxJvxWj3+HAQvti8l5yj9K6kcQZAKSiuvWvPwuG7fATP
PTF7y+yg18QeeyOj79vmJegq95C7LrSYLvo2O/7vsKmXDAOqzItg2inL8B2Ka9l+fo+cjZsPVJZh
wBPKgqcWMkcpeC54MFY3VYTHQleBQBaZJAVrcXZe7GvvQqYVR5iRM7QXct9SmcviorTGj4VMSzvx
zIfeyuBQ1bI7H3LQxA++A1jwSxGX66qOjGyOWuwNCed+M9NILCcnPBE2pVtH9waJ8AsY10DECXFJ
RvRbPLNB6pMyU1UOoaRI0xYeqU1Huskq5OnbXnBgw/hQTNhYo0HyLf6/2zx/hMCNup5fVkPL7sJk
9os1HSZJvYixpXB1xUAEJLTO4BFZvU44sGYeyVO/HY2h+JW1ILM5lDbXWgYOtTNcchql7zJTXMYG
ttgBbHmiAJIj3YNHD28EQ7HCN51P0yLZ7sYtWVjLl9TAtYng+xrQ8rQC10zzQPWJRf8lsSOYd7gj
gChw1gd5lbq/Q+i9D/XeuF1v3ya9NycYGZOJOCt8I2H1heOGyoYEzcD1xjenNAfHQ5HlElM0TV7G
YHvOWIneyEJxdHg3KZoTDZLDWmabSaEPXZ2vH0eZIrLxI1A3rb533tfBh87pik97Kyo1Djv0tC6w
uQeeReXZKhRPVyFkMzFjrYvkSr3YEjtHWEaEX5T8mhGE4gnr/1KX5NBIU+ayE0LnoScekbE48hQB
oWtyUVjd5u3oZ+r9opR8oU7QNkUzT9ns931mNiRsYIgRaEXfM1Lfcf62GdMFsJSmkfcH6Kja4xFY
N658t6I5VP1PCZu5727cZR7SiUo33JUUL/8ZBN3V/b5dZSN53i3Dcj8fVk29WqablkQo3KhfPfyQ
uBsKcnSPmL+TEdUF89Jri3anxcKTNhN7WRVxt5qTVALs99E4yVAo64ewKAY4LJfL9F/GP/Dhrdfn
mY4650qFUWBZUZ5x9cQ0RK3jtOHPT7dPUBQRCiLckY+y6qRA9F07Ojz5Baks6L9nt0NiLh5bbQ0D
OF0ObjIoaNH5TpcX1ydmgs1lMQyBY/8GWBTXuRZRl59z+7pwAz1iwjUhZLWKBbNwnQKnKeneLg1B
GsEKplO4umlswQv2c6HQLiM3kQfoSU1Aqw68uHgZ2thR1KU+oIGSOJqjo3XUFEbpkkZkvkHP/BsH
ojlvT536oo4INdV6jcLzyLerzjEjwRXEsOH39wjcLYLZ7Ts2BGSeYqfQm1CvSF/Ue+rnSMMTwFqT
1s9CEVeZiSa2bXWu3H0j+Z3Pyi/xDM4bZJW64qm321wiNB1JgN90JMZn+DE2AxZDsm5QD0brQeU3
VLUn5D2JZ++ET0yBRfFUl7dum2R7oLftqLhPvgPn/2mCYaOHGgxmQjxnUTtWXV8jegrt8aRdwx2c
5EacQ1eBBmAB6eIdEEgYdUqpaYRR8moyBdqVOHk+7OJL7irIkZHJktRHYVTZLXb3mBCNV+i9v6/f
RKz643M+PKDGep7b4uYaz17fOooGfjaVHcaQoU8vEQ+DurokcAqK605QhFeByGWpQ6fzZjXbgiKI
fRQHvmSVKx3IRtdiR939UlFLs71YyWcIc0PY145tTb8OQBYlXfBhDVIisLlcelmbN0B8a5xR+0yt
IT0SLL9L+k6Zo13KPsCQVIA0IOaf3IfBSfEMEWEnGyTMrO8UYE9k+QIHfZbLeVtogp0NVXY1+R6B
jmYDmVureCBK8YlwRRrCK4GZkinSGtVEID+c6fWe+KfBndecGGBPxSYpAar0EU4vFPQw2hoxneAj
x4/wY+njnF2q5qMGnkTYshVKA5o+PMMWWafoEUAY7JHoNPmxEp1ZRD64k3DY4jZl5/rQ9tsZ/30I
xFL66nqv1h6IHOoKWCBR4rWH0J4OOHeX/FNlVjSQMbQoFCO4QHj9ctvplJTvR36WmssoODTh19GC
+zzZi09gx+y3CeoA1wLcI55RbbYa2hZm8EWIChE4mb1cwn8vwblCvHx1i7ntlmq1ZDJD2n8++OgK
ldNDnKKKsD8zFuXKHNVzM1ruJyjlIBx0cCjUusHCc7//baA92JKZlbr2eNjmrv5i32AtpbD6ag2L
kj7kBEMh/s6PmTPahdOlvJuodFFwrtMVVBFVb1bKVrnr6s3xc7lOVKaQwKFp1pvlzKRtHBMGqW6M
+BOl3UiIDVKWjEiY3L4pXGMotH1EmwC/RZUaL2GmPPi56XHQHkCBRLpA/Jl6L4i/Fb91pHjs60br
1wfKQkTI84ZbUiPEtbQsh/WiJ9iJxjPch9UwtFrRDQG91fL8Y6mBjOFltB/zQ2JuLvp8Y8VwY+wC
I2NnUFed2maI+57bvTNQiwzJH1cpEvwGNaCGHk07KlzCLI4kdmnnZIZ9E4zRnE2eBigzeGpWW+iE
tUWWNeoOzDjHF+uf5YIHocFcGnEgPmGBo+7vJFWSJREdoc8DHeIC77hPBpI/czkWQ8CcDvAd7/zk
HSBLaQufH2tytwM80lB+dlimy+Do5wEoCP6zNYuxFf7bsCR9kNhd8yfJE/KFOBtPk5/3kYultI6F
Nd7czV5izbxlQI42y+/GOetazeswmxd8OYrVA0JZfJBXppkK2VzCtI1tPzpUh/Vq1hu9eaGbQQgo
GwZiOd99h9b9Ud2brv4GmZf4WPPNyr5xShkL6Hnv2MseYB83ZFSiItMigvpJxdBNEiIFH/Dbd7y6
8jic4kVwWOJdRvmKHegB9lIm6T/fRCEIRAOnGoxknbAJJFHpiMdjaHyDrcjT3vokPlTFu9jsSxwP
c/rJWR9K3QLF9E70LukLGqMgxmhoOLgobLzjdJiynWZ2sBvFocDUAydo1syK7j/FvThRHyBAw7bC
/8iX2irMiOTT2dBe/LiWt42YffSFo9bYINjYgOxqzalzz/H75NpLmm29A1b3y5+qDjtXNrtP8Uxi
lfuH5+Y/PeZ+86mZtip8J6RH4eNH9DLf+Xi8RsZfkLA1MTz9pHc3nDz4nxK5QH/XOWMW2UCXR0E3
xgoCOunGwzCqE1kJ3RF9FK3lwXxqAG8SLGyZwg8vFSbqZ9kfmfIKKEBFl3l/by+jTBtF6abSvgn9
M6pivwVQI1e+/hEO1lKFuZr4bSXwW+rWfsmTnbZhHPRWueRRr4WhPLHrV9yjLhNvduPeCKwIDALa
eouQpL6DwNu/7gcCI9ywS6kj8L3BEsN7JyHHDFPQi7L0yb4D421/crUfz/U+hKSTlcS9O6o8r2i4
wCUHTRLjfbHX4xUqEc7Y3HthM9Bqsaxx+F75XGRFy9WzyzKWFznnoadv71FEFvJfGtse+eBwk7Xq
JFQZNrzZIlKRkVOpE1u8KQEd0TRNigJeXWsUCLsfgMk3ipFZzlpEkN3nDyzjmn/or9YcHYrxL5kN
IWvM1wN2+bGZ8RIzZ2pUz7i4JOQy1pL47nYReAewXpH/7EXkfLUIVifnLkqzzCleQLtHTDOuEFl7
XoAqmPGsF52Q2W4l293loX306Z7tAi8r82bRADvdz7Rh3WvpxR5+Gl+SNPOU+oQ+hVjVlky764UX
5HV4vPSVyIG2Lak7rgaVmQxVkV7uJeRc8B1KombmJMxSAE+JFx+5YAB8fGEyqKkdiUNj0ACPLLcm
mEFR92I7kohIN4JBN5B+lQZTs0CP9JC/LhqB9eTyRWKWjKUof12i60MBcAU203h0Mta9D3e4SQ9c
jq6HVabOMflG9cZDXJSsbpavO8nV0NmuAUYGlcjB5qYrwKmfipUh7J21YiwI04ug7WbtusFFKHcm
/1xUFPhuvN0+6wjEn4Oi4zs8OjQJQouFHaradjaxvUygczQ7793hqvZLjNb254x+uztq5Ol0KoJa
GtRC60628hne9xNfK0aUrYyz6wusqEV+EjUI5mF/a4tJYEJLjMXBHBkS3UOR+GKwrk9YHi7lQn4R
+/YZZI/Ao2+J6yoDsPn9ghR7oXRwAMvoMrrR5JcpgNSQddlyuz1xUS66PIPf9Dz5A8+pdTVcQXzK
FXbqwQAbVsSEiLjmRQV/kaFkpFKeTHu2uQeBr4lUvhBPrY1v9vfoZBhbtwYY9gd02MwzP4UW/cGf
rPeFKSQntQcjnfOPNmNKj7IKv07kHYbZCjp5of+QKGFTOzwVb8W+Vmzc3FNt3JlK5RjCUq1CxmXC
UVVgf28vdsowrkyJXOVxevhabx29KdMfTwxwOTEgIG/G7AJf52IyGFR+n7HvlwfPoFfEgc+XCcVj
EDF1ayrovQzMVs8IlIjl9jAjNrQPRL+ksBSfkBst9l+gC6nMKYneyZPcEwpdgFXKqqaT0BYY+1uA
DO4xbkFqeCk68Cy3gdSYn9FPqMWy3NHflj/hrmnyGVfmcLulNLI4jzTEfZXPCMSNdNcYeU4SiCxT
s8hnQkxwOXSOdV0wMglEoOr31vX7ougHdXJbCxE391aiGp1fDa/T8hYopA3Y5B7XztIc6ifjOzra
i5MYUp3O1qly720b5AtlTPvI8YAOqj9KbS5rfGHBF7T2tNpUdvGv8fB7XWFA+aoovvBC4xWq1IIS
+ZvxfKjxfoEzspVlENwQQAYT+brfQk4Ch1VYjfZD2+o7QkXOtqmk6oBpFTj4xgPafF9ImHnRReSe
Up5KhQTOe2vXqdqNrIDWkF5JO7/oCFLcBvWGmqmWcLQCqvJI5w++rPPCpJ3MdzkGkAcID4pQ4bLw
01sOEQPkOpBVXO/85t4WzsNi+aIC+th7H1S4ZzeakmgNzsaajbllD+sgt6q3Rx73RtpMvvDFmvcq
buxIfDxTIRipNVJVOKzDGw+2pwSc3Q8R5ZnZEpImTtS17wNM95x7MohKADOpQQEWK3/93C3b1Ofl
ice3FQYH8QJxfqppYnUhVdfWpcHt46fB5iTnaEMnMvGcnFSkgmjoykoKjxkFWCQt/2IjXk98I1sT
EUtC0/Z3c5GWiyz3KCyFZvWoQBwvpg+31gXkXsJQ/z7cbKTfkU2i9DbnDsqy6RtyAXHV5PeufFGM
TQ9p6igHIWRs7IY+X7YKfccaKre5D/CGTrLHUVUOsQdzDmBFElEDpewBbA8Mcztw/ApIECtNQa1V
6dsOBY2befg73IIIXBVzBhtZ2xUk2EknRODNcOgM10qmfUmN30qZLj56DtMxZxAWBzkSAUMVVDVZ
vlzO8KeUt84/cAKQt3PET/BYuEQzg5NDNXzmEIHmZ9nolS482t5F6HyqCh0UmpBL9FnGFhmhR8th
eJdt7gRt942XKj8+7ol50iBC2zrbBdYiaUiRg+lalmh953HeXvySLZlBgNEK2xfjHQ4ldnfLfWn7
Kf9Hud/woebg1i3Ibt7pdESprQrrVDrf/fVBJItcayUCCAIl8i1b3aW+H1Ay0hnoAHlIAYnybxkz
KHgsretDfXaF3jIe9l3fQng81xnvmm60DBXyIJCSfeIaOaYtgLoTviSF97d7oEQ5w7TKYsx7Dudn
dEYF/QPtPSch4uhj4ZqYrFHcBFVyw+Ho7ebHB+dZ/beAVZqzNTfgKP4bHnUIwweiXRxempm4Ngxr
D3rnAvgKBc5lO4QQpNIkcBhms8nu59qOcyheKmh2uPLQ6CU+9qyjSdB6hZOspUF1TR/3b5tMbLkI
/6dfUZVajHo/euIFQhtWHyn5+nPATuzTjQoXzHh7OJQjPe14utRXAo3Axc9PFd7nTmKVU2uilRLW
guBrxkx178dbY/6H7peyyty2JXww5GXzgfB8yQ0Tfu4ieyLCDD7W9GqMsNxnx2AsT8Q2TOTmp/qP
xtN1s4ZoHreARRviNTMk4r319qA5udeOk0Q75wOObVnu3vi5bf86LP/20MbWAf94fGlFh1W+owSc
stTyFFV2shHmjYV7C7oJhpLZMkwvgkXOF97rObwUJi2d38HCQAZY39aN4C6hgYiB3aCieEQVFPEP
/houNSHGBPSjlRam1XGwV7RVnlK+Zqvs4Fxp64U6VQQWT2u0Vk6MQC5dg0JcTcu4HYTLwNJ1+QYv
/yajwHARWP0VVgXnvRLijnnqc6v8jMb67/ISPaXEUl1XMOoPmfNtwf8D2gsNCd6Iv/A382sWMA2E
+5FZ4Yt92hoYRJPEBp250BjnjejS6I8Hu1DvHsdz21Fo9I2+nWfy7GFI4PkeDV14wQoXDX2RGb1n
lV9vogZLvZbNlLAGoQY9g+5f5ZsgqlncDtGLUNScXJjzO53lfMjsZbUhMbWBSfgctqtjUpjSwBEL
FuJqDM3noo4b2iQCVsXsW93sG+ZIukNLfTEblTFxOr6QfS3lNKCM4BsqogqddrQJPmihZ/ubidL3
GQMSH6LXATpkLX//8/DZYgp/akkUiOWytApj3Mwg1rRR8876DqPKL3iQPhqAzKqdQnxipgpVTJYE
nxirQw3YT2Q6DMFXh/Ie7UIsoMYsqycANt/W5qIciATPw8eRxjM9UrajgQiSg0fzTyvjJy3ZaDbC
pD57QkbxofGbCcpiJKZ3zBfNNEswWK2EmLrKiIrL6Oa65+djldvqrqRzy1QVm2oAU/7IU4xOQQ67
XVE3uvAZymKGr4uEaVxl2eGM67qXbWPq7xv4crgqiVYb9qIUbLUQWmIQ1GhkVN5kr0E6JnbI+Xz2
ywmFhrMPLI9vgVFVbsPIxVhvlpiioptTn9McpAkKQGPL4HGgVDjFF4TGAQIfza2NKju3x/Q7OtgW
jRti7IoH41xpGnE4ZW3oNlQF7N3HQ1x3yskP/PgNKf1qXgGYDd+FjhXgDn8MH1oDFjzwbbwwvkNG
c3w0q2Kbjt3VA0zy/bSEo4gYS+P/MfmWOrZA7ynX0zJOoa7dbNWEtRw4sQ4EWJsTFofhjCUsl/y5
vL7kGnD31Sx42w1DhtoLLajTMS2FjrjMuDEl6xLE3hSXTwbPi36UuhlW/VymjLPW3UX/rrEFdMLu
fVcZwg477Vzc7bk0OBzvkA7UT+Z9ptDFzDJTYEB0+Kvu6Fz1pox5inBe7fPUGzZm9ohctJ/1UbNJ
cemm5NjdqnBhZlbyBgdntCfCU8c6f4IEO/hFyIj1RDJIyd/RrUpToahST4WT578Ha567/85fsr0z
pzcg/T2lGg+yDucH9m0VmIYKaxVCmW+eb7mtxzf3z5KkDa1vzOzRrkOGI3zN1hFpH345ihqQF2hJ
985faeLzQ1GyC3NpAfNQR1d4zmywelm0nsHCXTUtdhLyRDpKCcOYj7c+DKecvKnUd8oSx7qshH+A
XuVuyOP/Q5nr0EjSCBZpld6whCaytCcUcr+JDCk9jmEH3AqZJabW3zUlAhnkNRGlT+xANM3xYJLD
ESwrfHsbBRSip/GBiITmdYzQkClEhjfSjalAcII68dNIJQ+bI9nNbWZhfipqbZx1DyJmDHNXguv8
tk/FwqYTEADm+UAGfbN7wf0T/OhtXmmR7qihehBVG6amGjibP/ocZjO67yO2GQUP6k+Nt7qOa6Wm
GCqWA8bbRubRtxxZ5AoFc/DpB1FD7sUe3WdiKOMnnEggsZ76L1csQaasfD9eMT05ybDJ3uo2tzQB
0u8oYJvD/zL3/8D2uAzuDAxFXruqtqaVx8Wcfr95dEBUGhHMehnSpXoHiUTzMrha35rBbncWB7pt
ws0X5haqtesaov0sznU7/OR7rJsYLOGcxsAfb7icPOL8coqpRTGk67BTB6iapEiSlDK71GVFG1ch
85+JZxpojfYADdv4wcBoFM4yKja56MfOAsugfiUWRdlrOVgu3RAfx6CI7zP7qVO5Qo8XlBCEmN6i
KSAvHLOeljxIfUzVqDfNxP6dLjwGYiCYI9LHgbzqazBdcYgd2gAnl8e2hqCQ6V6lkCZb13ptwg/Y
PcWcW0zdx37y5gnQ/0uCZLZ2l4lZfJftiXJLdb3yL++2Ufck92++a8ojhoYPXK3iuowNiCjWtFng
YS+7hAwbbtlxDa9UHMbrrmIG1rfsRoq2K2dZZQQ27mkD4e6Qii8nKm+qcEvBrYA2u1woeyESDfBd
SY//wc4IppYk2jMTGfrSpeKnZy8aKinMqY7Dh4NV3kTvdQX+aexLvGumkQmuFXHloz5Vl3wp/VI/
Laa3HdgDWIKRvmzOmufbR9lgzP1yBU+UHuYp0gmUq4L9qcHY26wW6bb+vIpHUxU43QqWDC7XabVk
50q4kRXga47naKKm+TFiL/2529Lzs857aMSvssaVERpWJ78zakZsV2f5/hGeTml/Te9GEoj37t07
g/RnOlhTz4kr2SiyInxyDyaOBILqDcH5kwKkbB1zfVGFEfjLZjymdggS09nCo2z48Wtokncfy7lu
CZXjkLxC5GvF5WmBShyWdVJ6Rifd9Cmsmu/sxVSGnwOkHDITWDmrI1YpqMOQTsPXaBjqDPI7ScAf
q2qEUQK/isvs+ghdjw7mkAqjkxIgYDm+bdhmHV+cREemGErO+BQGVKutSIuRPk5nUxWxhdrZQIjF
1LBbnNEZ7+6TD8tOpCBxNe2HxwNbSz1tkiYGrY/SMP0LPZwswpkxEJE2kZzgsQn7wixylHkAdXGn
uhGGGe8Y37pzQcl06u3N0STegd9PXVBK8yM56pzvHxbRSJL9KIPMYz6g3xLrHqRHpZTC5KN/yWFh
FnlHITiDNohF1aMFJ821iXT3Vl5E1mWSsOI0PAcIIBpD94nsWuijPJ8zj5+YYuLEDpYu4yNDYA1f
lgtABTHNlQN3mF7iJMTnQVx6xnVF3dTCb57Jg+GdHY/ZSEuWgoETk6HpTWNk5IVZ6nMI9IRJIsjo
7bHKaT3dMqHL4lLtAHk2WStArHFZkXnn5w==
`protect end_protected
