XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o�_s��h�sC��C�������>�B���؊ �ڿ��X�7�`��8�;�c�̽Ɍg�b�V�U��gu�l#d(J�d�h��3�-E�.e3��m.0��, �i*�z`ޘ�Wr%ϵAa�	pl�n��W��'J����-j׿r�]"��gdkN�;�|�*mZ!|a���Q�M��+
@o����˄���8��K��������V-��ĩr��P$�qX���K���^�!ת_��([�Ad����k���TK�5���4l�T��o��Z�GV�A�z9*>�]����M܍ҴF�J�<ڇ~������G���V�.h�.t����F�^�T��@�f�7C,��(�H��+u)���B~Ĳ�˖���)@��.�d��i�׷X*��os�zF�c����%�����*}�����~������>�P�%i&�t4Ч'S�r�4������j�Z�YK�����	�f�v?�j]SB��"�j��y�q]e���Ȏ�;��__\���O�w%@����f�a#6H0\�U�H����QH=�nmav4���x���aXM`y��xB4�v�������[咩�~�c8���Pl�$W�  ~N�e��H�s�jx1`��sq,�[qQO�9<����C3��0���)}4{��3�d>���fs��B��(Q{T�!�"'=�v���-]f���u�WWڰ�	,�o��w�v>Qq3���dBY>�av�Xͷ]:"B��XlxVHYEB     400     1d0kE��jo"n���:� 7)p=��y\O�~�&�R=�$��k	Z܀�0&1Rӟ�7Q�Vrw�����>+��N>�;mzܰj�87�xcA��/:4���\%'9��[i�f0�Uw&Ծ�6��˛X�����Oj�Yձ�V	?Qǐc���|�6E��CgRt�wY�>aw��LL�S�\|#w�޾�E�Vm���ե7Ϗo�o7��^��x���%��o��_2[�63��;j]�H�-�	m����+�^�������L����n|��C��i"���`�a��G�C|x�Л�I�
�ڿ�|�,'ߙ����M'S���W̩B<c�9˭�΍���M�9:o��iwy�:��U�`�F)D\�k�������+!�X"�N�,�G�\=q��d&�� F�ڹ�WhX�@���U�^�kP۬�ޮ "d~���B�0�pHo� i�.t6�V.��XlxVHYEB     400     160}�}��8�ˇt3�@��-A���@ӫ���Lp�dB[>5e�!^p�� ��+�?.,�{7'��d��X6�]'~0�E7�.����I�t7��T����5]f��F��g}���t���W���N~�۹^�U���2m�j΢��a��@�n�6$� j�8 ��X��47X���Lt�K�a�A��\��q��9VY?��ׂB��F'�^�{���s�ys�7g��>G̞�\Ѹ��I4��s2���f�}L!����RU
�#��.���7f	�>��-�"/�鳠�U%��"�,t��hI�(eC��u��B��)�c�S0TU�M	�K��.+8
LG�6�eu�3�XlxVHYEB     400     110 ��|w���EF�ۢ!&Ka&6'�Ȇ����� ����f.*!!l�k6>�}L�o8s(V���]���W��f �~נ�s|�d����1��!����~N������G�HGv���>���*IЈԢh$�'���-Y��?��s�`=9@}�p�xƃ@��82������n�"D>J`��v�ʷ���Cœh|��4�3�eTj���'`5}��]Yb��ʠ��t\�
;��fN��1p�ݞ��~I�j����i�ɴ���ErԑX8�G�zŁ���Ch�XlxVHYEB     400     110��T���ޖ%�5z,��c�cЂ����$t1
�(��L��6��U�j&B�CTO��q5�I��}�2�QQ#�4�6����X�uO�5������Ɲ��ƾ��5C�{�QD��U&_��ܩ�Ofj�L��A�U����[�5�Q��ѥ&H��Te�j�2��j�l���Ds���jd���*.��HxHNL��P�����E��,ꅃ�5J5z��)�az/�Y�X��x��m ���0G�<.
�+\�1�XlxVHYEB     400     150U�f�e�j[�I|h2�c�������� �H�i�<�-�1!���Y�^'M��d�-x��ٺD��< �gquB���9⧳���̦p�
mx	\�# ��]�#�!��S���Q�ճ�*����X���	�*�O� ҈����i+~['�,��R\٪�y�h˫h�@�;�I&J��=+��r
;񘇣8��q0���@>�K?���ٷ����p�B��%T�O�ವ�F����& ���)߫:��#�v���M�P���È��Ku�n�gN��C�x�ڰ�2�l����|��4Z i���k�����;�I�������v�ͺa��,���XlxVHYEB     400     190�[*���_O'*�hӌ4�ۢ����T�֫�AP	y�z}��qf��/<��Q��	�N`��~�>%�dGs85PSӷ�C���9�p�d�FW�,�iNw��Z��~Gk�/{�P�7R}��jY�҈)��{�c���%e�n�̘[��/m+��V�d,���?)���̠���4)Dk85���q��C�����?���\�miI��z�hG�49"�I9�,�8v
��Mņ;Oa�g�%�R{�˳)���k?�kӜ1D���W�[��dt����Ew�#\�3�T��'���g�~K$8�^&aCt|=Aӏ�^Y�8�pr��<y���A7��������M����Z�Is_��7k�Ӷ�����]ƥ�zd�wc䴈��АV�I�nQN�c��/�XlxVHYEB     400     150<z����,�j%�"At_��{I�{�
K��V�{�8�����vO��-~R(4��Z�Z�l������N.:LW2ԁ��̍]F��j����%�hs"���E�K���y�����|fԘ�����V�D���F����O6�C���OϫJ}z}�=p��2]��-�v�2���R���6N�#߭V�e;�e���4��xLAea�n[��� d�_m�Ti)�Q�{.��ԇ&<�AY�!��2 k��VUf���I�<�o�9��ׄ9�PU���"ܽ�}1�ec���#����\���F�݊�kA�d��w?5qޤ.V�/'�I����,�wG�)�6�lXlxVHYEB     400     1603��A0H��;�����Bec��6�BЭt�@8�i{��-Щ��� `��$A0�l�n���9^J�z9�H� -{��H��N=GM]��U�|����1£�W��y�YǢx`�,e��mp���`*4@7�3:�
f��(�~{DQ�pkh�Y3
�� ��=��F2L=�����'��8����J�)'���3A���!��͗kp|���F�ԣW�(Q3:$0��ݵ!����1�h�h�fi`ؙ��b�s���C0f��'�h����Jn��s�|Ů@Ce��T�k��}ȩ �-��z
�X;/�)[X�fp�:)��1�C���K5�/T"�䝻b"�*�7���XlxVHYEB     400     120��@:��]�LV���]�/_��"qڠa��q�tO�v|�"vL�f�MQ�� ���?Gբ������K�iy�5ߴVZF�V�>ê0%�/ŎB2D�E�U#Kg=� �+�`3 8�V,U�چf�t��!q��b~)c��j��9#�7뀜��WT�m`�l$4�-�.L%\�Ԟx�A�� �,�UE�v���Ї��"$on��ϝH�����(\���\�0���1��I9߾>~O�c �28ۓ��U�p�@���<��=g#k@-Z��XlxVHYEB     400     1b0m���ױ�F7"}��k�[�������+ռ1��ވ�U�-c;��$b��:�Ќ=�/"��,�r]�S7���$�˧���o`�o	T_���->�����u��!�^k͢Lñe�h��W��!�,�v�R��PEj�b����E00{���.*w����5	K��p��^$�iS�V���LAenږ����t���Nd�zA�o��g�WO���ٯ(�
�!+�F���&�)���ԏ��� ��oU6����i���UX��W*��L�����)�Z0�>�Q��g��������}2[H��I�{��cFĦm�b����M��K9(�M�r����QN��9��O�%}I�>jJi���Iw�/��W�"ǣ�h�fa�w;$M&���Z[�|4�~�L�ަ�u�Q �Z?���bQ�>�^��E�0�7�Wqa�?�8XlxVHYEB     400     1b0]�&��{����6b� 5������SK2C�d;' �@/���Ći�/u�9By�Wk�f9 �|���A�G�D�����j�&�޸���W�������r�6��2;iB�Ac"#�}�+9a�ؚ���"W�-�C\O��a_�m���vظ�}.u1�B�5�]� �f �F�WͶ_*Ç�g�#+v�au����?�!����Y}!f�6*]M��]�R`��p����dG����SL��dwF��>��A}{�^m�<~�*m�|[���c��6��uF6p�S1f�"�e�h�P��J໶i����L��H����0UO�y�HV(��_j��W�{Y��8D��q��v!�� �r�n��f2�r��#���Y�O�l���~<&�VE|tLʱ�-��@�݈��a��<���uIXlxVHYEB     400     180���(m�gQ:� ��|��P�9�����:FJO��˴�1�+�3J@à-L�Y��l�O�a���?c�
)Ǫ��?U�Pq�%<ah�~�c��D0g��I�l��$.e%Ar��*^�"X;~�@,��e8s���"E���������������_8J�WՆ\�J8Wh�������o i��_�)��_Ԧ�9Х٩�����	�,x-�GXIu{慨�fp��XD"N���ذ1-E�zfw��������dK-�͗���� @�k��۬��w��7���'�EM�� hi0\���p���X9#uqӗI�[X!�K;��e95��~��;
s��Dn�8Y�U��݌\�=���$����$��˭�d8Ɨ_��XlxVHYEB     400     170xv���nY��SBװ-����:F��πv���|�~Լ���6��c�7�8�ƲOBp��a#ྶS�F�E�W�ǔ�v��򧖽P�0[ؾWߧ�A�ߵ���b'��A"�a�f�ډn��.�RC�T����fs�ːf.��Lq7��!,W��L�e*0�����d`pk�0)R �F<����X�TO<0d4�b������5�b�D��%������#�4)G���#����
��Y�7�o8��3S��+���l��Z�t�]�StW��l�N�O�L�RW۰���\y�G1��/ �bR�D�v��y!(Z��Gu��z8ǽ�\�J�:�wb�W:�˓@`���\i�XlxVHYEB     243     1004U�&)�Ѭ|��42@�r,�WKU���LI� ��?7�)FԄ���B���d)�sΙ.z]g���Q�=�����u�좨÷��ѳ�8v���¥�$EA����Up0��r*�z��n��K�ʞ~�ɫ$��I�1���q�N�,S�ݎ|������׀�8t�:���X��Gt�קp!'��8
/q@����m{������p��n�vN�o=P3��Q�n�E���xl�W�͖�hh�M���/ǌ���o�fg��K��