XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���/v��P�B�r6e�v���Fd!��"����`(¦7����UU���� �K�n��#(�*�h� 沄b�����?�U`��QC*�)���2�vڄ��p���O�o�bMw����O̶fl�����A�g�G��+��m�e�PBS(���vU9`��cˣ�f?�9⇛",F�?+k$�pv�/Gf��m��䚞F�g��q}�k��l{�����1�$����>f��.߳�l>�8q�9�^�m	��V�ra�i�O�F����b�:�-�O����4����t�a��2V��p��������g0a���e���T�¸�焻�hӥ�ri�W"S�;����DSq(?�^RS����yc��2q�;�@�8����܀����/��d�
�'��E�<��υ˰���H1����`<�=��@<jȦR�;��y�g�Ʈ^Nq�BUQ�M��R:��#�����:��> ����2��0;Rpx�#Ƥ�i&;K�����9�-�V'�!3d^���m�Z�F�n�6Q�
{�C��f=�|XW�m�B$94\���Q����<���n��nJp&k��"�z�>�(!2�|��7)ϰ�g5u����e����BL�����{�J��:�[�����?do��MM���}@�@{2p2��4?s�\��.�����8|�������³��~�n(�8v��M�T��f�F'�B���o֖�O��`��ftfi�y����7��}�m��V�\�ό�&"XlxVHYEB     400     1b08��C5�wJ/6��O����m)�&�_��=��D*���'�y@�X�ƣ) n���v�b��a���E"�vkDa(��lO���g�˟�'�aSݿ��u�6��w�դ&}~���G�A*���#f��ei�̝�v����<Tc�
�_\(>�)���b���#��tA�*v ��t������2� dϭIҁ�  ����XR1��[12"��ٿ_�}o�oq�.�&��V�ƻЁUѓ0Ᵽ;ԃR�%|�*ɍS����R��	��'`f��W8����|Ɇ���|�N*�΄dW�C�yҵyr���	$����\ui���e�BF{�M�Ʒ���{6�V�-��`�R�`����hy�yh����W�\݁����~�v�Y;ĊP���ʯǯ�Y�4�?Uso%e9M��0]�epA,ՐT���к@�
+5s(��XlxVHYEB     400     130�`��_F��o�`$�`�����FeMF��9;���ׁa�xL:��?v�r��&������d�ŗpf�T���W�_�jS���榚<�2堳�ea�'�&�;v4C]#FqM��۩f.�1}��R��U(>7������(�թ��̀��Dkٽ��������0YM!Ya�)U�9R~��/�D�M�w�gZ�[U-*�o1F�w��UG��� �2�|;����^��ぅF���[�&�YM1��:�<�$��R����j�/� �1^KR�@���x��î��*[J��XlxVHYEB     400     120K3r�/�,��$����<�z�~�0j
�`=���.�k0�ԍ�|�������S�Ԃ`��y�/�!1���u�W��1������By�k.�D��pB/_ݑ��
t��Z���Y��H
��sN#M�r�5 ��f~�H	 �X�u-o��]�q w	��(&"���k���	�k��V�9��hDn�� �J�tq�MWe��wA����J��-�S�3����d ��t�ψo	�u�{��d�n�>�8�����͊{������.��Fj�������P&ZT"XlxVHYEB     400     170������.�6���:Į.�x\a����<�e�����"�5� {	�7��R; cĝ�x�lX'dd�^Y�e��f�p��ˑ.�C_ �vL��aiK������/��(av/z�"/4��!n���\�M�+���3"CP��q����$�QC��ܰi�a� �m�ո��;od!#;�/�G��+r���C_	Jڥj��^v��焈��fk���V"�h^�.�O�H�]í��ķډ+վ*���Ii�BRj�m@u��G}yt�c�N$��0�dϽ2O�t���Х��.���/���8	�r]{�WZcيAc����mɨ������B��0���ݭV3d�E"R8�d`�
�5/P�XlxVHYEB     400     1c0���`0;<!�.��4���՞�6C��yX��0��_���^��[�$~�U\o��(����L�X�Tѱ\
�U�<Rޒ�u�S��0���F���v��T(,�
�p9)��g}�_(Qi�t=�oտ�ռI#;�>
�>ƛ�c(�Y�˹�ޯѹA�j�`����u��ٳ�~�`�7�'���z�+�h�F����d
}�j��!JH�B̙:��H[����O���%%OGϖ4��׎���lH2��w&�ZT��Qq z�J՛��3�g���ZG�4��8�&�C��]x
�Qn$m)&a�4Ͻ�:Oאw�j�.300<��Ɩ��	��\���hU+��)42�/��'�kq��a�$l����~^���ӷ��v�]�:xQ%7yH���X�n|�۝�~��˗�D=��g�CAmȖ�[��-�'��-O�D�c�pXlxVHYEB     400     170��J�pR9II����	FV}�N�2G��W"�<�=���D�-z���!�y�aY�Ә��zB�a��9�T"�.��'��Z�Y�lo��l�`Z�j ��T�-�JY!{=Dk�>��Ϋ�&K>H��T��W  ����h4&˲%j껈Cgv�t��Y�/g|����Ư��`��3�\���F����.hFy`r/��I�"<3��n.���+i��� ]��ɰEuL���'j�MƳ���yCՀ%=.H��C[O��Jf�k���8�$�J��'�8�`>C �ح���8 �!��2�Yw��F?�����=���c�?��G�a�hy.��˙����ď�"XlxVHYEB      5a      50v޸GUp �T2dC]^=4�P���1q-0��0rӘ%?���c��kπ2-�L�>�{IIr�2Hj?:��Z�,Z���*