XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��N{Ŵ4����-�$�Q���q����좱ܦG���4����9y[*��TL2�I��o�Z�x�3��^��~q�'6!�w-4�;��	�Pެ3�og�T�����"7	������+�}i��9��b�Ne�#������d�1���|�tw��LA�Y�Y�T9��ͪ�m��O a�Hy�k}�\N�t'��EŢ����I�����0���9��m����H��y�ۥ!\7��F��� Uj޹��,��Wbg��E�R�}��d0��� $����j50
���&Ki4��UE>�+)h�U�X�ۃ�f� f�O��Ca:"�mǚ��l�郓g]x͉��.M?���(����aڱ���޴y�ךº��P��D�m�x���Vdb�����!�#9��P�e�u�Fs����u�}h�
����4ְ;A�~N\M���!�Z�%�?�5�*��^�S�As����ў�y��*�O�l��Q3����!�������0� ¿*�m�o���w��O:A��ycl�RX�b�,���gxF:;��%?0=�M�syـ7E\�;hJL�''��{$����WB��ʧ��N�O�ϐ�3��1��s%�=D8���}�Y������kz�X�~N}(��_L3�m��F����y��F�6<u�dsJ��]��z�z������ ��j�iS��e��=,��(�^m����{�瑌Y��h[�g�" ڟD�� �4Gl�pԶ���ک�Bq�XlxVHYEB     400     1b02�2���b��B7pr?�yc�9�Ɖ!BH�z�����Q��r�bֈ�N���Xf��K�D|I�N��U��`:�_D�e��w�]�L���e�-��&�2��y�Q���2o�\2���R���?��c�~tD��f��!l�vF�ŢM��
,�Yy��L�/\��z�=��`�������������ΖyҸ��Φ[5�����'�j,U���Ʋ�]<9����M���n�q�8�B�%�Q�6ȇH|z��2��d�����|���j������*Xޭ��+�������*$�M�h�o&8~�un��zC�H�������E�9�cP�a�t�|�aċ�r~Ò�B~�� BAP�>r4(�?�g��UnG�P �_E�l.��:�f��(tW4@� >%���>�"\���!��4��I;.�u=XlxVHYEB     400     1b0�����"(Ԩ�ޮ+p/�m���֏�#�E�����#�2��P{ζ�o�b kS�RS�C���-L$�ñ�4qLRvp����ހ@���%�k�����X�ã�B�ӽ���_a0$��}�V�]O�U��K���?"O�ŗ�B� m�Z����ʃ���3�!;N�u!�:ױ��&}5�Jۃ�Y4Mw�����E�Fg=	4R��2�{@����]J��͘4��?��@M��hEϚ&�XظgR ����o7K�I���]�m�R�^ϼ�+m���Gؿu�}zQmG~pI�S��֗;�q@k�#�G�WR�'�n����5$��7.-HU�T�>!���f��m ��i�$?�yd
)����h��#��OUs\e\H�S���8� �X7m�o��5�P��a1��dP��Yj� �u$XlxVHYEB     400     130��b*q��.BPoz]�#*�F�["Xn2���a���_J�?����5��I��P�M3�2U̥6%Qt��p��[Ϫ9�-G��u8#n�c:�����R/�wz��ˊU2�tY��0���2°�]�9If��@�������m�t ���r����/+X_vl���I����7jP%�nu��� �q���ƻ�K��s�O������{�^��@��f2u���>��k��0��a�I�,L��@�X"u3�>� �d��,�2���o�VU����-AS�mfeObʕ�m�����&�}+��WXlxVHYEB     400     190\Te�+��)%�}C`�
���o9��Q�da=&�1���ϩ�M�{ST�'�J{@�W����+̐6�W���-,{S�W/��OqTd6.��p�}a��#r:��_1Ӭb����n̞q|��]tBh��7v��D$(���*�Ǐ?�"`֑U�\��k���F��� ���B0��lH�Il��ڻ�D?<G���Y�C�=�Om5��b���� ����W<$#E��/D�^���~sR�Mr唱�0�������z@���Z���#֔=1���}�$��ɑ���$�z3^ �v�sLP�vUc�(��N�5���Q���~\Y�����qZ���z�[0�P�mXݢ�^̟�|����c��q&+��޴�3�[L��*�=`�U~�M�qXlxVHYEB     400     160������6�޴�eh�u
�nDa	��قUe"��n�0��g��Pt&�b��Y%��6��.'E�&�T�:�DL���H ��2�v�㧋���U�s�����ᱲdؘK��sa�v��ukK���w�˦�]C�˩�Ѕ�w�n�q �nI��@�Z�����Ӊ�Iư�,x��L� ���*Ms*�a�+	��9>��)-
�U�ӰY�t�<�T~-Ih��_��<S3������uΌ{��i�仅��nF��Q�����7������$@�=��p� ���?l�GO%�vd��0�~�D�����o���� �x�]���Z��="�]v���XlxVHYEB     400     1b0?��R���T�t�=?�2��J��z}s���m�H�|�	_��S��g$��ert���H�_��w�}��+�!�_|�;�ʙ�� �������Xd´�w�&U3=D�%dUn��֪t������g"Gl/������˯�V���*��X(�v�������ix����|Zk�e����xG�b�sI,qѰ\���]�,� qݺ�ɿìPg64R%�<�=��)����L@	�B�*��2MG�DX��ap��M����� ֻ���F[����·�>� Kw'_��rϴsQM���n��j�����J�4B��[�S����S���I��-�Rz�*W�@R�����4��u��޴
�ugϙKB���к[���1���(�ZU�ñ"ubrv4��l�s��9���W���r���R�[a���3�)��}r��]xXlxVHYEB     400     160ԢiЩ���?ĹK�B7�^�v��)��FQ���]C�S�2������껺��ll�w�j��:.�s\��\'�&%�Ъe^��\j�=�;�=ޘ 3��_DFZ��%��HS�h��� �� >BQ�E�:�p�ҶW;L��2M��6���DuE�1MvJ�O�	�O��7DQl:��������T���Z~j�gT���Ĥ]�O'0��zB���e�����`�	/�e��`���\�)g�	VDe��fߥ�t��Lls��[�r�����\��� ��-��˔��a-�S;�l��]����L��rn�ξϟu����&J�DB8D��~ʹ��yXlxVHYEB     400     120���6[�>�}V��y7����3a�uM(F�e�U�
����{C�/�_����<�p��7ή"��0tE��g#�+��*�J�vu���:�ݙ0�^C�"����+�S8��9Β�N��O��S��ο>_ZH�A-R���V��ȉ厽e(��3�'�@[�kK�ȅ�zP����87D�G�y��q�MHS���-y�R*�]��#u��ΆyN��1�+�/���6|*�g��8g��Ǖo_��Şz���Մ��S��O��,{n
�-�=*�7D��L.�$2ZS�U�պXlxVHYEB     400     190����wk>�X7��t���`�5�r��@=�O؜��)5�61fω�fDS�7�u"�u#Tj=�ѲZ�+�V���}(˯�z�8Ɣ�6��0�o#����KY;�����q�����a�t����:ǁC�N���u�R�:�^�U9��VvVP���KO����Dc� =\0�����k뵶+���{ki?��ߚx.J�p��e�8�dmZ�^�	��q�A�/gY������}%e�5�R�s�)�mA�%��;��)S0Y>c#PB姟��=x�0����FfH�����T��8�i��˞F��kzY��,O~��C柙�;+
�[�U�x��B_hֱ�cI�����&Ùb�UU��g{������S~}n:j���-� ��<�x�JR�"��TbXlxVHYEB     400     140i�k��ڜu�k��ņ_�[��:�%LXu� 1zq�IE,�J�;�|�>���Շ;^��&@���u �?�m���EE>��I9PI��n�B���Ҫ��V�#Z4	ãf�����u�1���;��.�
�H�_��g��q�ͻ�T����%�G��f���r��F(�"�ڦ�����oy�^;To
����#	�/`����|]���9�U�[�=����hu�Ņ-1$\Y��!,�٩ڊإΉ^F�b ��E��O������J֔���WY����so����5����A�q2���h���9RF��,����wXlxVHYEB     400     160Eka���f�$�;;��6�/S�f��^V�F�_"��
Z+��E���&�K}e�;�h�G
*�@R�r�Jw�Q%=�6����1 X�<�̖�U4m��77�r<�"���2l.m�o��~��Kr�K/�H�S�iL�.cyf�P�A��V���]��1��ce���!���aqJ�FHܗ�Tc�z�/�N��p��Jw��B�?����1����g����$fZ��R
�2X��%����r;L}*�i@�^�>V8٭���?
�,�ُ�r���$'l�*��J��϶A��@p�6�? ��jUO�Dr��uJt��s��0�AcI��Q�L?�֪nXlxVHYEB     21a     100�:!�u&Q��L��s[��IVm�6u���Hc��[ZiIi*��ޚ�_���n!63~/��bS�ZW4�mcT���v�0C����m�z��&{<�>j�ۯ����0�Ԑ��:�[�[oz��x8���x{�����ǰ�����Gb{�6cyS�G��]�x�]��Q|鴾؎�2E��3J��|�b;�pH��U�H��z�]�i$�f?�H<�e����2���|.0nZ���������A�(�сB'�q��g�B