XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����h�l����n_^Ӵ�K�~�J1��oyZW]}KI��i�->�p�e�c�`F?�h�_s��$�+���y9��A�i�%
����.����0��BLTW��=�p��t�$��r��.9:�_,�;���E͍w�cևW�����<��4q�6�
4�� �8[í����viz�΄�".���HR�L�½u���C5��ç��kz&d�
��~*SӋ�]*^ǉ�on�	�!�ڀP����i��V�Je愪��m�ź��8��L���6�if}&>�e��؟�_��,{��ž�v�ʂA�A�E������v���W�ۇ�!�G0�Ν�����6E��.ѐ�r>�_��C">��)p��AM6���\��0q0�[�bJ�d=�ie t�ʖ]va��Ԏz��HQ��x���d
�5��c�t"Nwo����˴��ʭLA0C�T�7Z-��{��2�s�vB�8�Z�����V�)]��Oa�!�<�:���fK;i�g`�@e}*�7�+:�"����>���:W\���o@��Ӓ#��.GD-�[t����e*U��v�Æ8����(�9e�>�8�䒴# �vo�� �ޢ��m�	�f�ߠ�	@=�瀟w�����>�p�	�<qD�#&�nh�f�?�_��B����C����3�.HR�;t�3��줱����܆a+o�A��z��[�]�/�r��70�o#�[�������ߵ��Q~6ٓH򪎎�L�daH����O#�G;]�#�F�07�l�XlxVHYEB     400     230���2�����HК�Ͷ_s�Uά��H��)�D^���"��\�3?!o��TՃ��X�Ӓ(�>�[h�F�X)����T�l1����
�XG��@��Q�@�s_�G�!���&�ׂM[��f�3��w�J�zs�<��Ǜ�3j����JE��j�����aD/ݕ�̿N��P& �T����T�c%2U�a��p�*�cW;	�p=�ٶ+k�(~��p�54����UW.quNC�8��F&�3K���ـ�*p�p!�~�K�����4�K�0�Q��MZ�҅�15 �������G���jGgoϊ׫�no�����_���698s����e�!���b����T1z{>sA�]������]|�FF�+�>Hܫ:Ͻ�T�7�Ր����[���N�iH�n��"��$g���-!�פ��p\����m�'\�3�W��ům�C�.�l��y�������V��qs&<~/0O;��]�K���f ��ģ��w����!6���g8�q2-�B١N�THOڱ�N��L�j��� j�%�%�����XlxVHYEB     400     1f0��u��Va�G�ע��0����w~F�Ü3�0�c=jCa�X��1VF��=��jx��\ˍ�����,w۳.=^����-�@� ��FJe������
��$�G�g�,X�oK�D��Ɓ�kBd�*NCq�:Etb�D��uU�;��[�Lgx��kl����u+����A7�
[��V׊��f���y s�6�%�}b(D�i���;vB�,����]�����Cؿ�A��oeQӑ�R"�
��R᤼v����/�����cY4K�EX1����zC��cфX�b�^�G�?�{p�7]��&�g�G�B���"C���7^���L�M���\� ���Bձ�=T�fe�I��$/@X&I�����?�At膕~�i-��\��Fuk=]�&<i�>r���MGĚ���[P\-����[��ĘJ�<h,]M�q���
q��:r5�����˰�1IpÆk������ߵ=�D�Cn�����BXlxVHYEB     400     1b03w��2����u4�ܑ��nWT�5�2է/C�ε�}��F5�=s�F����lSa]u�њL����'*����_����{.y�ᑥ�0Z� �S�z�RFJ%w�_e>���qAfp]�3."�F�����MM� I�O�SRF3ޢ}�#9.������?����[�:θ�c��a�h(gq������T'��7Cpk:�����C���ݦ�����I�P�݁�*�}
׉��N&���� x�-���ɘsTv��Z�p��Lp���Ph[�cuCd�(�qU�i��F6�xe�C"��F�=�	��Qfe��\��S���2d&KQ��p����I�j���'�����h�p�x�j��[�˹��^�d|��zbV��ʋ1pIs��:G:��酉Y3���qH�P�fuXlxVHYEB     186      b0����ծ/���h��5�&N9�G)�>S`��Y�5�c1X�����φsǧ�����?�<�k�q�DN��׺�����4��;4T�9�{#*->3�g\-�R�PD�%��6����Q�6�.�\���	�����03B�l�dC�8ež.sN�$[���R�a���