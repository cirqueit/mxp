��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���s��s���L�2~rM� :�e�r�t��\�z2��s�ps�*ܚ���2�{�H���O�����6�X(+��C�a���>��Y.������>��M+9���?a9��Q��y�=m冉��1m��sj�0�3�}S���!j��_�	���Ti=&��+Q<�i*s��I���$a��Ʒ�"�Z���l���%�PY�_�yT2��v��	^�o �q$�>y*M�TM�,����6X��,������4!{�^٪�5��0�J�E�����]��ib�_l�^�c?�"�խh�^���h�K�6:P�XQnos��j�����!U�w@g��R�3Sm� ����Q#5:�:�K7#�S�p�z$^.���_^:��-�mD#f���M�+�F�-B�HZS��x\���|ˈfFvr��v�osn�PV�z��@Dt�\�7�i{� ���wֱ�4�Q	j��R���$1r;$�y�����*���f�ڒ���}��R��c����!8y��O����˟[ul�0p��n�j��I�%��%U� K!��L�]�� OF���<�.鬐�K_�ς�^)j�_.�ѱ��(����8&J��.!�Ŕ�BR9ȵ���_Io���R�r�����v��
��AC�,��5g��G�u���!����a:���0��>R"sE���(:s�Eo��C���Vřo⸮>{��W<K'f;����Y��><���
>ǎ��]�i<��)�_�#�R�B���ϕ��λ�`�;���Ƹ0G`P��{~W���1|߿ۺG��ړF��d{�d����� B:�P&��ǀh�6!�C�x�l�ࢽ�cu��,в�1k��؝Vz��f��_�����0g*�����.�c4�;�������Qε�> ʫ���ƿ���P�� ���*-V�):�Z�H�z3�q��]N�.o�����C�%@�ؼ8j+�'��������ω&� }��>l�@L�w�K���%�����"�x�Ja��<���Pa����U>Uʣ��k�cQ�5�F����N�']zw�?�Xt4�X"d8�>��Zqx�LD4Q������y���{Ժy� ��ӹ�j�\��R>�K�@��	c$�e�ơ��	2� Sω+7?�ζ�kRý�����q���Oߟ
s�/O* ��!�S�N���p�:�A�5 *��/�����xPq�%�\�֚%Ҝ2A�������Z�J�J���Ćj�����������?P�ں��M�aZ�$0���I�gr�Ȱ��Tෲ��1Ð� '��M��4�}�C��"9�����#ᵔY�QބDPZ�댱���U��y��n�eP	�V2��!,����GN��X�%�k �5���X��h����@��	�? ����_U	/����ƣ���.&���1�a�ˇ�O�����?�~=*�u���'o��񞟷ޛY���d�װ���iH~8�D<�J����U!�]ӸIɯ���� (�4�[�҉�6��tq^�2�J�h�/U��W��o#��J+ak�`��kk��6��5D�$DC) ���]��GHym�R���)N���\�w�	���Q��ȋb�SٺSr�+�+������,���T�sN,Ԏ�eŵ5�`T8��{gw˩���R������<Z���<���'z�H+�����yC���U6b����K�������|t�	��m���*֬v�W8�k �^�J�m1�6��I��^����W�Q���_�)шX��Lv��$7����-��Ӹ^���D�֝Q��|� Å{v�<�NM�����ކ�_$h�z��e�KD9O�췏�(�q)w3Q��	Y[����2Ȑj� �M2��L�k�Hua������v2D�@ce�r���^�}���_���zApO/�$�z��D�a�-�س�l��s���/�9u����d��-U>�R��T��7
��`�BC�GKܥ �۽:Ce��)�����\1�0m,��h�(��[~@�Q��$�X�NOE~]�|�J>[���C6O��+N��_��y	�������t;��ۈ:�����/T<�
�oP���L��ܿ�$�K���{��v��ϒ�U�l����hB.�g��Gx�@hWյ�erJ��x��
����1{���+��ai���A�Y�
���"xQ��!=\,��;��eކn�!b���!�[zP�	&�א�}.�Ӹ�a<��m��#4�잕�y��l�3>�h����(M�?����]�:��Euf��պ���0h��	�ka��и�F{5J���k���o���t��ƹ��I�����3�-�!�`��]����/r\Tu'�w��Se�����v����n�NCO{�9�C�4�rƫI�;�)V~�f�=#��^�,��=�`g~^�GG�"���|����eL�(
�k6<\h��.l1�kK~, 3�wq���%����[����},�ڨ�X��nN�ƥv�pꞡ��^Xl�${F��{�7w�š��3�P��ު��&���V��"zu�Y~��\l���@F`��9\T*� �74�3��B7����?�����^��ei�������V�S�TS�W���K/�~�Ӹ��#}�g�����դ[�T�fD7��9^R��`����3ѯ���~��r��&������
�]���/�[��Zl�Q�́g��¿M�R�L�Ɏ��+�6tr]���X� ���M(�,��	m�8��~_��_GC���C��=���8&Z��z����;?;�2���>�WL[%6=䠿>e;���6�g����/U�������A�	c�5���7&8���#��O"���@WE�q�9: �	޴W�&a�ʪ�=j�u���+��_���Vz�*���\����B�'�޾4,�l9��r��0,Z���}�Vs��ӻ_�������8�����K��Y�U�`��zVë�z�Ǿ���{R�~�q��