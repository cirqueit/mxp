XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����*�-dt6'uֵ��_�h*�S���h~�]�%rGIM�� ͜���]����-��?KϭV�,M�N�,m��9pb�i<�u���-�[��[q�YÄ+8���vb�&��]��0�c%S�n᪭�����	=�7����(ӈ�֚1R�6d�00�M����E����w�~ۂ��"�j���$jg��U�DSK��j	��PbW,!�n��_ٴs��s� tf��Kb̋�C�T;�ӻ��b	O��/�����O��G�t��1H��1�v�05*���pϧ�q�����a�k��t��\)ŷ`� �?Q�h'?��(�:]�����:�d��u����L*p����	��ē�F�Т��K�]݌ޛ�[߀1�&Tj�n�u��R�p�{��/E΀�/IN��hCmR�����&�Mc���$��s/C�;Y�i.�HS��O�g��}A�W�����&�J��=F���,9l�j�+�Ν����[�ډӯ�����=������U�CuӨ�SK	��@�����&��ՙ`E=�Ƒ���z&�Fs<�߶;��yG:`k)���ݨ�ŔS���vrg�gb��-�4+=ޡy��j8DQ�9�O�ӎ�~�k�4��C�蘨��Ѵ����2��@��x��`��J��Us���Xz�`Δ~-
�k4�Ű�p��n��mI�vGd��:�	"��Y�Y�ee(+{�f����)֞���^}�D�,���2_�nm���1]��f4,G�鈵Q�̢�;XlxVHYEB     389     180�U9�X�b����o��L�zg���X4e*��;��4gز��=}��rP��8���wU��O��(�_��vL���#�N�x'N��Y�C�R5�.�(�$�a��}��QC����hקfk+}�,��u�ۋ�!�^UE��w<�Vm�&�p׹�xp�F3�V��q�%��/�@�u<�ƾa�z'�3�C�fmcE:`�����
=�0h���9ԅ� 8<7��
�|N��T�䟾�:Ϗn;X���=�>4�*Ij
T,�@l%��և�C�6�<� �>����}aN��|%����3�yX?,a�u_ �~���DH�;��h���E��]��L��y��玿�^Z��I`DP��+\.���I]�dЦ��z�