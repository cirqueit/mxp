XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'#?̯�r��o��,?�P��<��e��"������rdf.��PI�qu��9n���0���_���v�&��v���PdM��ϊIx���c��	�6	7�3��D�j�blZ�r�e0��)k������G�}�ek:h;��,#�A�޴Y7@[[��n��:�[���~��'X�ӕ�[r|V�?+^ 崽���Y��!#x���;��YQ�|�t+DX��?F���0��ݞ��"���J��������M]�PR <t���薲���"=��.�4�ImA�a`��f�y[�'Þ�ń�>��S��(�gz�hԓ{��!ul^���L�*�1�k�����W��̶����Z�Z�:�I���k9kÞ�hD���	5����M=w�C6�]PD�4=�8N(�l�z��iD7). �wV�@e�&���I�!���,�d���D���bT��^�)�`���|�vd,K;���0�񱅓<1d�����̪����e�qV����2'��U+N�o�nө�(��Rv/�nݏ^�d�͢Ubm��z�p��[.�!��1��K���^A�Q;�-�w��:k2snǄ*)6��AZd�$}Y2�|P��`����՟d���a���ĞB:lǞ��I���vp�� ���d�{���e"�08���jvy�?��c�2ɬ��$RMb@:H�k���Ų0W���`��Φ�(����	�n/v�ƀ6�u�$�y��L�� I�{36����.엄7��-�.�XlxVHYEB     400     1d0د�5;�C��ͼ��X���|{5f׆I���}���6�җ�Zv�ac����i���wAKӧ�r����]��4��fG���mA-Z{��o/LǲOa��j�/�ǣ�W�wRm�a��CL�ډ��Z|I��#�yg1=>�!<EΗ��gm���� Fa/�?�J���p��o
��moA��{�FuA BrQ��Eoq�����$�	��|�$�tc.�:L^���Eb�<i��zl����6�I�&��e�����s_f��%��&�y:+0�[��d��}L��'�%g��^4$��ל��487�.$�;�_��ס���$̅�),c �V�7�.�v� 07���|�%{W�*gK%fz1zKLH�W�s����3uO*!a~qw����h{�a*֛`��;)���ǭd���? �]k��&W�`7לyn#�!ī��("��XlxVHYEB     400     180i�*)����Ҷ�5����@�����X��*���.�g)�g+S1E��>�W�
T�A�)�U�:�4:��f�V�x�ڳ��~�i'�ep5`DM��3�x�����&z;���ـ������6�����xl(���|��B���!�2�9�[���h����V���WjE�Q(h��N�&#f�ܴ�mL���"��^
o��#���m�_D�=9H�]Ï���fN93����������
����Z2�8L6��qf-��E�Dsi��q٘�IL���P��/8^��4�Oq��������Q;��k7�&��A���=.U��z8[{7���Q��� ��8�m҄{���+��y}��$�� ���=�I�XlxVHYEB     400     140q���iY�yr.p>�L���Ky�O擹�`o돫�~i+Ǡ����Q�2���ҍNџӝ]h�.�#�۴�Db�K��S�����;8�]G@�p����D���B#����+K���SZt����Te[&�Ra\9��R���
�Q�囷4B��:�g�,��w��c��%}�#h;�����,Q� �u�|�wh(��)E��$�N��������E��Q�^�$L�	w�<EAq�<�q��ֲ�u��Rq#贁�a�e�L�R�O��"%on���;N�Y�G:�:����Q�dh,u|hb�I-
1���{���XlxVHYEB     400     110�=�Z��n��&��
tg3�������d�u�#<t���5l^"��c*m<-�I�����_zkl2�3H�סIk]�3<��)��?����y2�g��X	���y�����j��2dc�����I$�F�&����o=�!@9���l)X]�\���k�
�B����(TrVa��~z�#�� d�,��_x��o��f��������K(C�`� ����n����L��x�:��G��yy���j0o���{h�5�G�~�_���XlxVHYEB     400     130��r���nIav.;ƈ�k��$8���y��]�l���E*%.�ƣ5.$��%{͕6�I ���`6%b��pD��d��f.@-���/U)�dlJ+c�wQ+����}���	�@�Ԅ��Lݫ �j���xWhx�3t�##Z9%�`v�g�d߱V�`���;�,����	Џ탁�m	 kQ�Y�,^[�i�����?�-(��O��:,Dz�5$�^u_ ���L�Yw���-�̡�����zq֯�a��wB|2�M��G
�X`��!��A���'��8R�2�X/��X��Z0�M@�:�Җ'�XlxVHYEB     400     150�����*��颎�$-�0��3;Or�V�_���J�!�t�ͻ8�Z���{ͮ0�W�Ѧ4��|%.��,ϸ�zA���i 9�U�BṲ��o_ʸ����P��Guas�f`�C��̨��a&��h�}sٵf���\k͈ ��� �Gk���A�B�= �>w�p��[@6�j_�o�swD�y���|���^y��j�Ϋ>|;��p=E��q~�2D�
�c��B<�wlp��wn>�Dh��tά��qM��e3>���M�D\u�/�mqq��;�XI���*�����`7��'Y
�%�썞�A�$����ݞ�E�xa��?��i���!g9XlxVHYEB     400     1100�aک$ͅ�ӊ���KA+��W �(��Dk�d	�BdI�-5+�\VI�V��޴��W�-���F}�(k;���V�`���*��`���fwq�iF�;"q�tN��^��G�l��.�<��oB
��U�����߄j�`��e�X��Qף���)����!2���n��օ�v�#��}!\'���C��i�+���N�d���#�V���U/�PL={����~&a��4Q^�;s{U�:\�"������E��.8�c��y�q�����XlxVHYEB     400     1c0f��+D���6-]v��-���朽Yo#��eX��/��*K8V�/�_3�B,�� u��-K�����>9}�f���=gć�j?�P���r��G~9�qoLT�����%c��u8K������|H8(-�z��f�d�Q���2z}�U�b�ߋ 
�	�̅N.�8�NL��(�wȁp-N��_���^�He�*j���֦T����ގ3yN���N�Smrm`��}�i�l�4����m�Y�Z��,Ѯ��%`�.��\��8k��1�c��iM־7�YAbo��ZAe�0ݧ��n���X��.\A�o�o&���*!��,�"�m�6%��H�ca�ι��<���v��EJ5�<"�S6���Māi��p1���o��/���2�����s�x�+ÞC齰k1	��[�Q*�������FQ	7�=��<=�)[<_|h'5+���XlxVHYEB     400     150>2 �_�)'VD�1��;.�'��P�=��KV�vP�˖I�R?<K*��!����#��V���h�b1̔���2���L���mG[cW�![�?��s�rgOs����IT��^�o�p��%=��IFl����t����o��h�;�[�{�K�!�u5���04W.շ�Vq�R��}�A�IӃb*�B*w�B��n���B���#TU;��������6/
���?���"� ّ��0���=p��l��cn���� ���KN[(^]� �����<Y�n)�2v����U�R���hB)�@`~E��Ԉ:��1l]�V�#�3XlxVHYEB     400     170Ξ%�s��h���Zȹ�l`�0J�9I�^�~����)���c����]���7-tW8�9��Ъg��P-*r ���:��Vh욽�W\�i;���oMb�z�� z�L��{^���b��J :�a��i�{��9�ຘp����Д����G�ۙW��҅��L��X8zhN�X�9��l��+�^����e7�F��Ð��'��9�ϲ�i��A�'&?̢�bi�,�p�?3��v蠉Q%���������]^M����d��u�y,=�U�Ov*6#��lmU�(gi���2����ٶ6���>�ZxD��+d L�|�g�,p�`��l!�Q�C�>�2Y~��� wtw:[XlxVHYEB     400     170±�n$�\p��Y?(���3�߇\�h䒞L�e��ST�0S��,`���	3������^/��5�Ly�9�)Va(d%aL�-.��!��1 �D����nd�B����9������1̘y��z���S�d 2 �kd�q��"��bk����f�����-��N�C��W�P����K$�w�i' n�͎�Rhc�}:e�%P)�z�wW��-�!
��w�e�:h�`m;��!xO9��<��(v�����ǻ����
�����쀉$@a=�m���a0	P!��ɖ�ez�K�j��I��E��d�A/W��C/�|�)噏�Yҽ~n��ͽ�{��N�"=��w�C\3	]���d}(?g�~�XlxVHYEB     400     1f02�d�{����{3�øPtȥT��@S�����-<2a-����{��������4}�މ�O�1���q��j�|"|�PI�޼��"D�TK �_�9��N~����q�C�U��NӇ(�#�Xɗ����9���)�SVӶ�|�^�j��8G��'�(�c����/�K���	�j�z� E��V�֏��hdF?M&�T�F�xuI8�����N�� ���ּ���
�����Tz�z1��*z�s�����$q�����W�>�!-����G�b�-*u� �ϱ��<$���8��p��9S���}�%���g�Y��,g��2;&��f��LİH��!����EF�2��B���IaG�1����=Qz܀~l/�0����pw�V��ǵ�+�A�c�F�8��#[J���S��U�-�l��^���K�S3o������C��k/_�i��K����#���*��G�G<��:�ژNN����AYXlxVHYEB     400     1707&�5X���$�2�9l6��:zF|�&���яۆ�U΢i "|��T-WjaDsJ�|�<�����GB��; St.R��ոf%Rƒ}��E���cz��a��>x��2�pR�*���|����2�^�]�X�l6�Vq'�z��֛y4�vBy�y��	(.�L!�"s�4@Z�Qmjcg�X��*0�������ψ�L��[亳J�f��CD��x���J�Q=6@	�?�d��6���#���;E��TpG1O�w&����qJ���!��K��C1��M~�bk�i�(�2R�GF��g��<���%�.�cNE�)����u��m4�-����E���'O/��S]�)*y� Fp~!�;bH=}�q, 	=�XlxVHYEB     400     190m.kQ�%
5�b�~ho��3S8��a���i�X,���rnx[���u���%#�}��˰��M�4��'v����hJ���֪xzgR>�G��Q)��p7�_���ۓ�q��ށ>�Z��}p�<��������u���1a�U�}Y�_����}��
��W%�+P���M9VV�	(TCbD��ǁ�ø��Όy����Ks�� *p�T�!g�B<�Kv� ��Vf�Í��C|h-�����X�G�M,�3��ro9���^!f��!3�J��V��ե�ɫ�a�v��I0o�ud�u\�P�H������%�:�H�G��a��^j8��0ڕb�}���0:	e�E4��P�����.H������U31˱�,?�9v�RP�XlxVHYEB     21f      e0c�~tL�E�]�#���3�Q�&�����{�7L���.��*�V1������}$���{.�j�+j�b>���
�g����=7�8|@��Cmmo(���f1�>���0����n���f��1�3�̠JI�����f|����ϡ�ai��U1��%Z�0��G�gj�L�����E�x����+^XU|�-��Ja�k�S���T�$[�}aX:Q�