`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
3sjK58DuYzSQSkXORRzAuAa5u6FNe2KUmGxs0YOIOwTJUtnoBragbCRY8mPV77eXWdy0LVPbnDWx
eBujrf/0hArPl0B4SNt8oKbtsBWdIS7O52l93aoAemVp58LF8eoU/IA2FsHBeg+noEXpAEZz7dVX
ms/gX+HNdxJve5+Qy+1dEfuJs0mEw7wivMeqifSffRfr6+joh/dBPb4puKKY8JApZNZdnhAmbto+
TOm6PA9VdHp5QJCY4wShW3P7pvEuXCCdosVe3tHziMpQMHL8ssZQe6LDrY9It4CMvaiVuklNXFdE
SXlzvucqVBSNDSqMMsqomaEmd3kdqSrjbI+tmNJPEqo4A3D66Xo52xSAwDmSq1llPVT7dtA2aQX1
W7nnEwDjtcMPKmge/fQrFpKTuiEkWmN2HXHx1bO8MblO575Lm0fnjDx7WXELLFFL8kPETiv/li6n
NClM/5u1fCUvlpAVM0CMR3Vn0v67KJCJnmr1v9bm3IDmjIuuggGOc0qyTWBKAoR1tOog5e1ZJhKH
kxf+Iqvb6ET3JGMUQFsMwh8WkNHgIcLolaQU5UZQA24hGMy3CiHPmepP+COjxkE3tSWK8WD9O5Jq
sb6gjtTV1jp/JaOzTPOj3P/5ofUzeUBiHMuNb8wkdVgAZMsYyrM07BlWqI3ZWF+2/0870iTctIZF
/Y4z+CI6b26O0tZiAykJJttAJifRmTu6K5yckvdRTXlzEyvNjj/i16owFX8buuHbe4VVQfDeuCUu
UpMtp853e67Bg1Z3RrSx3BIRTBtV2blPBVtduBQ4hlMF16w25g33owv05RaA6t5+uSnTg/oBnwPA
4FahCcyO4Ip6Pf15AaFCbRpBZiCGLVm+A+Oqi1wDcLbeAqZ6i1SyqX4bPeSyRzpWSwHTKT88ikEW
gWAvcNuo6bA1rxZkj0X0k4oQP9f01bzdSEFyr0KzirUbyCTpLA2CxO9iAv2hdUh6OZYQyC5YfO7F
cbcDACRIEGmSyrL+vS+o63Iuzr71R5CuToxMH/DRvn/ZlNShsh0oTdCmdCbxcI26euZsSuuiRkPn
3YZZN1u5WSp+iZkW752SNbiUPPFTwCGmHux/qhjuBTa+5LQZ3z2Z8xrCN676evJGNTrmrdquV8bX
aF65nrzl2WQo5DtE7vjapQoLFkA8aXdJTj1aDGFjX+ns5Og9+y0bTtv0El2AjWjwYZpaRzsX7ZaW
4BBO/zjOMouMmDsQoccsCgVedAHs6KCc+ECHNrao3jGdh/QaKdMTHgzmX+07DKquIzUz2HC2GPRZ
BzSQVyKzA+vKQQ9GAndqvbCmFaoADD8pZMd28QRBbGPy389jO01P3eVpFAUvBfj+iZbit5bF9Awq
w2JgjobnaTUxRd1YWrOBtfcB7DBZiedMW/0w4YGynNNr3wpUyz/RTxsC00VAspFmzK+10HxbRIOJ
P1kGvte7VgkNHBicrFFvxO9g729nbp7bHk8Aewk8hwsbYmD01YaY4F8AeJ2CKVVgS5g77sxyIVO6
LYH2qOhN/jvd51jpv9F03mnT3D7GENGZjWMBI4aU6E9SR3l+/ELgmeytpuFjyeRuRGWp/om80ZSf
Np8Mti/thWmSJ5rGuiWf/Y+cjX0vog/0M4245UPqky6MLuNpwqfZ4FOyGEJfFBx1PltdYUbSDghH
9EjQsHVKIzWFDmvl8vkze9HteTE7vP98avhbMjgY/+uZJnT0ufAQIN5oIHKvHmatjLbc1T32bVw+
CEu4aaZhgWeVoj17iviTxaY/iOY5Kr8gALYUg1GDxT6JtRvOmTiO8/o+01e/+S6cFp/txF8xF0Jp
+lIbTAUrZYqqYuy39Ofq7kZXO5pbhDHj9j0gUPThc9JcxMrftflqkq/2TOAaQjJJmCoWiwf0Nua3
mKzYhgVXgHSMOicd4rOpHu5w9PpzUl/nARnmHm75McPEtFXIfHjzpSovpuJf0LFrcLijAis01s6N
ffkqR6I5YAduYEwWrVHvK1EeztwLOfamfNB6CiOJ4H+tz/asSu07B1NEBUL2Na3IDNcsmx4Lt465
HgNwBhP9UhEWtIZODfmo7Ky5/OLYeLttVoydOMrvRmotiUxMTNDZSnxXPPTZKE7g8yQf8VjKaJqs
i5APXphbatEiSyV0h+s2wHAYnoIByhjC/j9UE4ghTFybR4FVVjwNNwg0yjdb/nqauvwBCt6neJB5
9JHPn4UuU7BVcPs4ZNxWO9O5OmCMwq8TBMQ+ajT6+xR5xT2xqzI21pc/lS4zofyAgjeMzHI7zVIG
IW728MPUCTwkxgcldNxu6882KQzQJnX/au+fNlKZmC1fDIsJMJxKr4ocmp/pCNVwYFs6iFgQeFM0
quID6TBLpfjJEtlVT8ACge8n6iH3nzDT+yWWr9+VWpy68Ie+lQ8UQ/n4fWNg0LU8VYYlqI7ziCZY
3dPHpflogsDSFVpcB+MNKRaxfZk+dsEvbIWvYadKM4xLI7bid48TaGoRIpZrHrdaB7Ct1HfA6fie
Cu3WRcs7DPI0iab7la8yyFksIHbT7nV7RsBrPDfRkoND2qLdKz/+9qEhZ997DEyW/N9lYbIhn6H3
JGnWrnTzR9EwwoybIYc8nSgSlY6ssTvHtYIkSTeeJiZiLcqEdfqeOe12koqZ22IxiE4fBDmz43Hz
SeXLUOr/ooKWtM7JWSTu0zo6x4kIc7MUn9Kuh5yqKpSphAOwzEMo+0CEIJ6STC6niyfPIECYKe9t
qS7tkGAGunIffp0ETV+d/7AXA9jVzW4g9D51ECdRWtrYD9ey1wHPDBTyG/pqXq+54cDjzhc1Hrza
E7Aj+Wvs7ZVQ9QctMwY+r243m6TbKDS85c9uk9USs3XKYIZj+ma3dLyUQhdm44WMCAoHjoI3Vmup
agQiiCsj4DBj4+CSo/Le4CmFzokXGDzFipZORWGg3JgFa5Q+gu4cGiLatL/5HXsHmQTG3qLXM84U
aD0GJtrmp7cE+hVEkGahFgEpuldk+oFd/lciv4mHk6fo8vZLSIAdxdhJ170z7tt0kD00ncZrsMLF
SEDxcwcjJ5lOUuoeLZt8m5BweY/xxfgD1Zp3HHo/6fQfyQD0iLv8DuvDPyDwDaPYEOsT2UZDpmBq
FAZcxVbeUJUs0pnUVgbsk2kQI7LZ8d+ifiRvrVKDCHxi5d2+8fDNrBQ+ocrKhKFN51rE9aXQFuLP
O0Z7YkJdEce0JxWG1fL6qNzm3FOvBHu+grCowGSfcRyTEFu7P7J4c9cT9eQzQPfR/OIirC66rNPF
YM5Pwhoe8wgzT/QsW+eGRtwNllnVEfpZ5jmhIC/8MuDHBklnwGXrwzgaX5pencOIP1igEcj9EnG6
eYO88H8V7Yea0TDfM9fa7w/Y0Tfds0Js3esjCaoL2XF0maAt5m79LMmS4gR8W70ZV/lpwwNuBHaI
SCrFtZ1FslmYe66RwJTnfNNPPpbj17EPyNFVAbyykQ6qqToIZYSkmzHxKYRaDPGqKn2Cz7q1wb8J
O0lISCHzLXR8xMt3/3wUmLE3qgvVXNs8OJOh2I2srsNW4thTsqeBhx+ZWmFP/f//HMtxwp+vbPBx
SLIXJwIKVDFnaCRp93mmr7faRUTQqv8YgFs7a2xU3xRC/LDXIA7ol8XDot0ytnZ/0s9QFXBWfQur
6hMNi7E4B+B0mx4VSPIRysnKnHrE2JKkLgMWibrL+WxrM+LlPYEggnoR7CRnn8K85nOtIeSGXXy0
BJNDVl1cQTuxkr+z/y5E5YuqVp7v5r11HBJvMRxjD5CB6q+zfhh5B0XbWTYfqFU1W2A1HtmoykY0
9CgiyasH11xHL/QAfJ6LcrTMIsDfBmWL+vCvy7hnk3Uks1E6nRLA4rSiN3dU34HlsWNcw85ctQk9
uGc74XpTbWkR7Sp8OXkhQX89z2/noDgvsUFyObMAdcfBqH8eX/VFB6IydEUe22SsF017ijAI8bmV
UQRKdb0cPhYkB8QTZqtCAk2jzxQdjALXY8HthZLFxpAUFEq7M5Y2tZBNp14g5F/hghaNj6YXsqlZ
7bdO3hEkFDO76UQFxujPsAnlG88g3/KjLjTjEhe7upfpFt1ptC4cImZzz48UIM/xlTBKUsSa4hlM
O+Vep8R8Y7RwLWG5CCIifVNj92VDNPmdw4QIOa3ic3vtrRGr7hA+g9dEueMUjxTmF3mPOUvlprnn
HXJqzpekIs7RYYClrgMcGeQaemFDJF+rPplMVOrtzISjbc0Qb0xkMbdglrm4153spD+LwvMDGhNh
dEaf1Iue2xFt/LmSTLt90zNAVABUb7UcpwKLKrhmS+0n+5Uy1jCEUs2tdcf6NH6w4ZbqvixA9V/d
npIWLVbAhGFq8CNwYQc3s4c6lr9hH5e1YqDu7OJaPlptS2TudU1OjO43cIzmU9RgDmgRxg9GHYWY
oXHZXg7Y12MBZ9okcj6HGhj3aX5L2buu4DzSvUFoqaEPuFJseLZdgZGi27b/3kSxThXv0xJEnAPr
PKf6B9QD2v/oKWzfQry2NTtv3p8+V4cvkTUrvDMhHRxaCBnW7RqSpSrpQ4zcT6Tf2nbuKkn6EZu3
J2ZnWfhFn3AQ883F9JxYJgkYAlMbZMY4kXHSSR6jsPjKyxfFnzsq5y+gu85w8Ud27+7McRyNUbjI
y4yEiBAly1Gl2tquN/GLIYdnu9PqfHaDDZtL0DVfKOMNKogGtsbeU/m7/R1KSAhQW99VxQ61yH/a
1vn6a8fy69aqlq7ONcudaPhGm6Pvh4eO+/fe5Dx49PfdlUy4mQVdNiicRLT6IlHsE/W7IaLc6pMS
bmb5USreFWLw0RSIjtsJkLjPn6ddilfdQ8P2AkiNlcxMYov7P/FykF21+515xTCVBKI0pidKKEf3
CdQhSTJu2ALFyzCW6XyIcAuCuw5EcLSJbh0Ziwtx/QaEkVqaarA74Ncp+PKQIAs3aLfOqJBmy6IU
y46WEuBaO6N0g+NuWpav8ESLA7iZkoM2WR6w1owIiGi6Ouuoh7x9Ikrb/qZF+r3Ty6bSH8FJcqP8
HaU3Wfrnl7uRlugps07ab6r50ssQYqziwufPiDVaGuNiH5VOUllkB1geq9zQQm/ae0la0nt6gyS8
bL674xdXX5PPa5tvGgFxhYuctSI2TU+x+wrlor7BtXPfAzzlGQTOtf0xj+urNsBmjxUntZ9fw3oc
/RmNmAao8JD0xennjC6ktRU4P5TqLMO61v8at9EVPAvCfNeTA95D8ilv/yQzAAOBHph0A22ZcOGK
/JatD/JahMvZV6qaQ4Q4XS/bX6fnMC/7BZLehXGVsW9wovIJfMCgQ47LtRGiYZcaF2RW6TBRW5VN
78F7tTV1v+ZMpsB2WUBpo/lAW7e7E8GnzGI5FDhsEh8Q1G3QjqRj3u3vS5ExsczYqytx4FB80dhj
nKfXF6K4HYwwGup7HaLKY1c3Qk3aa53nhyFjrbL9JQfNnOg+r5OTjbCCIMjfjtAU5ZMIPWNMdnNf
mMI0KSj2Xiw9PmNXqQ+VpUJ7NvS55jio7mHXVQ/rvIZxlrb5+w7gU4rrmm6KrW8RRvlcUPjl+Y2L
Ve9R+msA/TJEnajSsMSlbrrTPB5kmUrolnkjRCb3UjyIeFPeh5emKYA+kdczRH7A0e8lGUorWGYp
Fi3fOKm+9D3luZ6SvSAg7LuN29fnMX1quWwWTxpRAHAbk/eyyi8q9idtj7vhQYx1O9HbxpXmoRPd
mvXsiMex8cBZWYQUeEB5gzd8AL+US1/etd2xuAGUUFJGlBS41M6WCkQc8fHod/HgKHzVd8yij/9r
klfIc3dP84MLZh3MvwASaWvXtjBY6aG0GYD8Sj16muqAayKXNhEqOeMXygNFaEejfgvQrhn101nH
2UC0WcvnJoe2VQP8Ds82x9zZQmJI5Fpe8NzHrrgPGe69ZdhJrUBIYshELtJGkfuDNWHP0zJfR6HK
k+19KetHUzPvVsWQctubDiFUfjGDVTEhk7LadcCc+SWzMuYoHqV1oqcJZwbf+q5+rbWarjmHwJDe
fxf9UW5N1r0pYaH6rxLlloZUnAkQIJFYWbbJOtkROSr/4nGTpFoEwH00FMipsQaPcaKvmekoqhTd
TR8wiuNEOZRgdomY5QCWEAPQDp3SN2FeBWQFRHMtiHQ9QOzJagRHklDzuvkTRpANOdb2gQ5EMhWp
deMtxlimC9AvqVR+crfUpQN5dRRTuHL6LauAJvZEFq83Xon6m+yrSD7zfVE1ILROD3N/T8n95eMc
DnojwF0agUzXSKrYYhuO8EEicWo50HtZjCV9cT/HF7MtNFNmz6VoiubTpWN/3JfyxQO5OT08jXZ2
9iQAg7PQTnxp6CueJToyByvrubuKYAEkBLobKgnhxz6soGx0WCMsIWvqmsLOOf0bVKZPW61HV3sD
qIE8yFg5U9bJWt1cqppgp9iIZOthwrIXjMad9kjlJhGyhTkVH4BI0G6RFTMy5NYDqN8GYut+5zbr
QfYXaAFQaS3xNevHB9uhooZZRPdH3W3NiLBkYIk48o6FugXqOr/053iuIzFytYREr95Jietecvos
QHujT1qmwEl6MKk6Xow+jpdZAJRWTNs4frmEafoe3IEOpGvQjOeDJ+JksPOfLFqwcg+lFBcbDFFL
8VZqLNIVu7pJc6NQII88aEJZ/Z15QZba+SynjbwmDgG/xBoUeiMXWjUdCliah32rnb/sGje5MpZ0
/YIQ+VUayfbr/hAPb9myjaY5KlZrZeCZMDrdiCr5YxQiV4BwAon4Erpm0+LFYccj/XImwLv6tSoK
dgur4wpn+RTrGvQxOGMhbcx3aIKhdeynjDuMViZYixV3QdmB/v1JYLf9phlhy62MG1SS/8bZMDbv
mBezn35RjcPuXqIXWOMaF2jyi8nSZ1R+5h/3qFp9CX11gLHROqX5TgWWC4CoryZCyyoL87DU+SgI
bmqv3kTqdaGNEegDbGVSwCCr4VbpNHt3D3gDlTE+AXKvKRj+zsF3RXzeP2mDHkyYDnQTw/2jHyBZ
c5wlph+nktDzqxcQpJAoQhOv/XvQ8Nkj7DnDe7R4ORlMoFOc5tBako5gIWi2sqeM850avApW28Vh
3hQmBJV+tRehz+IPYW3PclQuq5m+KpjVdWnh8IfLThseW2HlUP6pb1WPaybkzRQ7Mf4U9Q6mA6gQ
1CDBaYZMMLwRd7tG4D5usVtaS9wp/8+42fklxzzel7OigqyQxGsAhMxt3VJZI0OnFnTutq78rAMJ
CPG/+E6Rg9sZ6znFmVIh+zcyfL+V05To3ZuFR3g+lDtMgbqGHB63XjQN7mAaZzmInKQ8OkMVJTWD
35kr4sJz3zkik+0OB5B7Y96iRvEKr3lBj0nkBlxpMG3q4w+xoeiNlKZvwN7Q8ECpcI5xT9fsoBKu
rga0SCyKtK7cmIEXORlRcN/VqGfuWImBUOWj6NO2l93ByQfg6gm0oTfBt3Szk00W2yrv7Y6YknQq
mb6PQgoNTSRkiKNTw2wVpb8zztraeVD4S6+XYBy1YxlfMtBcX+C43JLIM0P9vOv/bD6Mnwzi5whB
xhmVJYSFg1uElkBABX14Rq1BaYO1tmN+IL5cD6ROhynE3cOSIQntmTIAekjbquvdx3bfzHyid3v8
r0t8wiIUEI6TG3bWVYhj1sU+iIm0kWP+q5BnrpaULIUlRTqItdjDdiX2h8mEoNbpCVQnZtYlTcOn
nP/tqCom0d2m2lZJU/DHpkPblTuX0v9oo+vsYQlmt8SWa/EaTTYJIQBdeqFrlCyDr8/9jT4OLTFc
mmOfafck+AkG0yJK838i43RjJ6shuzk8oWNOMHHhoz9biBHZO3jIB7jgD980dnsBB7dfznQcVx9F
3wNDMyOhvuONcjIbuARxEMALKIAxJXrqGZjGZo7f9DYURqsUuRAO87QIOtKWqH1g2GZu7b9MGbWi
vfRi1H7vL2zHV2HeJNn9+XiGNOw9sETkJLBJV1+25G5tn0NoRXE+3hXoX96KSsjfjRCNiChB5ts1
eLJOwB4X/UEB847pdToV5CXxmJg20MD12J/Xyd7ZYvVIygkLjDRATiL/IQWWmk6P3xscKnsRNjVn
Yx34Kq3yrfhnQcA2gbYq+B8DGbxkbeIVU5Nr0CyCv14vM9bKUe3jdylzeiBPXsAqx2Zdm6a+7Hme
P7CLJkn+kXcJLYjncVUxQRyKQtCUOa+dRHESc+kYY8GFsZuNyK0XaAIWGB6xvksx0+Vwml3cEfty
esVgkG3D5blbwk+BPiaqbCHQUEVK/8L9nDFQ1Y5WmmpBQrW3dW3njRUvC7l4MDe70PfMlzjW46J9
1s8VGKIdaYIRiY8oYt2KqhvVBWQAsk36VXrlTBXGuGmxXLq9OSJRyGEUWw==
`protect end_protected
