��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���ؖ�Ә5��1�b�0�Y���xǪ�(]��W���3j||
�p7��b���vbk����L�R��[�'�a|ɞ�0 8K_�Y�w�Џ%�Ɋ%G�7�^�F济X�\s�)��Utl�7'�l�Lm���%�?�9�o�"���F�������&-.U	&�gCk��"�>���@��zR0u2�i��T<��=�n�_O��������mI��>T�XX��_Gx�x�q�=j'
����v�|h��vB�� �"~�����/g�r���\�Db-q�V#�ܑ5�`R���	'ނ�ߵ-g+F�(�)�2��ɛd���hl4�ME�r��,<�q�(Ojx�mݎ���d�D˚���J�F���s����+ �*�s&���?��l)�}\>h!�R����	ukTaW>/�ՠC@E�܇[�/ה�T)� �g&���쇡2^t{���Q�8EJ�`WR�g�j�uq�� ��{�Ȭ9�6�>nL�S�K���̓��B%N���M['<�LrބCw������#��f�ɾ�S��A	K3ZH�#���#���y�crUǱ��<(�N�||�k��c-��9ʷD�[t�b�~��sK#�YI1e @�㛈.�uQ���пV���j��lyY@"�
������J@�6��ҷ��{D�K�2������d'� ,��D�O�m��,�g+9����B�H�gJ����T�qʜ�qC���L�+���j}�l=��^7p�sw�O�Ňq-�����n0���l`���&c��mF�UU5y�+�xuΌ��^���Y����c��W��	����YX�o'9B<���f�U��ݶ���7��䵨j�t�{��2����e��Q����Xqܤ�4�P���9�X�k���7L0rXd�#{:ۤ����¯X���i=��f�D};�F��w���R��):j�G#� P
�ͻ<t�&�I��0l�x	E�(t�G�U�7�כK'(�����a��Dи�"J�)�����.r��Az:$�U�>s�jv��E��."N�N���ً�lA�	��Dl�����2����9!jP��6����͐b��!����L� �1��b��G397Ye��Yk>Ui�G}Q0��i�Э�{��;��W?��D���u�ߵ�RG���Sjt�L�_�4�Pd7�uDt����8�	ح^Zr�n��6��>�0��U� ݣ?��3�9���	w�9j��{~wKO�'9�Ny1���\(k�^r��P�ɬ	���m���Vv*6��c�r�������#�n�������6��;�	����jG�$j���rMb�'�%1܊�۾K̤�#�[z�AZv�xZN��!t:tAfgچ�D�F'K7�9<�2ǜE�{�����m�X�:Jւ��@��ڇBNa����-G]��0��]���4ᑅG)_��=�n:a��d���5��������.�I�ͅ+�d'k�jǙ
����s�4O_��3�=w�I\�B%�%_����v�o�ٓ���_��	ӕ
��(&$����n>�����I	���ow�����={pl����d����i͈��yzx�}e�B>�]��Tm�3�z1�UDV��Yuz�lǡ�&�C��*�b���vqw⾾B�y���W{�8���Μ��o�1�Ͳ(��h\��.�_fʡA$C`�7��Me���
8�X����Ssɨ �w�7�n�z�=1%:����`H���1-�.S$�>f���W��c1�0a-
G�%�6n�֥��=��i������By$�$���2��I�G��Wf�+P��Nѻ'�x0e]ݪ����@�A�hgw�O�+Ջ�ԃ A�~�m54�����Z�J�q���԰ks��EF~(%)Kh�l����.5�e�'���vV̴fW*��}�����B��C�ܟ��K��a��FЂf�E?~'�)��xCg�1�k��RI�x�����l0�E�SC�
�u��
E%Ӌ�ى�����@SS}Ta�X������Y�#�])b�J���ce�w��	�����%t��o�]F���C�E L9�8(M�C�Q?</A��@!ʥ�q��}�ź3��C�Ͽ�w�c�.�-
��-���<��mKI@���S�1z��z�W���4I�����`@b�ZIx�������.n�T��T�iJ�)�&42�Dp����>��`�q�K��Ϳ�h� ���X�/i#�����*g�y�]e�4�Å43 �~�%Kj��7�*�6
G�
i!�2�'�X�KޡD
Լ�D�G�%#�ġ��YuA�WZS+����2/:�tj��q��Ͽ�ƽ��Ta}a�-ş���ACg*U��I�ztq��.�Z�ygUg�p�J�
�$~�	-t���gT���;��OY�[>peA���Ζ�^R�K&������ux���?���p�UH\A��4��
����|���ƞ�$��:gro4\�N���~Я;����K�J��)A�\)bD��\>u8�IVnj���k���c�����a��d�]S�~��Ur�"�<��!ǥe!�w����c�}�Xh��$�����pS��<�hu����8ӡ6$>fUz�x,Tq��[o��C�q�}�0�Ď�&/ͧ�[�O����Þ�����@��)p��<�!����(��_Q�؀a�L�o)�M��1��٥�+ƕ58P��pv	���7�x(�3x<EFذ��P$D�"��K"!�5�8���0�z���߸I��(%b�V̤�cغ�Ԡ�҂f��%l��.���zH ���z\�ğ��jk�Wt����`����k8�y���kc���˝EM�X�1�S� ��}��N|@>ֆm�Ȃ|f8����1YX{���e%�b�]G�@Ո��.b��O���f��ǲrF�1��C���3�!v;sA��/3�[���Qe��݂� �H��1�:lp�p
�|3T�)�aU�͹�;ca=k��v�JY����ȹ�ܟ��P�����c��(�rIM�Ƕ7�OH��i�$�3
��n��νT�b��_��'�_���x
t�:^�������_7���R�4l 7~������A�B�)줅���+�ӚZ��� �qy�U|*� ���0�aTe�ƛ�m����6���{Pm���i���i:��5��(��Z�zA���1����th�*�ԣ��|V>��o�,΁��و"��ũ��Q�֫c�/���l�4��fR ���chѐ&;:u�ٸ�:�?-��+���n�:����fЀ����Ôyq����O�҃i�<���O��9K���aH�����I"T:�X��\�^�AR��;�<.������>�_�d�_��ǐ����f�e2`ۜ"z6堄�Qu�yL�k��B�DZk�"f�茼��B~'�ާE�e�<����\<*�tQt=׬�u���(΂i��Gአ7�d/�
�,ejC.6� �+
�Z�o�{���{N:�S�K+%[�0K�P��jI��x�hӒ}3�#$� �.��/��ɩ.>�����^*�
��f����u7�4�3 �=8V�q�ʭ��	��^��.��0�Y�����[���C���ذ������~��<H�&�b<s�U��<j�=�����gJt�=���˲�q�@&�b^��&f#��,!N�E6��^���'�|��D�F����
c�v7�^$�@[�!�kؼ���BO�N�<�|(Z���8Ճp~�0�3�x�-Te�6������'1�L>�H«�Jv��WP�۠L����^=�_�͢d����(�S��d�a�YI	��E�'����P7:���F�+�8���c�n����;��E�����v�MC:��W`�6D��}g"�K���] �D�5��)��1��+J ]�(D=i�D��~z��<�OfgGr'��rpѧc���΀��0aכ��C���������VQN��X6���#N8�$��r�-@��8:��#��R�$�tȼƕ,�C�z>�B?�_�HlMl˹�X:%��Iᇿz��/��n��Q*�Z�n#b�
�L�ݺ�ל.�?��L�@��t��➪���zd  ��W�����0?�44%��3�u�k�t6G����� j�:������}R��Z�-z�ru��Y�;��e����4�C��"��6��Pժ�6�:5���O�µ��Cb{t�NZN��o�����0Q+&�=g>Asa*��PQ3����a_��F Ճ��dw���{�K��4�#���������_�O

���@�-�=�[�9<Y���!����EͩqR�	ދ�¾��<
Ղ����n�l��I��\�e�y��l����{�6�Z���Z�/�(�p�u�=�t}}��~q���^d��� ���@�p�:4�jQ,XAߍ��H�f�����>y�	!?��=F�3�I�fp-/�z{9�F��8�<-t����k��������#��m��'�/��ݠ�C�����I�B!Z����Kؑ��N���|��!��k��H���M�h�$��P��?n�A�*��0�x��Q�9��#�஁���VE��<&�pi%���3)��J7��D�O�:�^��&�++�;���b�|X�X��K��)�?i��q5�s[���vnǿ������EX�fܢ��]}��"�E0S��+\3�o�g�:�e5�-Ј~�U=��/��Nc��zvȶ�����?�Ê�+�6�9w���!6����v0�j�?�Sb 3"���:�#}�HN�Xb�(����8��0����-��������j����ǻ �-��l�A�>hS���r?��)7��%�ZW��K�:,�N
ʍ�������a�ZU�dP�^+I1�I���*���f��wT�7"���M���l�Bڡ��փ$�8���U3�)(�7���̄�YђUw0���Bm=t�4�D�u�9��⒦��K)�Vh����M��g�{�CO�(��b�8�'Z����qZ\�Z+�vG�����m�hwH���2�k����A{�����ol���%GZAYPP��R迼ؼ�����?B0uqp�̸p���,8U`7�vX4�@��8���$�2FM�-j��� ��K'�Lȯ�?�w���r�%����Y�p�+�v�7���Ղ����u�oq#�A�8�qG�zT?!��P��Fg�-0���A�G���gDw��R��ˁ���&,��j��_�h�ݓa��8|�OR���$V*�.�V���
:}�^\g��mA��>:��JE�N�������`%r�D	#<�t�f47dn'ML�ţT�ZF7\�j@�!4X�[�H��i���޷��&�:�z4��{� �T ��D�I�e)��<�-��7��䪊p�)M���9Jts�a����*݆U�/G��KwM�6����b_�5�L�ą]\B���s��9���'��)�4�96�{�V�����ϵ9�+�Aj],�}���3�k���/N�m~�D��1w�]�C2hMT�@y�{��	�5���-Db8d
w�� lcn*%S��-�$T����7���x(��U�=~$G�|�-<�y*��g�A�WR1�TI�+k��k�h�O7YXV�ɤ�-9��j)"Y�Tc�sQw�x=X�v>��R�ߡ���0'>�>����0��_X∃�p�'�n%��1P���z�)���<~�[믪�۱=���0F�%�UN��0���?� �ϚB���	�b-!Dku,��E��5_���/<5��X�,�e��x��}"�=�%瀵��t��X�0�:Qv�f��'ik��Y/i��� #�#�(=�������ޛ!��@�B��az���xw�9�ֱ�;T>�0�&s6B7�Y�{�̣���bz�����sC_�[��q���5�(d�	o�y�j�ά6�C���<]>��s��f��4+<��EIP�Cv��{�;���;�@&��&✙������UfI�A�]}_ �br���=��=��|+[�ؾ9پ���lNZ���Yƣ��
czۡ�����p�6v����Ü�-���9t��HB�KY�8�xLlf1'8+���-�����.��w�+��#b���w�Ul�K�3Q
�����L�O}�����6cQ"��l�����1����f�j'�6���Z]�5l���"n��bŸ";�=��EM��` ��썜_u9��݊�n�Q���D�yG&#`T��6����R��-�L��_d�eERk�q��ƿ��?[$VE��Y��<Ty����a����r���bQ{%� �}`���rɝ��B�p�P���9^�E��]��>xAw��}�U:��Ɍ��°�b�'~T���4'�O7��@T�_�|�dgD���{�U�k\h�U������V��)�~}��b�	N>�z_�b�b�;U9���6��Tc�:q��[�\�M�8~�  jk;m$ȫ�l����Q.q�O�� m����_5���� ��v����Y|Y�~-���O.p1WBSj+_�	\��-3M��TB	�o��En
����Kc.��#n�Rk��;��A̟�X6Ģ)�?ݣ8z���iNݤ�b+�H5~H,TKU��y�"�t�~������ \0��g�D4��:�V��:��L�~w3��̚Ec~� �3B� �Q/(��Hn+ޯ�`�y&-�������cvZ���
�}���I����0ď���u�r�D*��S�o�X���29�&������(���a|	��B�3J*g.�1�B������k5M�4oW)(�N�?�p���^y[7���,�@1����^*-���rݢ�QLdc/�o��GqOu񚦾оA�ɻ����Y�8��ՠ���,����-�������w���X�1g6����q�乁��
��6!�i���ˬ���b'ԨSW!e�dڌ�v�-��f+Y&ӭ�A�T !%D$p�&3C��j֤�"G���],J�D�S�����V,�a�m�,6L�:��~���n��	84mvB�X�Y�q��'4���<�����j�t��y7�������AK]9ګ�+r����;���d�j�k���%W�w���|��//J��<�����/��ճ�{|$�b<C�kfO�N�lD�ү��d�y���K���5��n�K<Q෫� ��B�?�#;;��^��He��>�M�K�+"a�*��C�~�X��sYp&�w�b��{x�|��1��Z��3�M�����\�$R��.ZN�U��_��� ��?{�6��h,�����59�X�"aPup�sr���as<�����O^�F��@�7־�,�&�L��Em��@���=��3����^@3����zo,�v�������)�ub�pۂ��Tf��U�<m�͙�0�$�����)��Aכ;ǧ�v`��`�Դ�ag�+�����uZ��W�x�����>�4��𙈎/�[�	X�^fPN��.h�qi_|�>�	�Hꡕ��+F��һع�I��&C��{p�m����S��/2�z]9�a���6��V��2%%���	�g��P|�B��g��:��.%�]��� ��3�>��3c��������l�l��h�Z��^��d1�:��*��Zwd����N�M��v�� l���.¤6�$��w&�*ݓ�:��p�-��|p����e�pAD�+f�|3	�G~Z��?w��F�FB��<4kq�M�xg��&�?�m꾰"�6�ap�m,̌z	�= �/�K1�\��qK6�4���Ҟ[�DN�*ឋ�!��4��3!��9eg����%:�g�2�ě�t�u��*->s	�ݤioo8?�,T9Ш	��>�EfBx�I� iH83�J o�f�\^md�o3����~W:�MnD~sT�>٢�j%���Վ�f�z��k�g�2�tK"6�%��n���2*����&��ߪ��cD���y�I<y,�w|���˶w젺��B�+ِ��u���lI���}j�W�^?@*�}��Sk�^�ۃ>a�� h����#�ia"�g��i-%�B+H��8u�����^#}֣~`g�wR����ף�pCi��Ҏ������'��]�6O�ǵ-lm�H|�jK{�<c٨��p�׷N�L�}��#��+��Z?wzc�	���@࿨
6��F�w�j��ж��]\�%<O��@� �(��6v^C�
��=6|���X�|�nv'O��T?M�@��22��a�ld��$<����+d��x/'��2�R����v/�[�c~Ɵ�%;���tg�J�8PdDJK{md��t@�}H.(���;�g9�[BT���O���[�q��(K:?|S��:e�HV\��U�;���rX�*���cMjV׈������o���Y�
pN��\�P*&+T�]�%$f&|��2�+C�H!o�����	�p�0 e��q���/j��?S/+@9�fz�n_����|�x��k�8-9���5���0�#]
�HZ�[A0�A"w?t!c��]CP�Ա�3)/��a����P�e��iƬ}Q��ĄUЄ�}��;m)_RXl��dH_lض~�{]�Ĕ1\�J����%���z�˵�m�E��D�0-�}i�V�E� �M ��1�x'h��j���5^�i��̜�2�Uu�SRy���	���ġ�}x��Ɖ������u�w��:"<��>Ϗ3�7�:T��&��������dѦ��(�q��Y}n48kHPǝ��K�����k`y�fb���m2���d��>�W����E��/F�w�Լ����W����1��_h�v��e��^jkF�\+C��f�a���8t�\��o�Ӽ�q,�y�ɔ�Դ{쨘�Ԝ$P������	I����L'2f�D[���錃�E7@�����Q�zv����q]�ti�����������Ή!�
��ٸI�.���d� V�H]�4}Ra�Y�m�.w��UiH����X���q#�
�hۣ�f�9)3=i�D�ʼ�Y����	ix>uD�@�Q`$�4��k]4ד�
��M��,���!F��W�!�4���Y�����ܻZi�����BY^��Wx*�h�.>�Kr�1�+N�@NM�V����b�@�`���j���)��_�@E"��Y(�e��̺inA���-�*�$I��$$���a*�"��sӰ�kN�?F���i�

��9?��F��r�+[����sN�K�#e��Y���<�ׂV�@���������Z��3����ԣ�F�k]��8�dM�Ա�\��aaQ]�����_��_�)Ӷ�(.Y��*3f>ż����r�G0�C��<�yͻ��L�s�b��� �GPL�w"=�78v�fk�zS�t1��������gwR\2��S*g�f���/�r�8�ß:�9).�O��Wq�P|P�ߊ� ����c�V`=�4��/BS%��l0cWѶqC9����/��|2���[�J���k����6�/�8K��6J�Gq�@��կ��<s�
�ˬ� ��9/yT��a�|P���􏇣Ģ1Ul �Hx��	V:�|?}�y�t`H,׆�1�X-�_L���&	)��+�4�u��-�6]�@+.����@��p�� X��t��2�H�	U媃�>�/��{���Þ7F`��`���¶Yw�Yh�2w�h��4޽(̔�8f�ꆟ`�[!�O:�4R/tU ���������h?��P�C}���I�G>�C�p�\���H�ܬ�5'��o��k[b��*x�I�'�5T�$��$A��{ڸ��.��;$�/�9�v�L������r9��� �H!�4;��V�fP�	���I�E
P�7^�L�r�(K����Xe�H���=TM�k]V��K����p&\�Ph�	�t\i�=��nGkՋ��^ezT�J�6 R�ö��:�t�[B�e�w$���$��U7�A�p����Ǩ(j������w�7�J��:��;]J�����&�|�@��I9�S%3jЊ�� У�H���@�l�1.c3�F��߈P�Q�h��<'� N��/�w� �t��1]�dZZ�,}΂yKBl�Q�����0�l��1c1�5���m��F?K��#��PK\�'����H��Ե��5؇�N�j��Ŭ_��ω��XgV�I%sS\�#����m�ۚ�y���ijav��\��םs~�ƙ���(�B��ޫU^��:�卓�~ֲH6TI���Ֆg��\E�[Q5�	�BLq ^���m�o3�*sv�1<�XP'Mּ.2�d��վצtU_L����������qzTO"@N���Sz|�G'̯��N�5md���:`���uD!m4PA>}T�hZ�N�6�؇�[�y�i�L�WDX��E��ņ$N�+m��8���q��dl
Af�t�?(C/D��[~?l����5=��%)��K���Y:-.�g���N��}"����e8tf��zg
%B�9�K������ �yu떐�� fc~����I����um�1�ͯ�V� d.�Զe��&��=��FP�i7��WP�u�J���X�Y"R��z�t������O3?���|Z�a1)��(���cJjh�k���=MXU�u�qoz�-B
?z'k�N�GZ�^��<�_��-�����41��>TQr���RC��+�1�l'ݿ�MvQu5Qfu�9�//���ର���i���H��0v_8�p3X�Н��Q�/�l���X�K�)�V}�]c� ژDå&�UeǸ��΍R gm�X�x*$���g�aZĴAw2�����~��1��rʥ_�Q8?�?����PZ<6��a���a9;([l�����<fa��c�&�U���jE�j�����p?h���I�-��]�4i�W=�?1���q�q�9З�Aj���c�nG֖�.�ĆN@�X���g��ҷXn���W� �ܥ	浞�e�*���o qd����$����-���4e��ƋP�N�p�����4"�
A�����~r��#�����������$���v�d0-ܰ�иIs����)��:?�����"�����'���d��〛���+Ւ��b�X�ЍW9/���p�1�G|_	w�1�sP	����^��a��U|�������K����)�=?�$�[��Z�K`����c5��m$טK&�D�Z�<�Z�r�屌��l!��=b9
)�8���Ɓq���Fǿo�j�f�r��S��Btz�z�t�"&�\�>����TV�y/�A�'��=�en�EFg����߫?����b�5��A���f��!��D;�˦RJf�`�H��P�D�oS2h��'�H:̿���R����\�r2�I���+һ��W���������@��|�V�]��1��Q���p	�X�y�5��p���}�z���a���P�['�a4���Ğ��$�"����'|���շ����-�=/EI���;�g�I�� 8���zr��d`؋��`Xߨ���֮��g���-����#pv��[�0p0�e�I*��I��X[���\���b������g��H]����3q�G���5X�5+bl��ԝC��N�01w5��19}��>I���� ��|�Q,�:A!{�$���'�ʀ܌K����w�Г>�W���	�E��UǾL.M���������@E��	��5l��F��������º���o��{Q���I�(s����5�܌��X���f�7;���p �����	��uM���_��@=`C,o����U���AF�lH�.r۸�z��z��?�ssW�c�z����G!B!����S��-,�g(T��)�.��^�K��h/C�}�h9�jH�������*�*���瘝�ѣ��ZW~}=��VX��z���H��`N�U8Zp��l��2�KQ�lp��4�h~".r+n�olW.��)XK�>���|y ���lD����ڂ�4�;�X^��Hm�ѪVt�"L�����<4mO� �;�ޟ�~n�1 od��J�00�N��hD��
��	6�>F�+� I��:`�9ԉ���w�Jчn�<���梐�{�&x{���;J�l��[�@|�1	�N˧*�G��6�}������=�3�y��l�G�gy�-v�枳?L� ����<�!�j�h}i�g�)C�M�|cG^���xU��E^� �ut�����`n��=�&�Y��Z��EO�:��Ĝ���� ���<:�}F��[MMeM8���`���	Z���I,��\���M|>Dd'��X��%�T��M��K^� ~<�Jd��Lb�����r����w�k�W��N��_h|����k'>��:��qA�o"�4�77����@_п�/�8�g���⹀��`G:}�g�����5Q���9E
��w���t\����:X���nXW%�4zl�܄�94�W;s����6��O����z�O�����Q&8`<�w�L(2�a�Yq����qQ̔�<�c}l�~��s� �x�ߓ� w�Qu�V��t��1�HHb^c�}T���>�ģQ�! _����S'_.*���=���/���DIJLGTۚ�7K��!����'����Y�9���S�.�Z�"��F����oFB�p(�U1��q�}��]����W*�'�d�ސ���=�i,�y�=r�Jx�qbt���P68cv��C�?�}C( ���/�H��J��9n��W�ǉ��B�!J[EP��f��*U�GV�Ɂv`�3j��
�����u<J����R�ÓF��oP�h���K���w��W�x?�i��Q+�i�8�@ZO�@�:�#Hbw\ށs��$�\��Nc�̩�]����jh$��Ǳ!P��g�n�K�#Uƣ���G�{ԗ�U+7��sؚ$� �-�_��&jo��*�?ӧ��5��,K�Zw7�Q�m
�Ít�2�!Y��������JEWU�`ԗ:Ȅc��0A���u���@NlS��Vh f5���G΢ާ�=e�>��x�͡I]��f�54�}�ꒈ6sl�`J�V���iJx��m�����|����ep�������E�q�6��6��T���l���J�׬�L���/�����ʫ{���/��@_��~�ky��D4�=�`~���m�&Δ�)ǏV	�"pY�p�����-[!F�X��O��^֍ѻ1A���Ѡ�D�M�ڀ�W7ځ�SЉ��Q�ɗ	�`p�<8f�$@I�Ǣ܋�35n�ٻQɺj� ��K���1V�5��H��T:�B���n��cy�|�����}�T�`V��ye�bI}�������tL�Q�݅��)'7$	- �r/9�A*Z�Ƌ$�7Ana������_��F���?�݂�P�ߟ�F�D�M�m\װ�S2�b���Eպ�� ����	r)�PRΔ���(w �/�1�h���S�š ���F1K2�����%;���QD8��<H�T�ΰ������j{KY��Lq�2v�7��ܩ��cM/�Nj�8*	rPQiE6|�p���\{��޳�`����y����Y�S�"v����=���0�K�%�\�~�N\�����Ė�{P�'�?���zˇ ���}5��m78t!'5Dn�Ǒ[��V��YR5A_ZԶj|��.N����� ��5�>��f6��^���R����m��n�)��Dv^ܺBr�&��`'X���͐��rVã�$ةC��p���X���^��dj1�5�נsyiJ�s�����M6q�<�e�#�Og�p.�m��Ĝ�17̬ ALS+�#� �Ô��HA%�����(s�l[�]@�&����*8[N�O��`ezq�H�C������Y=��s�udw�>�@K�yvM�r�_H����O��k���w͸u(a(e��`g�����e��D��)���܄����t/��DW��?����Tu�C�eU�	lw5����7�{��iQ6UV�
��Y����1hYbm,���;�h�.|�c+]�B�~��6�MQ�X���T)�p�-�ǿJyr����a�S��}׌��3* ������3�R��������3⚫���T�V
Ֆdq���?s�Fap�8�	������堥���ɦ��l�h�T؀U��Z�g@����~u��sn�83�q�>&E��k��ɴ���/�ݞ������`��<��A,:�?���'4�y���,4�U���֐�B���0���)f~�O����v���y�,�����8?B���t�E.���ȯ��#�H�lv��MR�o�]�l�6��c�`;���ޤ� �EgP�"�[d��^
$:! h�����1*+wuj�e������N�%Z9��oUj膙�_%�{#	_w�����4e�j��}�3�������S�ԥ�A�4�c�t�E[m��`�5V��x�Ɋ�\�X��"E�.�F���2+�R�^/4�9��}G�o\�8$�c���'��an	,5Q���
[u d���P�_��d����s/����>SX�Y��!>�r:��t�L|�y�ą�Oh���cˡYz���B���hF��<�k5b�-�����c&sf�Wh�vslP�W�w�9�����[d�����4�H��ӿӻ���-�q)H�v3pfxoz��²�$=wף:����� ������&�PKI�wk��b.��<��'��D6����@��@.����#��!�і��<�/�"���ƍ8r=mJ~v�]B2"����uf���E���I��C?��?�����'g?����ڏ���A7A��^cw��:��v}IY?�tB����"�5�[��#duz�.�IG</�������&���J��/�{*N%�I�����Ri'\�(����E`p�ST)E�A9#'@�I
����dI�Z��"�мH�E�Q�\<4G������UE�{kU�ٜKz�6� 13e8��/���*ynv ���m���Y��Lt��@���l �fy���×'�arE\�w�L!IT ����0U <�]{&l�R�t�Zy* >$E�D���3�_R�&aL)��n�����.����i�&���rGq��d/����4e���%�I���(�ۓ�)��N�kJ��_�b�~f�j��@�ஃy�!�1 ��,{��;�i����7a)R��6t>U>ܹ�u=?	O����&��Ʈ��/��<8
�F��)k�yn~j�U~r@��I7�M���az��ϰy�,q�SU�:q�c�i�׿
�Mw�n�AT�n���>i ��	����^d��TXr�k|S.����X}� 8eA�?cb2d��*"=�~fc{�+�љ
�ӓ��?R~5�n	�7��Ms߆��*ږ������U5h�nL�a%�j���!9x7n_�6p`��LT���
Z�yYe�^%]��Z�[��8[��@z[��t��yS9`��D���Y�Q���:бb��6�5�P���#"?셡���A��sG��D��oI.����TU��+���Dr\j�r�tJ���t���E""�� *.>�OE5��Ӛ�&rUY����4�JM�Ϊ��� [X��-)�я+>s��o�l�׊�o�.�_�4�<�5:�u.�<�x�8�'r�wu���U|�'$�����=E��(����iy%N���ѕXH�2�"(�%�[T��C��q��(�a>�9E2����z,@R"���¶_?IlQ䎽�Z��tI��/k����
T���.��W�e��a��m�Z��Y�e��7�����< � Zn{�3(i���:�:����3�
��7���Jg�u)����(:�_�@]�����n���d��R�@���̷�}\����L�
������w������%^�܋#ۦ�o�O����d��'��z+���B[?Hn����<�Ӌ'��<�{�p�pդ�|��&����45��,�W�e�3��2��I	1�a�~�����ه7�� �G��-.G�����Ʃ?kpT�[���8���%��x���']�hxa\QT�t���r 	�ꗧ�-g��I�q4< �� !����ۀ�
E��Ku���QSg*ɫ�N�x�B�NZD�h�� ��W�d'�����;}QiKR�%���*�B~����3���ӭ�q�1Z¦�����s���C����Lz�`�ѿ�f��T��KX��g%	8^y����j�����H�I����<TQu���X=m���}���}��k�2�3��̘�s��ٹY�J+d@�F����%�[�{��%�^^����k������G/q�6w�����cM��䜎7y@��z�|{Bbԉ�Ca��̹�׸g�0�Zs����G��k͏fNN)���*�CG�"c)�\��M+)����S9�i��"<ހ�,�3-�z�
�մ8����^���8h����e�j�s(���#9���f�R-3�Q�[��tY,٨a!$;�.��[ֿ�����W7�>�jnH�/�Qfw4���EM4ep�3�u�R����`�L�0J�-D�ڢ�1�ʻH�t�D��P&n^�ּ��
��� 2�nT�cB��Xw��������}�Jlz-�,'���'9�y��k�TVV��m��r�C�em�T	Aj#�ky��1P݌q�iU�P�b���F�����Rs�E�\
��>��c�)95���
|����|�P�*��wُ��4��[��95��U��g��1�@��8�;�T�LP
�\dA���L
���-�Ԗ�L2V�(�d�b:���鵤�	�5��%5�&ɭ��4�>;�B��-��h5%��O��*RK��}(O��(�?����|�O��6ҐN����Fs�#�ih�r0����n��H(ɇ��Bal[N��j"�\k��ɏ$l���I��n���������	���6�k�C�º�#�uKm.�o����mW��0`$X�qd����l����ϳ.���vP-��������\�}/�]�O��-lh�$UH��h\��Q�{J�[��{��(��	ɬ$Bϋ��LS ?K��E��9�w��\Y�<�h��3_�r�?�h蛢�+��k~��p���r��V�K��ezYN�M�y*�`���`J>�6��=��S݉Ω�.���$ U(P����O߇3V�yy����3�'�BI�a%UmխNi�MH�7����4&ӑR^W�_3���csg8��B���������L�j�i%ۨM�qHcD�L�ZO�/E��������� �ɨ�.��c\
�X��!�#��5v�
7��U{��{���E`�����\Q�y �\��ơ�VȌ�ׇi=�>�y�>�v\Y�I���X��8p#�mq^��ti��x����?-�`f1a-�uc�&[uS����4�Y��q|7���-.G�qzB6DOH�4�� )���kR,՗�
TW`�J��_��f5�X�\��F�l���}�<����|�	Z)�F�͖�n0m2�G�@,[_	a:�x���4�Ymc�K �$��~��;��ʋ�,��k�E~=SNUd�+i5.M"�.�t�|��f'�OH"�鱜�{��B�}e�y��5|C�(��W�j���<��Y[�Fj�g�}5����<��U'�C$�@{?C��� ����#�}��A|��	�:����8*%����4}D?]8U�/�D?4�{ ��۫\W�ݡ�:�Aϣ�"g!>������u\�h��6�g2��~[��ex|p|(�C\{Z�σ.[�A�!=Hx����Ia�+Jzg��޴���;Ɛ������~��[�����N�����[�%�?��Vq&�i#Т��Ɇ��l��!������m�R���!���`b��vx�g�������!���/6$��
� <iF\�a^R��i��\V�,E-���������m�b
Fg
7O�fnԓ�.w�@۸� :::��f�^���)���O>�)`���Ύ�2�Z	�YΗ��b l����$���'�Q��:I�������i?
8 �:�QX�#�#��
ϫ�lhz�T��V�P�8#�v�Ug�c�"f�'路�W�n�dМ�O�C��˅�����=XC��b�)��jt��T����;	�ƕr+QKt.���Y��aTg]a�����3��p�G�[���if�8��K��jC]��$����tѫK={>���['M�E��r�{W���1.	��6�3j�v<�/b�|)n�{&3]�ɢ�>w�x�[�5��A��_,߁�b"�_I���a��H�q�^x}䊤��� �>pyx�vq iyis����u�-��Cv52D�h*�ƣ�����>��S[
��+��q���rn����P)21��$�.�9\e�|�_�U�a͚�`������T�8#%|�&u"{�Ǟ���F��9 �� �{b�3��a訩�rV�j����s�V:�q%�҈ބF�+d��6�?��J��̼y����l�g���HB7w��4�K�0'��'.L'�?�I����Q���D����7F��d4_�R����ͯh��f����4�1��+�W�iE�-:��݅��ey�@�v��<�X�f��͆�8p�H?:�G��B�+�7ݴ���{H2P�Rdr�If���<s��% �+�jM,�5�����L��VI��������3��J]�y�ҍ�� `[��p�%�ꧣA0��aaa��&�f�-ip���� �	^�Z
7��<�������@ۮ��+��ك"��h���n��(��~i�G�#��C����TG�|P���2+���"�}���v;��%DS5�.��v>��J�	���=���8����g0p��a8�Ѝ޷
x*���AƉP�yg��jZ�shd8b�
\���-* ���e���hU�?/�o�]4[	�0���ڷ ,vP�b$�p�B��	q�oX� 3��N���W>Xu�Ч(�U12lM�C+���|��, ��yqH%������s���'ê��E�W����P�O3n�T�t��N�^I[!�窺l���Pv�^8��z=��ޫVh�m�2S�(l���m��C�P���J��P`S�U�����B
�'m.�Z�Qg��G��۱��f��
�~s�+��1�,hB������%	�&�&|�d����$����!��b�`����� �i���q4��+ ��n�I{a	��"g��u%M�� &��OK�Fΐ�yX�C���A��w�������^�y�E��T7GK>1N?�"ZS�0���h������R�>�8���4�]z�[v���(d!ٿI����CRZ%~ٿh���H��V�\�����$]�[��B��Hn�?X[����0u<����3U��@�˩p�g1!v�fj C���MUj��9�h�
�k[<I���S��}"�Lt_�2�Vfq�T����e����dU����xG6�j��!tθ� m_�T�$.��s�rS��\ @5l�O��#�Pw�A���Q�-Kƛ�J'�����h�x���E��|N.Wk��M$�u��'���y�l��b�=c��#�>Xw����\�#t�n�+��JVm��4���j���)5/�	��I����(}��)�Q��n�vF�'�"�L���(}9Ȫ�X�������&E�$G�jX�5�I����7d ��a�Z��4��`��w�ѱX�� ��bL�؂���[kɃ����Y��C�?V1����Y]�g�����F̱�?Mdb�oA�1���Y*��b{`�J+�62 w'N�o���N�n�__��C��%2ho/#\�.��e�S|(���'d���Qf�u^A�z�4�F!B�����y�����p��%=̏3 P ��d����9M��3#E���	V���.�=���-����m!���TC�' �\=�vC��Q�ʦw���d����� 칿6J��#��θ�6ŷ[�_�!ĊU�7(�1����g��F����_�x�̦�	po4d��[&�����(#l��m��Oz�+Z&0�	�<�k�$��{���o$�3o�^��Q���?��H��3O�M ��
n��YK"C����{�M+�s�/{�%�$���8Fy2Ȝ|e�L*X�iƴ��$:��Q��v��܇r��Օ�H �l�>��iQn�f=��Y�`1-�FOI+��I� Y������s�2���9T��럁R����}�AI��]�FI�ʅ�a�yt�#K�,u����A0��=�d5 ���ݳ�x�D�o|?��C�ʜ�¾�I4�?���%��3���6��*�n�T�Mm��:(ƵŲ�WP�����f�u��$)Kc�n쑵�0�L/F�h�~����#��h���
��9��ɇ��=�Ffc3�Sk$9D: J���"Ys;��n�b�M4$��<R�/���Y�.c�*S����SS�t��0�<�e�E�CT2����p?�2�X	{��dI>`K"�6�ɋ��}��Wb=�2���a��x����0��Ԗ
��\���l���}Ľ�?�����}̹�t�zh��HƞW��o"j~�c�<}6zbs��ަg x9���vt��X�a�vY|�����Yq��_t�����8�2P��,��;���(������u'݀҂W�D�L�����_�7Tϯ�����%Ik<��
6��`�	�E q#�Fo�f�qܟ�Ԉ�a:�2+��hVM(������Q�g`��Z&��(��&��ڀ�$���{���h���IF9?DI��ޒ���LH5�X	zuF<6�Y�\w��3-ݨq`�# ���x�ϻ���_,�^�u��K��!"��=X�J��dZ�XF|���*�1E
������9	#�y[�]EVh���iҙ��u�^�s�F��ŷth���|�g�8wWC�^��:8K)��m�\/�ap�,@�{����#���F���(�? �uqR3j3�������}Qۇ5�g~
'c�R�?6REp�)�XT� �SA0���qaB�g��I�!\����)R ��o='���U���#SB�M�T/�\d�G�|��`X����z���>	Q�uI��l�>#������Z��L/����5��.VWd�����oh$��U5Z�qS)yDyK�I ?q���n)؈��O�[ ��#���u{aph���sdRx���z�T.�'#`�Մq�@0 �gu���y�pњ蘡�˃��a_&N�Kw��YKV��H�-�*8m�(E�~�w�;����>e�5J�SY�Y��+�:z�g��ƭq	ӣ���
&�s<�|�Y�+I��qc�a�a5+s.��.� �g&X�MRc^���1�k?�G@
%.i'9���\; �����'���X��wz�_���\3�9��L����A��g��,������H��0�1��ɇ��E �����r�${"v� l����/qq�xˢ -�weH�b���N��u�!c�$H��+��>p�t��8��E��\�&v�̩�s +�+Jv�IG)r��m��؀�T�HP< %�=P���j�� �x�����{5 i�|B���㧢�;9�<��0f�d�I����i�E�F�r7�.
�@� &CuI�I9>A
�`Sp��� )�">u��ד&x9�A�-ȕ�U��Lo���8 �s�:��0G�0]�K��%�S`m�^% �Ǯ��L��"�>�Y�:��.ˠ�ۧ���Ԭ&����	��<H��j�6��\Ge�W'�2l6�+9p��Sp6�5�N_hOX����r��_��F��D"����E���EC��:Y��'��ȏ��.'����Qa��m�B���ZrY�3�*���20V���aѦ��.�����F�M�B�;�EY�[Ȫ#Kc:nX/�4��n�8k�q��
qU���[�HÑ��M�)�VR������Gi[yH�~L�0y����%<|�T��mh�bɧ(��ڻ�hH��j$[f�hR�3��[��7�"�(\2��;���=K�#��=]��9?�qW/'9�!�<�Pj?ڼm �~��5�׻�C���d�v��O�,�M�^׭��W�pZ53~W�C���2�^O��J��4���1�FA�D_��=>�4v��N�]9���mW$�5\�Ꭴ�7�%�O=8s+uHi�_���r8._�oX��}敀�%�Ԍ�:D�7�d�����iIPЧ� �e*6:�]ځ��PxKBà�-ɘd�(�~Z�d��i��t(:��j[�8G��۟�a,H���hݐ���MdM��ȓ�%��J���z�Q����'� hn�9�ۧ,�7Mw��9^�b�у��9�A��xhm�Z+tz�����4i#4{O-G��X�o+�
D�o�6bv���Җ����wX�15�|V�d][l7�D���_�5�YK��X�Zu�W��"�O�B�Z=6^}���E�r3��R�Ayʃ�65�QH���
�.jÛS�iv%F����*S<m]9�uUD�J�n��%�;�����Ρ�T�	:��COd4�@�j��]���Qc{���qɴ�E�C���(�(�>�� �s�M���{/����m�1���Ď�O�6��R��������������7�oE0�#+�)I F��G�Tqr����8E�w��8���#��3d�5H�p�'�ň�%�־L� �1�w�Y���"֓�dǊ��|a�����=�8Xm�71e�e9\'S��?���)�XƼɔ*UwWVEWqĽ��&��s3N/F��^���O+����T����=eP�b��r5��IE��augc���2�wJel�׌;��8�,��S��}�A�Q�3W��kg;�)�v����?�������nU6(�q���~0b��!o���~������2��6�qq�)���C��5ؕۊ�]����p�Ƚ/}�_¼㞋rt��`�-~-UuS�9����J912�}x�
�DU�3ni>�*��/�ʜ����]�@	��f�ӵ �(X��:K� >��^mij��l�b
vCєpc��nOuu�X�h{A�F��3��Q�of�`��m��~0���cw���	x^?�iY/v;��rg�=g��%��5 ��+:���קϭ%=��& ��ꔭ��5�����<�d6�>h�L�����{��RR�V�N_�\��I/�󿤒�_C"���s����Bй(J�x
R�.�QPb�,v� ��˥U1��v���Ձ_AT}2����^1�� ۺ0�+��������A�����JՊ�3�wZ���(qf$�v�����P-݂����e�Ѷ�U�rǏ�$�u��z�.��( �����V�k�`|��7����I�����n]R�+2��洞j�
�Q;
̣^sI�F�8��9o��>�֧FrK�Z�a?�B�����.�A���y5��f����lc�^O�Ů�ʧ'�C��fy�k���8!,n�0qtv@��0�%H�l�D�۸e��@rc!Ó	����-���M��X����6/��g��
>|[q���3W?�K�u�]�:]b=��J5}�9�ş�x{L4m#4�da�]���b8��Y#���E�����_� r���}�����G����E��	=�xӂ��X܉�)l��^����}x��A ���F��A���sXĪ��U���>:�����,�#����Ԣh~�����S�ܣR8V���]��Zb7���EJl�x�Z�L3�������F��i7?��1×<>E Ϫj�pFT ��-�
�U�$� �6�?3u�!��J(����Y������X��%}�P!�unN,R�{�+������1�w�XM�I�����ߺ38%a`�g��]vÞ:X�����p�#i������H�1�a����M:��O�<�Vxyɠ�Wd1�*�W�-%�53]%R0/�����*�E�m�z����AFT�&,<­�@ɯ̪�y�}qh;�Ԫ9�J�������j`�0e�p.:4im�Jn��.��!� cR�>C�il�=��_d@; m}.w�̕��L��s��Q٬�&����9�K�Pq,��/X���0}p��;� k��V�����kKũ�LX6��`���nGGʵ�
"��P���'�!ޣ�
5A��������3��X�.T�^'��������)��j�g�*����ҨgF����x#$�f@3�����ځY��`;!�!5�������]k�Zn$Y`iX��jAT[��%�~�����F����d�?���/�1�B�Et)*�C�;qFwS�s0���(Md� C��VG�1������%� �f�*чY�����)>Mr��S~0TS�,x�:Y��-��"_L���8&��%�Cv���izT�=����FE�i�2���r;��g�IO�V��|��˚�����B��nGWa�)�����X���M�ᱻ݆#���*����L���4/r���|5��p}4?ʄ5?�H�K�n� ���1���$I��=���"ߡ=c�[��]�
���s�z�`���EC$?j�Bj5��,��'���}3H^0�j�}�έ���z���Ɋ�Y�J�!ج����v�|-Zo�؅�&�vj���Hg���b2���v�Z�z�n��W��S���H>Q�ҷ.�����$\���Ε蕢`5����-��Te��}�8�;��ʌE�,�Vr��~څwȸ�'�ǘ��v�G����pǸ���xe
#jޢ~B�K������`u� �.c]�pWO��Ǯ���m2a��zHEAc�&�{?�m����<��[[?��e�՘���}A������`j�W\��6�;��٨�9�l
�������� ������c�K//�	�)�}P�j�p&���s%VV��λ�:��ĸY�����7�H׬O����e�6����88޺�����>�^c����"��F�,<D��3�h~��' ީ@�3�H�����r�B��rEx�� w�y#���4nURœ������1���OYw�広>/{��RLC1����Za$����̨Ԉ����V6�)Ԇ&_V
Wn���ٙ���R��J����j���*g1n%ƛ1R��>� ���C�.�u����Lo�ѦCR�Y�˚n�]U���!\ϟ�D#(��Sz��&���zd�m