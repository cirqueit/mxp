��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��������wTP�QY1�M��^1_��Rrz�-fF���`bq���7U�i�]��f4����p$ ��ҹ��>��dsuRYy�9:2
�2U
��FO��2��ւ���o;�3rl����'h[��z�&Ln���>��+c�����4�3% /���A�vB8�3�К/ژ"T��` �-�$G�P{�e��Õ�\D�=3�x���s	��c]ܰ���0�kȌ4�!xkZ�M)���.��|���x���Lݔ��2`��,�yv���T�E��ȞB��rV��,���^�
�!*m�{s4�j�QPP=
�58��3s_��rGS5׆��H�B�B��{����#�����X�>8��4��~ig/bYwj���r8
���U��i�!�u��&8�Z6&s_!� �qh���A�1Ļl�VW�ѓ6p�7���ɤ��'������f�<�v �cyQiDls.�	�ѧ�gf6`��ny��mU"��~w�:�~^,�{ i��X3t|�3����^�s{_n*��Yg�c��1�>�r���|�z��r�,�4��rT������*���4�B���"�S�,�6���8g���Ɠ�f�-pB)5��edι��1�[�e�p���r�+��j�/���A�N �Ϡ/�G�M������;�;O�[��	3{�sI%��0�|��/#o�m*53B�.���Uix��լ�CmL�/�x������9�\]�LQ$�~a{�`wD'��/JݕZ��m�9a	q��xи+���{l;d6��ћ���F��f��)����:]w���pL B��rthVOˆ�4
�_f�!m��՚'}P8.b � �a�W�<��9�\p-��}'ʥ��i�6N��˔ � ��o��D��?`r�M�Ċ�Kj �͡�G��K��%J�>���8$H-?���9�%)ڽ�ݵ��
#m�8�qa���y�<RRF�r4}����r^Y�vu	��U���ϥ�,+���PmŒ5��{T�g�30��җ�N�?��.T�I��̟i���q��G �KBƋw���[�8҄92��h�3���f��j�'G���_gm:�Wv"@�z�\L�2}�-�.�=��-Di1��x�ƛ�o@�M�A7x�����V%*cvs=!=�Tq�:�`R����3;�r%�ŉ�|1���t�ˋP��ōgl�>����d�u3Y�?l���������d��_��]���:B�'��q��R�Ȯ�䪋MH^S�GSdɉ���4<f��AB���p�j�0Jg�-�]2}�Z5o�B@��Z)��ll,�T�&�`_�Yyv��c��9�%���W�����k?m���VP|\�us��g��)����-Ǹ�
w���ދ|�/Yg"�û X6C��T�m�����07q��)���i4��{�}l�����t�]t>㺍Qje���ҫv�G�6-fy?�9-Xn���a�5�b�ڣ&�IT��GF�Ym4Q�'�m�Ā����9�ʰ���/2��o�m+�.N� ��Q�d@I����Ne�/����E���	˷�Jr��q3}?�Kԗ�Cq�	Z���9pJt�[0�"'�֢���3U+Mm�	�N]�/H�e��ua����0�xt���rW�)K>W%��/)݄��~k	MV�]���.��`y,x���&|<�/L��4IK�p#�g��0�[�Vνbޢ/�;��!��9��F[ ��Z���"i�!Iq:m��I~��Y������u���|�h�?8���nH�x��'�����@Ը�����*�R�ŵ�ل��@�S���1�!g*bx�S.g ��:fIjz�X����}�ā�'�3ޯ�<Ex���/�� �2����u--�[��w~.;��y$v��J��76��� �uJD�9]��ml��(��Zz���x��=�[��h|���1�|!1z�}����X��`?�\`���̆�-��?`]���;^\�Ĉ����R���'���T��u�;7Q�@�l�8E���f{�'\6V��MT�4����x�Y�tO�C��!��4/�PP��=|�yA�{�Jd%��$��l	�~�;�Ө�X��6������M�+�ٌ�Qq��1��7�(���A�q�l�}f�o�ɔ�z���*�w\��t�z�֕�`���2��a*��3Pt������	Э�-\��X?9U΄�Z�؃��/Tx����4�*�J<���=#���7�h�
�h��́Q˱�Z]�	_p����hq?�?��И�yR����L�n��k%�/.bT��f��Ah�̲y:=�L�R�,UL���8]��u�e\�z���x��&]����ل1�T^D53��I��<�xs+g�!�3�x����L����i���"��9i�>���2�w��`Fm�`t��#g�u-����_.��2�9�f�+�a.����w�ѥ�D�4���B��*~�(��S�Ph��hѝH�ݓ���|���0�/=~ƙ������z�n���=H�q4�#ل��q�a���ыf+k�<_τ�b�xl����4�α���=�<h�{�!�@�����Ⱥ�;��ΫJ;Y�H�ق�
oL�E��-z�=M�۰[��4L�
��"�R�g�t�Z������A�d�$I��&���,mĔ*Fbj��.�ΐzmG�qi[��m"e��ԃ����r
�; �^��2�A"P7�$�����.̘�Q�?�~JXWu�����J�`w jL��RU��sq�v�f���HL��<�߶�"�+� �fҒ��2���1�� }F�[�v
�\�a��i�~S��3�=+�a
�w��I绁�+P;��Xm�G)Oc���/�t�'�c�7Npw�� %p֜�d�jT�s�)���7��
!����q�k�c@�v����|b$W�wHd�>�8���#�Q����s�/-d��v��ÏA�D�S�ۇ���ꙻ\g��@8�5~rZ��f�_��Al���ɭ��b��xt�j�@�2,�/�(��fE�	3f�X�f����$~c~�ː��M���gr��7��6�\�~��Q@���aeO8O�S=T�W�2�X��EPV��ɧz�
������k�+�t�芤�
�~��,�L��s��2O"���	�3�	���-�U[1��>��C���R?�
Ƹ&�
ز=A�6"�1R;R&SZ�o�Yk�RoUsLdq����튂b��k������]Zts|[st<_������^M�
�+�3w��#C�3�퀖�*XIU��Qd/	��7�8�M�����k�H�#^�kC�j�|��Q��/�Q�1��Nq�_�:y�Sh�_�I�M��k�P���0u��/F)`wj]]���E.|�m���4ԏ^:v�H//�:���{�V 2����?}������zuM�y�>#�{������r	��t�s�XTJ[0=0e(I����q�
���d�~t~!)�ၒ�S�G�=~c���/�/�}`�[�l�F �{�yX��|��V#yy������0>�1&�)3%�l���j���wE)�"�[UՀ@�	*�C]�ϔ��*k֫Ȣ���� }�<�^�A).J}8����aZ����a[z��{�GuO�~�:uB�!���D����Kx"Wl49�֟�3e��1� ��R)ԔWFh�G<&�Y�$����^����&�C��\���Bm�?��![�6CL��D*֯)�׳�����v�!�+g6G-w�������"&~�aJt��P����-��b)��ݝi �3)BGj	�@�
�lʔ[��`���H�405*k��r���(4�"��f�J��i)Ј�C��H/<�W\6`��)����;kWq�
��G`�Nf-�j�v����^�ypx{;g1�aA- ��l�=��W�zW��tD��,sCu���������qp�3R^S;��1j������F�g��"�#���JT�,�dF�����^��s�W��#���7>sOK���eK����%�t�Y�o� 4JY��]]������c肌Ɂ_>+����-�O��f&2�E�z�������M9���Mw;�6�f��:�&�q$���'Jo@
���B�N"&>��IlhR����ь�\wߨd��B����Fsuu�W��yM�,V���f"�A��r��>�u�S�C�y(1�0������C�\3"v q�i�)$�B���7F��,3�����/��̎��$��X����5�mm��\.�d.Z�M�#>��B�s�e^���Mߕ{`2����N��=��g�^IeC���B�������YV��&�ȡ�:.ƹm.�e��6� |���Մ�kB���K����蘦q�D�&�4�S��
~��9��1��/���5���1Z�� _���r�����4�� �C	r`]f��]�g�5��Lz�U�K �6�m�(GC�h]��U�]�i�@��5}�J}:��.j��]7�6@_1b��C+V\W�_�|vmsЬK�>(
�R�U�@<p����J1���]^+P��ϙfO�_�KJ�*���lEL���DN���}$��������m���������� �wR�E�bbp�P�hvx�8�k�)M�Ɋ^vY'���+	��kg�!�:L�ns���of��MK4�RVx�*������@�n�nE���n�L�a
w♟�y�B�cB������&:rs���Iň+�&Vd������r+G?���m�5{�����lڻ1AHB�FGZ�k�m��QX�VCP�M����I��-z{�3�rV$k7 5�ʚ園���i���c&#�,0����E`��_�]Gke����հrd���K�U�JS��(txG�@��J� ��*[ٍ�Ar���-��S7�Y9^�j	��پ彉E�1�an�-�X&�4�0���<�����<�l�%9L��M���Ǎ���J�t�%^�� �Y� i�\�),�*�s��]��)�����N��`K��:����;L�̵@ѫ���峌���D_��΋Vc�%rNt�	[��),��u�K�����w漃?�!,�?����7q��x�M�e����m��������wXՊ0����#��A���g�3�H�5���W�U�kѨy�{� ��.+�.��(��J�_��<rX7�M��y�ԃ�aP:X<}�S�T�C�7�#Z;n�P�M|�!��������w%����g?�q�w�>�E3�6������-��B�Js�3R	�p��Ƞn]�)d6c�;�zϑ��Uv1��*�>!�v���}�V��y���W+��q��-H�+���̦��ۖ�j�h���n��E1'�% F��G
�J�S^Wu�&#�����yٷϹ3X���p���J��A�0�.r�R�O��4o
��z�'nS>�M\�����W�����G#�Sb2a�Ǉ�d#�g���k�.�Cc鵽6�--���}��W���Ұ�(�DG���vi�O�Q����qb� :?[��a�_e���A��c:ɰ��W]����_��u�1��jc5��*��ל#���S������cT����K���b�!��3%
�0���"co>9U$wE�3�}>t_>�W�߲�8,Pu2� �I�W'�FD/��|�gE�@��:&y�V�\N��}�|'?�5������'[�v�1$��8S���*o/|f;n�V�r����Z�'�_��LE�"v(1�R��8>*𛅸KG�;�G�v��sA���u̦nN���o�=-S�ؒ{�fϩtt���M���k���<��BIU���D��������?��z���aV��l�zcQ~�5?F$�^LS��Qs�W��Z{���q��)C�?J�J�`�%R �*�=�<����N<~��g��o�������G���p�)f̗���I�r����}���PK�j�Y�Pj�����>N�S$)�^�1�[E!��H�.JY�