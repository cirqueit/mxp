XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���\$�%���SY�՗'��q1H�u�E�2�P
��I���f_M<.�)�5V�>���?z�j�,c�"n?,o����>��ĭ?'d&�ZZq���C'��q�gi�+Oas;��ҵ2PÏt$���8�'|l� ��Ŭ5f��;{c�����4>�L��Y�����+(s���\<b>��Sxdy.���8���e~T�f�H�E�M���:9Ly��62i���\�V�YCR��sܙY�|�J��:X�3����C�5�$���*�/�1��������PĦ�`�Q}�t]���{� �8*���L�0�H5>m�H%et�t��;9�/�/��ڜE���󙮗+��I�`�JQ#u��b��1l��'���iX��%��5=�"'C��td A����������'�Z��N���n*pǑ|�|�.�i>C�QD�,�Od�n��g����a���pNA2�nJ��V@s$�'���q�S�!��yر%��@�_��;��|�I��W�ahcZ5��bM�6��a|�$�S��W)b�J u=�g��e�ub�F~���J�DM����x��-���$g�ŋo�r����)�380�
8�]-q{�fOe���ޫzr�ɘ ��6ۺ�TI&���,Q�p,�ļhr�/���,e��nh9{8"�讎�A�~���Ckx�[31�	)�Z _A���J�Nn`2�Ȃq!�;ԥ� B�`�՚1*0¹v�8��_�m�Q�4�1��T���XlxVHYEB     400     190"���u%e��"�\�δ��Q5:�`�lq���C����9��)�������w2>��3�3�=�oP��.�hD��,?�Roֆ-Cbk&㍔gb<>j�"�)��rm̖YĥO�8Y6�j�ȤG�����V�
ZH��H�O��L�x�=�Q(oy�M:��%դk���@a��Z�rX 0y<y�=/2$2<`��ֶ�+�5��k�@��h��y^���#y�5n�����������MG�I\De|�O�63����i�S����d>	i�u����{e���S�6�K"�Y����$	}�/�bϗ�C^�\��Q��?��S�ik�`8�B��z?���c����Kˣ��F鲊q���@�*��O��?yIeA*�A8�yZo����f��ր�Z~��XlxVHYEB     400     1f0�3����y�U�H�G]��?�M�P�C����K]HK��	pq͠x3tN2 ��'�����4�g�i?������H �-���B�@��E'��b��q�BgQ!��ϩ�D :�����S��\�����e�F���M�@@K����-�0)J�٠dϺ��VG�%�i��<�N6G&A'�	1�� 0�4�)56!&����"8*�?
jN�� ���͆����~K��|��+z�}e��8v�ng}oOH�#/���`��H�67��K�?�������v��Xh�$Z3����۝�52�ߟ�S��Iه\(m�s:���hOb�z6�*�k�Vn�|�����k�N:S����#���\&�!��ڢ���ᄿ��%DAaN���v;G�@g6�r�+i�x|ep1H����"a�=���e�ݗT�3O�k}c\��Ha�?0������M��,��!�r�E��=�s �$A'Pp<���8�Y!mXlxVHYEB     400     200J�6�	F�R�@�2wU�����GO۬`�@c�X�pޯ�
�u�!X��d�C`�0��Q/��A�~�B��T#pj񊩤�p�$@�*W����8_W�/ל���
�V���1�]軁bӇ��E���=�QX�Y(��.�u�J&��F|��9��6�fA[�������dQ7���,�ݜ�G�Y�h�b��<N�I(a�
��d�c�7v��^�;�Q���uk�U�O1R?�����\\��Ē�[������?�o-q�Jδ�y�>��.�	xa�s����!!
��]�p�K��д�rIixi[c=����������wC�)�,��%~Uu�=����a/��[�ѕ��Ǜ�'���GBr���r&���E�4B��x��_*���W�1@��d����d ��I����2�G)��DT��%!nޢ��8X��#��R	-/j��6�iDĢ�����	�} B��/1���Uy�o�M�f�cY�����.�
@�a�n��ՄXlxVHYEB     197      f0s��z�wFw�b��C�yฅ�d9!�B�\��>	@��^�b���"NW�=���d�@�@�
^�a�:�_�~|���+�HcP���8�%�a���z]�O6g
�S4N4���p���`¡��p�Q��taP���W�#b�L\(�������K�I�5������tR�!dl��BRZw)�O���v��WD�7W-~<~0�֖?jb0�ZfcP8N�{mSꮺ�E��IK