��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��ЈQ�� }1�+���E�����u.�,� 5�	���@���E���zMj�?����&E�΁��E���1{%~Tg	\��/��у;��W�������bgx%���̜O̦jxŗT=e���ƺl�Π�]G@B�2Yu�){�SH��P>(����*av[�c�J���&�:M�J��M���ItEU�V��YC+�m�*�T�}��<� "�H#�h\���C�1�VC���$��OY\_oG���>�_d"/��d�& ��F@a����}�3	�ҳB���C�<6��/#�o֥��\���+�g"�2P�m�E�2�G4 �^���`�k^Y���ld$�f�F�a��B�B]R��5��\
��ܷ��Dc��I�8i�2sΡ�V�p�9 F<+�:)	,bj�}���#Ҋ��Ѝ���T��f��Y��!_���jK\������~�AK����00ͫ�"P��ka�����Ͻ7���d#���,z��*���&$g�n��Y�P���ٮ���?3�k�����v%��q��Y"V{��\ئ_�!D���5/ �����xQ�ʦ.�y3��5�P�v�j�&�3Z��<�����B?���R�E�)�r�3��|l���c\==�n�v=f��\��!��ҫ%2QbбV�>Rr��"�e#d�!�CA�>�E��I�p�矅�Eo�"L+	r;�{h���+`�#T0�Z'�%t�^�7~����W�V��{����+�WT�M���Cm��N���n|"%���S��r7H0Q"eY���{������n�2r��Ԍ�d�^��z��䶕��ɐN�J���/rC�1���@rZIYyCYxT;�a��TCe������KC}%�����(uT�<��31�Җ��/?/bv�)`��ZR�Sq;z���������`���rȈ�Yy���j�x�GD�oMᖔ�����{����4��AvS!���d26Һy8.�"�s��Y���q<�7h��9G�֎\����j���Ճ�Ç�����BF���0�����������O�9�T�u�0]���tf�IAU�HF�D ܝY�qP��W�L�'7�E/�?��#�l��u�> �3��_�\�  Z~:��C�K�3f>��E�n�f{;�e��E		���Qâ�\3�J5�U�O���&"�D� �O���7g�^ㄠ�'Es(��j��Lc�/����?!=��&����0<��� ��)�N��-�r���e'P�m�ˋ��h:"��g,�\��}f��m����}�m`Ӏ�:��"=��ɂ���_h�C��Z������RTdщ���i_@��=��}�Ғy��'s5�Ү�y
1�!�����0i���3��%91a#�g����ķ���Xsg���6J5
�� ��m�3�@4!dh� ��)ܱ�&�|�Ybu����#L���|ݕJ�X�!gpzɤ�w�(�`q��f��5z�2	��w�0a�t	@�k|��r�SA�&zш�i�Z��x�vsZKE[(�9���B�Wp��$� ��)���H���+��\�������?In	�hH~-D��2T��]�2
G�$N7�f�Q�Y#m��[J�ey�IR���9�1u6��{��|��Y��֍~f~���zE-�&�\}��\�V}��N�T@�\B�Ã#�T��r@����o1����a�˳�?�a���M~�l�E�n��Ԗ��I6'��e��-���'x�(p�=aQ7r,��/�ը���_�ֳ�[A���#�k)◗$�S���k3��e�Ė�H*yJhظ}na�����ֲ��f�E5���0���4�#�[��'�ĶU�m�њ�)�M@��C&?V�����Fqۚ�>ެ��1�;@���H豩��h�����(�t��32ټU�^���琾z������a�beP�N-���c����6��2��"� �����q���O���A?m[7q�AoμT���Qpu��E�+Ce8��G����dO�,����zy�J�*��l���Q�V,���aZ���%�!�x����=�r�����{�[*���������Ӈ�ç�!������U%6�#��6�ns�T$SE}�D��rM�S��f��S�z-9;��jĦ������z�nT�$��;����2�姀U5>4�h�0
0b3�]�o����,+:�>��	��@�#6|iU>�>���n����,vD3��`O)֏�*�g�p+H�Gʔj7+|goO3K��1��YA[d�W�U�q��s�3m�S���/H�Đ�ָ�1r�"��?�[�j ����fǁ���3�{�#��R���aO��@Ԙ�JB͂H�qpM��K��G�6/���q5���Y��#�y���E� ��͓��gTK�6]�[�'����;	nV���$�<,,/+iɞO����?.�"��E�+T��:J��YV���*�p�}z��3��V��i���yM]su ���ތ�񣄼��Vu��,�'��z,�+:v�z���O�~��C�φ/8��Ca �/��M�l����b/�"-H��l�df�kIȽV��H������K��,�zB^^���haL�����#<����@M����TC� R�{Fj���]̞b:�*n�uK�žs�w�1M/��٧v�]���dqu
nλJМ�}�6S��AD�g��Qt��|E����R\.tS6p�<�AK'��AԞ)?�̦6���<�V����t��l�bX���?���!�O �4ŚZ�#�̔����mdyLt��Ռ��e/��j�`���11Z��-KwzA�gK�2�]��3޽��2}�(��������2�uw�Y1O���'��C�p��E|����s�K�O��f�ؖ�؝���{��[��e�ñ+�w[o=�G�sI�8�y���0��_�w�A���G�4�B��D�ۜ�Z �/v2��Ք��*�S ᖓ5�[k���c�,��Oh���k�؎f�����B�_��vᮼu`G�4c.�9���(;���-�������/,��jί$� ��;K���j��I��k��y���^$yPVr�tG��.�)E�̟#�5�/�����J��<��������nC[�b��im(���,����JH�j�m\�d�{lΚ7�k���|BF���mDa-3��^;=�8�4�/�c�S��$���\�<��Z!�D�̗U_l�h����x4ڗ��"���@'�Liߋͻ]
nc�:R� ]��� ����o���%�)��pLj�z��}���H���h/���B�a(�T��EOs�+�WK+"x�.���<&z�^qP�A�����谳�6>�Y�?7Q>��8�Sى%$��T�^$&��\�Rz�@Q���L�=�oL����-$�F�e�7I�L �ήm}��+?������3�����IC|[�W3�]���I[���`���h:$I����R�	$~R�jp��ؚ6_���!�L�K�O��6��!������ƃ���^J���MR�ٝ��ʨt�MT:AC�=���0��I�	�Nw����S���r͡�l�=g��a/�{��Ѣ)�#���WZ'��E�G���N��*Q'�����]��4*6��j\�7���7e���E�k���Mb�)NEV�^h��u�4�ɗIQ+J��z��'A��:Dս`�0�#-F��y���+�>�6�����R�3� ��9���h���K�����E���7:t�xEXQ�u�����l�f󆓟i��՘5!������Mˉ��nČf��Ee!��S$8l[6�F�Y�� %j,���$�N�
�ϗ�IB/�C�')����`�mDn�¬z�^Hj�
�Ժ���΁�hm�;w�%�'>��_��)�� d�����J
���O����z�t����#�F|���auҠx���b�0m�n�֍Z/m��04"tK�U���W��@͢!8���d�$r!��A�)�ͭh��i �˕Zs�?���H�11z�#:g�6�Y�"ӊ5(g�a��˺�|mJX��Ā�s�u����Y���곢��aOJ�4a����wM��s���y��_����anw��/<�.��_��_-%/�񗌊������okQ%�ǘ��=X��k4�e���7�t�P�OE�GNȴ"��1��;�[{����[y6#��W��|��sO����WȡP5��ؖ�k�l@�e��*`�]�b���Ս�i2K/NPE�� ����HX6F(b�����H�3���,ʐ�3�[����Vpԥ��J��6���3�Ժ�pi�3)��=A5��{L-��ŗ�r��i+�`[U�a5߉t ��f�EO�#�����3M�I�w��@��m��+H�c���+czHP�յ�[�'G�����wBK���F�0S��W��Z�Dćp��N��=-�~�F��d�LR���!�Yg��O�������<xz��_��Sy�A�����\#NL��P��*��$�Z�K$���2����5I3�b�[��>H���`<��Nf,�1�"�ǰ��h&�2>���Ic�y{bd�-�c)-V�u�`�^� ��Q�C�h���U������2@���t���9���9�h��h�����6u�ԇ��*�4�]���LH�v��]���1q�	`"��lZy��i*�x#��՗��M�:��u�(l�|�b:��w��K+��`�</Ƚ��sp��pU�jV��!I��YG&0�<>�5�mf%m$3�F#z'��a�#�Z�����i�?���:�Jڠ�Bު]��T�)K#��eEL�����Y�����߄#�P��X�3���=���Shl!�YD�gȺ��$�(#0�BSr �e�[�f���:����%MüE8�Z�hG�;�����b�Y��R������x(�����aYv%T�^��NN$�����lԙᘚ�vM-M�#��0y�#G7�^d�j����/]�ըvgN0s�E�����q�\�FB�c��hӼ�@��9(�ЩP/ac��#�K6R�T��k���|�J�Y�b�RX�Rf�W�k�튔�nki���^Ջgk���{U��0��uu�j�>5������$�͌��^�o���sK~a�q�`9�(�i�l#t�W���3���>�zq΋� �;�E<���5�	�r���ʇ���]�̹1Ʊ;���}�����W��#e�x��Ҏh*)�Ǔ�(n>�u���/�>�7n���e�]Ѳ��_��T(������3�>���ɅL%LL�vE�V�FQ�g̎I�z�a��!E����?��7�3��3��4}4��c��y��8�J"� ��\i�)�\#%�-��,�+�cf�H��&�TD�_�g�G�c��ǅd5i�ń�87I`ۗTc�*����d����Oں�͚Յ;B]�$�si*ӯd*^��k�߉u�.S��r�j�!`�y�4,�Pw4�u7j�G� T�b�B^���� �Þ�j�ڦ�lhc��k��f�z�I#���y���r�r�c.�P��RA���}�E�~S���zW���;�-p��K�>K6�� PF%����[�XO]$L��f�?u5�N�:\x.��K���#�����qۤ�/����$j:O�4�.�M��ښ�T�׿�@,���#&s>O�3
;\���Zs�E����X����ږ��G���+[�,q�"�q�!O�pv���;���IO�ǎK��9;�/�;f��IR���Wk4/�4I;��@-mMׁ6��O��%W�I�0JM��> gv#��%͢����=�lAc�^�9�m��bO`{.,�^�W��|�[rHd�N@9Ϣ,b����?�V/腜�%	�l�����S�)���yl�%��62G�����#܁)ͥ`Q�֕h�`T���;����ha[��a�U�@rp����;s�j`I�P��)�g��V����>��[1���� ���+����ÊC�@Zrg_ �4�O���@mS `Fk�b$����7D��`���V����lM�OA�$�%������R=nS�A�2�0����(2�J2���&4p �qǚ�0���:R�;����\j���zru����$�@s��+x�Ձ,�b�T�m���5�1�3�dW=�N�ޗ���/�v,�#�	�dS�n[]�e,a���y�Vyv�h`�*�Ա��L3f�+y1T���Zz3ƹq
&��>i�$����B���K�	��n��m�F����]���^@ʛЙ�	ud%/֏�i~d���.��QK�b#	*���uc����k2ݻ�a!P���&|�-:E��1�?��i�C��q�*���{jD�=��e�����C��Qx�Yuc8j][Ǔ��}Px�����k��C>����ӹ�P�Y������)�gYZ:4궓!��j���N�~V�ɾB/7\�O9WQ�.��'����C_>ǱP��5���). >��Z�-5G�O_�a�������C��6ĳ��cIXN7��s��ɝ��2�'�9(:��1ի���&fsxOʿ� F_CT�;��j��V�^�\Za�"";
1F�54r4?�°���%�c��Tg�#"h5�;AZD��b�
+/�*'%���_e-l�h�i����tU�1������*�/���x���(hH��٤��Ñ&ޝ��G>_��d��'g	�IKA����f`(�45jY$"�l>��Ep���� �9�=	�`I�$��&�
���7�j�@.'��G�X��(�v��X���{�/Nt9�EĒ,E�/��Z�@A�UH�8�>�VԞ2m����2�Um�5���w�d�t������̧�Fuv����]�0�4�)IXK	�m�bG��:� TTP](,�>(���/�|�$Y:��ua����^2tUQ!o���P�V���h^�:E��.O�M%����֋���Ֆi�@ͻ'\h��~��+P���)�8�X����E�%���ͫ$��m4�{�(�q *e-@#��{E������[��a����#� �X�>K�3�
��2fOQL^K÷ح��ѭg��%ȋr9��D�w�^+v�&�=�m����R���/��o�g=��.���hj^�r��!��"�/�9!^��W&�ٿծ"70U�>Y��-�[�� �	c k�&�m����Gk�w��	���9j$�m+��n�3cz���V!i�<5teDd߆���g���<p{u�1
@�����*B�R�$�d��uֆoQ�-J.~��>���/D�V��k=�1��4G�p���ُ�B���JW\�84���*��Z��B����/]��]
��E>LyL���#�}�~$Xє-Txe�d�=�ߘVk���=o-������䜋Y�H�#4r=�p��Vk�b��;E|�s�~
B`l8����b2or��>�F�g�JV����#���4��]g� `�U�0(�[ �.�<
����j�0&������PRSNk��0��XVg�%�-�}��ӭU��_��/�-�p�^��w��/�#��������+bc9�;&�e��$*�0K�x�*���}w(�e��-dG?.&AR����0��pϱ�D��!��h��Lw���:��Yˎ�Z"Y�U�4������z>��	j�$:�Ìr/V�j[���r[<�k�_.__Ӹ��Ds��|C��H)��>�:N��K�e��Kl.	�Z��B����:�Y}����NX�Z{�=iJ&��)jI�Ӛ�n���N`�+܋�=�J�%����0n˂�3�e��Y�'D�Z�Au+���&e�w�(U۞�h�c�m�2+އ�M����GSC��Mpe%�=��O՘�ucb�6o�/r�yl�-�� L�Ɇ����|P���=,��޲���C��:}�T,z�6ܸ�<k3�2��zn���9H1�J7^C�u�B��j�Y����s�ݼ^�N�� �um^c1Ƿ���[O!��T-0�u�k�z \�9�[9Mw*�51�v	\O$i�u�v�5��昞�P���!HL�Rlo�\�.�ս���p�����L�E����6�:���\j2:>g���5kЩ̅Fb���e6ڛ�-�.��Ύ��d=�\�ޢ����˥p�Mn�\F�u��$���QHF1�����I�[�Y��Ǝ"��� ���Eeڃr��W�}%����U��D�s��J뵺�o� t�G�l��(���\����H�̮�*��o�7�S�ޏ����^a!���Q�@%��N��y��/�(׀.��d��/����!$��&�i�l�z/���k{�o�q�p����UW�z0%qԾj3ֲ=�ݬ��t���t�&'h	,n!��w��VL?�%�j�:����.*�^����5�����(kՓ|���l^�$�2w��y���0��Ɲ��(��Xlm��%,���i����o�&4�Jou�Դs�����5��N��G����w�`叄�\A�n-�ofQ�E���p! �辗���;��g,�e�f!w�j�v�E��_��0f+.s�K[zSAjOD) l<�#ǳ*�n˻O�P!d+�VF;JMj�OY���	԰;nu��Łv�%��މ1QS~Lv�G^��A8@�΂�Κ�K��oe�T�l�2�ȥq���r�N�"��+o8n�Yy���н���΀]Ip�J!�ܔM����X�tx�KC��{������&���he�L�
ϰ<ᦚke'���s��,�M���a�XZ�� �
���p��:�<L��J�l�,g��o�y�D{Q�;�~��J�����aW<�!�������'���Ì
[2Zb�N�?���Pw�z}�� ���v�_�g4u���v\�sI7�s��x���q���I��-Dۄ�s
���q~�yyi�]��	A�'�ys�������, ��7���[�&ފ����F�rr�
�)_��dN:#?�[����f����5V�(M����6�i�w#>��gqc��
�P�`m����-����l}ºj�� �<Nn���!n��xOi�3ɼ��n�i�I���ϥj/s�+�9��_�p� T���	�k�-�c:i��Pg�Pn�a[�[F�W�+�*�49 4ܓD����@a]c�։]n<��f-��H��#z -h�A��RrRQ7�������G�n��ro�X� ���V�$�bS�qQ0���C�a� lY��Qh%F�6nr��+L�L��w�<�ag�;IE��M<x�0�e!1i+��v����1։ș�ۡ�S��Sd�rd�:������C�\Iu퍌n9K[��-ۿ���j�Du<��m�����m��=q��A�ż@�y����.���:ŭ��U���H���g	���Q""+o�Br�)J&�j�0��)Z�`���1�owY,��(��Lu�H���z)��؎yO���<�����
��HI��-��f(d�T�����I��'A����~�h���k�7�U7{8&�L�b#|Q?�1��p>��V�<ޏ���F�ܙ�\Ṇ̫��8d���.�s^3M��``�h��	��7v�7�rQ�!,��1�J���B���a�2��/\|�͚ϔ�D���"���'��3,�"��ƨ6��R�8y�iM~g_��s���"��G1�NG6{� �KB���p���*�$ޫ��+mcN�7��).Nk�9'�N;sźD�h��"ā�h�?*�1�(���+}l\�z�
��b��D9�vD�X�d2Jm�ʢ_��v^�^�����.�M���c8�8�%�����`g��^���`���^I�-��d����E�'� {@H��Pƻ�U�u��6M��/	����
#��;H�;f�^vd��-�VOm)Xc7.���Ԗ�ۺ۷~�,F���(tBp��d:��J�.x����Av�F���[6�Ф�/SPQ������-&�i�����Cat�]Dw�5װ�`��t��<3�Z�c�,������ŗ0J�
{����6:�;��`�"�/���,Cc�򸓰�_����z8�p �T Vh�W��0n2dmt�� ����']��b-��%��_9t7%JO��* 6u���1LWȼ�m��\U��Bu?�ߨ��ȿ�v#��=Ɯ)��ս�+Οi)��^�s
f�����]x�u%�!/H�eJ�C��v#޲�N8"nb�.E�
 r���� �˵l�`Q�O�H�b^��;]��C�?����:�3+C�K-��;<��S��PU�g��z�^"�~������l����ĚZQ���;�^�ue�]��:���@o��P���M�L����J���wͮѸ̄�%DML��+9��2�y<�k���.�%�ZϚ����b��,�H��"7G�1�}���A��G��єQ�@O���V�W�/�6�)g����P(���{3�$7�+�_X��	\0��#�'(��G�m��NE���Ox�����G-���G�
�R L���~&c������[��0L_Ɨ�3�։9D���WW�X�r3nS8e+�N���ٳŘ)��7�/u&��Z	Q��W�Aʌ���0���A��g�|r������%FfZ��{��Hl�o3���e$��T�3��cY뽯���v�zb񈑝��� )�d`�>�|m�*�����3�q� /*ܼ\���j��-r9�t�%?s���"��ζ��G���������0��JZ��F�L�&D��j�|����5$��s9��Ik��oFB��R��6R�n��vKriꭘ��,��Wb2C�R�6�P�]�GS��Z�g�}_}h�r/Mg�+"@���;���"�������G,%T?Y�oRY��V�^^��g�9�Ҟ��P�x���--$���?�����w���Y���|���]�5���NSe*�����Q�s�#s��n�ǜ���溭�l:�[�f��� ��>`�B��_&��sZS�3r%Ǿj��֓���4���Rl�C��-����"<���۫볜�*�`Jv��Vģ����i};T:"8x�Sȇi7�3F�����5���)Z^�ou���rv:]�V�n�/{R껗#���+�
�yv'GY@)5LިY_[�[�'�V����I�b]��=��l�>�p�1�M�3Ⰻ�P�i��ʾ[����6x@�s���l�m��ߕJ��d�]��ڧG����B�����Upi��}`x0����>薮�]%xU��[�D�q�Z��P'"GrY���!]���BХ���*���/��"���Ih^����k�ƴ`7����b#��W�� �Fu�GcROyM�uG��7���b���W���0emJ�����{_��n8��铠32��"�?�_�Kgs�� l~Z��%:��j�9��I&F�[��<���E���*���ǁZ�8R��˽� [ǫt��d��)���<��^�����6P�h.��J_pa�]�1�D��T
���g�G����j��q` �BNO�!��4P�����,�>Ȋ�uٮ:���Vқ�:N�޺嚐~�V��:��@(G{��j|�i��T'-�_�y��PY�dIt�R"�Ϡ���m[�>:/�4�-T�$����I�yl��3s�|���*yr�