`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
x2oprkgOfGq1Iogb8qz6YfCa06HwNuOwBCHwpKCMYfW05z5d7qOMx/3HApR4xDXvzLAD9q4ZQwDg
W/37xWWwzNbK+057ddm2Ncm2VydzrIsTI1jFJTyC86wM5O+7JUWqZ61QY8g6Uan6be6tf56VkJb7
MCvwZczM44PMxjewqetjX58GGrncVid2CMeWcKqM3Gz0oLOwotjN6EqBd9ah6m8g7B2WGKio2Yyy
bATZAuYViwpGOn5/opT0sXjkhG5fTSukT+QC2tCS7qfPgFgc/3vJvwr01LoMeDvdTkIq8t4HY9sM
MVvfyN5e4cxRzmbcx2sh/PhuwHlqUK0vwP17onPD4zWlLsc08OOHmhqHeWFPLUwWmYfUisiz4jkZ
t19hMTNaEKk0Zg4I1ZnM/6QNmXB4oEMlR8/q6Iezgn3K0uA52bUE2qdI6l87HFmsXJ6VuyPiIZdU
CI44ARsBD2xHC0lEqEiKf3chxZSY2jc1seo3iMgdDzcx+FGB+LBphZ6pEbELldzr6nrGeKEyM9kX
njmSwyOK1iXvLqnfTwqIYuO9whXgx4YWIxvyIz6+SgRY/eT71DlEbgJQyWuWCeRj9ow0RQ2b3uIC
ychJHkvcdduFE52k3p0qgSykkKB9A1kw+WEwa/XY/w09kM6k7wXZvi1VZ/iOVZGy/A/cPmruOif2
HhY7Bq7IlaCu2z+XWLR1ZZWw1GVReXWqA4ozaePctoC44gYGQ/C5D1NMmfAHnEFocaxYbprIBqC7
XcGRtD7OMx9sHSoAuhmF35jBEBxj3KnxHDR0WV/bFso2OrBStk+TN7bZw/JS1rg1hLY7E6pW3OMN
fbd+plSS+kkSzZRYBf4nYhvLnM7aIrCuN5kBdDhxT9rhJXS+mx5Cjx5YLjnmLZVgYw+i1YWnR2ty
kQOcoJFio2CrMjSNEau4JMBTyoZEV4CtR7HkR2DEn1uls3GJojD8H3VloWNwqBMl4WhTbF48ychy
vm6whPfFFaN7WFfaXtwS1T+F70K2Jc9sSLvwxqW9oAKfjvIhZwn+UaodINKlF0JyRXSRXPlH6Qyx
3vmMWXXZjoL3OKNP6H8J2UXhKVCvbgaq5Lh+TmQIJBJJBMwkELqK36xdTiN1SLH2gAt0fK727yIj
/xP9eu7B92Spjb3eeZhPsCQ2S1z8w08rclNM7XruQz9WSnCbCq6s5cWR5UKzeAZ/C3nWVTq0Ug/v
YJ+OMcJXdrBYMrwqT3KFz1aJ7HgZXjcezf4ixR+3a+KqhevP7xq0S8LEnS9HwKfRpHc8SLyNIOWb
C6bb32yT/PBIDLUcWnD6yOKJnEiqGAftPQPamrGp3cS8SeV4UnBQRoIHakYnWwtBzG+mo8x8KfQa
PaXyev3jckPN8csEmh5OX6fPO9sTrncIdIKmgcTm7hCK6JkTBtbkA7lGmQgaeqr0cNDqs2CCr+jv
PQ2tvO5/4GwT4IGkStxgWrvZpzu5SOb6k8ZEG0NWmdK6uoySWxE1u4pMvNFPFh56ddRrequE81ah
Sw0dVi3FQt8w7DJbvBWAPjvkujDiQQ8AEY29qip0mk9KI0IG2G1GdTuCNMZhViS6d4yDuryKeWlM
A5yn8AGyvw/3sg8u21abiqgZkm09yCm3PYy5C3zQJtsPag6Hk3FqkX0c6RRi1sCeqm4etcrhW246
NNbHwrrUlD3Tj9AHvloCx7ZeXas7rpP/KkiZ/g/4RuvidTelk1cAOFPPGAUBhNK+PbSho2p1q2Pa
Yxm6cfA+cFrLNqJ17PXumd3XP8mKmvkjHaTg9262gTny0Shfl13K3X+uMWAZcdKgnPEJKGWgdqWD
kI6Rhrl0PtzdlUsfFrzss/wY0c2rcqY3Q7+jpQF8kDxxUZyQV8FtZLxfLpm3cgoZsz7Mr6eBW6sd
A4903JKYZ1dPL8IIxVz7QMzfurBQK06EfvKbXfIqi4vkQ1OtKEnySTh7mKSvwMbXvOEZtfKF/Yp+
WvNjXcFw0/UPZpBGlLGTxQLbuSwutRMNymsQWOnq4LJk04JdGN0a8EUHaBOt1DmCH7LdHW38GyjH
rYVNSZjb91hR53qluuYGIXeL7AvgWH31ilK5cMC8tD1IMzljFtVDQdS6UhWAZHZSGtyTZKM+dc0u
PVBHEdfjwhiPwSXTalawk5t6NpMvybsCfbiYzUYxAS3pQMh2MC9lehYBgovOSCYYU/Qnx4OPQFpJ
Ey1mjLmONxpzJamktUwPzX4Uq1uioptAqR1Lk+v84bHkVU+q6UVkLTU0bEYCNZQjXpTFdsqZNfax
GJeXdP9dXZX2M4Hf0UyeWmqQmPsNtbTvdx46p4bVJnyfsGWKS4GVBRhLQGocCV2kG0M8r9W1ksZ5
etxPC6M1NotBpGiXbT0b238KuDOmLnoATXjtGDyxiNxJ1+D3bAuA0QJAYgTmmpPwAE6jhGStJVk9
lrlWoY/IG+Uqx0US2weao89PHGAlPVG5VlNPoBEnKN0SuW3Xt58SGIwRifBxp0dZ4T/aSHBYozHP
S+72zBhym0FWHd4ZmC3NnVBGoCWy3UW+JGI6P3fwM4OXCXQoQgdZgCwIHMYFHbVikmkqEJ72XCYc
pssEDLHRnUIBytvHsqe+qUK1szNWP9lnAcu4/m7mdIAGHeEuuY1JBRBTCoB0prPQ6ghnoZVIBF8o
ItLbL7qk56WYB2bc0XyJHJIu33cir5YrBXCGQLpQwncQAP43i+U3bNwWDG9EzeF0VLtByxvIVagf
ecHbOPlVNKFhNu9v8EHUXNoJyjIWvaV0dDCW81yjrNF8m8ZdwAlHo1sJ371ODsE+vK2qiTbbNW/u
bipiRcWl+t6yTMz/14dSNwODMfzCO0MI6CsTfsPirP8Zc1CYWZa9Vu4rt56lcstDU1V8dZ9Pm8TS
LUBaye9n9aDIvMAe3GXjt3md98J+wSxZeelpI1nQTHcTkLNNoX+2netV87oA48wczuyKFX67491y
VWLhj8yk2CmHH6KmpPZTFPkKim7oxUngmVDTUq0ZzkXXR+/bNg83PqkDgljhAloE+eyJp0aDajYm
iHEQQMeAqjBBa4KfY2GEGDHfhA5nuhdYSgz8DuS0+a2c2TONQz1faPmq56/dpT0j0DbOwqI469RI
UK6QY6iJwyABMxLS5+PHMU+G5g5WSpHN1r34HSlpfg==
`protect end_protected
