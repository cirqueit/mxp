XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���z�B��!_� ���N����کt���1�@��.񃬝J�`~}�;_���^0s�|�^�����0��1[1�2PGA�SGu���������c����꩒�*��FO�O�)����A	̉��T�Zz���y���(��AI��ċ2��	O�f�^J�m3 +�!G�25�9�Ѫ"�l-�����X�(*��D�e���QZ���C�3�03	>�YRm��l	j��Jn4�WJ+� ��U����(��z��̊�8��f
���{Ҩ�a�K����$k��ž����^��D��ɷ�K$��հ?�-1�RF��=�]�<O�d"�xx�)�mK����+��҂�]B;0��-��nj����;�L�"a�#7r�������/"��a������)?�U�&�PY���>��w��6ta�J��'킌���+d�w�۸��7a�X2��y0-����k	�QF�5揕0��F�$���cek�����&М�1��FO�ϻ,s\;���K`����W<nʈ���z��f} ,�@� ,*T�<��|��!kM���^x!O1:��>����wz�9C��Dsr�0���e������FA�QXo�������+%�u�87
(&�v\�n@�0t|8�Y�:.�"�go[̝f����0�|e���˒{3�?A��t���9��)KЦ,�G!�?�?
�Q+)���:|�>�DG��x�S}{ɒ������U��O(�G�p��j��$3�X��s!J}�q�`���ᇲ �{XlxVHYEB     400     180G�`�M8k��f�y�ɞ���ǩ*6M �C
�h���-�}P�S�,%��i.P�CDa*���4� S/k,X.�ȿ70�D�E�u���E���h����ͤ�@.,���~qYvͪ�"����ь^���V"��v_Q���E�D�%P��9:7(����h��)>4�����u��o�T.&�}0'Oh�N�tW�r!3s=n�-�ψ�	{4�&��9Tok��`��[o���{&A5>����㯀ar��iI�4.��J�����0�[�2g"F�&�\ĕ�-�F�J8��qN��Y����Ix��(2�t퉺x������o`I��C����f\nU�/b;�.�~��%>� ���^�T\�����\CA>@��a��0�͕�%�XlxVHYEB     400     180�jDYxP�*�U+<\�)�ޮ�#�G���dcJ=P����Uw�ޑI���d�A�Z$f�֖ʾ��V��6�+��֓$�\�LJ����tt�*m�Y�,_ �\�"���%�s�׃�Z��N���H�U��%1T��⤏�״�!0�fٝ전��%�?mKǟ`�VHU���!]�y�$�J�c��C[A;��A� y�ڟy������>.7�G]�Ƀ�~�"0~��l4N�I~���'��}�Ȣ�튃�9X j֠g�o�k��fR�/��r2d25�R�T��� ���O�@i�?C�*�2��O��t�=�����+~���0&�ag2fh0JG��O�\h��C��v1�'4�ꃝ�ў8��d�5XlxVHYEB     400     170��8������|SP�����m�$[i'��3�DS����6�{�+dS��. Բ�`2�i���W�p�����ڼǷڝ�l/��r��X׊zx���H[�I 
ϩn|:w1�~2�򏔰�@B�O�c3���N|_�����"���Nd%џ�t�|QNS�Ն��*�hE�;z='���uB���X��b =s�a��2��G�]$wڼNZ�$Cc�+����9�� À!q�F	���I5A��
b��֕gh-���[L2�@w�>�^O����^e���D��#F��c�L5%��������6�p7r�Î���!�F�}�^˞!�:���7�����kU4x�a�f�!��sx^N�Ϊ�g�XlxVHYEB     2e8     120��JZ��֦���QΈ0���3��ԣ�*�������Ҕ�4Q����Q��ӥ���Iҍ��Tɵ-vL���{0S+5`l�6��F��lOv���y����!6�\2������x�
����z	[�ɸԳ�9.���al�2��(�S�7���-��Q����+;UEQ�ͱ>I�ux�I�1!`@X�ވȦH�P�	̯}�S��;ɪp13&{�W�:�	@I��lf��zP�-$��	�e3l����j�����d�:��w��a�)�F�\��X�$�����c�(��m1��?