`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
q4L6c8dy8aUdT4yxeYQa1S86Qm1WaWdHHgVhbs5HK+TW9ixOv+8Fhg+Sq0MB7t/8qO3AYx0aTc8k
I1ajlLO7Dc6bIaGeATKxfy7ThEenBtaLJUity4Vrjut5X/IpOMveX4hoSEGAuRIPkdTxSB99kVV3
/MoWAf7pXSQKdORkr7wxI2BwyHtjXjvmE1hoS9WPd7yN/Q3skL+t1MS7So6PsLP5O+1K5/F7nMhJ
O0whp6Z8cFpCtwBJScOk62dIt459/dgEGZSywI6VDNRiSpKaqDEBhdRrGIjbGx/9ZDVuvdGaVLsA
U4ZB6hqqwLV5s/q8y7fNgajmSAtesLuQxfm/txr/sTGsgZlI9g//Ny9b+xPM6n5GYrRP7lnvxyv7
qfjhJ5B7eVS6IQorMR6jHZ/hdNvY7x8ZWt3W7fBel00+Vu88+QU4MmsIfMXW4mgvrpJXi5vzVVic
Xob6sF/pGknhE9+WP9ujeSZ2iM2YZAMySCHobyXPA2NuxIbYXCEX9tW7XXhD1IlsaJwWTrKoXq/f
sNY4xEOPIPhUjyWmruHGzf8WO+uJUDMe9ydxLTOzgUcE+E3OGzebsLleYdVRVKhtewrWeNFIlvAX
6eAWzRt2SybvOOHdwDLGjDO1NACAJwRAADadlDf7XAWIcncuR9iMRrcFHSNn83NuALCkljA4LUdR
FEo3EhKJUGkjDFiZ8ZizeuBxmgJPYMigT8v1RNSzrYQMDcAFBMpqWZBcvbhqIcVvz1j64ssqnV7r
A7wzWu7Kx6+WSt1t99M/8b+B43ATyRDxUnERqf5YzADOnl7ECTHEV4x4nb2m+p0x02GH+mKGAWeQ
c8xIWapUm3TQ+TyKFQniWlGF3K5xuSKQ58WfeXJnY7rlpPK2YjTm+JU3mYg1fcg+35yjmmMFEWhB
bxFVKKFQ0+3kuEn2coTo/RrGJFmYSz1pcugH+X8sOzOgpOE5R1yDmYaNFgzxM2gBcsWEjYBtcefw
q4QvW6ErKB4e1zq2CvIiU7xTVAURVmy3PI85m1j7W6738zQd6wyPPfFYassYKfeslUqJHqIrL+QR
59QTd4amGKHa+QXKBe8i4PmX5mr9eazI+hhzL1P+kaqKt3nsNryu1bp8N4TPGhwOEmlUG+RJkajy
tmNmQODVSyfwgjrju1x7X/N+vlQt9TqL27rzuKQjksBTXtwqCSBBPxxp7Go8seDWXw7BgUQjQjzf
e6DdE5YMHJ568mAsShlXKz+lPZFuTwhddz+gebfCVl0LMAnLGLfW2+m/QxE4gVKBiGLSGdWY0Uot
6cKU6bFu1pTGrMVOvuG6Lpu7iZi28XEcbf7WJ7zpWftk7mMUxLZul2bz6IAevGFeLgX2UdmtsCyM
yMeiHFznhyM42MFpRvEr21f81paHezO6TNOdLtC9vfBDR/rBdz6qtacxFclN525kgEdM3mOHQTsE
2QFtsrpn33Vw/oX/D6qTejNZd3lI4A3lGmNSA4TrEa+RcTmWpXe5dGaU+l75cNZI8JHsp+pNRe5H
YqnuWydbzUZP6pQ1lL18t2ErpBAmIzGSk2gA1s/TqUbOI9qGWglL0fQIZsAtzzlyBy7FkJ5R3eYj
PY0gfOJv0HfcTjV0wwU9lpamINRLrDs+Gd/y1Cbqbsg91JiUGLRsg1vnkNPq0ToPHSO6hDf5T4iP
BNQVGUTuZC+cb+hINa5JAFS4QU9TQF6WO0LEbjSyFs1z2e5oAczgqfo+4vluL1LgHYHRPLUhM3RU
edfdEssTtcVz6K+TRvlvsp3FZ/XDys2s235xHk3MQgUCo1S+lvgO9EQVNGHgq5FxyicuLsf8dXzh
oqIS3slYkW9LdGZea4wtqJLnOgv73wY4R80kFy/tX6AJU3asrpAOfkcYN+ynEEmJ2GoN90AhjW5/
uN0LbXK4hNcSyl7SO/ZNVeQ4Nf8W5HgJbjIak403UPWNMXuL5MlxPrxE7KC6GDRtiMmnK8pnQsDZ
1HGwSNPWIvESd8Uof4DsrCcrdIOd6F3CoyKTLfvaelEmIEufouMWT+DFgMG917Uiq46gcfjkAJEy
CoGweVXEPFUcPX7VyrJ5IdiN3vpUYCEVIcoPJ0slyfjOLwW6fWvQk+TP7e0l
`protect end_protected
