`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7104)
`protect data_block
FJEKbMSXyDYdV9lZ9H3XWMRR9vz1GooJ5pqfKms03dy5R8yzJQ8pslP+F5vlkmmPoV3gdnj+ItKy
Lbtm5aKZnzIAte4BejkoclyXfEBfNdNlKf7LzgSQLUbeddnWf9VGGA/GyVuOHHPW6JmpfKEfT2fU
UYRMe9FScLmHdJPXlejBZa4PkXQqbs/SKxw3uZ8wAvTpiYITm1c8UOraagy47k8dsJUkVhn/0kZ2
t0EYhvnkiL4KRpZP861qYwzpbpSZm6IoSXxJczKixkzABngKSkFfiQ/UUVR7WDrD9QWkNp1I/gWc
gZSYcaNqQjWstrvQml8NeKtOcB04emugW32WklC/Gu1TJrUJONZDAFEUQYtSY0s+NzLDKbS62R1g
R6A4ujyjdNp4T+IuvD3tVRazyBJF940KmvNaH74JK0fMxF3xDTEuY0jXrRVlJk2Fd+UBzN7Pps3G
0CF6gTO1LnpbrAKXMGQzGelInQkPabGFHN/6GT0VmNyu614ClZF7CSrxmHWi5VVMpyiapeLES8+c
3Lm2bsJbkTht6m2yThRDVMmvvuA9d1vm0V/QgJISjwaEc8UXi6/kUBPGkJXFNzJ6m3HOQMU/+7S+
E14LI5acSCdpmeWFQkLvBf1JaD0mrQlreNRXCR/eV4lfFJqQLqPeUMnCGqOgnQe9S2h63Th7ghU/
+x8gSGpdUXz2q9p0/sy50AtWW7T6z1wTSvoN3JHvLYmRb43k6rKk9Cp7rh43Ct/h7SuTnISPBM/q
bG2W6Jng2g2zp9haqWEHfMBjcCh+AbqunqVRq+LEMmqMXvv7RnQy+A0NOEITz+cfng4I08vM6evK
QxEZKqiCpvxFLKcBfTmyWVj1YS5kR1H1jHMJu+6Gza0tTT4Y4oSJOl5Sl3m9wKNVXj82uLzmGDnp
7hsbC9EmR00SUCmsXTCMYHRDEGDI+EMcFiH1WYny36hPhNI47+Lm7mf2YJUMr7b+aJbzxqpI4jIn
nGNVQRvdVi/bKFahB8bpygTHeFePpdNHgb+9/dHYsYFjX7SQ8KysgKknlpINUPXpsjRNXow+plGv
0ZgEm5JEE+NKl4RMhys5HsAkkFV71WExkWZv+42tv7ATbCHxwXlqTFnt4QRhnSk6TMp39VsnhC2D
SQjZjNYG7fgkGeHpoBkP2yuc5N6H37CpYD30fhGMMU62EORndFBsppiEAZ6bV9oIhtNOInLo+13q
sZrHolQPlVHUsA/+l94wd2sc8OiP4yHEgjXkXrrO8XYqBv0F1M3L6Oj5HDWqGZGu/CgpCDnuxt18
y77Qb6oQtzcGQN+93DV/SkcgDG7u54rwaRiars7CAwEne3MU405jI9K42gHnX9MI42q3pLr0IDWq
aMI1q+/mNOJjFYb/vpkxj8sPJImhoJ8Hk6L/q051T0ikkENbWVdWa4tcBS28qgYGgExaTbJZI3QA
NDve1nVPUv6lyvzpbdGrByVPLk4SjYAW5zEZbx2bLCiHTrHgxO2q7dRPeW54uzEwIVB+hnyzVUKL
0OG8ubWnWkUi6kuKUrme/oQWg2X7kg1w9RPRCXtWlU7vKCPwgEKrRveJCzCA8OI8dmviq9ZPwGvF
ljVjGtgHOyQ0nVyyXi/D6y0TDnfZntdV1KTV4qmqMHWPsG8ADVfSMjDNXVpgxAonXjL78PaOHS/f
17RPoe/kJMSt8tCrPp5sAyWKkW3x7BF20lHPjYKilOas4koQkPkjkkczunuUtKDIM8wgPmHfWF4Y
i8sjscnfbyTWvKycVoWwQd4v8QDQ45pLPRkAPCIVtzlb0KgZ+70lgJWYqplobfJliCaKoAEt5UPY
R8jbn+G3TdvdaM1ek7DD/go/iYdoA7KKLWuERlgJvtU1PCcPflljk5qBSPAFUDwoxVWkAlnY0Ec8
icv0HZXqKYTPuGgACSiLTiyue8WV1d46d0d0tPiWfNSy0v60IM1G2+0u2G0E1rhdYm7yVzvBGHbt
lnv6sNBrSF8nrV7MPN9S34VZ6ICXsHbw7f1XusGconG8m8y1KKk16LWbea0JGP4Xw+5I0TDxWZ0H
s2MoJNeIJi83Pn/tk9XJCndd3DiUoJIl+5bkGhEwa6rcyXFk4uUqVpTYU97fJhQEpXpQfCvYYtlo
8gSZK/42X2rVjOikUtuY7WEk1Z7KznJBSAsF3pQ37Ko1KTUcKHQXXVeN34WrFFc9CStxPkzP6jxk
QXbrtBsMqv2Eq4/7nb3cLs7yxhmwcOvESjd97VhfMmHU+z1K51DKMM18fMjZHuS46CLSMYrKHSRu
NNos+sKQRxlqph3jiskWZoe/L8pMs8AvlxtcPa/Py5KqiVx1PkjbtDXbqQmKzgixLA1F+yxKPXMm
p4IRbLn1BeXWazcWDZxmIcKYpRueFSTzHxb6X6Hi3NEqkgcqoLZdFMRj571iJsMbmFXnl8uUkqb9
AyV1QTVREDzBlJKxrQ0a4yO72z5wZP4z062KUI5ykG7OayEL3If4YwbWHO7a8RQMCM5QhkRvo1li
HGVhTlAelEpm6u9g6D8uyL4VN1HJ4RmdNNIexovAEaZRsyYFl9N+d+dxOjOVS8ARr4TYk7JpA64q
IIIAz8uZKbdQNYO127TFuUyk7e5cfCqF3raPxaiBO9IH1gxcLVf74TbVo/452dUq+N/VwHGf3U9w
5s5XEs4NSiwslxwNFmEE8tz+G+9kL/Fx+M4feTGgNmLrnjoBAMjJ/djAts0SwbIIChbHKDq4FReZ
5LHB5eLHf4hpFF2K5uwmlbOHH/HG/tt+pJysZ8W4vzaMEpeqfVlN0ZjW7Yc+ZTZmKuJ+S0xAWhug
3ZmBjCmOfFsjRh7atFH+OVI/LgQgv84J+2dgZ/8T3AUqdiA+pqaI024CPeswHNRyGID0WldnRNNc
DvXDxO1CiQqbQL4rMe3Pl6JMP76gB/kfKgzZlx57hxsxhgGUC4psMF1y3EgX1Klw5Ri3oekTtHwD
hwOKTrYgifthetrpOjj7pBh4r9g/sVoWI1RoBM7B8tdowQdEMmBAzy186bQxVlThrWbUPekDwLdN
zW1CWcDiY6lh4wc8+W2KkdrcGN39mhD/5p34SbQIAhHZ6ekjdmRhTFdLevUeag7CGCOFwgOdD64u
Z8WOAZ+1yc2Z49rYT8W/ZbvnpAOZkJf1IIYu2+Q22GkwdUI0H2UcDVw57sDQEZlFwdMr0gXerTsG
CbTzq7ZbxSbMJWs5Cw7zzB1tzHEPbueI7Xaa6Rjsl56+lPESETtQIoK8V2CySUcCXzMGUGS9yBCY
ZJcOGS6qGjXBdMuJk/ElKZNdKv5/fQp09O62pAwGsrA8kil6MNYt0DS+vB2RR8pJWnXELUIhgQxQ
M6gweUd3Y2X96lA6ycDjATKHCEzj3mhh+uc0Wn345qquMsZ8thTwUyzKWEVKRxbfpfJJfZSDhmkH
LAl8LbHzW2MCozqIuT21vsvEFnGCcZuKFh8ucdaqcGN32OHvb79hZwa2v5wvUJiLH3XpCJH730na
fOvw6Rjbg8SKAxJ7YFNc4DkB7P4Zc2DIH9xIZ/sCjqHtgy2qp8/qnWfgzhAamrThjweLbd1Vu0kI
aFYLQ5jMK5pegNsH3ctTV6YqILnFq8TgvE23aG0MFrurO2EYqAQ/RY/dMJjDEW0Y04cFU3yYLQKm
mwr8R6W57rJy239DoRNrQHB/HWkaNXIZ82fEQiy12/0COg4zV3P5CeNO1s4wtmqJXyfGIe9sfE7x
CIPanQj8NkeYomAyAWNAHFhgI129ypUwiK9pQQU4L26e3KZnCf6sQu7c0zZg46nPk+UQ7Gr88tVt
Cz2Iarr2Z3te7crhteRQ3y1GD3PNcN1BqfSWnnviqPGJHhnjfhOQz5z97HfGouiaSRR1tGwvzJ8F
FY4RL5ra28B4Y7jWTjMTUDRVtutnwu/olXrU/Z9BeBVAH+vUqdcXbR1FgVl4qN5gxQ0qKVLoqWxK
Qe3FKJgZ01N9nTyR1CGleIMutQaxy7ENiovLjYln1Oe8GKAJseL2gXYtRorw7bj83M1I8u5xq/4D
6aWPQRhJKzvQvzJCtHDBCezzZ6XN5JKWFBAjHcIV5lGSTWt1wkqQgKrn9Ktb5cXK/e9SwqYkiXCd
Z9tf+Yyq1KTz3al9WwCgJBHu31TmAHLfcwxqQZeKyw63IbksPqpeATCxa2GtpJgpO7tXlgb981JH
9ucMTbgdzVe/Z8PNtNq+J0kHKsmCC8Bhkrm4ci0/p23uomB2a3mjzjzPwe4sR5c75ieEgkYD/6of
A+2dj2RITTcO0WxG0T7qazDVh345cOK0v4MiZQXiNJkZTMrCE5ZTx6E3x3scWSddJ/kKg/mmqxga
b3Xd8s7rYg1ORrBtMoXFJT7hdGXW8yUh0Zo8hLVf+Cs7BjrUvl690HZDS8G5qMvCrVWzz+2pfN4N
REBZCzmHkeiwPsc2IjU0gfhv0Fyw1xGZJmt81XmvsVjUJlwNDNNVtE+lo3l41s42fbPABO9A/A2k
6TwiwxFq2oAj/PGcivxDbTi9rmCsu+WjVO6+yY+/wE0Vay4AmZCm1/WE6QLfhJ0kjLkkZnJhKcXu
n/z+k2zDwKs0svxEWbDea1B8As8yBkQfQRM22krJduB/jiqd5QuTQciJsT8gA8QtKTgwtxI8quYU
a5EqfacqpDFCbluVGPfFEOAGSgFe6H/owPftr5muTembj7rLn5GWDtKot/fsL3CShU1gLhJdvQ5k
XD8s3NVzuu7zCnC3+Dc6T0eyds84dNZHmUk48kd8hRssMhWruWt2ULb+mF4cKQk/eJpKhu0BVL5G
Qcu12wejtQT5LAvLbDZokDg0vWV+3epoUjnf/dqYAw+QHlm0uEqjSBiuAVJKX4fhDcARcR01NUpK
B4YtX4BL5NVunrbsrJ6V8S/jjVMU5ffeFIDNqFXGAPAMMHeS7IczDwidCyDv6g0wHYBYOW0/8Lt5
iOJ4XyMqqUEhnBG/Wgs+8R+UFEQqH04M36Ls83Nj2fIt8NPrvHTwm8cws9nO+fS+rS7OTTTvsWW4
yBnvr3bgBg1HYvv442DT7Ame4WfDwK4L4ghmlemvcOzIyO4GRjwUUDqYn2BTMKP86egOu41Rdeur
LcIU50YrlwBLF4eSr4ENh/GswG3gQNuKf7tOxMHbG+xFywEY9+JA4xX9oG9LQF+wK+w5TDnun1zZ
zArtsfrsAwKHvB9Zx/03/A/iaF8iNFc84fMdtj8WeLMNFGx6g0e50y+xoFKxdgHxRNRux/Gm7l/K
2eZMBSN1lUe1f/bXXULNFGt6nqVFxXX+P3Dig2iGXJPykGI+wKgf0Re0wxUkQ+0djvPf4DCF6wEr
PExbT6hwby++t5Vu7dooF6WiXYxjk+FCc+IVejsPJ1ZRb9S9BAkvCl1Zt1woXCDYZ9xYC+SXC+Al
kex3hMSuS7039rMJleJljfZIPnpSLr472UpadNnJKc6kZvC0bTlpuEr2DB/pKbFTOScz017e/dX9
qZT0MtnMBlt71k8Q/t05NFjpCeTQhBiQkJOXETRz2Y0qxSDNmjzeZ1bqQTd7kplMvObOpW+TZrQz
konqtWsA0QZTvEYLVr7mug5KyUpFYJHvmRIoC1vNrZhpisKovHtnW+z51qZHu2t78eceeq+BULzC
yGLlkOTcLsQqD2E6klqoXnvpEzoQDPf34DKFEe5Vi7gsA+hUHoSq9sGmIx8i7uomhPnGlPMjP1+C
jdRY8G+a6Ls/EYxv+p+K5ngkREECA9R+huf4L/JkueZEcIyZu7/2/pFig+tIGXpbhlUdNs+t2kDs
20JLROJuJHmuLsbgbDubn87UX9oKm1NXsQBuHqoIdmZuAW2anWnReW3tPsoyts4S/KuFEd5mD4Y0
Gy083zaSPlS5Xg1kSoKvekFzYlVJWPjTCS5fswrm/uU1PWZYo1xVKubjG7wHd4FJ6i9BIfYQygb5
U4hMhU1IotcnVjmTRyKMEUBxnX2uYByvo4a7FX9SNBd8Je170y/BY3Emsqq07mpvIOtsN3Y+LjfT
NEErbjmyNlXamyOTdEN0mHFAox0f9muz12p/a3fy/yFaII3VhqtXH56aimOcS0bF6L8yWucDcKi+
hD9oQXOyKhscKKNAPZrjC0fOj1iXWV9avixkCJaTfblwZ2lhPBKr/UXB5ynzYYQRfZLTRzBLvJz6
5beGiFaeNMNzmWALLj64+t1u2mYPDogf6z2UOVTSAQF6vYpyJOesqnpS3g/vLqCL37QukPAROJBH
vr+gE8r6R3FvDJ8reFDlXyVidhHWmozd+L8xhAhXLrtWQbHYqn9A13DSVw9xsBlLF+BeaERJtNEz
vf37ZqmLboyD7qny676OYRcgs1ASoq5oAbbwOH/6j/EUwyiO7v2hLqpI3FNsvf2buWLLGx3aOeOk
OgEZXgLR/F8hjiPKIhVI60FdCINq5Y2Zr4L1ARimT26H0QtD3PxGNeuu3YuTeh5DSnYm75Rqn3K3
JeoolXWvgySjTsQ/jEF15fHRym3mv4REzpJBf27RBbgC4ZjzmIHpUxMNXHWFZC7fEP5HGHW5OR4H
5G7PYBJqA2qjL5I5CqDs5pyeEfTOf101SMdvtk+gMZUCYniX84dbhLlo8CBhq9gMnLEVcSTHVxRY
zAEj08BPTzEpTDNFN8+/yvW/S1z8cjdDgjJ4byG0wyFevLl0ghShIBPGz+CQHsyIFVp/44BZM/Dg
B3FuvomKpGZi7aKJdyNLaZDjN7DrHVKOFDs5ticP1LkG4rYdZ4H8BDqVECB87aWbO4zr3ubAzj4S
MDd0V/HetgoZOVvdQ9eS3pDfmks/BR2nMG9vT2Xe2nQfb5SxGIlMWGW6lH5vf0QUVMdHkQKeFOT4
L2fkYlwPM98pxaLI5o3F/w/YEX0442r5TN01seCMCjcqQsYHsO2JFZrePkDX8PCR2cQ90iQHd0+k
qzx1mEf0VGXJvmB882tv/Qa+ibDl/IDt10yDNIGSPdH5/3ohGVntdaSxOjowLHRdWkuBis5rVuir
su9wo4jSUe8SKdgr4svXvNK6d9hzwot2kEbFJOTrd0twpZp24o6yFzGN+WrscXQR5BXHm1DmmysR
yGsm3vXKZVyvrM31moraLRMX2WB8bq9YseaBRi+paZEWoT4eNXyNFG5ABkvfRAPOTUzbaqaKkBrW
4PfyC1hyHq5QW/7iS4jimUM7/3fejJQ7UeQ4lEL2Js+plB0cb7icAuENY6bGJMAmgXxdYyeZfDLq
AmVVmDCE0G9MVb/QuAR4SZqeGwOVXXao2ZTsJ4/VWlBqARGDYgA+aqJQj4SwMptsgI8qEpfyua6k
Yyw/OfdHbrEtZwhHrM1megarRx8kz//pFyRXFX7JKudIQsygNXr+YU/+GW2/8ZPDEbpbp1FjXvar
yR4RtAihQPvjgTBsFTvkOmJu4bufO0MIBJKKDaW6Q6HpT6zy4lZ+8rpTAnmpPz+s9TnfB8ZeqpSR
l2ylAd+mq+xC1nc6iap7o+UaKNSpHEeCGgkm1sCNuANhCwdHX6h9sQhZ++Zb94/hSy3k46tx/LhM
K0gky7Ih/v/pLYIlB4MGa+7fY98jB9WPbyiqcQdG+MNGaicu8NPdzu/S4j/jQ1//8SOEx4A/jNgc
4nex8mr7swzqvE+6LxElUaqAzsIFbzAA2i42RQ7DCgQlFLxilIj9Hs0THvG0jNm4Qyr9qnqqApM3
R2trSC1M00qkSJ6enszpYrwDS3zXdpRNElyGoTaz/nlxP/KKk9+Os8gWf0to9IihcwTLtKs7rBTZ
qogsPdcWoI4jf8OboCdvFC3hQpu0bRfAZmcmYPResOMbjJWHU54lDd+tScKDBZ2DrnGjvS7/jJN8
ZdjcWkovf0ZB1VTr/a7LJrocpMaoA2oaLn/3YyHqmoh0X3Cftut6wd7I2R06amk0HmY1Lry6btuv
FwAqMVWXbZiUCMbG4phYYypwrIZfbxkRP4cMnut5WdVrs+C4J2FVXi9IeH3rVKkDdVdrQFxznzJG
sg9pQHqm6p4O41csEBMdpZh+sx+QJYPiZZKEb2N4IdTtunvXLcM70bF4fr83pWIBrgqMoGsNlc2b
EbMmzcjqVG3AMjceH1t1H9f97K4OhLBqABNRN/bCJDBrxMekDMnYoe4wl9uXZnkSHRDr4ur40Km1
m0XAhM4EGoJGucho+vim0JHCkyMFs+gJgTklDbGzGrNiswa6Z2rqRRznwq2sznuXGK8lRZ4BOwkP
ze/P20ibNVXzqWU1vY/KvLnu9tFlyh4KJjlZjKTgqlY4P2+T4dBy/HAnjS6JDtoy2+WBywn0HwVJ
isdaq1fRJxqR/9YNOx0uIV5yXnQ2me0gJYxH8veU5RAReZL3XXAxyc1FEsAfPMCp7aLD/lwegUpd
8Q4SEqSQ0Ew97rag7r/QpREMR7hO+nJqIFndXmXA0YnxNu80D/BAUPupl2jZTGr8c4W9xAVI4h6D
6Z1Ett0t8XNanMOt3CpteuqVGWeLdFXcwtKvGWSQsOtPZ1fPwKC2jHBRM/gnIPbJxqwyP0e55XnB
FK9OltkCNif+57NPsQJDAFSribQ/8vYDOU3C7yn0Do0Iz7C1TGF39tzQcLbroWQgqRWzd6zKPHiX
O4PryhaIAtBGz9IanbYfb38c9/jttiy5qQC4sidqq7beo9ELIgg4Tp1yz8Xc+bCNZWeuYObNtBi2
BdYl9nJwph0CtWXqzpGmZq5l3xEbhjakXS9y5wRk3bYpDY8b0I1A3WKkEnjw4YS9L1PJ4IBloy4f
NYhzhaTc3SY5sPB+2h2nO/d5DkpDd7SSe1FmCnSAtUQxC7PgWgUz7paHdeJvla1lSE49LnzvCuSH
d61tRCFG+2ZZNnCLJ33IZCqsXWKmX+/yZAyHKYyQKn9sszn1h5n40WiK4p9pNXMDUOhvQTscfUVQ
7SHzBEKSBIWnUhrZ2kmC3RY8rZLYUcZxfOiVgNNEkSp30U1Q6ivxmqCJuTIardmKLZnSXPceXLCE
FcztO+qUKXwq4JcTuXZsibFeE3NipG4B1ZJgULV1SbZT/6MPdy2pinHXJjr/Z6wTp4okRpFpPXe0
1Xr5ZkHR1nIUguxG0RzDH1001iDXdDCs6Tckg7thGf+CV7+7PCqEYYJk/cLm8q+oOwNbKT6pzgIk
r7lM+b1n9XALanU6Fk+Wk2UkklbHeoRx0ByRo7JadL8h1kMEQun9HTa44k6THWNABk714FkpUz5c
uYGJAaBz1S4w+pkkERa8UcTOdWdQsiRtlEvvSCA+7GMw1WpQLho4j/KgqoK3CRPxLJdAyMTV9EmO
zyn7hKaMGiFW6mLxwG1g6J2nRAjujvxnuBgjviANzfuI+PQ9cvhSnm1JQOEQIBsNqRNvMKJWeizH
6CeX+o68nRgW/CRozdqfy8R4QxS8WqWKqB8Ui5PbqHWTsbU6tePBKi8Uooy1lxLdxj2mEZB6mrGJ
zxv5WBiiJUSY2jM9Ou3hW9u43lo3dgq37DKFfytjpiICKrOK
`protect end_protected
