��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���T.��%�9HF`�Q��$U�H��q�7��|��J+����j�V�����8���[�p�ώQ��ka�k������r�(�;�Ay�E�0�,l�d��2��0�9�jn^�tJ�%���=5�y���K��
�z{�T��aJ�b�?��룾�o�c�����tXʞ�G� ���s�l#% ����s���O�^X�NY>t^iK����B0:0���O�c?��N����d+�7đod���P(�՘��hZ�sk;�}�:n�q�k���"������ۖﲨ֌G��'���3^���Q��_?�2������]n�W�_{f�0v1(jj�ؾWf3鸲Gӭ˟�X"�͎�.�s�R��S�X���W4��;S�o��]F�ɷ������X�+0Y�g��U�ž5�o��&9Ք�O��k���6.y��� �f����E=9��<S��s��q&��d����\FU�,��A<�6��;�����h�b�4����+�_�|�.ݑ�Sn��v��I6�x�f�v}6�}- �5�a���Q&�l����H�]�>H�T�����?%Z���9x�B}�t|>?��kE3ḮN��T{!���PW��aS.�#� ���p�Kz(t2|��iU�)[V4�Tk$*�Z��'ֈ� ��`7����,sG�P�2����η;}������}��O���jZӊZ[���V����3����f��[dWN� ��(|�����?�� ��1Vr;!�jP��*�k<��ŗokr��a[�&;X㼾4��@���p�`R+�S���UY�P��wV�	罫�]_-G���V�/$�6���k�qO�l��i��E�����F\��WH�:8��i���&F�+�ƀ�O�d9Z�|����rn�V��s.�y:�5�V��$�
u�ӛ�U�r1EFn�Wq��Z�	�i+�t��O�~'#j܌��4���:����H(U@?�a'/b����~�i9�6���fU��^=�Љ�j���/��^̋��2��*�J��B��y~�9>��^3_���Vm��97~���T�z��ÿ��UP@ծ����,/����w�S|��4ʵ�SA��I���76F�����Ϥ$��px�,�X�]2�5����`��Y���!��B����P@r�S�!��j=;!���sB7l��㱤7�w55�M�3��Շ�)��TR�9����Cq{�&,����C�*�\L�/�N�7 ��g�}C\���Iɬ�o�2��fM�H&��A4}���HM������iF	h�EhX(cQ塰2�I��#���p��;-����Zf��y���-E�7�Y��D�6�ƈ$> �1�.��8p��Nx�g�BwDe�����w:�'A�h���:��x���w�����ռ���̡<�l�~m��$)�wӌ,�ڮS!�S+8�ed	�a����E���d�:���!�¢��y�v����)s�&zHK���GE�\���چ�.Y�N�)����n��66JM~=�,Y�K� s�іI[}cM�geU;Oj}��`~�pM�"���O�gs��i��<xk�Gn� ��ϸ�����I��*�͵���k�we�|�3�4�z�T�_��(��������K{D
��jŮh}ǭ�-��CD�M��W��եcr*�oOiQ�=���A��a�\b|i�`�|��T��4�����Gt��t"�u�6��e���#�K)�+�&�b�H�ޮ0z�`}���&B��v`{�w��L1�em�]��=�F\n*j��h�͋�/�6�)�鶆V�Wͬ{�����V�Tr�����ε��H�%I�y�w5V^���~L�� ������_�����֠1i����ל'Ē4h��S{+�Q���'&p�����]�ߞi����F��p�;��� Їv�D�k�����D��'�����#$o共G}(Gٴa�N95񸾧�uu%wf˧� 6�Ñ�L�m,��{Τ��:>����0�a�c�1g��xR�;�yp�ݿgM7w�[ �M49��� ��jH�v��'Vj���!����ý��9i��#�j�.X�n��n
��y;�8?�yJ�u�h�4���8��"ބG�6��<R���\_x8��Kq#��Ɓ�WTo&�9��o2+"�}R�E%�u �k$2ܟ�G�{��?�$��%4�9�&cL����UL��793������:*��+���g�6�|�ƽ[��0�p�*�+׋Q���(���i�3�N���Q%�;�>�E�����ug�8�X���)$���w��Ic:?��p1���|R@�*��䗁#�v%���%4���w���I���D���9�Q1�q.��v�!�i�蹇V�AFO�N�`�������h��\|Ź��s�4&�k�Pi�7���E�#%�4���������Фψ�N��L����
#R(ץ+m�rm5">1�,ق���ʚ��/;�yX<&i�:(貓#F�\�W�ݏM��m�?g��gT������s�=,I jK��� "�?������,M�ZS̆!�-Ѿ��N�\�����h��{Bx0C�D�ˌ6�%P�r1�"�,��|��w[�%�M3�j{.����M �p���&����X�9wc��^�7���?�����I-ʳ-���]����؍+X3���]��6�Z��@h�[���9��c��.I���NQN��Qux����T�G+0��� �`�#�W��Gi��/ʧ?���zOB)Э��>Ӗ�I��V�(,����5Yd���st����|I�*�J
k��hY��e��kcR1�9I��=�L��w�̈́.�2���j9�'"��4�Ll}�qw�:�id�GRQ���:�Q����)����R\O�;��|E%���L�;[��r�_.}y�>9���?�W=���!L����</���6����WF(�MƳW���-ȡs�*.����k�-�aC�t�6���Y'��K
�(4������ܰO�@1#<���{�	��� ��*���,�UؖaDJ��;[2'�-��q*6��Z�l#�).��{�CȄ��U�e��O\AHŋ�`��7�����[�/�i,�q
��<��X3P9�ҷ�Ycٖ1���x��vk��Q3�5�}�E ��N�)��v�Aj�޵�f�*���A���"�a�U�[��э�WF�ʞ�.���n_��b�Qs�v} ڬ�Iߵ�Y��J2���*ar<�v[9!�Ԏ{5&��N��V�wD�*Q�i~~N���EY2�PSuG(^�22��l/�-O��,6�n�]��"s2�=�ZZ�0�q	3��1]�Tm�������0��%Env�t]�O������1=�P*���Iص@m%� S&�����W����n��'T@7���������ü�*�#�`��d��`\9�
)H�r�Ad�L���1�u?ND�|s�SFm�v��y���R�`/�h�y�F֏�F�-�Ɖ�)!|e���e�����h�*��@���0#)����`�|U-o↿%|�ɾS���0hƊ��ބ�j��~������ѳ+xfyv,��:��^�7��IV��������/M�ˑQ>|vN@tV����yJ���� M<�$	����
�sĞSsvTͅ��b(Ɓ����~����k�R�P���MF�\����Ӣ��Yw���y��{a��`���m԰���Lh�\��e�L����r�nA�M7?�~��^�Nڬ�=2���wB�}�c��	���e�\��y��i)��y���~�V�B��B%�esdzI;#/��K��JE�ͫ�7�u^��(�5R�])=��v��8k.�u�ҷ���T�#��������;�÷r�8��1�K�L�:.�\�}�Tń��?�"�H$�Zʪ@��G��w�Ќөv��L%ǩb��}���ň�nb����ѣߎj�9q�$wI�PĞ1?���]
���kn�6yϖ����LO�Ծ�G��p��pR��*����*[At<"E�FiՇLXռf��>�Qg��W��x�%'�)�׽<�v�#C�l��q�$��5�(�M��z�@{�xdR�?�V0W*�:�F�4��������Q�}��TB����@_��5�5n��ӰM����i9���
E��=�_�<{L��qp5o�<H2V�)�Q3k6�l3FsWpJ؟��b�/9�^8�_�S�e(���)�J���VҒޫ�9�kY����S��ӶP��w�(!>�;����OV�~
���m�����9G��\I�Tn���eճ�S������	w�yc/3�_�Þ@=�����gO5�B�˜U-��<]vSX��h�7mf-���U�'u�=�_m���4W�mOhN}B_��v�^�LV�o׭����C�|���!P��u�)�OC�<Uݹ������p�*���
x<�T���(ϧ1;�R� ��2܎83ƙ��X7���_��W�֨�E@^��j�t�#IV#�'��d�-��vG�^Q�帲{Z�1���`Y���o<g�D%�����,^�~?�v���`m�Ð���!�R?�s۔���?��̭�ټ��I�/8�Mx���;udÅV%��Ί�x� �sL'���:
dd�x����Y夵�LS���2�;6�p�Ъ�?�<�W���~3K1�-%�����Eڳh����v�g� �;��Zf8ȿ6
�D�2F1ץ���ȠGk�9��>'wA�����R���g6}є�=g�m�NZ�����Ax���z)t1��e"��3%�5�-�>��ioFP��@��j�䗪@�ܺb�z'��O�@����Ϋwj���sOmJ�$3�W����-���$�?�z�����՜Yq��z�>Nv��ȩ�ݎ�1�*�Cͥ�V���0⬳��s1�h[|x��H�聟��B�]S2��V��r@<7��F��b�����&E+�]��p���?}<b��F �R���+89	(�w��d��d}���
ge���Q�J�@u_t�J�V�Jt��/��Uc�EJ�{�1}j3v�� T]3����pJ���k�ץ6��N�H����+�gF��g��i�� �:�'��@��0���U�I�#����>�D�b8��п=1��5��>��A�94c�Yb��h쵽���^�`���*;%�C��I��1�>��'F�J�k?N��Tt��m���|�Ĵ0[��O��e��rq��z1�Y����?�gD��y�s΄!�A��2i<���D 7�S��A/�k{��OpuMtV5,��6�L�Z*�l.��]A�	���S��-���ΰ��:G.������������`�b��~���V`�irگ�8�s�%�9�`�7X/2�k��2@N��%ֽ�M��S�:N�O�n��\\5�s�� �5"ȭ�7��OO�qA�������������/�C�)9Q,:��v@��n�t�I����_#����%�>}��(��p��7���3��eQ���f��;P��b|�H>,�P �p����"I���f��H��a�D������U����澤W��d5�Rݪ$3�XR��Gȯ�q��<7oc��5��GmCom����/������zL$���=c��o"�,-͗��|�#���2����݀���_>SXB�����嗸��^PbN8Y��M�E`J�� ���!_>:,���0��Q��~.���]����q�f���CJ����(h����7�BƷ� #��@��j��Git����n4�O1���$.*)��BB���&�"!9���]�+l,�P/�6�����zPF���X�Z�S^��	X��"��-�R�gӥ���7^4��pv��^���t�������li]�RصX���~P�۶�Ú����� �ԏ�\���ļ��&-,�"��Ĝ�F5fO��6�T�!M���q��D瞗G�<�}�D������Uj�ya�K�1l��Ch7�^e��~�t�T�x�u�s"� Q |�Xt��iE���6�L���gI�F�j���Ҵ�J�����p��<`l�Fws�(R�`����C���p���c�e>��v��U쓴��J59(4���́%)H�J��G� 	��N|�H����)����&��Xc���dV�Le1!�ߐ[�Pn��K`�<X0:��(�?����P�iZ���`�Ɠj�n�Z�q���~G0���D�X��v�����kP�Tj�n��@)ۛ-8�0���d�ᐷw�t	����s��$���uri��w��
iN�ޕ���)�q^WG�p�8�)/ %��L O����|�O�[N�j���,�'b�3�'�3,�me��R�7K6yR�2(`j�I��8'V�mu�l3�gs�Xw�����HUʸ��uAy�Z�eS�U�ms�
�]Q�u�@ϼ����v�ݤ�r�����?�j�b�4:z��
Zk�F��Ipc�G����=�(�?M_E^O�V�����x�f��I�u
{y`��(�)���/�����	E|'m)2�7�����bQ�B\Mu�ʍB�0������| ����|�7l4���'�g�A���hOQ'��+Wk�x2w�䖏1����Fm�t��i����{˦�V�UI՛�7+ݍ/v��En� ��q��E@��eQr�"�'we;ǋ�cX�If24	O#<lK�6�Z|2Ӆ��&ΠE�Y���}��~Kp���>h��ju ���M��� Йف�4�\KI$u�b�*A"���W�l��f��T9���+3B�Բ����fH��<j���5�2�� _���G߈�eU)��A�ָ��PHyO{Bj�1��J�y�I�4�i��-^�ǟ�ZRw���imNVCl��a�`�*��k���>��T��'����� �D����7�0{�r�:���+��Yi���p�`�\vE�MpYn[��l�H%���=Yk��"%o�]眩r�M�p���k,�g�ڜU~��I�Xt��5/&�t�Y��_�]sѯ���~7�����ϕD��j�N�΋4�8Ņlt�X������he �N����5�d}W�He���9�Q!c������l�]F0�i1�|��$��@��9��ws�\ɛ�[D�V��*�]/X���#���Q���a�TXZ�Qu�2���2�|o�3�ƕZ;{�ե���N`��D퍻u�;�k��8�B~�Ѩ����1�{�ݻIT^\�g�Ѯ��8}��ޕWI�J�[F��U�?�\���V��cIR@��z��Z[F"v�b�3Y��/�jx���|Õ'Vϟ��`у����1�l�!�rh��>%<b��3���X��E���B���F��
�;�)���{?2�%���9hcɐ=��K�C#��t0V U�(�b��{���O�#�
C
�"���*$���F ��M��6��)[ca}mZc4%PV��D',�*��c_�4AE�?�=y?w?�����6=�6�����{ ���i>�U�խ����E��3��#�.&��!R�+*�@sN�XC>����,�@|���b5$Cx毮`�L�c����[�ET���y�s\���G�^��!�%	H���U��¤��Tkc5�Me�җ��1  ��.ڊUN%1�Vw|p&r�u� #+��AGU���r��F�<�����>�YG����Y�jR�H�&��ben�^���E��1���I�zU��|��O/E �d��Ә�D��$�.o{�&y'�O��K�rd��J�gw�!�S���D��(\2�Ț�����A���ҥs\����_�����E��N�+[vԅ���>��2M���F��ee>7���P�w�̗�R�>/K�Ldo�N�D��3��ض�q�a�q�!����{����&x���nܒ���4�i\���w�qg�7��	6�+���"u$;X���_�GX&h�\ڝ$7���������2�kI��.�+�Y�:t�
lS�Rx ��q��������Yj���7��z�����$�z�s�F)�l���!F~��=..����a�!0�"%�n�B�m�u�K#hU����ȩ��Μ��˽"���cͽ��sNk��J~�]N�I>�d�IO��KBaG���Px��S�p����S{���
���b5�
��F��W���H^d�k�tu��S<���������b�f�j%����~�އ�/�Y�r�e)��4�m#8�Mj!�&j,��<��U��D����"�Lf`U�B-�e3� ���2�T��c��WV��qA�j;���0�*$d�N���<oճ����*��-H�o���"��)�=��l��w�O���ZNT�O���38N_Z�q|j��s�����|�ڴ���64�w���NA
n�HI�y�/(a�݅����~�ZF7_�P�Zo1�x�P�����8�}�����l�Sj_�
�XN4�%�t�*�9���hK?��-5���N���j��7L,���J��q�:`��j�_'�Hr-�?�:xTƔ�LQ�c�0^p^���]P�����J�Y}��n���\�I�b_x/���0!g ��@?6R�\#�8C����6t\K.�u-Ha����q�y(A^��?�&酳Yz��9���pvxD��n���I����"�|�����B����/KG�~����RJKM��:D�y��kRhQ\����N�[�X*b�A'�2����ߏ�������A�W�pUՁ�H�郉��;2���ߘ�/W?�� 'j�f�'��_�(>'�p���j���Pm��h4�
O.�s�Z����C~�wYx�q����4�k����3¸���N��LJm	��B'��8$Q�����w��p�m��������g��>1uZ�eD��B��!����W��
����ɜ������C5V�;�$����ԺvOw�dd%�NW-⦉�����'�,ig��d��