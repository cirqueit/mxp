`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 100176)
`protect data_block
wLh6Vkf3mrP062eUjXIblNAfgfAepqxPWkU8zZA+osW5OJXuvwmTDZ6UjUSuxf86U233xiKTVdgT
h3DnSxXOnSVppRp4pyWVvUX3p6ahvPBQADfoe1lh1cJcjnvspJEvZ74I/e4WAV9PmxjrBtgP0+Ho
eC1BKFiXTANlNzbl5Nft8WT384rYk8Ik64888C0h+//cD+y201U/kyq35VnQkq7L3/Dnz6hfJs7T
S8OP3KnOV43ahT3KxkYrr+z5oqiI26xSfHx/9A/rycYTOeZ70cxFY5WpO3t1e7mnpKl0D+4IjzVg
cDZBm7sQakORY3zWqbYgZDDKzjVmK23f7mg7DKtP/sOfjFxwtDsGJ3e0nyowe74XYmshbV3/1i6O
3IHFlknJnIHo0PyDOo3meP7ehDlO1XiedQPJTkjmeY8hUbzMkxsQ4LiJwl+B9+FBt6uUey7CtriJ
m6f+6ehZqj6wGUISgy6t5Y+F7IUqa1oX9cNBT/9n7Fyn5XG+y9BXfIXuavOT3KmnKJMJCFcWIhT9
YwtWldrBx6VpzZN06e0+AhgedkM9pfOqQ060+FY6gEjnN35lm8RJspaawGMFIClsHSo/P4CmLDNy
Jz/64kniCmCacR2dTEcDeKBiPJ7gkBz4qkFrL5J+MRma6froh8+JmoUudY5b1uBChp4WA5n6C3ym
Tt+wJtiEFGkhliNeTrzbWOF2DAZVxYijfUnWmpf1MpLfPtKNMw+Vl1FJH4Iuv8F2aFo1gH8yyuIo
a60HmDHuSJvrYJOIxasTMb6wdpwGPRiQYPzjWQ7lsgz+EvqYCeDFvZ/anbwqD4gT0Pj+Sn+fPaHD
QjEBWHUgcJcafd5R2aERblg9qHscEH7CLFQIpKGQlpS4AmW6lpR00Uf8jNN7tLyjiwIzbBna54JS
/O5Nh+sLjszDWGNgYIpfLQ+jnvBNYz/gEz2pcQMp4oQq7q4OvmRaNHTm1T31mKiLxeyhuiG9bLRd
UU+AiW1IlokOWL4GY5MVE73X1Nwgx/8p3bfZ5i+6l0fLexfis03HhSWJj+5aC1AtsQQvw4sPDkI6
dJPbOSDoX1XWKnOv6fN2GxZIPnwfecQmwBIohPAXi01RPf1KX9m2zR0sWN9DdX+h8VylzkghbKZu
PCEoRUwnWSw5Y1UjlREDtbIPeVpAx0K2XbSAvP6LtLSbbkxKttDgUgwq2ER08FSIyZ+L0iZ9pYOM
SgrNO03jM8ldOdlpW7cxJr5tX9gyXt2876jZDquTTit/1EwQ1Ui0VOtze9bRh/Im6XC1tkuqilcB
cdMicTs5ifPdSArTRaNifzTybC6wfgKzExXrAPFxQCz2fXsF64o6mpI2V6DNmW5KQtp4HffhCB8Q
DDsL2JjULFGxtErENNApozcnDHsnR1mYqaO5AFKJ2VJe5rg84A5HdZCskVdL8+lfMgHswYjWDVIA
d2fJuZh+gvmE1/u7i4ExejYXh21U+dH5JFFXa0V9K8rHE1x3VZWmctS5fPEI77aDt1rIHmfgaby/
K4kpexcQEEa7el1snEZU6kCc0tVcecqRNBuoSB2vQFHOhNXEd7XnAoxg/NkYv8eLvlhgoXQRaGKX
n7BlLCitOUi6C/D5ipQezuAqqF0Y+J3w5yo857rO5C6vlB4Zc4CpQJWjtNKIn8nggQu/zpsbvnxt
Trqfvq2t+s7ZAijD5HZhZe2agw0DVgLa0xyPgRSZwc42pIejQ1CuMj4Rr49/wiFab6pKUq+BsHNu
nP6rrIgetMf497LxLt5svvVG9X6b4eTWo0DXPmXCQZhk1PnCl5Q1OXTDjN+ybjCJoJ67EYNRwkO4
ud8AMmqJ/NXj+JJCje14d7bKnuTFLVXFak8B+JPPdIRSURMZxME0RymgOP06CmXrV13W9H9EfSAZ
C97K1E1Qd33a/TT7g8hEOq9Q9DpFKWTlsMymdFmRNDad5XAToTwm/KFYqWUrWjCzpxcNtzmU6ab6
XZvpt9EM4annr6SAbX9Vk3BZfF7cK7FivIPsYVJC/QTQY4e7dHqVIJslqFsjFydoqnEq4EVBj0+i
RM5vh9i4eeE5X7CIz1Ls8+2I6Vj0EY4N6z3PDhUSGq28VKL4ar6gzx92HcoEp5Jt8oLpKHlI/qdE
/MhHFpCaWfbz4m77R99Oj5j3oF2d5lAAQEVprFSy57cI5+mehRT28ZOxM0lFbUoSSuzA39LYe187
6J+11aOE3XdlhUPFjkOvBnSvp8rQcm7y+W8BGYNVnTdi8qNbaZh1fYTDYoVS6ybtW1idr7L/lxbn
1tCWSsMea/vdb47mwdc0xUWAXGx5ym9kCxXv+T3Ju+nDLDufOzXyRYOO9FbYR5UVelqSp1X/7Euf
2WpHmjHwYt2HCsVK5ToZLBA3EgYowXwTYRhqtsyc+yXyvtiDTI2Kx5F1sMA+iUMX2Sdo27GtmTrp
DyOIiSh0FBZ7xNnc2WS8c9FREVY77RaZRZayT7MIQavZSlBzuOli+AJQW00iT9g6Rt7LQCl0bJgs
ys0B3rjh5FpJPXABwQTyToCmlmZ9F9LD9fDQRk7znm3l7LnTCbtQf/Rnbt++UG3yUe8JR3YExVsH
4S/T77ft6EtTbqPlsKXeUDUfS3xfZi+9WaYUOKYQHBKrbicThmNf+aqg74bkPZ6eFsJKQJ2mqqPy
+ObQLlas8uVRefp5oCWcm3T2MhtGY0ideFxq6GXV4zVtCFvrnMUU2AuDp0Gq1z6inUP3quomdX3V
NWGG0Awq1Q843xp36lVhR0xnFxRa/Fi01377AFQ2OlewZjVdn/RsFnKj4DB07LNP7vX0VTaaisff
rM9z8qLEDc2qvoGE8jiODXB85fgPTTzLwgN3HroPcxsyw8KOoyIscPV1u/fZB0Uj1hpI5U9U5ES8
077+Bx1WEUSMSsEi/k6I1+fpCofNuk0L5lq6x2TbpJYLOSo9VrP1NMEOEf0GMT3i0yKM9/Kh9C35
cFDoRxPmaYAF4bwqj6v57YkICr7xHH1I700daA3AzBM3eo+irRnohs2Jn6pZbImGzKSfKwwuIWIb
OzFgsua7/tZiCjsU1ABpM6gCc9gmW/+7WhC3YL/i0JxFo39EuVLwIb+6CdkUy3SCRCk/d4F9j8Qr
K+EFwiWuw5gyfmbEjQFXFsYKhkmI8p1EOlqeCi03QeEGRcXJkjIp25EfOQwjFXX/8BheloKR7u0B
aY/qtqJ/pCHZQvOK90MxWiHCDyYImVMKMXIdhK4aAgmzLYk6AnPJ1CN2e3XQnpLct22Qe7zevPIQ
TGVuGnvtsSI8n+oWCM8bJIsdUviGTkgBNFOVjtgA52YPuMQBrU0bZ2VbsQMylLh8K4cgZw/GFDE/
L0itvs3PRa/pdODVbDne9f3fgmfnpfHmigaeF3deK4vETtHFTWcBXENca9ey6IwNAnVdbth5AHVs
cApti7ud316cVKT/unn8qO1VQMpy1ttphOxrHo3A2IlMWeQDnuYBtTj3K5oDx6Mo/tShFmi/koOJ
5V5SjK8cck1L+eImxFoy5twS3arfxB3XK8JIgkAbSRVTO2I6MchFreHEEsHiWYtQWObhPejwuBBi
8Fg1EtJ9i0+doVqmsiPyzxBiml4OziUx0QRhCY/TEgtszm8D0RbibLWnpotqcKEw0I0nNPgkPFSY
3dlbqdDya3WIp4Pii9vnfADYAYvj9mknEYNzmLCKqUHq5qWgQGCUMHO6Yf9TPMK9rn7B5tlVkYlW
dcuBYPZtM85zY9ijGXaXetnXEkmltRxE95vQJ0Yi5ialuJWmZSMlPnj7o7bdV5lWDgqTxEnRjWyQ
2YNpkt+jEtYP9t2RO3rjMipQvTzNXkSF/WNz2tx80+SkUtIE+7qB0/Ggh9+/9k6lOSfRxmQkriLi
THWkXUHQBOlr1dLkJPddwcFOqq4ladJNtdLAxGqfg3U7iyZ+YyY7DY1c5VKImxf2lbZI3G4IJ2g6
ovSfemf00fAyJo5r3hTbrO3e+4PhFDZnEuXzwwLHnosEAwhAVP2qAmyrAl3DfuhS8a2ugymsZESy
8x96Tf3MoJlCf7q8Ua0oMcy8tPk7i/z5nIIcfqDH10vw+KKfTvkrSSoRtpmoOwCKamvI5jLbSVvX
E0pLunXLzoGYwwx3DazFYxcrVPpmKTE5a8+AyPy7L2q1ktmUMzWM2bYxnxdcUvHPK9fKu1rNJvxa
ifPA3uA6VeAv4xVwGkoRFB1XVs8XDc8hSKAw6TqQcepaUkIJsuE5e15QeXr+YklYiiLi4FB9FcJQ
2w1wP6lEbKbxW3Y75pYhfWg9Ya9WqvTlB0c/HgD7UPAVsCRjPBs0PWV1s5ReZa6baFG4Z7TcPxSY
egOjlY3uYCPZZZwtI5r6smMP3z3xYLSi7aTmWaXDQDY2MDe11/X5wsyzH2+jfHk4krCcMOUMs6Xm
qQM2uIe/XgpEKDPhk5rlEIKivAhxJolm+fH3Ku+vbf7u6+q9rozG6BYgP66RWqMgagDtYO4BK22u
T5XO0r4XAzufxYu4oAZmfLn2xT0L7EVJWTD+DFWkiSoFWxd1dWrlSuruORWWxjFdBOADszrz9rDe
0kIWlvIbt3kn3HVCAbHE9wLT0mes8Ol8JgQGMnIdJhx98AvVElodQYV1BV256yEd7qUALTmgc2g8
pHWhlQ1y2S83bGVjTWwx+3wI4KpIdSoBy5lh5wMTyQcbTSYBJZpZ6YTJMd4rk9Fn0Dg8ENSOIMGC
TE9q7V6YJqY9ZxQXtdIYeJYy4obUSg7iguQXULl/45Ijv56q6MC4y5nmu0Mfm68CxVUdHGrurwAm
qadGFOfIqddXQX0jjgy+jKyGG7MM4SpGrGrgZBeGztzhqPX9g8gTkxXR3PESKvcxsvWxUgakZ2hX
Rz6DH0cxzSusCU9gB9WH6Dku1mLykj4iJILk8R2b+EpN1hvqrVT6domGyUGG46P3NEuKQDaelKRE
0mcKSB4qKQ9FFVn5cxGp2H8FFQ7k8DVj45LM0p8vBgFxnMo3Wy0KrXvGmCThnErcTb9aBp/c/D90
cX11j+wDb2vqDhWcrUin4bMUVD8Gxy6CFWl+5NnR1RRxDJt2vFCepkMgfusYlZJf4+fuTORjwf6/
l9FbUKV1V2r7fcPixHEIDyWfH2XDFwnP76b05JeeZrLN1c3um/tYaunqOhdwn5QO4djuC9H1SUNT
l/WDauNp9XJy4SY/21NdBM9EsCOHSSCzCn3y74lu02MPkPWkESOftVV5vKRtyjVKcwZppJhFzgbn
2DNk/GjNfnXCmor2tRrfy8CZM42UxUsUBMH8vZqLIME9foczT5Ub/Y9QnX/9wigA8dn+TXpHyFIF
zP38L6icR2turbt3NJL6jSiPDEIQUZmr/AN27wCAOs9i5enkIgf5SofmnikYO2N8Qlz8ZgIs1CHp
OAjdBiN5TfmP0D827jHAMqL/qw/gAWibd+10Ut16iEiJd0b9Y8cD86SdVnsP4ZQGMZQBSl56z7DP
7KDS160mzjbDZi1xZWtYMJx1VpMkikoHuIZlZJAaWs7dh2mUsqh++aanPJ78x8q3tGogN1n+2cWZ
tjQZca5VkbNO6FVRcYl97zAPfJucPGmqdP33OX4scO0IRi+0f6RJVkE1yFHoaxbN4h33g/Slzgfu
1OxdCzhP4twfkTcRRbFcETuvP+BC1givkGeUsDpynl7yI0bNSOVSwGDHliV7IODSEqr3JxahfgBW
g0Ot5J5pTPoTt4rm0VJ+QueCWXCnDE0142DWkLTDQ0TQsA1hwc4Mu45Y4h5T4ypQQAeh9u2DgkNi
0BxEkYOasNciYY6+9uHtx3kHjyuXI+Sk2+Tstb57Bku4Ng/dge5dmleqBglkJdaz8S01M4pot7Ks
kuQjgW3n2zARqzVan+MVU/Y7+3+6EQ7oMeQ9YmLmgJsLS4ETFV93OjF02txxsoNBhPUKpBB4Aiw4
HV38jEhjALkARHCqD4xkOKOex0pPdLFm5zhBCwAcHZmX2duSqI0LRujg49N6uevUs4UKA0u+U67a
NOtaNK5J1BEUjyoWPZ5+6YKMkPzFVCqWb+tgd8vtUoBo7eO3J/Z1m8SvZ0BJ2WK/oSv5/y7yzApn
GT3EGeYXb1cOwxrlGXSe+pSQFq0/PX1PmMG/mwK1NolkgvYW7Fh+pZaTycQhA56hmiE+gpXbIRh8
QFPFjiBmaCdZ3snfzzohwWfLI4VRZqdE6mfJmdkVY9PfDEeTE0q0nzCT+KJTb2c5ZXJxtN78iwkM
DMNuXtR8k7/LiNu+7m+cEM7RaEXhQTQ0TvchncDnkGE6wuGlrXxySyeVunxQdk1Ysdjxr2zoew4I
8WD14cuzsL/qf4OmmyqnK1WsVFN9mMDhaOI33+2rgod/7jyPJGZICTzDctIVGFO4I7DOvrl3necK
Da1RKYQNRnNWR9mWt+smwKzxTA0TKA9XI6sE7yxpwZL+iYTsWI8QKm0+tUEvV6R5nrVj314YMThf
MgF4gjQRdUe71AhfIURByiRV3KLjZ6s70ETHW1GoA/u8FgoDRe7HYoCBPG6+GvMZGxn7M16JfrgX
qBR95jo0umryFSDZkuOBNOeqwQBmINxW6XPURZ5Aiqak5//s6bcs9tHWxtTs+8zkLXqvNC6eF2gX
lXIH7V7su2pI2fJAW1VGN4uAHpe0Jx1nb3Izd47oZrE4axYO+AWqKSIXa40dgfrI2trEVb4O6DxQ
VH0xNuekm8F/6hOyH1U7pJ3YRxtmXT2/lvG1EyykhvSFNzA6Jv59F9mKu1eFIokYLNSDk0eomGEF
lnlGxi/5RTiQv7E+Hnu4HuHUJZoEqIBTxUsdbUGsF/yiQFXOJZnymPsaokn67yifoIfVSeLbglWl
9jllTv9RTAQAtrdq/3h3JjfWlU+oqCOHA5rCteKMVBJx0919tb18q71/QQm36KXKSOby7ANnVckJ
Ti5mC2CqMT1sS5VpbAPLS+NB3Ef6+kbfaYG+Qgd28k6BNKOtNkOyodpHAs2j9oJa1jN5jc29fjt9
OuE6MtSv38HutiRPKvegdepDWbmXv7PaDYENtc7XTZtFl9xVmuCdsD4mm/lAu0GBuGAMBE1IYgQu
mq2Ni/ipVbhpf9nzd5KAxfP14LU35J6dNG+imBEMVB49J7qwCIXnZkv6JwYP5hDQTa1e3IwfDS23
kKXPKdRgANw15DmsELuNuFvOApgbe8Dqyfg8sTK+K0oQYUmRhyOdrRVndFDpMev9CKkQ6yyN0Q6E
tyXlTHDzXNZPtOBHixb3I2YEaxGVQQOfCYUfaQkKO2G2NK9Qp5KEXhR0v9iyDxZNeQRFn386ZNXA
4c3xFukF35W3/PmVaPB0TGz1ll3GCSoRZyCTuO8spb8GgGwC5Fx6L8rQlPUnAS1GNlbtWvMYpLnn
r9h2HCkWMgPhVI7eplNN8hncxop8v7UR+Lz8FJQm1fv59p/RSsI+2FDXOKsqEOW4hOxjSdToBFmR
RZ2MUfMPvWjUA79jLqjZMMpojLg+UEhQU1i0aZ3U5XUV6dSySb55nSNMBobcCq9H4WbuyQIVpjCB
iK39fMBjv40JC7sAV5osViXnzLc9wG0bmdICxKgKGDIv99hLPyN8NghLmIRg7hp7vlcD4HTNDf7r
TigR/ZZtHhVJb4N5uRt99u01gLwm9yLpGqR2fQCP0ZpCbyfCvuO7UVUMXPfuFN6hgJoousQn5B6R
gwXygNMuVHWy5zKqOxKJBtxV4bMoVDttOh5P50D62KhH0wrg6GwsnLnG7ey19VqxOCFxF6QVSegv
UA1p89joc0W/KWDM0CDGDA5VK2r1tH2AJchEJGqj+EUWE0PeBe0bAsZV2Sd3OpQcKvMzy09tOxN2
DL/YFsjYyZ8Q/ExE8hbMLD7USuM/bEXfszRNRSnPz7rqVNJxhpsKKsY+88yeKhxxlVcBBuLPbveu
tBfY4c8dGQGqoN7ffVUqqN7tGdUbwasjV+pUbUtyis2z7wv/hI2ksBL27oYhGHEe2E3g0dTL4y68
X1cDo/Z7XZscw5vuUpl0auHqe7uifs4K4StAKeTM7Grzohxo/CXrSWVLIm4v8pgk8ZwUhUfCxZ0P
KNYLaWjq7PSTPRWIuKggS8OfF6PzylK67jNmXKuIdTffXkrBW+NKCYo3ck7aeToJKmmASUFIIV/s
y/bc2Ii+r6we2tmamxdmJ4VkpP33DwmAVpxY8ds+WsPMjPGMX1j8Nj4U9M4v+s8VUuD5kqOSly+U
7XnQLnOfmuFvW6BzaSylD4goNjET5yVf2UDqUImwMb44YJjdG117VO0ez2EotD2my37hA8jituKD
ytmqT6sNcVO+G1dLov5ezjI4b9VJk/6Ug8hZui5LFhtkOAtvh6x7zjMU3INR4LzMVG/v0Z28lx+t
Rm36pIGFAYAbe/gAeQn1fk2SDx1kbqZfmbdvgiBjWNBjWxjt+wYxtqqroGvRSZ3TxhEARUzDqnVw
tSpc5waF2UT7nrwtAenkFofVsZo/SebTDRwD3YOQYFYPEeFWgiTw1Tp4bHtTHHkBTwlGKVMba5BB
Bp+nOG8eiA6U/zm9qWF04D1dEv+hO4gzFSd+6nodtUOy18xVnXOfhVLDFZm+mklVax5EofH+hH68
gzFE+6dZSG05w9PdEtUoGiD+5c6IdIYFhVunuBf2g3Sm/B0mLOcnEEPO/Rtd9PIaKmlOtZ/4Mrq6
eUrUDIyTQNR/WcgktwyASTI5wm3I+g3t4sdjPCJ5H0FyoDlu843HHuPQyQ70GFzpaVZZ8NSypJPq
aRIO72VD+Sgk2rXJDS0YXsVWO4uZubbCnW2Tg+sJ1+tBr0vVGq180E5XcJY5wCvJ1XArePaYdGYO
PJ36m+BS5MZM6WVjcHjQ6NY3cR7j2/Hb0SvcCG1OMr6ZnGfvcIo+PYUq+wWmmd8CrmYu1jmcoLFe
I+remE1rN7G+pMPA0tDmFsutG9OZI49qXD5XGgm2v4smpX+78e0Vq4ZjuKn/6hoVhwaXUplWOiiA
1cfeYCpCL+hjzH43U+p+HFk9VuSdPCEUdOEN33bht+NvqmJkVR9mT4FBAjnEta02l9hxcb3fAa5n
4jmiDvuBKewazT9dGbKrVfqZZ0XTb1DePrJuUlHU66st5Ez13FfU05VKloRkiLc30aHKCXc2Y0Kc
qrI1xMJEQ5/p0ugi088Bre8Ud1fYyIQHEjmvqfrazAdWnvrjtE7gNvCcd4HQP9nGP8mcwyVFMd6Y
XFuhdghy5UjiEXkqhlGHIQF6i4OUp4g/vSGF8BEvvMUi4mYAxet9CnK9UlG9/PlQHc62PFOZHxRN
R+pf+up4NjEl02w92pc33q68h3Cjb0XMY7V8BVsOC2kcUi3RVfx4lYLJRBrJTL+NA8eSfuw9+YvH
Oa58Z94LFf7lGdlzS2zUbQt7meIXb6Hq64OnqutZ6o/J82VxXRD6OuCtQZ9l/FEwnHhkwk13iMgN
vU1446TbbvyFzmZ/eodVajDfHn49WXO1iL1EmwT5plBGkdcehp1uuNAH+b7EEDS2EZNm/S8KI3Oe
ZXfMBDjPVaF91uUCr60I1xTFqH5iR6XFkA1nKpsSdCPByFPX3j0jNBY3fkztH8ERihTBS4kVciUB
cE9O0shcemCt+eE7aBAakKgKy30+xFrsWWg+tItBuyc+S61QcqXdi7acQifMrnxbNs4FVdYT3D0l
yluBtnq3oKqrvoSRLxessQUelMvGGU50oniKuhRRDw7c4h8TVtwnkPTBVPNnHmxNKdMlc7yJcKmQ
b5NiF162DFX2s5vC/NOn6xMbPtZIziXkjHrxthRC6AiMqcR/pWAd65Bg8u3FXUVCXoI36rG8V74d
wTDyfsz03ho/l3jbvIVTqv+PQGIPwT1HsKiJC3yjCwq9rr95iZfwmS0mV69thEjQmGWREed15ISn
4gno+btTc+/wrdWKCAsEq+IZtZbkYNYcp3D12dVmA9ViAqz1uGWYv1j4Uq4YUz0wVnzVqy5BJEoS
+YqDwdA4hy/BSDRe1opO4p5/QnS07/7AC9jDneTkMNd+2yWED28F0vTVGbNi83XJzJMWwHXaVtYf
XOX2h8/ef4xiCMsvxHSUeEWbJEwvsVbp7PpTFp8xxM6eNb3+Ql1kZW+I3qZophOGsHkLjJi1J36w
CUtZrzVgmBMp1P0xECcMNwK2o8RPmfmlzTwdTtDeZsvwssbBwDA9CU49b6NP97kaLmgMBrxtIJVD
duJ+TnqrzEP8m5r3hUDZQRktKBnht00Q8KAoAsDA/MBTw8fpQ+JL4f9B+Tu55IiqFuM8itKdNO78
VR1g9CEmCDKJ2CDcMUeFJhkbf4CKvDtS+50A2KpQWfpqpDa3nKhwmd1X2LFiGzKWGwlj160NOcWm
Z40Ag8jPkN2IhTP1wX+kmX8095I0dmwCQ6+zLbaLhdkjIQcELXJGk2MpIlBkrWznxjFd4dQyOs1k
rBSSJX+PC6fuay8n1JbI3uWCArgtvWqQ2tZVfeoWMTTNF1EURF7HJvGO6zEL3kV4cnFavsOy7C4B
Bp5EIgq5jrzkY+H0xl9BPs5sU0zMgk93gpDaPIjHs8y1AW3ADFrtR7r7wpOuT/Y4hdZfLW47bNEv
H01gtmxIVdUNe3j7Jd4XoliP0Iz889DaQwxA/vtD8OwdhBA8junpxZOCCzKpB+7HsGywB9X7LZRM
eCad1PpGN61FX3oDQgmrIlP3zEC4iQU7pM+eqpZysspmDFRzUJsLvVPtVWnIiFAl7Zr9Op3dzZoo
7rfgBx26/9AK6sV1hDh8IQqLL0yILrmNr8x1VmiBACdoVYnRh0nBqPqJ3UT41K02RCNGpy5mBom9
2G+lbI0ykFznf1aKgc/Qxm2CgpnMytuourrIyLMJ5aj4TPG3mY8miZ9AOtdV3LpUVc+6nDCZ1b0+
/7p2rMT9XhY7+61q6UXIyBY8RFduNzV7OVzt0fGemgET0GMm0HAmcl3JNiOYvc7MEnf/9ib6mj39
8d1V2TIbzB8KzvgBJOfKeD3B0c1MBEnaK+q4CZC0zZ2WmzeY3zoYTWXxRMkBgohZp223mnx916yy
NPudYVcLLGuW0e8kRRgh1ilh5BrGcPFghJkqavEHLMtPFhWr5v6DaC0IpfqTmovejxpMVBcQW9tR
82tBA5MIJHOJKLAvPewwi327BK3LN+wbNv5We8E+EStnHMIvpKB967z021MUIIuIY+dpNElUhT7I
QMjPO/68ZhswFR6aXF4qyEH23hTGhhsYL/ehQWY/FDtlS3EbIpj6oOKCLpN39dxP0RzzpzWkRhXx
ria3zUYXmy8HqpyZ75Dh4HfWvUQcl1aD90iJEk+icnMO2q2M+ycFaOGO8y4LAwzcuORqf+RjOf46
sN/+ZFYID531jpCyasYJsAcgmMD1Nfx/qvMu96xS8iEiRH2AhqCje/3/bB3YL+s6A/iD+MWhaXUP
onm+LQcig0oLPgmjOCybjlMj+dqr4Sd1LcjpG/4ZG2AWHmUym3LdDDFTb1EcUzt2l6V8mWbTGRx9
UFLPPIlGBjvMkQUKyjAdYsYoUFhZBCXYwIqagSdSy5UfFjkzD1/dtMMsyypK+1m/z2LejyiGYcLL
FpWdKJiV+BLAVhMyxRGtCkOaQAC6GqPSG/I/tGRhclE9fYPF/AQY5IglkkybZMTLEpIy+gmkKnyC
SxRKwgpBauVgu8b55+wtYlnOSsPJhJzlg1SQkb913vwwOoA29+VlGYDVAW67NUkua8oRka6XmWYf
pgn7SrJnbAWuAABlyBg6nLA5mlpUgWvbU2wT/bVu5RdEV90XrecdUoOf7r5GwfyqCoFcxYXGLkdb
9rMZpUBbKAF+Ta26RQDwIZWn11EzbUs/YhDI1c9Cf6asTuHBkhgBQZOil6CMx+LLwLpyeVYAlMCa
qShbkaMmjJD7L5/ZDlmTzAtBj5d8/tStQ/qWBIa9TCGkU34jLeLV9zr8Jqo4PGRk1Iw2BXHM1OJI
muAuBWtDPSMrwhSLfoJGfjNGPDZIt4yODpHaAFJf9I86dETTU1MiF5oAef5i3LrXJ6LUMztHeDLw
plc5Z1mOOaHQBy0n4HC8vnOUAMYmWboicv0Wqa3CeHNL1JCex1CP3/Y5msc/aIOzx5DJ09gU/JtF
+wEwAf3+rF+3RgKWZgeSbs6FKwnWviJLX27xAzbiASIAFExi05R80P9yT1MVXy+Rsfefa+Kp+/wS
SffAuxcGN/2pQzRNVdW4wVcK011J0l0METiMaF3CGemUextd2HoFiLC4Uprq1eBrI77Bzk4J25KT
abkN0LzW4TS/TEIiYHL9yWxYXidG3fEvv+XEy4eP0SV+BR27hw8S67+eoKu8Lj5+e5lU4v4Cp4vy
aSirX5cTc6QpfnwSLR7vHnFYvUIkgoZEbcimX8jJGiMmSlSeqgH6iR5aGNts/Ax5WkUNii4cx/Ig
2FhZ0D9d9u9Z9oQPzg2cb7kxu917ZmSJTSPuYUPat1nm287P7WnZJPQ90D7YLiXqRBcUfUS55dPO
lQRiy6kamY6kbwMxqaYzDcEu8971UNwfHm4OzfzEP2Ad4eVdV2n2gTHeMFGwttANvUo0fxTheb1l
RlAkCGIDwCGOTXYDiMPYBUpepqgjJmMdsIGiusxOltV2OoEIlmN2UtZcjvli/RfdxZ9xiOxKEMeV
0aPeGH2N45i+zyW9N/dX4oATgzQy/2JWGM3dpBBo/VlRGHn9Q4uZWa9eVzz8Ikc7JDdY4Y7Nmn+J
krPxASK/0a9Yv70mWEnBHuLXMKA3ils79AstUq7qqUdqlwr8jbA6MgaQx9hqs/82xxHhFvEo+86Y
tQ+PpSfH/rApf+5RpG1fv7K0CTFGrJ1J1StldHYgPjtW9h+cs1zPvZ4MXeFkDLYigLV6RpGAd1Rm
7kOIMjx8syEP6bkLlrRPH2iWsP3auoVyJq/ESCL0BF/bzBRrj2VYJpaCMCS8ZS2D4sGBlYUn3omd
dAv7N6S4woi+cjcL4uw38rFUeoyIVn3REKDPHUkWYKtlPo02oUwebYJeE8He7OOPBfoPoDZrGxpA
1P5bD7/h7uUw85Zmwo7zsX6U8P5xdM2Ct9Flddu72eDUYBRGud1MJ3K66+Ju1oBdpH7tV2s77aqa
QN5SChg6WWKeffPtiVmcacaQEj9AIh9IHNyArjuvRpX/KmxDDRK0lmslA2O8LpAhYcAgDYKVJk6C
3SV/kCPyzh1raSIAtD45FM7N865DSIbafMdrYI7ufT6cIjCN1plpdRxxoAEmPv43WGnaalbPPI9u
kS8q27dO01LCH6DFtDkPcpZMIKcv7y5YQQzM4E9tGGWa3WJhezLnMGRBogCaa7RFIfzxaZ6NLx6n
CygYEJf1/7WR+qfoabt1QlAMEq9WtpZhNXtIfihSbAB/jHH2zDDAUXC+cJ8vd/LD768r96Ehsbim
EXtQuz2kQdDCB6jMYvzSfWCo6C4y3gezXKX9UPYc45wtkl2PUSlpgIdndtUqqAE74+69YQ+R9ufC
EhScgr2XYSu38aLgSybwUSeFWpzfv0lXMyKZEvAgicNAFJXA3Qim+6xHngXv1C4M4Ebl2ZTfw+Ns
zb7MxsSWy6dViniQ5+au5nuqm9AgNQth3Y6XXI+gD20UxSbRMWxIKCx56emnMRRZZySD8syyVsa6
bQ9EKFzCqSO2Ja1ioJoBKYMubu7DedYe7v3thlueM5lYZAjlPJWHwA1dJ+U6Lfd8seOMrPeG+FpO
FZSOvDACiIoGF4qK0PbJEdoYKuaxDb/Sr4zSMYWBMOXZHDXeqc9uhe+vB2eu5g+3I/tRNx28UZfN
Yone7mZIqRiVkMcODOn0HPZU8Ck3gZJR7H2f+ivc40nzUPVWZanNU6QbHBynqL+exVpUXgSl4Ex4
bqA9coi5a9GnW3YQYFpOz1F8S5udmzxuTRx+05jayeQbVRVNRu0KBthIolwU43I5QwfkXubQ9l/C
nArv4qUk7yygY4svMSmt1FawzCfUuUa1/NriLZzt1pKeTrNKnM/zX/JyQKLxlxwFXk+UG7gSntub
s+hGWyaZeIi0aQDw7O7l+zQTS5mI5fEdu85DIMVYhgT9vEK2BT2pKIZ33MfX7C1k9Lq9S3O7ORf4
q7kMlsWT0BV4/lfAhPbQs5LNHPWsL3+1CXlnuU3T4Ysqjek8LXD0xs7DJNxxxqGeWw044ya7VwK1
ls6mC9x8KllghWRB7RoXA2yZ8ol4Vbjt1BbCm+9yOBTCiFvkUif7qRMaCOf2d8mBjuuFCA42SQuu
uFqJ2egbeLe1F3HKf6OflbA566wc7YEJHtXzGQY4XZFEfyENSbZEEPgbKgS4Kz8+r8GkRXiTz9B3
bGDAkB4mlKldHTLHjK0iOGMI7Uj5eSI32gJZ7rN3DlIBWGqVZlvYD5ourdRZiRUaphkZ98Pp+6PV
kOA0Mc3HHcdte0TbXufQB93RpcLXaMV4lUH7VfpLLJhAM+PhpLTg4jslw0cZwnqxt8rV1Vm0LeOC
eay03TZ/L/8EX8iJJk65mcq32MuorItPYCfe8yU8vaAy2IbFKtSKuP9R1d5H8NnVVFg2pKs7zQKU
JwMCbnoDubQz748VVxqmdJCHGnYtVoPJlrRDXtXMArzBCLzYy61MAGRcnIo8N+yboIdD8g1sRjeA
rgea482tVmXfrz+QHhF6UFhCZbXhdcytF0MDIiwkH2wbtTRAy8QTIOOb/l0L+iwdixXK5z4TCh0y
bc2KAWNoK+ziEe1lOu7onFfgkj1MvwOMKE3TSNs73x8+Ft2YksnO+LKM0AaMFeq0BlKuMlqgUXAe
asA45cUmB0TqA2Ns5k7wMBpiSNPTUfi4gNtGIK72vzl+5yTwfTnj0Y3WsYD+XTyL6bQvt3T/o5KI
3VbP8PZeWY3F5tyurJPHsShkrev1net3kBxUOyPmDPWd+j05/8SCtHDGHs9HEWp49Q0XJmHZyB7v
R00aR3OAWm4roMzgpUNiVQjIsuUW6rmKiAwaQl/lWlnZlMjDGqd4zww8m7CVZhoY4ymaFL5E+fIa
0NqufI86/fIfsELkENwlB7IplN2Gqit4th+O6VA7P8C3Gh+l3YAufjuw44OwTXLDl7+DG18jrjBR
fRu7da1HKEYpLSxahBksykv+bWlzX4URlzs3MRlxeN/azj3zVqhq7ZJvK0dm2oLA9IVLZUV0oxRf
uBKy0cxas6aUANye7yf6Oq0XcQQUTav6x779WRFgcWa6RZdVPjXcEytdMfkFQJYHTzftIDW3wTmY
xyc4QhJUHgJBJSAER7YrgUen4Rn0yY2wI5cIvOR0L624h90YGQDARETOH0dxRcSt4JJdnQNqH4vp
8WvFC0cZzbMewG6Whj0uTYh0WE1Pop/ftbHLRh32N5o5FpAohypa9mbA7YH0wyCyihs4PmVaheyd
QwgdxVCIq20bDRsdcg9cdQTxd4UG6ngQcdBXgacL/PRBCCEwmhzniU7jYRuKfnx3ReDMEyPbonHa
GZ/Pkqqy91ZlaVh6iYEeCc0ZqbXWGl2VETXmosWvR9ZSIPMSYM3WLQc8epgMDqFma248i0nC5tJV
8CUnNcpoBa2hnJPYiIdf5K2OtalGy3Q0Mic6u5YY84T1bxPajOoN7j/JVPV8U30CMXULUXBjr7gZ
29TuQDsgzWvPZpZokdB7y2dbhbDVWXr9wXLqI/h8MPoqpSddQnjZ8rx2nUNNQV5EJIuNot+AbvJY
ODa6gUlmwUXKZaYqPljq9vQL6RjFMOikHQVp7CNZkPiVZjZUIR9vVLVqPzN2mW+aZAKqjLNG97v/
XMtFElLc3FnWZtuIFi0yDmUpJ2ajF+EelgMbK0xDaw5jRo1S3yqeCP0/sU5OBZ8MavkStqZhUfyZ
TDkXR78Vs4gfeJLQZ3SCd442g/HqJREwtVSrUF9bJirzF9eVop4LMHkrpbzdjXvHF686IJm8nc12
tM5gVc0O3vZJV6OS9R5WBe4WHmRD0fAIoX7VelBWAo9Xs9Bzrmr2zCEPqHRyGT71eMGiLDpAHT2t
cHcahVPE+uiUjGYVuf0svL6jKvXW9vxFl4wKuqUBXfSI+SzuwBY+YsPVGYx8/OF4brAYCFdqDsp1
402TBuM7jZnnpqVtTp0aqyX/SnN7ogULk78RtD1er5bSYobwewAbLkBMcEsCP3KrANPR7Q+d16Hw
S+QQm+769FIAAbJw4vk73sDahhmODqien61X30n2BnH6gpHTmw4FTqwdgVbXt0PEn1jSAuW7pEbV
7zG97eCK22urMuBcsmhoA9ML+GDu1JFaA+42Y3dGn5pE/XSYUJIHs8iq+tOzpy2arDWjcghDzy+C
cawSnWB+AlwgCkeRTp4m5CL3ku0PbOjMMwSVIsHZkSJI4EHDckOhPsIcIXhvcwrxW7ZPegJoFHC2
j+/90yG+Dn/XhrQtvuf1eFcR/3RKl+fm0DdCY37sQ1DzWuYYy3W91iaZuMWcYpB/iHJ2izWuqVfq
fQr71bUcyKzCJwHr0WBj8xwxt6Mbt3RJZOh96bLClygjVyRpWTqy4DjuwN3ovSrsnbu3TSoAtMIb
vtEliLWvwsZ9QGUNHL9ymHU6JIv01W+2poGOaPY8ZVonpr8wzLiAp2wR9fCZj+pWPcgQqxBfSTh0
FsbVqfPmCBVb7+RK3HGA0dfrQF9oHaR2qOxSMVBNCee3P6i5GjGuzpaa/ljrB5jkRfhdGZglY/pk
TR3SJquJSpgDRUCarJdX/aWl9mKGGdBd5O3lVUPINBZ94++zKRinw7RNTAeD2SrWA43o0+vEiC3T
iSAoezK7sNCUPJLXHWph9JuvCHdwgwPT3WhKTz7vzfOS7QogPPpfsuXk1I6wQ6rRTltopqA/i1Ze
RFZ5HrXXuoU5JUKLNBWIl3GSL1IevXpvUOnuekia01pWJRCc9fmoistC2rTDGUEkdvV5Ke/E69EJ
3DGxu7sb9ASgUkvOObcKKJUieb6tBUTSEOc9iQMq5IhUFsGK0oWmZBu6YW0TCQW3rL1tgcpCK07D
XGq8Ygp4gPy6ufxc/uKo2mf+XoBUp+5wfVQ211Z+J2gikKR+W+yfnUdv4jXq49jufCpjGrTGDH8u
N+cBv512eTxc43qzvVD/hTUwsAHNaxPPrQoe3fwvVZ2AlsSjNzykoawEUBAH9eatrSbcCKU7vc80
HTCo/Uytw4EVGGh3hbt0sYAcB+RFNB+vvqoDOqVh8xgb+JEyVrBr1+k+lpOXSPKjtd096AsVa2QH
r1kOYMe87Qu6IQhjw5UfDGZOxU+b4pbKzqrnTx42e/ntI4vG4hV68shMJJRA3Lp9rVSAfumcdp8W
g431ZMpwTaAxtoMCeVax+UBW0rOUr5NGzWUp9wxneYwc23XGfHGMWjVJ5mCIDq3oU2RGa5QvXXDr
8iLJ8PHxCL9Yhtnto3XnT6ksniGhu39RpcJMyVU9iayliPXobrMmGwB/xsIEt5Cvx5vvfRihSlQz
hcFiLRmQWgCA0D52yG8jfRL9F60F3C42bSKducS/UL/Iz2SoFgAxvi8X4SPMMXouXjBkt+XX0F/y
vx1F8Bq/iitidwUCETvOLlLpsclPmWpstB8aKJUu2lD9gWLSMtCVubOAh1F9K6na0G+frQT3wp01
wctwOJuHpB+tYwbN2F74rjItstiWih/KlE+kA1GI1mxWCUejMKmqDYi27UxL9gjdOFfNue3bTvBD
lFVYaMHJ+IKhHulAVEADVAqDwtLX3kZLf42yvz5wVFLBFAktYKg+UQ2EICDUdRM4uOWRBvnel5+X
AFUTnuK5eWLs2hpgtFfZ2d+7k/jivJaswkL0QX5b1LHyeRjEh9CPt2BrytKlfMmLLkG9ZJs4unlZ
V85nCNEEKkkvmWr5MDW4hkWLOS1CRUQpULuFFo+C/ed2azaYjrsdwRDN+Gc/iqcdCADAxSnVqrmP
1junyRczHBW6bZmEuNDc2eyC8dFgFuGedF7v42HV0VvSf3mYOIoGeO35Tly6R2HxZJb8S610WRKz
n7yP/tG97f2H01FbzYLIXlIbLVcVYDgf3wcQe/e2Am7/12zdieeTT5A5cHios5yLCTVlji8auYpw
tnwHW6rir2tFrDIc7rzTVp2ZYu0XWxNJis8T6+b9jHgY+bddPoAfAM6W0fPKaCAhzuznOR7DGQmI
6fQpRMbJ31dIk8DqAAX8pNnAsUEP+8TuwBX4+dIaKjpXd6O7gUYUtl96qHjpluxGHjLFrBYCvKwW
22ROJv0VLhiopI6lFDFnaaQ1SrDZfMNbVYZe2eFxnRjm+k6rjokqeMUKeQRY8008TIYJWRL+xH5v
sOzU5E2XIL0ctO2obLluCECOzE5/dfVp8Q18zkvfp9EfW4HW5+2+QmTkoAj73yu/SjIqoRH1+Hnu
WvC3308ERCvnLgI/POl7RVxISPw0zdzbj526eAAWISO6/l0KU4H37s9XZqRgIq2qG0wi6pueTg52
mZTHhzY1DAH62BNLK2LTFK9jDVy0THQ53UHIe0p3N/IyCfJRxEE6k9CUnafxvJgImXEJIYruAF5g
M2Cz0scA8UOl7Qtekah4cd0tAs1PkCYnnkYXZCqanMAWyvBe6JrZwGvNidI9Npdg+0mTVhqSgA5l
fj199KFmgfn5EnvDRZcPTn/f+GAC3zoKOSR28cNIrddkpGmmywpE8t7XL4GhZFb/4XNf0XrrfgnH
di5cqGOe1LyMgb1dXRqH0xgaenSC1rZePLszfsOYPV06/pT3d/i22tkOp1/VjB19TK6PDQa3oKJK
tav8PIm27hLshhmJ0catpfX2UauPed/GiwR2BMLUaCld9ZDSCS1njS7mlY5jI5kXsUmTkcF4FAeV
SUjqONqbJL2KNDwsaUZzSApTbeuQ1wYnavDiMp7xfz65KC8XaJVJIcUKsMOiUKW/HuY4H8D+mgqR
y5CCz+MOffVJKd5J2wYUqUWc65T/dEliclXiRp0noznTzqKd1Oxx8kXEB617ZoltT8l1sari65CZ
kAKamBavI13jDh6d1PgXi+fQu9LGbbcsy0fRV4UkSSsIw45KWr744zj5KmYrLIsp6F2ziJnSwcu8
zP+UhZB3K9jtHz13HAaxuFJNDX6ZNpiwrGs82YLpmBBMrXORJ5BtyKbcJaT6zQL5a0Ua5ahU5IeM
wvHDPr+2S8jKdmbVaIzLmg94q8NFoxG1HXmQQvwElQpwERNqC8mbfvxobJ3eCs1goibbUVFMI+tb
J5QF+sQsUZMEJIaZ8ab49+iXUdQndbET2KBNtQAAnfdcPMbG2TiqYV2C81FhVLfRZqqNaTJh1TgE
M3WAom8V1UUP1Kq5EZsOFU1fqwoQlr/Y0kloV3mJQHBDPJy1xPDwbK8YPQsUj737sogNmK3xZK+v
6cZYsB1tfy+PvPpAp7ymhvE3471khiUHE0nw9HCklETuWTBVCyDx8yBbEzDn/ug1h55cPJLtyD+m
3hPrvTdZWyZEkbSq/Dpz6f6QI93HlYN6T8zFXJQhLxz8Uf3UH/eVDXq234TLGBnEbVi3pkbd71qx
zs1ZrpWTA0CisyC/ZsnR8UZDoHYvCZ9k2NOtFkMhdwQWWNLBvvHTor0xcxaLTtBz0MLU9f/BSV4C
oHU2mTw6rBIq6+Z+Nsiq54L9jtKTeB6oq2a2fQv9XRrGtIdgXVM+BpgEy5wSqvwgFBNPnxc9X/ON
JvTTC4vp8VgNlozdSNmi0qP4Ob4qp1NWXEK0IXhlDWTmrTqrFS8xRUVJt4v0CVzq2nX52+R+CCJb
nX5+fEwgR5xJsJviSI+vWkQTpK/PKtxDcK6vTnTnE0+8DpC+vgK6+CfBXBINfCnFr6CIhOCTdJ+l
TyVwXL5QZburGmnoaRTft3oUlF/K6l7ObxvpQJfIZqoZ3uO24TmJluoLBQWSnEl9+WSKBPeQu8E/
+q/dZpj8dYamSUG+ubucWbXIBIAxDLqdjtQZVMs3iTJKplrySHkE5X8I/4ya4CuMvCn2uxHJ85RS
mDbw9W4E2Te0qjiHIBG7dLfcaxof8NOOFA77ano6A+8l3vR8V1z2Q+vfzXZhU6vq5Dg8OA97Xt/s
rey1DISe793osFrRXTqCsNXx4SPNqRkaLlLb65fLRa/eca5gzDaOWATDDiXLEAByETjB6v9/DYas
WJqDVEtx2aBZM/+2lw3fmNe9FOcz2f9BavYIWlEnC+c4vGevr+3xRA+9vams8I3kvKqH/REW/OSx
A3ScbyZXxpoyPYVk8HmXX/86QzxqgEWBDoY5Byz8PXdpy0CsQU03cEuUelZina4Yh89bZQfpJH1J
veDQLfKx46aVVbrMSJFXj/ntazyHhOD+IV4DqWLQVrZeNSNd7QhtFYc5/+RKWGlidenSLEWLJQVH
ZtrbGKLRBuZrNK+7kFfDu3Ra8XfUWOnGb7FOZ8QkFOAUKUIrIzSt//TskUDMoaFYvl6IfEHrnFn5
DfQecyMwjPGNXhqChTTJUPDnxmDlYSratuzlZykik5e11pdYwVNSg7XMg2zmCLQWtMyXgZCqtYna
ZNZYq+ccQxwaH6CnKBanAqS7Gbk4q0UTPl21Co9XBIVYSHMbxq7F/2eJJN4Zx9ECi9Dt49PMKYKg
M1jQxFZMwnbGOqswesG+LL2i3jwnZaQdLUmPA6LHYQZOaM5mCpNP5yK3IoiRxh6o8fcDGUiLuSTT
Kkjf99Q7hrHWvcbV2pFECynFjMjhM02Em2tDhplF6WJiE9oZUL3rMhxNpKJ6ln2l6b6bmWt3kbxs
n9tDIj2OTxEjzBoaKTtW03GYfeA90y3SRd7MqeXe70EOibOdg8JsPLpMMconJoDwoLQUdGiAUBw9
qQQV32GMWCe/6SVRvxCxQwXdSJiidH1qs7I/S1wep2u2ihyL5SCXglbxNfmKTRFFNs94xdVyaqE0
JBPgvHSUu4sz+h9UUSHfGn7KzIhnCxLPMYMMp7pXy6KLxj/jFV7dvpgCIchjf3u/z2k4l1DsRvg5
2xImoJgWFIbMjXhBIAArYv/AI3U1FXaI6uUhTmEmufVmBOmjuqE+SNlCtC9iwAB1E7Ne11gbMRt/
f6fqEYzHqtI0IM91qNAqEShvktVO/Gp9jFIXQ1s6uLOEKvhJUxlBiM1STAiahpav0HWvJVaNQLYN
lokPsvlt/CgagKD0jwH1zYVyKKbAgD3rY0Cd7aDVfbrwLfTfKheoCygAndhM5UEG81+I9pI26RCQ
Ze7hokzJzIVh5QebCndqyESAl8De3adAYGeHXfeBtFMDaReNVXL4FZJoxBzOmv7sKCh93hAQQf77
uLFfqv4faGX7tBbFbvCWqLFByHOQh7KLWtJoNVStopgDXKZQjIvagiCgkXoY32vb6NeXhMXZuMOq
7SDzZDuaE6P+2CGhKNJrJlSnJszu+8qoZ96cIMWBqGL27KYHGe9L7MJB6Y/H2ePzewk3fmCoy6Fi
9dl5i/kpkSd6eVJIZ/QR3KtkeTVwF7YA72gEdbqmZVEMjmkBWVIr4QLGGjydbwskjJ395WNoffbs
h2ynzznNivwSxEqf8NLL8YB+K72lV4E7Gf6rAU3OvNGOtAPuxZZFdbTKIPVTgPsqoiy5Q9PqzUR4
PCXOTPhEfm7ZH2QuaDpAY/V4bZHX85X6oRWX2wwksSLDdnobwn9Zkd4UpRVavBp7UycFqK21ItKo
wUqt3IWHNLJhiVT0MRqH56ozZ2xrn5bJ+gFLfRVkCOmGx/jvsS4HNKeL7FEQ5ceRwpKS89GuKrkX
NpGEhcq7ZHT6NyPzver54c9FSpZ6v2HNwqDvWW/q5nNTg2CgFY0bePm3fz4xnS04/jIx2BxTlm/b
iPVbPXF1JGPN5XPv6sXxOksbe8I/dT3w7rvj5d1nDojcMh5WRcxUwQcGEof/m+e4Zwy4t57DT5zS
lnLY2NfEkf6Uf5UhhByKpdOiwUQYhOFM43rlVMTxMufa58qrf+QD4mOq5Y6X7EsbEngyVfWvPdB6
V8ygtXPu7F3hkl8uPvymEMZKRxe+sjwa3ZWrOGTZXfnPGPPAKzyD38NbJn6fq1mBpIlKoizClekR
6piMCJrrbvlGG66Ts+shnJgj3Fpof0zrOWDvWjt3S9CLH8dLhZqOpX1vm6Q5Xj7ZLl09V5tjnT7y
hucCA7vEAmCEbZr2W9UzGOdeJ9d2+05UjWn1b01FXxbVOhBViP0ogkohG3kSENeplm7UPNzEB+ho
qEFMJzsiGYx+00y277k6ZIor9caa9CkH0WnlfBZCgYGHGxX56oFSDitn54hOWQSWl8coNKTnFpoE
gozoagu5SXaJ0tjXSUuaXgeVUbgIpxKHqXyg/aRDFj5x84h0jwYPQzYeyxJeE0/D53mnKE3Snaig
ZoYhUsxchOazeUjuVccGvQuRDKNKm+Nc9IJTSIhwL6NKccTGKPJKTp4/S/Nc50txkGtULduoWSiX
XRgaCdpYB9rr221AEL7ES91ecskVYsNn20A/VzyQrWoR2JNftrxO8UX6wF+UG7H5gFd6GkmRJGH8
mx0gHL4Batvp4yOBDC0FM1221uP1Fj/K5gIdvuyQZsnP+wRWKQp/BUskcMRY1J2VSCQtpbhMpqRB
XUYPH2k/wLnP8DCtvbqLchMY1H+4xGEDKUooGK9X+MShjMNlaWS8RIwyAUDJ/zNBDRqyo8oFo5xk
OsjxbdNb6iWn/9HaeS1Ic/YSnxGdOKa95XbQVVO6wV5yhuTv8Ox4jB5L3/sX8sKwHsFYqSa68nbp
GR6DO10U6UpnKYFiSOxTswdWs9vS/SBL41SiBaBkRV0ZqfM4v3e60nGd14sAv4mb2nUA0qzoiN1c
vAuSWv6JONZBlGzZKrdN4aJf6RcCAWdoHtAJeJT8pZCpC62+Ww6vLSIynAldaUhnwxdi+uBtIjoB
cK78Np6YsUVNcW+RGUTu9g0pHAvovHnWkkxMG6cnYD3wpZ3c8XAGkDHLLgm15fVC/llQbo6IRErR
ndZuk+qfcaEydtdZu93LHgMLsufypGbGokOK5OYnmHSsA5xxOiQStL9sL3jrN5/PVfhKT2wUQI7t
Ency/BJmbgW7yoJtlPNymVQDgcvy9eYCLV3nzCtzjcQzqzyXueY9JCDCzypC38vBiSkmHb2hIVsC
na0mUFjRAj1cXc06iKGcsa80xOkZ94cDsvB55Hr9avI41Y4ex8joTrrdIOz0nI7NZavJkQBrLDIn
T/yyVZ7EeingKR3hvYGISo89LTGtoQyGSr4iR5d97QXv3A02mhTPVlfN4xMfYH2yr+wHSSxRXoNT
2xPR3AGeKp/BmQ4C/lLpjVYBKtoCp4f35C2Hc/sEC9G2bTRTgC7HPKZ3nsEGVkPsXK5mdHOgFY9h
87P3iHsoF79t+QKPzZcvL1H8fDeYY1ZktNUjEWDCCq7J7nNd0WNg2suIbI5CrsGOLhjdJdy0hBIY
yyzss1S704V2lo8k+MTvbkgAsMVguihpj1YQBum0qVnfSBphgf1QZtt9Eb6jlMdzC+XAFEDhsLiR
qZkUz6MeOz61NvO0xtNiFYKeCVuIePTnVzzcYd8Hcr55coPTmL5eFNLZPlif0kJfcF5yLRC/yXvW
rz17IlroFwPHLTdnVxT7zkRuuAA5lo4UDbFoHbcco2EJEjcpQ6+1NkYg6682TH8UxGnkH+0nALtZ
HV8urB8e/v0oivHdrdA4SaZDMSD9vf7HFELbbS7iUMswdQ8oWrFsLU1bwWReDeRmDk0T1OC7axLJ
/DxSUjCd1Ob6EcGcmDzyU/MaN6G6jzfAAFz4NQaW7B6tf1vYHiGdM/1MbzvoFxRBNMV5f6VdVIe6
k5B0WtVd8lkNz01ccmDb1u+Hw1J7DIrnnFqb3Alc3xwwt9xTKWig7yn9RnpAO+IX0znRG1fhfrum
nlGuPkGoAgHR4zIAgc95wJoY6Q63vcDGU+nZL47RzQYV0EcTQy6WMARdZ05qPEk+6Ejjcta9BVu6
zurENGxK8UMXMATf+gkFJEqdVtHYUOiGdk5Ap+deUuU2a2L8esR2aCvUUpa/fwoXJpTERga8qeVI
GmOGhu/PJ1GdKJp9Sx61krQQ32MkbZoHIlztI4VbPakJN7n8qNW65Opl2gCpikHN0c19M5e7uuF8
AfQe0TfdToh5QK+iIPlMz1wzevxQlrrIUTit/PSDzASTnaWcYpSwg61kyFh/I1P0gBJfh3N08wpQ
NBg61MrimunY5uZyw01AgS2nOpoUKNKxUQWXgJqnwu9Bb1Rkiu6a+uP2PwPI5obdGhNH9TC9Q774
fBqdRiMn4Mn3QGs3RAK9esWD2sKYKuowlwDPN9E25+ER+7juJtSWUVOGt50wvb0kulGYIrymQINO
hl3fmAPZI4aGpCCLPBUyl7xy28z9jo6hqnbwOPSzlYJgtRTgxqeR727jhBT4Vjr1y7H6Ec/4FIMl
kHizt+QJFBNFC/jsEJmvf4vV+XXaAmYdvq/v8tiazH8ouWwKsTipnK4hDrqCd5998woGfbejbFnU
V5cZf/tgHPJL/td6hjYzX2aHLcWaIOY3koupMNpRNrTj9vPzkgmEje41Gdl+4/JFhtR6Uqn3S99I
PlfBvTlz1BNklJqW1d+b7cxs6ICjON8PUK2xFjat6tLAzZMIzuK14Zd/4yEP7jUFgZhh3awybLeK
92krOWq+wSCnVfPb85YByAN33iDTATwfdHDL8lJOprKjwPCqluz8WUwpksfdiARctBIij6kiB/4R
gIHs15wBInv/+91d/BwJkXa60sCf1jRZdHFkoSAcHTyAzSSYakmcv2QpEn56CUTQ3upj3vUx0337
pCaXi+AHBxzDuloHVaJn8VFchL18ORLZPmcqyM3lE/IOwz6AShT2Ft4jQt0m0rZkwSA++vB2p1jg
q1kx6vIK2q4dd3fyR6CFn7ixCiojQfhBafPPJtFBp6Q0VE6gfM6pO0iWjqbY4l/KVJUSjJ3duZPU
xMqD7XFZgGvLo28Ru/+QTzV19HHgBhPJ2zwFeVOWpD8/vQ7JnpuxnrzB/eV+5xwtJ5yp8Ql3I8sj
4XUOxIZPTeeElomtQDQb790R6tB5f02bRx+TS2MhqQ6Cjp6oEpJQQC8xPCJWLsBkMn3APJYjrpLz
oC7tjafJig2p8cZdWst6iA+WNuF7Gno+oFdBcoTSqnmrzMGE3vQD7xnf5LSpOeq+UOtV8Q4jBDsO
pdESs6op3gguGPRVIX4at+oByWwTk7orJV4S+PyvP+1rAwEpzYuLiEHjcxEPSfGE4cz2zti4cKdh
R08pWoRDGy9eJF5H+n0ciZSFCykjPm7GH5AYGGM/1QMRsVpMpgBTBe5Bbt7QQojwMiDwDtnQWU59
Bc2OBW/RRGO3bsTfVN6EYM9CsWX0tgKwlHfooSeDyfbNHAKpSfVjUAoryRgLdijRzEsnBkHK/LvG
V9PTDsUKohIR6SrES0wto1WGPiaZA7okK7J7HDamR8FZuejdZxCV4ptq5nCkchrLtwox3aRcQ43Y
WnWZuOX347J3k25F6qk7qz+PYKjAuCU7VSXcY4ruWNX7DvKCuhVOtUd9llnXBXiwvvrnGONo5NFl
gAOFYuQDIGGut5VeTsmMSRMVEG8BOR1/69AXKPLB05h++dJJ+wXmpw5OHAjRkdEfW35/NOWmI5n6
ddkFwP4v8xaR04x+5MNB0TQhIwcdJT9NzXKVsXvTkmBFq++kxHCJywfAcJor7ZYDb6RpFRdAKuom
JbEnvCUN45v/fhd2ggXvEzmB9I6+UXRlZ5aauc1Hr/Q7wZ2qR9UiM6O89BcKtX98le6m6TZH+rCr
OPerGIVc4js+BjYizoKsas4cZqr6bWz1ztu17bzR3O+KnlcPVL7YdBTO5Qt3omQCrDvvlrKyaWL9
u4llpBoaSueg4PoN6LEsKyrLqTZLXqCB4wnpbd0ahN7Im1wjuUE3xuFRIlv4lctTfPr8DdOGbimo
kkD9xt9vAhToXV5hX8hMCN8MZdmxTCLjOcobEySA4Fm1w0Kgf5DBQzKmyk5jqxnUkEnh73vADZTR
DAMveJRFrFZni+jXUL8AsuJlQq6BKo9qh1S8HOVm/jmBzjkmRFQ4qleceFfCeuePbNiKQnoDaqii
8v670TsR3hmSUfPc2jmcasyuMe9+9j3aHRlIlLFYyF5cK2vPjtyTFMirndNOzh55lkk68Jpukfgt
YmpZLPky2mvXmA2YhTSgC/xpDmKe1uP4zPOGrkw53z516+qw8pdg4fYgD/inDphBIRaNJNiBqDE7
Ue2gKSxa2XFPGQN7VHHcAbI9MTN1i4YCJT13FJ+pwWg+SvCWAtxrjXfLi5t/MKHESb18wvxH0gAI
slDrsZuBMIFgHvh+QKsxSHOxZVe5ck9XMv4a35qoc1z+mJecbI5t3x+ELQ+jsJIWcSOyVixBotjw
YrKuYONpNi+6dPYGwHHNU5Oq7RTPtqRcYBrfGrJXOL1cWfrYLe0KYuLMmVrRFvSOKTdIv3+VjitR
uac50Ur/mMFyER1QfkXsvmv2ySuHdrGn7H4tQABbpGux+zuXwwr7Fskygi9wBM7Os6fG6GsTqVdb
+y71t6rMsg5rglTs6t42qshjN7x3BL6SpZPGmkEDyqQJ1QHo2q+x7DetWCcGEoVyJyAi4A1NUKQK
M6Mvs6nCECuP5hVK51V0liAjsNt8nVET1PjqiUGF+zmRKsNvwXVbMkItKJnT6fwP8m0I2nlKPvLP
ZVGfodZFfC/8avfG5yarMv90ID6sFSeQYWRwp5suRigi5c/Ddu8UetY0eiHN+4U1qB+TvJlU1XKR
dePBmAaWcOLgJY5kpmMjPaES2FSaIE61Yq59XT3KoVp05XezHpYeZNMunXqkbuiZ213po778/gLD
dEr/WUTFr3YZtuPy6z7KjhiERYiR+iXomDnZPwLai7hYb2oy7MfzgUEuyozjj4P1l/lIZar8UK//
XZofNzXsgTwugQxieVaUSq6ZjFTQ1QrQ6o92ma0MYas7MweYMU+4vPoS3vctedMmKp5X0svFrzlH
h/eMwJFUyEy9dokrs8Zz8XgguctcwJ5XTh3bzACwTXASP517am9GDwDA8G97VzU31moeMaPcEm7X
7XnvCTSqAowN/EgQ7pa9Izpjrx8KoHEzQwy48VcWaOg9KehtVxRoH93AoSRhvISH6PrlwLkY4caa
FNJo4sWU5p7+Ti1Wfxgfdd0dT3npnIYcsCuUPioUpC+Ykm1bCKZRQFl0FAlzDCLj4lRIRrbYj3rb
SaT9Q7AUR/DjI+8xPxrYF9JqsE4Qvf6fXgXae3rUPAgr0VHatomkllQyg3RFt7xZov6+RhKUWC2T
KXFhfEAoBK3HFF6+Q2WYE3Kx7Wz6cc49TIYAhw0GEhFpdjwOrzYa0tgSzYrdNwgy3OYomxFLcVKJ
J+iY/4u+XJph1VQqF1mNDqmbH7utH66Oi9bDCNdcbH6K9IuM3kyWdYtxnnt/5IapjCVGVwBURrOz
dfqFKVrhL0Dufl06ERQtajkT/7JZGKG5/m/5CMofIvOzYOZuULfVJsGNVSrTnFcn/sPUJBgv5X7W
HTcZA3GV8E4BYgxoxIKJ4514eS0MoVg+8J4yj2JzQ82dYUKlobh5uQdY4uq0KldrKIWNbWllX8fr
9A3AOq+Klr+Vjjgi6rLMMCMdKPs6qGqjsuz2b0q76IknmPMUuuaIOZqRFzFweGeq9ZacCZGsF+0v
TfNeOfMs7Zkc2vwu1SHRd+ngJjEwOwPIvo84YTOTJDnRoDouV5kilaMRP6TSmVIzJNDcuRYsaVY+
d2rXpqNR9m/VhadJywR2XzoTSlKOrVckDCNM3SOAwnSiE3ROQDURKg7oSEUSWrXIf1inx9+botx6
zo6o/XImcR6ZsoP/4RGKb9ufjLIUcQfitjveqOwVGyLvo7MjCM/RUgNBfchjUiaVJST1/bfZjYo7
7tOKZx177SIqRFZfP+Uc8H6+9cWRYy89YPlbM3ZK8cCaLQ995rTcscE7iOGyzqnDsEDyrZPeXcvd
66JEF6fN81Yi8rUtgeHZx18T3KnoJK+FaegDdC0dcX+6MPYf+DI5/740Z9JZS24bZEEbbvQl2J/E
zuRstBoDJjzrOCZ81GG/XYFlN4JkjrnnkDI8LSC2fl42vX1SWWayBRgbJ6u+YpKzwKE6odSXk2Od
LZhGoKQkX2xwRn4y6ELhHPakmOzDlWxjT0mZ+Bc4eJOgwhA9D6MQhXlmVEHg9RC3dPv5ih0KMhUk
/gjgrfehGrfK+riFEMBauspuiE4QgZAcGnv9fK0RiGl6Ol9nQ49O+0JIQa1eByjuhuZljz7Wv4Ul
Wn9wkA1FqWnVACkHqN/k1ulunaQTsRxTb9yzO9lIfBOjzG+yQ/8Jw5YOn1ApO1fKw+fByJ0Iyq12
QB+zTOeGuR/ycPjJdEf06VwmcawajnVIJylXQ+LavUX1xqzbUveZFi2tOktMHiUWpiG9TTRGpDa/
Wuq6U8u9b1cj0BzG3qHSRrj0Lfs7msOYVet8ZZB/tDbXzhieQ72ZYScpiI+j4BDSO+4OLIrsYw8O
fHsTqXTDu12aKX5SIKlUyjvvpDQ7CyHB5CF6769G+yXmYEPf++A+S8QbCNJocICbnZ+xBmCD93+e
IlAio4tLG7CsEaqe3oHfKoloTt6s+M8tgaDFKCi9uebVZoiKmwbWWSXb4GD7niS/KO3usdsDpxZc
Y8yqN8g5F4SrhqL+c80/9brnxtDv6vpXQPNtaONX53+Ix7m+2JpLeWSY6SP2VLu8QgbGXd4AvU0m
mQZv/yGzK9gLPq6f5TNmhuQXfP4WdyUeAr042bWXQstVNCRvZDPwclayvaLs8lZElrrG+Q2qu528
+MS8RbWOW/XzLbT//Fa9vm91IyWiu1jG7zfJLnnZ/qKtvrCC3XV/YUDmEyTDHLCI40dqcfN97z6h
IjdnDilKSQ4pEYGLV9tjULk5a0hy+O7lzVrXisFuh0+iIG4IyWjMd273RFo+JZEijru3Uiciw3yo
f2OVY/Y7NEgQpZ49eNxIogBJksXlChrjGPTYr/rDDrQhDzoByIIxkuLOJv04bJd8LzXgynTaeJGN
KXsnd08N7L5J8/v7rNAFkO5CGamuiUwz0CcUb9dEI7StLeZeNTyLC1uN66Ltm2fq+5mx9dFy0hpF
YKvOaGMETjAO19lEY/am7lPmme8nR7RMu0lZG5y5rMwffIBWfxN/duSRJC+JNPYns9jrdOrjwh3w
app7pJ6PIVTU//X1yIlNAxdWbU4uGAB2mFqKyl3GeDC2J+QlhQ4Suc3jcCf8tmNznD+fyLmF0Nz0
LS0llesYXrEZpWt+zznoXmUDvUEFasSgyXQxX6Sjz2GnNLqktcL/r43AyPjbRZwvGN9BIchOO652
/7CUKqKDxGUXvgxlJKiq2LycY1CuII4gW9nAFjurODM+jGy5UgSA/uwGT1ZQXsxeU4S148mtX6wZ
YxdqRt/T0QHUXL2kGLRr7e61kMeZFpv0zjtZ7/hZDLy0Yl8MKLYLfO5Y5byRRNyBMVMp4qhuiXWc
vXGziegoBXwH7Y/khhnl+fiy1c3Ij4PY96QvYrM3UzrjPeY3gt8N5tDNivbofieSZeEjDVuyeUM6
Z1Mxm3bhLzX/mc/Kj47fVX1F5q3ShiTRLwllFf2vPxrjPj+oGBECpHuFLl+H5BFsRLuqgR65+WE3
vFXteG+WxAqym2tUwYIf1wOBFEISJYGvOo2VoxUYGjjZoo4WqVBIDEDbKJ+/N+pbRhQ/zQ0iEUww
a9CCd8wSMWcQykPMcoSn4iecYp+KBrHLfGxJNGSptFnOEDSgBF2lPmw8bm/I1SfTHR/WCKYC0PcB
tL0bgTHhkHa2IjStkhf48Sggxyuj/MDBim3qWaZi6hlXyaXM3JlAmYz6HBvtnhG0bEwKXl6pScjN
3OCADx+NqrRrgsyfF6AHrsZEGNFs9KOwK1SiqFXuZwwi4fh0HPp+Lc+loUzK7kBzZLGZOi5vyMze
c6jPFKXaxa7pegjxm+wq6CwVhH5JoGgMx9afwRpLNRSg8+LexZFdf9EEU0iulZTIu2BtgZf/ZLRC
TAfmbA+XnEz37tofnVNgcGUW2szlABCZezeo6TwQut9NWR7Q8VEtffOUIPZaM53rq0dB1ADDAUsJ
M0oRJRPXLjefFe/8LCXR954de8pf9NGXsTBKK98+ZDWkJhYd34Fk66IGa+UH+Rf3zuSH3QoWLZDW
WC94XZBr97ik+f37oLm8o92IMsliUPVMN8tTwdzfv4c8dvKYgACEmKKzN48Zsd+hOk1vxJ2kHbgO
c+144vmCPmrOFGvnWFuE8yMXj0rNCTpcU7ZLImqgxdiswcQwTGKDvt1KiRgbsS4a7SKJv8JB1Sog
4vRvgLyz9e2hM6gtZkP++rGQLaEJchvYCvMdExdvLLRi6iNtmFJj34jh7GkVYPSUp4CMNd0Vh29X
9VfbW4l6vcGHJ1okGieTj4zM8JYVELq/dPreqhI91oIZmlzux0JgBdchuf/Fry946rC5cGIeKT8M
XzriF6agPIpQ1CxmosJCDYPnD0TxZU0euliqs4/ByfJfVoWgviab8bgQoeY/mtOcI8jMFMEvf4zh
xfbCtTJdRPPfXKl6MWm0al3i+DtM9c40myEUPXxJPQaBHg+cLjfW/d+pe47/5yTuMTqw6LsxkviM
4G4JInXZ7G4VQNeXM1Gh7XS28YJMFK1k7oU4HyM6pMjpXdbUWzk0FBDmLG5kyudhXhlpBm1eCCB5
qfrRKMkxlCKSY94eJOhEs6rAADq8ZVYpYTvLdQbnEwp6MYc0BXEN8QadfkC+fdRajJ7q1tDiO2vb
4afah3ja9hgzeBdBJ2Dz9fk3rlxmZdG2Jeu9PK6+N4lYDer0jdV0JCNH7Z4W/yuzrB42CywyqSl1
R6po3qvoO1xv2tHEY8IFEeDsvolYYKLCaa8Rq3o8whW9JkqfDD6NgDotKCKpICH0+QxKKNCTux2/
tRH+uR3HUAXfybwim0nxORC8dzx3ln9B5WuLDIEyAin0pl7PWQFoGt2dZ1b7vaUt2PWpeBnm1d/d
GaPIH8+5KV5mnCEZN922I4YvgusxTwHv/TSaHvwA4QomZab3weL/207g8pX1aMT0H6Aj48QQg67M
HCb+o4JqNwvKvknvfH6bwfUhr/OiLlV/nkEqQjj2BnjzV49alHXgjhkcoerRaftZ3lkZUnZ2bopb
1Cj0ws/aQC6vavejd13MDyjR449a5meXATrVGomxZFB9Kn/eNe00cUmeU/L+fId6lCWA2bpmyZvZ
2R93Mmv20wCkd2n2T1y/GO6dcynWv5D7MlmVkbhNO8VqBJ+LB04+wh2omFDW4kqQHxpFChTLcp/f
IUOscp0kHDRsjNN6oEw0ArecdQLRQ0HeOoLUYZ/EZgdcpZKrd7NmCCe9EPLwksYnyiPDCGO/2oAK
xXeSgPWSGTm9B9kBzGWkNItQ0OloptCe3LM5gK2uQOJsmqmfa1DGLkPZ0lMNw4wB5fU1OSP9nVoC
FoffRxPsmSWfgXdKs8IIvdKEWKhqgiA78exDwA6QOyHKh5j36K4hpXR9lgi05v5qDyR//AucMhX9
IVGLMk2+CM6thg8jDdOYplx7XaPC5R2mdPbDeJJRXkBHH+rkhXx40QoY9FIx67B+0OOM/8lecLa1
kXrxJtmph+6valYyNknaEWrxLuF5B7pNgDGl4mZ7r3eSBvvwYMaag2ZT//6JA6a8W9fDPmPJtrlv
7kPVFgnBEunGKgUMnMw/T3AABaVQin8L6bXJzF8gBhQF7PErlgDrjZZJROUREqn+xe8AxWh2t39j
BTCTYFVVEZyMXJRjkcMak8O9wzIwF6ZizxcF6UvkiafRZe0oNqzH6J6DvzC7tzS+ZQ1WBOzf2gCz
tZlJrZbTnvXb6WUCC2NNucNHcVNfv2qZOWLC3DFegWSVpYYn08gYMAvgQ1lnBX067y5P37hKvC1B
LCY8aVjefvcvMqL9gzKnSBxNfi/IvdJqMIMzZbpTqPl5NEDJfRJlQ4ABDGhPn2EvmU8fsOHzCa+i
9rfuF8C3TfZJr81jt2DFz5F1jFys9+HTEIQsAXzOTb0QhXVaF5M8jwrVtjCzdPWOp0T5EC5zM22r
4B37K40CG6nvBZDrSiWAD6ZeKcfCji+fMya+1hHlcANUOuAPgpZuUaxebOf4+T2tm4Ivr6ccmnwb
cRhbX+RQdwXxGz0f/aJ1AAHQcrNthMY90brsVyNASvUpGU5EQxSqk0H3bvfmZ3aHjx81cwEFZuUS
2HE43f2FRL/lKBUERQe+7dnh7/cyoRo8CH+ekU0l+kgGvNRQ7QD+XJtzHcFibgXfHlO8YCI2JYZv
xP0rlQ0k9D4lwfAvYOZPPxLjsrqREmWck3kyc+7ThU09ZsV3rOc341jCW0g71g92uIl5dDeQdNGZ
iSzkpaD5dup+TQI1vbwkF3ZY/TNYEls07cPeKdnt8mRXJDZGHi+3GvQoTBXla2hqUBLzzGCeup8v
+/TM8H4Y5wlErViXknkB4fF8IW3pQvH+f9Q7q+qEccDs0hVQzg/DJTSwZJ6+TVXXvFLDr567/nIo
shCfRhL+sWC2aZrgcnfmL9dnD/DmPvDIf9KB+rmgODZ5F+uPhjcmbzFsjy0CV28REcG3V8tjxMxu
upC/kqT5QJ+BhA1N/quNmAUJ73lKL2iNvFhBpzkvW5IyTUPFLYggL/yg/rK1uLdpniCvbdZVxp+C
Y9UUTeyQF7vAPXX7qo/Kcxnz6gByZPOrB1rWHrzmfYSfTiD+bG9p8hZcfw5MNDdQ+QOvnfs69LVw
zb+G+7KL3AQQ1O8tuoSG5VY/lA/n0JanG4KrClGCZxCnF4DyPc1grDB35zoi7sdNBn9YYNXMsqT5
F651dmUby6+XTeYC1osfmY1Sirl6vJDxL1D0avisKw1rPAFsAOukzy3PfLa/AAZiCUcCRI/45xsg
UWWmwJ0akLS5gf0p2Ok4i2E9dQnDdijYfFlFMMGGK5y/bz3ixxTcKd2mLDSmzbHp0jiqcEFtylgw
GLaEwwy+1mQYN1chrklqGWuQW1bptjOwlfBBE++Z4/qdB6+LZ22VV/5+ErI4EW/azxRAf5USlrj2
b3SI0G02XtdaaAEyYWhy21Y2xXibQs9SYg+ceRUdk/vqKglAmdi+T0iHZyY3WsCuZZx2ybNvcSMS
dMQzON/toxHl9UuKH/sfKrCNMh0a4PyVp3kzcxfYf2SmNMjoODe1hqne51BFWpOg/CsnsVGoW5py
p+wXc+oLR0DaxSmlspaN2xd/FZHL3WvDuFor/XoZYgWU3bBE8cSd17IOBh5tc2RfgC8gSmQJbE1P
YUGafyCFO0Ygw71XM+1x7WmObBe2iCVM9exWV/jc9n5Nax2MF4PxRdv25XPeu6VNy8iZk0D+QvPY
WY5csIztdvHYHUQAQmDM/OUhW/g3+q/e7Pma14fd+UYv+l0Zak5L0zk4xLcCfBKDebTIcaccReIw
zHJqDz15MO3gCCj3tme+P6K3CvgW4bpPUxWajJHFV7fpMUgiU0cWVXFzgxEH5ANflM9duo+8S43Q
80QkC8qfi8nl9b4sQtmuY5vMuABjekwT7th9yuO7Jt99ENvcA8Ux8QZ52pPYgnQArTSLUhYmdVxA
qGbWcVbXkCusPYFg5/vVV5YWNF770dD5+7te2FYq1OkuKMJOEj462cltk6c1jI+GYMXoFUljxHku
ao/Uu0M/zcd30jJcrwdVLcpE06RFzwbcxO0Odh8yGipKdeAmgAgm4EXYAxQvB+eX5cAkgR4lGgdK
E25TVpEPgkWL46JvBrEgBUEZux4QPjsZP05EYW5XcmnqEr1gwRmFcusxFQQIifV5v6fr1PIdgWIw
oMHs9DyyCvz2mghliHEoNmpJU7ujc4ZAi8xJfE1eUCB85OQTfD7oMolI+KSeG0+uC9S7VqdrgWeT
IpPN960YuufwtGnh6SCX2lDUTV3JwqLMNfAMG8bVKvyOREL3TB3xykncz7+7VRdVu/biOl+PW+1V
TFJCkG365uVBuqKvclpKtsA3tAgeGJUBkwrCGpbvaCjWoaGIDOY2Ql5AEuIqe31qgvAk1LqFBWZW
6g1YP6ezj/p/zxze6VaRmPgOyWZuSQUGPWuBZgUyirLP9K0xNd/N9orYwhTrdvL1v0F5GnLopL+b
HVmNlgiSTfM4v26eruF9wYhZ4cTpUxV8IsnOuVw3pg9+Z+6BzGS/h0DXp9V3eZ2Vejusj6/c8dsU
MHZcTEVohC0Kra+6gbX72Zs65lRMXRlyud+lU/JZQFk5NU0YBw90yQbsd3MqFb1rlYZ/otPnhj3O
+NWmORZWtVoh44JvQ0ZLWjvf29i7DUCSkkjfhLedCGNS9gml2RbB1PdJYz4MatGP4U9QlQjzN4N1
a3RVnG3u6OAt5bciVxTU08rx5wzVNuCcFLsv3MVqTFH2KPtWU5G74LQlx2UFR4euHt1enOULSMac
bfhvQf7/WPEaM6fahFjoeSGFtiQfAybXLPlFD8U+hrXQpqa/khOiMEOC03p7CnbsnmktGAaQcmX9
tzMxd/Imsrh8II/Yljx3kQmfFRDQH5jbXVa3RN5vEK8SdxFqCMWXvhevzdjECqmLfYan1udVnQNG
lgCAotHiJEaxRPSJ0qi6xuoSUtzx78bOwXr3NRxkGbVCWPtRTyQPdszlLOG3fWN0F6aFgjEiUoIq
gBVIwQdAeJZ+7NdM7Jqw9BydzT7ciy/7RIQcupW3stlAbV3Kga1Jo3kWiEQqmj3f7HbUWpDQ8Pqk
GFzbA6IqWog/yROvFLm+9jW+0GLoP+Xx/NK2upUhTAdo+2ZZnQ6QmASonwyxmPEPPZXBt/gxHe0v
TKzIs6j057QU3HZaW2pih383VgI3dEp9bAK10tmrqTwQTj9rHzwD/4Scg+j/efa1GxZ7+sRaswMB
A/Kn27bYG9lSR869eXEV437OuLQp4qPRI5SzQveQ8S1tVv9pAie5bkBwcoj2fJEt9siahRoJc8qL
nNA3aCL9JlpnJ9jNxACTtwnDgXgLc9Nw1Vf/i+RRhiBhutb27Rp7ptZSlBKppTAqLSzdJIT9HM4w
v87hlxXshur8VE3iZHwEekb8xbtNWZC68s1Vu9t/ABilAhVQMT2+hY6fVl5FR851Rf9lwM9foST+
VJt4VbPLc5IfxTjaj/2id0RAwPBmyBR++JMBFk3+ybwqsXWoYxHbMsP7gZJXU91bqH6Z7tTpb2Q0
/IbGrr//mI9nGs53RsIpRdpRZKX4WnZ6+fX+iApMpoJfgsHKYz9OVnqZUONc4Vev/JPvrSFiw4wZ
HDbF+7Ht6R1MbFn3at2f+Tsqxa/yEIN/bpc7THCpPWRXrhUvhZLtrc6HO63029WkX8EJTxnp+9Ot
Me3/D64I64RqNbjNm2FyRlddcjadwyU5d7bLh+jLEh19nRbkCY0wsY9KykTYdyG47QXC1pTu7IHO
5hCfz3J3ODj8cW8UVt36rxOur+/ppSX8Xr372xzwrePlIZw/K3IzIl/Y6kwL9TOKS+ZE0ZO/NHVP
IcaphkzCAxeK0L+XW2cfej6T4gy+rPus4E6calLChFL7+6067JAtUf6B+1QBmKiQmOeTQbm96dZ3
DV1QXVywDzCthfH3i7TQp9mvZAbIoloI7N+s1M/E4spLD0ypIgqjTtJyUFL32MOogUTKQOfK/mMr
72Vb5g/57nP3n+2EVLhtd0M8IZiOBhrEVNN6l94Au+INxAGWvYAzdivDRasId/T5KJYn7UyMbw8h
W9G0s8m9/93UhKi0Sh0Lt41V7ATerql+yniTWxiGX8XVHPQolx5w6mqzKlS6hTNBHCmKqCMAAX1v
Hd+7jZ1Z9T1VjQJ/3ch6IvuwYJHLy7yiGUKuXoXUJv60EB//F09UgozgD8Knl4jDc0Iha3t0e8tT
AIFIMHD/NsUlwoFk0SyAea/mYuXAiHMctzzZpYXjUEPuox602wC/lap+k+4U6h5N0CYaVHBd1dOo
F95k5DCrQRP3ulhocbXaWIet/Z2lv5BexsNhk50D5iSDmiJnggXonbvbxQ0rCBmYuRyt1TtJ65nA
9PvFBn4iC6ekdJKxU/NF4mUXI6K8nKpATqAkyiQiMnqcf+Ig9plHSk30qmAeLH6nu5G7r3kmMA2B
cd6oqQQtWKvQPcJUwYF0FIKa/9CXQ9GbwsIf8sx9M3rWnuBxd0uJHsFnI/EuSrrmWtHZpTpbFkK+
t5CiXXicDBdyOzOTKC45Wb1AXnTUxzNRjMSXbgwZ23vhk+0GXKoEizNgTDUdlclSGLy1Gf1X69gp
mlL+jgXcyUuTSNdh+5KpdDQHcKv8NQwt1C5wC5hZouuwdy/wM3P3hZsIQWqPp1N9/JQ1XpO0JqPL
aIUE2yoO3V9Swh2Wlfp9vpSmLRcxgvWUGPtz8nEFcvMrZ4GYttDxJnL9tt3EjW5eF23G0k/YC0Tu
ApTkbNn6fkCmmXKs1USmIezLmiHzMIxI8gpsZ6ls8F6gmIhvAZfs/13nX6Frg8kHF/PzlVFaScQF
N131m7Tc4/wawJIpWkHJehT2aXkfhrvYzDFGieq+xAWMnvbvrhJU2qVnTTZT3RB9Rq6VaJrpx4we
iZIQ4jC3ti1LxrNf9J1EySSk5EtB82r64gtCEh98fjbqVkb0Ns9+zaRP0H02HQCJhDc/1w8IsGYY
3w1D1ATmiyA6jCmbx4kk1sPq2KWb0mW4I5CwgzisYo+XoW/cCkS5UOtRFtwElNDC7diMJuGZjGb6
WpUVSQPxM/CfUInBtG+Mha/ClUeNCsqYnYo7KTu6Ie/G8zR/YcJq7dblN/CcKlvecdKCGnhgNA5+
SW7N7tenTZ1RWkTuhcBIshX4/VwNdujY+vbSwn5kPbbLTLSRj0SvtmLzhr8/QyVRYicx7GcypBSa
7JlSDSOp6Sa8oHo5DhXGiGwARCi22hqW4cx4oymGWlELs7cGEENyUhfw/86A27R3qfxrVr1s5I6s
R8k5hgni9um+M+DahMUtHEUYoNu5scmosqmC2+UQJQa+xT5+Dsi33W54ZE/XsoQiQE7whEdEnjKo
lukqhZ/x2cDUm8KND60ibAQIvO8411mmAU7IHoapk94cs3LFdoixnoi6LAKNzrOrsC2IZbvaYpHg
E6b1JcqAwtCot9ydR2x2bBLaquDvQo86dSJNrtlvidYbMSEe8t8H8OLsM7av4FrKYm3sU8h6VGYC
06dG3au4cKQU6JplvsD1ay4NcMbTgtb5rB3Asl7pB/3pgqmoPA8MYwl9TiWIZGf+kS/MtUkYcpef
6Zk5rn1dWtfzz1U56B6wnPQXsMpuub7sdRCs3vC/HX+G2m0jANNdVE8nxoa0PFxRLPhhRS5xILFC
nMStLtmX5I192J7z6Vv6XcYuGu9CKDRj0bNzmf8hhpccnsfntlISpaVz8/BCR7TFp5T2yvkaMK6F
RqdEgt10L0RFQyLKftlvM9KvxgoscbktptYEmLK10h7ZUDeFumqkUIYRvrxAxm4W9HRuXYOtiSt1
WnANT8eRVEtK3BIT+6HK6EvWWM1Wml7SGllSCv2XG9W+DBWAJ+Pds7xw7isZgraYQTEmVoD55Eqs
Lfp8C/66Wy3s4Xl3RJl3R0f198Jyi06u/NkXjoG+1zeaxry/twp+36kDaqid1Dd72tCaTLUQQQCc
y9X7BZt1Eg2G3tHY0MHPOjyJ7WluLTolBPHIf8HKIvuj/OgBb6StNrx5EztNKFh5zXqvkS2rSpL5
hK/VjZZHi6ssxZ1QWmsX+OffKVcupl80r3fcRCnliG97cmgaMNtm5bWzrKtKUv+mEgDbQmMQX4hp
cc5n4wtJV9zL1hIdtOH0JNBX+yqWninqSu5xW+9VanAJNT/OXf5NNoca8+tVWildMV/32I13ha4f
nthunggReuPxgJiAuIZP7YGAjpgsZ8s3ey1GMYUd+Htw/cv3ea/JO+JOshwg+6nCcsEHUpvcD773
9J0DupJAwuYpZMldg4kCFI+/9NKqIZWcB0+abs1n7+MONmhyqztH0BJvR0Auc1A/xZoLVcUo+A53
/V8kjrvRK9CT5Xa3eu4b/QgBpUlc22N2LdV0kvjP9XvuoUpJzp7I/5EOwEcf07Q+PuCXGPAuuqt4
Ekza0/aYN9Jdle0INX4o/lI0XLEyeh8X/tfCHxtPhGSaGrvaCjz1+Xp0pmMcn0rs+RHVaOxqRghn
qG3zpEUCQ+/skpvgYNphycs++jIEBYkmJzxVLk6B1oVQHEc/ZF3SPbNbDUlvnxOw8nb3QkCKiyWm
4vSw8K2dVqRkeZ3h59nhiuTf9UiScr891jlIoNWM4J9KmeBEaAJR5iCtgEK6nKmYdw3uugL9wbzZ
ngAVAmqItTFurn7ma9qsf6NCNAYhPa6dK48jZNj86l2Xe6RnR4VzrKEeR4XZEjunKLqGk7ktES5L
C7oAvEojrCdwbTaJiPoxJ22pSahhgwCETNxe3ZuPWzMKenOZxoYFoqclp5kKhOx1oXJq4EOzqiLh
nxXBRkmyqs4RU773Opq+yJeW0m2H5fk0Oh2bvyZ2bGo4JJMRCkeULh+3sT93nrmjW843gepD+Hqv
ZQNKPha7fE88T7zrVf11igj7h02SAmiJa5S8WDntNThAfrdEG4HlVN/QxOT1gy8r29Mm9X5287b0
U6m/SmIJh22XipO4W+07y/OHY5xOSPLWLAB6N11UmNK1Hogfk15Zj5d5rV9TfVCPvlIQljb7gm/1
aReES5fjVgaYSisvSBt9FFq+fmyNG0r+zSNMnMVSXA6ZDOkdm9sBbQEZ/6iZLSAsFBdAjhGkxhp5
ghiPmdcJYgBxMn8STEfzTF291j0lXLQdaH+S08PVB8VOfFZoPOPeUzmF9XkkmtGAzI40iKpjm9Sg
C2nPvPWbc2v2hEr6jJSlaXO0RRUq18mnl86DBA/W36xVWm8aA8wXVcF4NRlvBFPnTbHUtL8vZmt6
SUadZjvenBg8qCVrTYdQgr/g1m9yLzodhtyzZP257WXUZx7uvLBkWfyJ4X8gD4beXrnw/uvj7YTd
XekT9+8GZJrscElftM3YKuZSGW5/N6OTm+TR+3/CfHJUtgkFKyA2WiH2OZpR3Cm6Xlhzj5f96WyN
rYwOd4AjNAIqr8WB1B2wUPIJgfwRDUuNUefjqzW7RrvzEl0FywirqPkFzxo2JdHe22VIPADSacDM
7MeVHkbUHopzV8rA25VJ8T7qH548NCQ89FddklzXjULpME6kAO3OmchYTamAZv+zwehlRb5uFx9B
DEQRXnK1J3IfJCKMc5iPkQ0yGK6utXJucajRXHEmNVS6BS1yoHB2hvOBPoMZ6ccsx5EchJ6+F5tD
kCgNAgm7/Xb+fQOkz77giMSrLTpBsBLv+XibzqCuVOI78LriPSodKdJSASItstEghk5DjgGQGLCK
hfHM1zig6ASXY4+y7fmKEw/zNnnT2fvwJa35AQBdbFYksylTcvyGrAv/5qMzDC2MNLH9ddAjHd8a
cY3Abj+q3RazUxLaENnlTWIHOXAAFupDteVc/Ox3cZvw1JRvRYMEb0vWGmtVVYD7h7xvQCFgD14R
o8c8QxVlBR9wnPj7PkZOi6+hPQ63ij9ok4p4n6wAxByrsamtyPeaqb5ukKKW2FnWAoLQPRFmqeEQ
NnBgLl/0CnI7tTxEP/JBDrDOPhGSu+GVGQb1m826PSON+UmD6KusAq6w2C59utv7oempcIAupsX+
MMf8ovBsgsY+AGrtC3UH20h8cm47/D94bvZDJFqxmDqx4NwSpsWkKSE9wgOSASK8PgheLJAWJev5
kaCIh4FsW66971Ia3S9yTEkMmDsr2zkJidzv1WruurcFT9KRqpQMtshVPARFzoQg9aJI2Aj4g6Wz
b5mqu/KXIjY9UhY27zzOlTP2KI+wbxyG6cmubz6p+3Ik2GtXmrsZQDApNqRQtVfiuoHpa4ng8jZe
fmfCniWPFGEWkVJDYkangyFvhanqhuXUqyhLph7AooRjXtPJTKV8X/o8ALQzQEVArzoF2silGRV6
fIpMe1to23/NXY73Ce/DyQUn6uqSqZFaM7XCUYTYfc+NfU0JC/ChFegtwyZZmrYNCA30QrJpixs+
nRQvykrhcfVHhAgPj4+TGEqI0pNAs8t0qrhR0pi2KztohQq8+0/xu9VGmsMhz2vvXKU+28k77att
jNI98ttR95i5vjuPRMDFF6YphZianO4UQZ0/wE642B7Ed2Gzmw+0uK5bdH/wlFqwgZ70tAjcPB3T
JftDzXvZlpEPGLwm3pAl4NkCcMo1zTg0WetvXLNooGOgMOQjhWtFY9wpjJRjisDWyWmVQ0siLeGB
DoQ1BKw4qCPUt/FLdqV3dHK1XKzSTfF4nRemIw5JqPisjql8S2wcAkwZWs9NJuG4twbJpNkPdh1R
kIPV6Ovy0ByG+3oaHuYl6BD3jdgJLO3ydSkN1bDe4bqVnzYGkW1CQ0HYW2UtJ+oNbiXSHQ0+e9U5
vguqUs53nT1ac5uk6OF2LXWPK/NVRZ7pQIQhBQsaeRu4K29n6elMCaWMc0cY5r/MZi5H+4vxI0+j
IeLFL1dY3Xy27mchAFdW3jRRo9R2abeo6Si2GxcVEAbdX6XqDGOQuG7Gc8QuX4Gog3FshvcTMuGg
kWQiUycyJJF+nkVzlGcyNju3YpBig8YsBrDgZ6iCZXUJmPUBWbAuC1CstyVq/AvfvUL6A1GWZtgK
1At8JMq684NFTO0akbrxcW6JoBTpAzN8s/3OxRMZ5c5jeArNXUn+uwnZ2h0DtUJb9INe78OwR7kX
7ud9+3G3iGF9GjOVJFzd9Jt8iiYQeucxJYHZ/K4kV71rbSC63JlCBFsrFVYH7gzhs+YgCU6zXwAT
J/1IYGjXifukL5x4vUth2Ez1lqKfDKVTRzyt0zTMDcT8kxpEFhraN4hXobuWojpm3gDnR5+aEeEE
l3z5yF3MBBhawqquln4Q/YLBQCrLEeO3DClwyIMW79F8msnnQSZNUWS5oH9PcVDQ/t5j8tfx69Qj
sCKWG3iCD/kN+7yVQX6L63aBTOxZv9yfcYe4eMLMANS013IKN5wtE05agK7qBcZ7QdwPTeOStM+u
9KEBZrP+z1XUaB7jbo337t1Uir45R/hACiG4IXIwjcblsxXpXLMPn1T9EwSgCFNu/APso+MNxJSF
Nvawknkewrwts9IYqcqHVSIYV4eQ+3wFylt3gKshEqP2GvLfQiOv60zSsuJ0C6mwBC08gqm+q0hJ
1pwRq+lUHKRAlJlRE1d/1X2E34g01ZQ9GaW+hR3dcjnkqBqPyKWfbqYNAcr6vO4sToZ0UMsi7Nq/
Cordqf2ZJDNKLGDwl3xvrZecVQZvd2pqg55iYV0JyVlJNMhW8yHvyi6/8q13b7Y64r0dJE1ZHWJp
Jve/Iblv7IqP3W0z7SzbUHhjd24ro2IcskM7669w8lcPoHJP4HBItHCBtaWfHfLsMEU59X2wgQTE
KjaCC4OA9HqgEHhvzqXVb88GqTluUntIq9L9uKHHVt4RV7b3J197wZv74OuBxjJWjttwT4WnONOC
eKpG5Do7GIBUpRioCXg+RfnfXLynd25MJqvUowF2jKCW6K9qXpX8WjwLKC+V58WlOylonA/mZvEb
N85p6zQ5xszMD73rJccMhW7YnA75HBbLUIQNl/beHpHSC+VeZHjOJ6lh+PZmOow8OXhdZdYnbWgb
wxXvUEsR2HZ6aOX74xqgjyaVwbVLWYzuEdhVMcmNNPjZ3B1EEhW7FjG6KUMl826UgGZBQWuB7s7F
hpTzOar9jT+uaZErohEctxv+Gxnmvqm/OBHhBbyY2GJDhi8s4ICEGeyvie1dnzvwr5+yayeCq5jY
qqn8f9V7qDc/xTsmqlQ+58ByMy75NL29qhCOikmKdlJWTKqSnGqCD60fCHuzt/yoRii3facQEsKI
OjF/SkOIzdleylbzO5jHw4KiI2LFG1gW5HWmltQrWnTuor882H85JCxyqYlPmKGVx9a46MDabvzQ
pY81Gr1/x3cNQVdDM3xb1m/0XihpgiVU6fT8/EZT9+pTzmbk9wrcX6fMBjgsyvzb1AzpaFiOIfM3
Je+vmR7ulYDo/9SCOxLHj7eCHv52miW8xERUiOJoBTPadXVWch8fjwVdu+IeNGFGsqMA77jhIq89
yDSlvQErX6xrZmeMFx6uWCliV7KR4i/wqMWE/g7MDehLJ+xjuAO23LPn//z0hyHPRZ6iqI7mD7C3
uZospAHw5xjaIFJnS/rFhsciCA6nCycAmnrknpD3QLe/UOVFh2BEuQCp5HTfbbphnmlPLCDapvIv
BiZ0NgIKpraN+H4db5DQhOylG4bWjoKCW5few2lAqqE7TsYaxMP7EGCyPnbMoBxX23jWdi9C0zWc
dVoEtUdu4gAi/Npq35SpR20IH7ZjSZARQqOX/dSR/sW1geSUhBxv76c91cbMyS9+tdIFLY6jSB/b
N+SDq8muU2zkSOy2ygWxDb6XvOkQzNyO8t3mPBaxWrk4eZHDuSYL/J/hozmQbB/18ra7FzK3YPoX
LOZ5bH/c5+0E/sPX/QH7nBF7ry0zcR4AJcbqDW1mxn779/NXCeUpa0y1XdjH94R7DFxJ1udunX2+
LqY95Whyrreo61F9vij3ktdJwxxEAQQBSGv399qrCRniCHRf7l2c3uUSM5wdfNR6YcuGVS93uLKE
Q3/d2ITRPFzmk03EPt5O7khlYib9nViuoa/r2jRPWZlHya6drrwydU0sZVYEVIv/dmoPRG+S9Wk9
84Mm6PSQmf4xFiOJpTk8IL9tNG84MfXJyKVuN4sOUTVjDK/CcbfgnTqkG51rOw3L9kC0BO2t4Hpq
0EYiUziZ6A9DZxfQvB5cf0SnpX9x225DVMZJKGU6XVihvfLxlSqX8E19kLNPIkC4wDgZSTdw0HNo
YFrXULBqyVhqEuFJj2NdUxQvv6NIFbs32d7yetJJAKlDznDhVuIyMqQhF4DRJtHDtbnMsM0qFWQJ
PSF9bNFFAupWZ2PJ+Io3unk5S06KIE3GLekTl5Y8tgiDfvf9AlcQJGOesdd1zoW2Y4Nz0cM90o5B
4XBhwIURN5XtsXhMO1kDVEQ+bUH4jBn6YQlGUbCiV4Z842sLu8zKTT0x1o6mOyOW8RO0NOOLKxVO
TmqE3ekbh+ky8thMKLEHTZo4Rmku7HUbMzgJeqaz8mkTTvTS8PbSKeqbnKVreeqY0de2kUVthV08
zMqHCq3ZYPExyf2v8pqeeHGU+WNKw8+n9YhKYcMOua2Eo7XK8K9vOcOneb3tpS+F6nEuO6eUHjXr
W0f+mQsu9SR70BJ/dis6BaPFiuZVN1dowS64OQLzyj6FI3GqlSBsHyFxmWFu02DJurqmcqkSxQUo
8mzRfViv7TKzm0beWrCrJGVfxW3lff8L34WrEYOdDOoMPC58LCDDJ5X0x3znnrsKN4lksVyEjLCd
tabxL8vS2g+dPmnWbdCiVrqCYRLGX6o3FKIPnbPP1fY0ZDc0/Dj1fJU4eR/pkP6paHCNsv/d+r91
+vaSpk1UaT8LJjatT4Ir9xGfG+7cV+tIQlMVa/CvhH3f5n+jUIadoIzWYCEFa7ycWpfICXEdxb2k
bKik31rGtO4cPWQ3D8K6EIErXKLmMgT4Ybsha9M2MuJachCvLaqjPSs43EXtT/r4vCTk/QZtWIPn
dGT6x/9EQtuUhN9aQ5QvX3rcCzcnaqG8P8DIgvLZx+M1E5xky/5sg1mTc7/T1pDPYJ61bPNfTXd/
wvAkx8CYLTPblxFcOYgrA27JyJoBJxEqNFMjYnlU0oSlChfjZlOYZhjp9/3fQt8AxNkhs/9sNAMw
aCbvRhpQokzWiCcHbDBbQNPWq5uhI6pLSkIURg0MWf8Ej4OnNEXM+czPF84zI7M9eE2juHgD5p5F
TEwA+vgsKIoqA5TMnxO+RLR9pGcFpknksbVksPLoFqgnsYVbCwqOGURVewPM65MueWOCdKQSiYnD
ikj6Sxgcj54LzNpOM9SclYX5sQQt3acIcP4jsjBTVYIfZmEDZQ3Cy8K5kPKLblY9qnUMQpkdJA66
zRiAsRvIUZ4FJaD58LOYfFZRJfTxlQOq/3pWc2LHkKMeV0Ttgvv3dBbYIYdXJPxj46f/3+MwWWLI
1wSpduKNuTojWAYXTpPKNb1wqKQllWYyI/P6iPU0RoH3JdUzx689Wju7A1t9SoabyZVLR3UDMRTG
PBgUaOms10Z4/HFoJYMeif9yOl6zNlupfRitDYp4I7TIeFiGUzWKFm0nySRgaK4P7IFitpGVEROw
A97bAdtPpDart3dOD46BNI22li2RtkZFlKKXiAgrdb5O3vh57D84RH1xtd7iEEWbqXQ5QQD2hzAL
vnFK98ZM/D096JX/RS0z3YVKrbxGWclX48Zw58mmT8g5xT4ZQv8seSeRkyTzWD1BzRH5729HfYzj
pKWpD0NBBMmCw11+SHcsAmN2//jX6sDjjXz+4WNJOPC82647txV2LnGQEs809I2HVExRMvoczPHk
ZjnaYzEK0fbA7VQPVgmwQtUDD0PfCbHN0MRU0AE9Z1fHWgeJnb50ALYB3W0jGzzBnThK0WIaw4+7
H71RfBYJDMT/gaVAvVE0PqQnSwLMeTBrpJrtb+HPsP+twPLY9EuSOyCIf3gfMW3eKBIt8gKf6hft
yBPq1yILF+VLmrfjme0ndz4NePS/Q7IoY4k8OnpFqdIctAczqSTnNIST9RglBiQ9TB92xXrNl5B8
RY9W6rto4GdN8nw/FqvITbC0wIgfP4q2hzEK8b4YKDHM93e2srv2JQ511ShLQqkger/Tl4BLUswz
gpT36p9LMdCzc8QOoWK1EtrkQeCIsuSkggBFfPtu0p3ajiHQ+2L/t6UkoUvuvMF2NPC444bRHt1P
d05JUeYW0CUKYsB89VXS1ZndFwEUQK4POhtQBi+NgILimXZ1RKvK/8b+J5MmgLh4bzPORzHbI2BN
nmWwMYLKo5iZ8VHhkAVTMBYMh6/mh4ChjoChCvzkTRminTv//+4w2JjfOZohzjtW5T5fqR97FSCZ
XDM1sXV1b7Pi2Dvb4+AiZMhekn35e9Z9NaFcGVWTsUBb/iffzhsamCJtcUpbnGqoexHeZYA2cHj4
hJHRilaHYEs6F0kx47MYJlfG9CTCDhLZBXE0DFFZm6Tb03XaZ7tJZVzgFPtOgtxz4pOWa+Mu8NT8
8dhgYYrcpOW3hVt8PFmPQtbfzWRBUuE9geTRxs1EKEbaIqYYaJ2vgN0JbCaPTgDYXpuuz1G2BBiM
PBW2To8Y4/5yh5nrqsURXIigongyHKM9QoJsEWe08n/7IHSxtnj2Y3ErvQJexLwZplOkd3iZv2QL
BpEvKOwUMqdVfZvWNIAaZnXxCdpNGIxhzH+P/4YTNSyvuussgHVpLMdxzGnugXor9OdIP7CseUEu
HMB+auw8cMRXu7vNLREBhZts/pb8fsIXuW+G2t0ggK/W0+7BXJLhEEm5wDFNM2AYugtkuO96s2/O
iBg5ivHtBrU4KA3lRYrW2qKoDgIptD07LhDS4RkwJcD9yv8RQpgm5iG/75OtZUFqjIIajseMmz2r
XL8vP49sTarcngclUwB8yy0GKUjgQIH/qz6iwY0e9LhiBbx3SIubN7CF9pJojBvZM0Er6+adSdh8
lIy6kWHL7Gt4/dX9iDoziPvvXXVYpTA8+jq7b8JCzmQFSsWNwwrLrBzWALwblKsiViB50Osi+yA4
t6i1U/S2G1d4/H4ZxVw8eeXZ9VnCQbGyJG8aE10dD3TwTyh5/hIqB+PuafMSTcmGwTKw82t16FOr
6llBjNhtW4ytoeY+5F/R5gKvlTfvWmURuSdr68ZEZzBx41fWYmHajFPTN/qIU+2G6zO6E4AKHBMU
7Mh2/J75nV0LMJ6m8DjctoNL3ZYRfMi23iAbqtkuXT1sK/LykmaiXJPtjMM+92WaBc7n3b38UB7j
2VkLrISLnI23Gzh2fUjJI1UY+W94lqdzZzbcGRUsbad76BH7bKcPArsRbp5EUh57XAJ5X289MtpE
I3gbpvzWqdA8vPEqhJJrtkSzOXpAWOgMkiY4qLP4J0TmVYvgbbROEM08FUrtvU92Xv+CfcdZoiSR
/+ZlWCxfwMn4/xCjWc8sN11gPgnz5CP5/WuJgcPkAT+YYxdK+UGPa1Za1nXJTIvaUGWd2JmBxmLw
azMGv4CwzYk5J7i6jGVKOtYsx0zmAQ+lsKUce3ncJLigp+5P6h+HDSwcUDSTDSgdbh0sLfOhOT6T
tvLXb95WrFiDODflJVnu6v6qLsjSlgUQY5bVvBnc95Ik1+22idDxxpcUWA4m69YJsi7uNzVzkQIX
pQUFM1hpcOQFuuOvzU6mpwBW/QD/aMc7LuZjeyQBlanUBMAxVfeiWLBf2YfdaCKuvM63YO4QFoDC
pxBqgwBoVUGrr4eGGZN48i0qsShysRyWFLLpJbKqv47SgTbcPYxmaCCsoNdI3Vqi+CRSPaz50/wm
43mo9Vca6CWLGwCDNxWbSeYESAoObMflE6Tf63sjywz6Lc/42Qna/XSv1XANRXE34vGahFlDyVv9
bu/4eKbcizn7TfClE/qpD9C9eXou/F3O4Hpw/jR/9mo6koa2VOzD+ItRtOuG4R7STh9gA5dP04Wm
ZH9JpYEvNysX3FgteA0/UlNKoUAvoSsmJ/RPMo0cSxVC6FoDrSl2xCMPJEvH+RM+DpHExPaGXCFe
Be6JnbZ+0Jpa91duNk8eW5mW23CWVQF8CTt7xqLDKv1UJotOjQs2Ar/m58CnXz4PkuCaQVBESIki
mNyGfa2Sp6GisP4GiALZTDYOJbmJQ18aufUMOgRv5HWnx7fojEHcMFy8ceM8+wpij7d+fVtLjmZ+
3DgPL+HWi4wauNRKVPY0Oi02mJ8gksIMtNw+eQh+KharHWdR5yUtMl21UdOYcY/8a1Hm9cQeZqQi
i/3AIh5/Qf4oikTU8QrprEkiKma7LfiKHcHzjQXIutDGJo6VS9regpn1heUIDZx+NY9zuRo9V/uB
DnLPqTiyMLq3Si7eywseNaQg5usiBvviXrcaMvHlQCIovBadi4BQb+Vbp6/jr+JvsUzNNpwVcCiX
6O5ooVbpNtmBLfXcWeKDoV6gMlWG6gRU6+OIttKR6V9XVTM+D9Mdua3kDWWdaDtlwCZZcgkq6C5E
3HMPxhHYbwJafNQaehTUzRkEUbn22TSlxPvPeRyTfqx2bvALj2RvXcPk4o4zfmg36IacY+t8rZxw
PAoHKOhEmK3kniP8HPqt2Tspx2rtV3qSDrLxF0LS6MK6jBqscstmjKeWyzW85Fs/mR5wS/BApk4n
Hc34k3skdAx9veY4ffFAMuWihHB6bxxopScHuU1QsZgSDeY39xO+pS4oZtoeJHMKs5Q9i3r7EtRp
/OgHxOIPL7eHBH51RAQeefOfLEB0JBXqCOj0QsNZOQ0Uw2TR55rORygz8haResCowFDCGMiMXa7a
eIVzj3l713RGhZu8M+ZGeuKhxkGdaLFWTlyL9YCqOxPoX9gkEcdB9BQI54v4kK/TELHngcZWLeNL
0gqWMvBf6gvy8VKX1mX/nw/IXiQBtZ5UJ4E+6msYkqdmJ3wPIBeRLreBinG0gegk2vA9XbO9zjDP
0jbkYIVVytKkXzG0lpqLdGM9RPQz9Ru0myQWnYfXQfodMQMGSnYWK12fPLaYeC/1Ydu8mspKcv8D
QbLRZ1z0+KBB1BPr2EtVNipKOyKBYmG8aNBZrvjASqWLu8TyPBvUpqnhodPC73V77f8qpZr2W9RO
0qYflYnGE3wBROjWGBTuTpIiZKRrD3rUMIO+plITZWCZ2o4f611wTZnpxyhKf+72Teolq55WNbvM
HXJvHopK6L4ZdRC9Rd+G0P6GOmXpq8eZO2Pt49Brj4HHHeSYUaO1iLNe4zXYfmIN+nIfEaF+fTl7
dZC8ovaNKFMlvQ10DQX4wmUGp69saie4Nbd9UXFAwryN1elOr5L8E/zAigl7Zx76WrCe+uVlAUnA
3Od4GOw10xmdxa5yuRwmwJ0DzKFJS0yyAM+ijS4+94pxQ0ffUpNO22nvmGaMT3b49NvTmz6YOk4e
O1ancmxEmoca3hIQkrluwl/EFjphNEbrhQkkyJtSYFL6yDuqnV05VNnqBiYB1svZj8ox1AATfEsU
E/6B0/SCszWNLs+/EbrwcZ/QuWnDMdGIpwaqgESY7BIc58Suj/GuInJJMbILDnmlWaVsCF9GnlHI
HzQfi5FkL5bTCq+BBV/r2kL8zproAUUUy3J9fMwVO2sDM5nrto7YPySsdZdWWoRAxkhRX6PWta4T
GixICch/JMcyCzWLiwKM0zxCvmcdXKHFqLxpcaq4N4TzbT9JjyKrxZusvjQyF5E41JoH650qnBLq
DPaykUVNqDkPT+5/zDO1SBDHUaGU48gB7WNOa4Ro57AELrGeU+xNnkOoaHyBV7MLwN3UTg8MNbX8
oGlb8HMvOpuRU1MQvNZq5WLRIap4/R+fR7GlwStFkK44Qp7xD7D/Ki6FmUlHftch/Vk9hIBqSzRI
ZA1Wka+qB1ODS4uE8yNK/KkQM5N3JQr+M8D0KhM41Pjil5HpaMJNVpPw4r3YkTWGKWhGih43/XLx
ESgoOCkRPdTNA204zTWoQZYYkQhbqMoN4Z/v6bkk+1QDyFoYMb2Su0PoMv5HH7wDdpLzK4l0nQfA
X9p2ZJ+6x46emww1FbAvJutWKeslZiIOTiDC2hQxxd+XUWCgbMqr7eMlZ5JgG2ydITzApageLjUz
DoU7cxjECj/1E1xvqjbdhkZWPiYZJbIiW108CCobTirkU1TOXuShQm0j/PUbEWnjf6uCodGLxz6r
AKUh+b6eaicHBYn5KLyQuspukgKNMvC1dPVcp05XxZfubIbKaTJljbCcKd9KUi08rOslZlVgYkIT
0McPPBHONZKC5EC+Eh678uBpzH9+HG63Clysq9YlnDYbyDsqz3aWBPxGYmOCY1W4lIrGvgLWZvfw
y8h2f4ar1wzq7JKDSgIHR1UTmpG506azmU1+pdjVXhztv4xwduwnmKsEzB4M9K7jxIhC/kxNO3YX
Kh3CSljtny4ovYjXxJ35YUbM6+GrYk69TI8wqCHKrA0bVfPm7uWbJqTBswi4TuAgOGfK7YMbuZYt
duTrmtycR05w06snLqZaZ1dySHXVJO2baJx1GYJs0nnlw1aAioPBt2cylz6MG0HibixdgIgInq/p
TWFMYgEmx5dmMiHCWyuyNDryxuvTyetau9OPbvPO2r3n4Ng7GICOSdXpW6kqx9xZjDhP/YmpCWxu
SqvnFnuGQBrXQb9InIIwLTQWV3jPwbikXQqqRGSmnBu3/g0RUu4qAAWm573rW9Mq+dJ6NI8Q7kec
ELNDGGR2mobEtrMYzv3gXfQVNG7A48VRB8gosCoNBYT/2KwT3e7y42MMh8eH56U7PrhTU+pcGJg2
UielpeCaqMdW6JFH4wo5YiJzB7Ml2bJ690GiW7701AzBRnFjd4MeuvKOu+GJau5uJdOUJXTi71S4
YD9Mu3jGJ4mjtuX06C76iFbYnI0yPm65tkV6WXr946vx9LfLpKbPwGnKbTtjXeJfJ4qAIDKbopqB
qFZ31Iru0rFgeUIJY6rIQYJgn2cIyb5IXsLFToAMl7OqmMXtw5lmRSchs0J3Y2ru2hKpj30m+HFe
+ndlSq9sBuA5X0Qpbgkf+NGP2K3qVkIS6Rvc8cZ7z03oGMv2Um6+smlNiSL0+c2q5rv8QXS9X+MF
A+U/eOFvdEV2XD6oCrcWaklQHBjE3XZ2/NTiXat3c0mPalNQJcW5OG7f7xT3dgL3tUaQhRjQSyeb
OCXvmhzDYvLJCM0z9gQYKKkFGaxpPp83HX0YxygFkzHG2bSYGt09yiH8I5MND5GEwyFo6wUGzTSb
TTSADrsJtjETj/5ZJ1xGoktCB7eD2A/LOXJ+U2V8C1CSdwJqfOnWR9sV0qohQMXvDqbSL/f/XkVn
Bz0uUwX90jfiKuse4DG32D/Hg1sb2hXgkpS0DKaQASd8N4fV/rliHvi9IqgRWQctESZ717CJway6
zjXUmTrL/i8ivsbG0a+V+Az6NrKkjY9FVA+bAI0b88UzPadNz+S73HWCrLQ7Fluw47B86NVcnnNF
WVYjEt1hvhjdvNRWAQYUgBC2I0I+lsnrPyrZRh8ewGqQ6lmC+U8jtarMOVGyapP5xMFqwyBz+SPv
bEp3SqIFpEQcW3e5gel+lexyFc8+HxtSBS8gnJ1rSB9ltYGLHPcOjwdCIUIGoBY65nigC26fSMKQ
bqmOfHA/SAk+JqvStjYGqFerLghqrXH5+61ZOggJJ/kvY+9fTXMbW0hFlhk7vPTVr7ZEIFHHfLJp
ADFl8MnK/Vx8LBRWOeACMIj2KOHRErnpp1M9+Rrz6tfWc8xQN3iCTwRQKubSqGomeEKCLz5ENJIE
UGiK6+OMna6XY1Veodxrp+8/8S/YdES0FQ2OV+PqLC3daN1EIu1Qd2aGhjLtLG6bZoxMIKjxgcl0
puLS6cQPpnAYEDRIFW5mJwg2dkChZhXaLCo19jBvKTSfBrfVs2NbZWd0o9E0jlisUKnK+V7nz5IU
v+80Dl78Nrljp87kKIBW0zUWuoBwmjGujsRc/yo/z3HPW/nXV71v1i3at7SPg82bPTy1c7tyHBYc
lAFdoKrApUfMT8FYFfTA09wOuWh/VrhKgAjCHKhEINJ8YORykMSDG2QiqjphgOuYeKjnV6LJje//
fqE/R+Yi9cLAv0cx29FP1cEXeAZVHMtx7pExmMt2bBKqTNybZlQlplAJuz6ulSzPiSAdTFvte2Le
/pqEjK2JI1e4ZydztxWklNMULnBI1XCIsUNOkjLTXzp8Ba7eqN7s2fppIYw9cQrQ41+MW5s5zscS
F5hfuJL0AZ3Cw1jigt08iVes+rbDR8QyRuCQrEXPC19vPXV54i9a9l/HRzZwz/M0v+FkDE12oh9g
8DmvwzJrPEDJp54wHEr1P3YeYuWrZHHRXyEhS+yURmXT9SyuQJvBxCcPw6PlMj/PtFYevWtDBewR
9zcWDl2hK9H0CIT05U3YIuTYkLXmufRC1BZ4AbefEkUXCZ0mpakQPjXoTIpnTqv5fBHklcNQwRd+
iauEP4JbMJdVjoVlCk5ok2+/Yu0R1h9K+mgSzMLt+NWFIaoydB6yJzbWDUc5oRgEw4vZV/KuBAGN
tCdS2GbX3MF4bKYuX3o8jmpACEjyMyWce48KpXuBpex4bY9CZLyBubHGUrny4+Jn9E/sdhl3GbCt
wtLNYSzZH6X1hPH2LYVilI57XAcW1U0iDI4nIvDirgihkCOb6HwvYrVcfriq15IMNkxfKhMC+NTy
OpXOPgCg5+RSnN1ID7Mauwwo5kHYayMi3xT68lJYQhcMvGYbJYCWtR0Z68UBIb5F8sZ8UCQ7L7VD
AZkrptpN87q2ACCvYowuo+BDGDk+jPROX/PwelqZDJJD6hKPCE6TJaKURxrrno1+vMLCeEffMQZm
GUj9zZI5JR5coKxWtSmWn9HkZGNPhGs6fAttRS+J9K/XedeHLI02K4dswxBP6M58yy28Sc8+y41o
LLoxvRaD+7cQB4pZIFp650mPZRFUbceKsff3kC3DtpcrrsjWFLkfoHjPgwPRdiPjoOb6Z+40LDRW
lIDFmgrRTXZvPhe2YLVwjFD1FuhWiZx5f1JEXjxPQP6EIEO8xzaUydKxAanZ7XRRpL7Pff//aV0A
eQ2Hlgpx/Bg0FcUp/7rHBhYr6Kh2Ndfps5dM5C3sFM7S5vbkT0x6LDBB//T9oywlg+V3s13ErkBI
3Z2TFIfVhPjS31Qjf7tTkQWjmtzsCz+SSNeL3+6NGeJXzKeNkeRwfYPGOR/a+k5Yih110XZ6brms
41WoX82e7Ktpe4/8P55CJwaBhkpUSx3px3ruhoIU99Yq7AMJJ2EV0ea7FlC7n64iMfHrRHDqMpUl
BtEd8dwBUtKUVMyMCeGyAZcokuBqteYeAY9CHL1fx2ny27wYz/+ebegKOrIQAuSdv5Z8uJf/3a2t
n/fvBKag/O9us13nJTSGtzOBcuyjiTYjzBqH0qi0Ol/lYqjEAlqLKi75IL7PXkvyc7xl4V9LHSpd
X8FWyvvFvwVL/Xby9zHeNi+sSMy/k2Cljg90+G5OnKZb096+1f+CFWn2iKkejPJX2clie3KzCQUH
vyIA5++5PFc6pNcy0YkJmt0Eqd9Q/I3jTa/zAb3kY9zeD5/olvvd3mGBuWRS0S1NsqH7CYc/8QVV
MCYcidmE1KZ8RwH+1ywfB724RyZtYNOXn/vaea5Pnvkle1Glz57a2Hu6QxjBlwHpRjkQ9oJv3P11
yPYUfb9rFiguz5VBed0vNDk4lbTVsP44u4xDeXBnTfIUg8OvgK/s0H17smHW7jskvdchZkX3G3tr
PInUDKpp10BH9W34E16UCqGMypQwk2b4lsHHnMyY16HgYrSRWEpwxKBLh+rVR5tbTspPqVJXrdCF
MTM+XEvO4fIydFyK1HjZDw7xnuY1+JQ63h2yG8RX7QC8U+AGp5i9BIY/bhNyIXuhtlvGyoux5lLv
3aZnydU+XrBtkmc9oWosuj0DgdYEUjcueY7aR5chXJvTc8eT+ZCx/bHB3wRQtYrPYpwJDVmvCgPy
jfdD7GeM+/BBuKaz8wYjfpXR/S9EuY9LJjIrbYGPB5BpndxxX0grY2MEJ4XrJ4GmswZlEpC6zMpO
mdoOe2vyJqijcoZ9DJRpXsYitIxTzCNnf7CW37jNflDGtogFf/3ZKDFr/QyrIXN5ZGGFkf0GC5vh
KVv9/HbybEopiTLAq+3NcYuHKp4qr1wHsRy2i6E7acUA1lIzAm8MC44WCE5VyeoWUxNpAiloPZ0Q
9RkP2s5EEuqV4PNHD8L326TUh5YL1bMLGzdCaJ9MTwHRCmRGKtmS9OgT/oM8CCKObwVD6EPpyAB8
Q3KxxeHxB2YQZRLxaDNiDu2QVa5s7DsanViQQxo9sNhrG1xLtgNsnV8k5YYBxO4HNjTYgV5LYxqD
Ug9YZoET3dIzqeH4aFq86ooO3ALxPfxfkIs2ntdhbkZhqahfizj6GSIKa6eGy4g0mLmQMNLZ6eGD
jNICLCG8/pemJoOPu6uG3LR1sEpNtjImcfGRtkUG5+RCXR5cf0RNED49Uav8k6BizMq4lm/TGDEq
B39+U0nAD5gFBnOhCGI2NCmG0YZEurtuT86zD59EgyeHG9Xrx3y3ifkll3D2xGq32cp27KFGdxY7
PTvrqkdQepM2jnFqzBkyivWJFfQ08mBkrItIQWrZRI5yQ/1T519j53ETMSX+YoFBUjffh8qNckg9
8V/HCqDDt8P6qJR/yUobktZQJ2Y0L5Ce3ZOO+cQPv0c4s/zBz8YARDhZCmRlSl+8WofmTAX3gEdP
2shh2LQ9+qum0fPvyT/EN0WOUkCOF7VIcuqFBfPrJ7k7wZpcXZRAQa+vPFkIp2PSEaHKJiVxyk7P
pKX/KEXgytIjxprsa6QMauJsJRr7A2CG4QwcHDczseWbx4LQULfeYyxE1gWnEptIXz9dd3u+795U
vKbXDzDgY41nW6UC+JQ5R61CelcT6xixx+wEJ6haHgxTqwdD41JUYYQvTyj9yq1Lu+uIpDBvZToN
2615g+aox0s1f4STfCzHsAmOQeyLqwukIGjm359LSsBmvP/4r2sDtQ5R0YGS8LKXk3qoTT6AWhK7
fRiO8q7VxJiKEEir+0nFFI4AtnD2kNrZ7Hqb7i3t55Vi9Tn/MqjZMRucO1QTKr1Sn5z7sFX83BMa
UpuEUq/6ScrihTf6ecWrv/MEWK1F5/ww0BEPFxJUpbsII4JZAVmvrvaI5aKQQeIzJFN+OB4rA9wP
JtiLnnYxVYcFSjgHMY28k1ZBD6Cw8TJioP3C2n4u36g2OnMx2i5lfQevrE1EDubzmlILcHTPBzhS
2od50WgqNc+XmhQS5E/WdI+6gZuo7HOWmXG2IFn4Cl+NYAcRZFjDfVWf2hP6pu4LHmfgV323G4/y
+W4cJ8/W0pbTMRRIlMOAADgYCKsJuDOLmghWR3Xkl30xTdyGNgSCP7EWW0ECaiJx6+1PrvxTrTUG
T9cFs6vv/x/KEUn8sPBqxODZGdsuzyKlzLY0Gk1vDmYFe3B6c8X16D0HlLtVFNimh2rKSiwYOEn8
8OxfpHyu1uqB3QKkRGTWJ2i4Cge7WTFyNcVftBvdORRHXePnG8ST1jiDDLsWr+C2pLR2ej+mQcWn
ZeSyQ+zZhdOEYjmhdcCU9QXDGdglOxjbErtDQN5ex/oQ8S5VkuZyHBDAqduNMEPu/J+AL+kSmf2x
MUkYvt9D1rmxx4W8097vgr77n3d65FRF7I3SsamwHIjbTZl3m55teYqa3t5ltQfmv5XvFQPifzhh
Mt4oHWwmcm0SvM2exLxAoqa1IDbq44qZWD1DqahZIUKHbfbZ06Fr1Gr5vFJIF1PPFx3JFlXoGHdk
aVxE6K59v+htmjph3WGVJT3oqpyaKr44KNRIEVsrllusApuNBuNNJql0KL14FBtyjbZ0W8N0E0RI
cBqcB0d/Jks7Byd8Y+BcFRHDhpKHDDekCG7HjfVOPQ2WgJlW4AlfbJREbHiGMOxcMLtjMWJ4Zsz5
9Ayy/Cl4LzAtKB4RwuPaYho31nBBh48HMrrsu+Cm2GqFJuQRwisSPpCYr0AnW2Eo23AdhlGnA6IA
i4E4WvXBjNhpjDQcP1/vcthE8vtV1KbYG3QoRblA7y118WgWZTtAizH2hqxKYZLuu1ERb5IYTffo
6twMoyUVnlLVK3bCiZD7PFn3y4JCVdHCyyprS4wAzep3F8mCbrOHH51JgzVMTrpjBhQKQokcJLKq
9D0N8sM4JO5zlaaY0Uttuan1lkIuG/KJvSCoHwQM0KXRw8Jm3nxf+CgbPV44XuW4x56JBpUhaJRk
n42IgN8OrplBFiEttj0C9tVmWDRsRBOw6mObbeOVi02kpe7mcoysAmR7l965Abax+WPIJKISUZzo
YOV7JThsTAqX/s8bu05/XBF83JMSapxA48HoqA6vWNw6KAfUB8q4twCVWCBOOk5nHAHo2xbyLnIt
Eai/5x8x6EOi4B5HUNmdHgaAapQ/vlrgcNrFUxJYOKtvXk8dvPnvQsHg17i2YaRya5bGh63hC9oG
p3ZJuRVwOQ5KrT2TOObBiYVOpqZTrVGuF5FlwBpERuU18X2zFf+kpsGVhp7WFDh8wAtD3x3Wyqev
M3IA5DsvnXzlSmpYQVjx5CoFa3ijpkyAm0dF2PqXOsVbFtdbuZByF6EtSKhy9CbjbIkytdj2v+CP
4/ougaHbivNOIshm4uOk2C2x7eF9sbcOMmv5XLRjdOaVnStFAGktsU9474aTBhYWqCbsDUt+USBr
WxFth003eBrqLDo1TUtDalM8a422Nt2eWXGidqXN5C9k9/SdIx0sXW3usWhGdks/SPEUDUUTDXIw
Qf6CPnNO4RTD3J+l+P/Q/MgW2/COxoQ634E/RguMVZdkLkiiRNSGg9LdElUzXrao4OiBVLUUUiQ6
GHoCyOJgBQ5r9LnTGIWvwmaNXWlkAiD6V17ZCwjPHv6AURQw5uOa13nmuexIP5IDydrhyTfaX6uM
fMxVnJdsOpxSIDSxFRQxJ+NFzX2F7T/W6fL+mAk2ChJyJI54bv97ATJT3Z+e4u2fLF08x+e+x1Ff
6C5L+5zV1dJ014iU6Wi3boIi580Frvt1AMCwA09mJWP0kZ0nBL/slCptCC8HA9otjWe+ZlaNK/UH
tHdxvkfsBkYjwVnJeaIXCTdr7Zu11+WBFYItQeQrHscjl1SdBuwqoyw8iob+xP9rLWMNW2yyjLQI
zVISNskQfUsyXg8LNI/otgh/HvTY8O77sMwuuaUC5B4YG/HHfI8IL6K3VjumJhhX2D5+xuyksceJ
BIT9megADtqcpSqNeWjLAoZZ5T1cZavnp8nS2K+xiDBHcFs5jPIfYyFhmzkqUvUlwL/uBbfJp8Q1
GAhopEaJLQrIQ9xqLYmPRxmKh/K4jbGxP3HNwlwfndiPtrwyQOGabGjCYMeL4ip8SAfw0eiPIqFA
tGCfOMlN9p99Q77N9IPEHa6FR9QtGOZf2aAs0kdidpyPfGkIvmB3AIcvTQpqmso8D+KNwgR7mcjn
7qLrybqWgEWf/CpkS6FAVp7GuLKuvEw2NzDQYkbXdTdSlQlxuF+kZxaC/DPpCL+zZsLxz1r9wIbz
dDtOpxzhY71xF7S7SR70wyZX81XuTYfjqVDBlzk1nUgUhvK0Mk09kAN10rqOmtEpyzsVaAOb2qNq
y3ZgrLy/WEI7qIghZJyZ2Q+aHqEfLeeQIVykiaqgdphq+LA/PI0pG95Z/0ut2nWVpH4bd1oj5qsk
6gUDaCwtnHwfcIhWK9zKxnnHFgdthlyNV6i/WCEtHbVETO2lW05Bx60YG0Uc8IiKj5WKLKorhiHv
GRcXAr1ue/PNoE+e37SEUdZgrWfevSL7xpPLf8jrlk+ACV4tkh6npuDnhZYVD3otiL17fbkxbcv7
Hv5eQONow92SxBhW/TwUs+g1P5or/j+Yo2/WoKNIwPOcUtC50BOYh42jQkQhCJiGs+U69uR3Uzlm
TFDexeJG7mSJx2t1/ceGwwVRxwhiWhref3E/qtgPAXI4UrVnJCfy0RhlcdzT6sKTqK7P9Htbw/c1
M7HXCOytH2oJ58khyb1ultQFLvO9dd1TD+1IBGsA7OjoX46C5BNzKkwcWGl9Oy8e+dN3ShL0kj6h
1d3rQ1krMY4oqP0E9c0oH3rety1w/QmUsAs6GPmL78UF8dsbZGlf7hpxiKjjJvtYxNuJ2TUfuDHp
lAHfZwnImFeauyJatEnL0k3AlsGke/RRxh+61FUeb1PyBjFVzTzTfDznYJyltNScLZPxoiCjFSBH
nzBfQZz8Veo5iEk7ePCNHJcWDf2NFzWKoVD7qdhpzy4v3NBkmDinm8IZJMHta+i4QRXnzsRkDeqT
Yhl8E454iMKpVySYvPjmPPszN1xCYqsxzvbViv6zJ2ctOVvWBsPSe0CU7Rw4tG2bckaVIYsSfLzZ
S/pfYnzxIcQCGLP6cb8ntJFQNfJqRq0rJUBPEK4hoyKShBLfwl1ltNHyDY2fMnjskqXWC5I3WLI5
ahCJhqzivUV/7VIoPyCLKDfDR83BAhwjRTOVWc8ZpVyIR4pzwvUy4WfZXdyP0xeq8fhlbhJpzUnp
Xug9Pbl8VCsqi8mdt1YSwotL4PyyyBX2AWNJBsyF11M5VaBeV+wZrUxVphIHkQEkR0MaF8SkNGC3
kgZvBJLwv1LOVmYrdVtqRQ5quorSrx8SkI0i+znpHpOcMwNZAO4dLJuHlrWxscCN0Zm+PyL2B9dv
OazcaACxGjZHJeOIrzm5PZUL+y1qT9/NQthRPCwaiF7/jiLBcr5WmtWja/j5FIspC+Rd54w4uo42
s9cPhNiN/pHoWGQ1VtqGKCYFPt3ZV8PR3OHfM1d21MwB3gy3AVtsVUla2dqK9D/0wKLafnL4hHc5
O22h3+/MvvRQPGP/cuaAw7rFo0dmAUIYA/AAqnLGPWaGXNiw47IU7bQ8WrmC5lbybvFTp3y3DoGZ
p8/ZdCoa4xDuS9LWzIz0aDcYJY84QGRDzI3Isg/xKUwUJozGB+aBdvGuffvMQAtnKNM2DvLua5Gq
u6cYus+WmFBlpBM6gXpVKHqLNPvM2B6RStxoJCfjwYWCrb5j/nrNd0PbuCNHCgiKHnc6SPD1Z9d6
8Z9WgRWNDBQZox0QFvHn2b7UEc83ZIvAfTFDweh47vLKH93eY5kM2CFDJGpzMj5A+w6nyqOA8vuY
Uj3sOEzEybbmT5PDXoQEcQWhtfvuP3CPMPYcSV2wyVDrY9cMxqIzj8TuHuPF/FgvFf0yRq5L7Bkh
/219KnUIJhX2H2WmCK3qnWaG9k5wl93cNdV3BCybuXNu+jH1+X6a5I0Job+ipdRzKBlvhuZXc8jV
uNQGMK0D4W/oAjY9sTYFmXFPTNtde8Wxgj1jcth1NtoFOV6rKk7mQ3lojEgBmwFRrO/MMxeq+Zs4
vj6gnlS3cNJEcD6B4xUPvaNaaZxb+9gecaK/pOlwRwZ9MjY/vl9ToArCPK1W149YNc0aA0ezgK4e
cpJqzQ59hQfEXjPNvs0iViRqndXky85ziaju6hUrdAOOZuvcosXi1pCEwc5mSETKc7GjMjAeelWL
u0F/CtTN/ZA1G4t1CujuRSM6NzI+hA1YQWFmSh9eFusuhS5lQL5BMY8m1x1pTmRqm0t+RlmSxMzo
HWXGAi1YpRPsRXbRKQ65IbelwKRbASHj23qRuwGRs21WxEFa4yWw5UUri1gDQiCCs2WzyWmR44Ay
r5Q0jEO0FcrrOlDRqocAfWSRZElbMy30nvL4a0Od0wmZA5foz8KEeJ1S90SCcBvhNi1on/ityxPl
oCGL0GAEdMCDiWrfwFLkYDfiTCOK5I4TzGtMoTIzMzJmU4IHkublCpxcUceTOdpAggTASKJlZ3gi
uFbz04RTkukS5nAnyMqZ8K6PKocqiOn5iywNkMl83hpAdxTlrUAZEKYZfXxo/23u2orhZA5HpIBU
UbXMF0w24OZcffxNJPmLX1TFvn0oKel7f2iziP/f4KrmFBAiYlbmt0/w3pbrc9GRMWnU8BBjbOfh
IyozgDRFy1WBX60DGm+DOI/JWD5bdP7rN7zTdJJSKZFEchZtuVIHMT5vpSWlBNQlN1yjREF7/D2V
TbQ5vNos/74uh02JnO79e6dXB3sa1B26Tw6Lw1CybfnOXZV9olQ2/dOPXKFhGXkebRbfLHyl1nzP
QF6BoL/Uk9tPzavR9yl30E1dWADl4O1UjkDxdY5QMbcxThB5Z7RRjk9F3NUpFMZKlbDUXuhQ+Xp5
TtFTkyk7tiUBW3Dx4iXtSUsCQAHNs8RB+M0p33yN1+93UHHeM8Sg+zrjKCNJw0IN7BtcgfKjYBEm
IhPfsL7U9Ap/OFnqpSyNQMPsHW118FvEVnbLrQHXwSmxFXobwNub+gR8mES0R9rEirJNoefq08j/
EqLUKfwEYcClveu+lLIn1trpe8kaat7TYi+NnWuM05hwJjML035ROOc/FpNZOsgXIFBBgX81/26b
Ev727d4AxD3RWJNsAOJY5RxeiOV8bmA6XhWqwzbpckLHRecCxguFbyhb7UkSKBtK9tBPF5DhFVz0
+lS9x/UG2zyuPozOZZAojHbonxEvTpaGTbuEBLgVs10Etv9RGo2gtq6nIOhGL61QhbyhfSKF5mrQ
tH33Rspf5qmA5B1zhAiBoleMh1UQ4F0N5+ToxJhqxSDzlj8ZQM+4kNqIA50YecR1Iwf4PDBMg5/W
rzaDYCKxNaWrEIM+yAssYCQlKnfbKtxl7RSSSWCpE+UwwAyR/x14VXFwh47m+1jwpkNYeLmMAC0K
7IfapVCMtcyqJEx/kce2sEKeFRXgRNcSG9OEJP9SfJaEYnTWbMEW3MWVNM7GXxVkr0POQwnbmNRf
SDZnfSaXbIOJTqacMu/Q3V9CXQkD5tkHHC9uHRK0YXGj2ztEYYmDHvKlhd+kjDT/rD/jpBVkkgSX
jlOfdKZo1v/pRE18KFQvGvs971mHOrnoRYZfTKKVOoE60n/ll/zuDltAE6EkfWTuTB8uacMo5pHw
lB/IuO+thSsleiA2yeEgnm06WRTEr2MQKQFNidKy327wt7HU+uYRFyMaevucGpJSrM33f0x9pbh8
pwrqYFDzqmCQHsil1O5MR0Y4kgFmwIEco43y9ToT9CDz6688sB1iXYfDLxcrsPsYf21TpPiCQQdf
qtstHMCWO3jymWWL9vLvkoQ3i7F7y1nm1kL4FppgnPW4Wf4zlqaAucYlb6+jfbzBp+RVBlyGvAbc
eqEyLKpRmO0sfqq30HIgxXhbuGGr+/dJea8RRD+OCWTOFchWxN9yXpJIKHdKJAQWwpzktahMBLZQ
aAH98tkqwETGnFwtgOgFwnQTzClscYY9vYM/hA9cqL0QdnY0QFHbc+WV+QfhEm4lWcp2ZGChXeAH
EkCiBcBa9O7uJXI8WduzMP8e/VbwoZHmMoWUH23F8ma100j/sFkiwbhJ09BEXQPjKt7r1zFAFOIX
Xb8q0gUaDq6llaXp2Q9xz8j8FJgxeXOvaeR/PE8QzDg7TUdedzTol6b2OSj1oOXFRlyGCKxerelV
Ajt8DkGBKpnfMeQfdwW87QG7yNlXOwddC8vyq5MHl+qEVOKCsgZDZQySLNT526YMetXCu2vyJ9vz
jgkfqHs2oHVrw7br5aHnOL52wP4vVU7KIB+U3yYaaUqF4LbWSHjs+wagSbNSPE3HTFZoGR2Kb2W9
XF2ldR7A3pVX33/ucue1/qT8IX7xsVX6OQg2DjKAtr39seZRId/IvDyCKWWiN1SAbetMl8okzhBD
jUfyEFJDeAO0wSE7+ZhT1NzM1gz13sC48LxZiAeUbZcyLVe4D9TgWk29aDuwJ/f+lQEOCaO3OBYL
ohgBKOMA5kSUveayGAfOsKUZWJIlZWRvNgnudz12jn7+0H4E3AG3UW1Exc+YtlFFISTevdsbJZRr
vexQ4qAekLXffOwG8xNZGRjCMqyLLb3KDkAgIDby8qiRxGjOHHXPK9dHex3DhF74iSmtX/ycTpHI
g4jSfP3aWOC7FNOXr2IHY4b/pxqANUy4BzleoIvCbgCKVb9M8xvL7pKwpCMbqyroX7dIj/gDdTK6
NNgzrlxSt6DY0NqumW5MkvIm6/mJUdrawTFAcPjmo4/A2eOy1E3YD8mbC2RAso3gy7g+GGi8QjDk
lmSL2YsrrzmQjOgaYdVyxpTSGQZ0rHPH/ZQtYdH3toFWf49jwH1QedOMohvQ6Onvf/NIMk48VLrN
9yxrcbHdghgmqOLVQ1i0nFqS4JRA653qK8QC9kCetZ1I+vXPSepDSCdJebcccUP98ZPuuhHIiM2P
yUJKNhvLf9dyziWZkFRiJ3mLyLg+bIkihtjzrrIGZN99/pJ1z16gyv5mb9YZqmREKM42EqSsNKOB
71zpklHkjTJetRiu+7En6U51rhO6Q8h8YaPE6TC86R/Ye0/PP/XR6tDB17XxbscI5WWVH755l7de
PG9vUJPZKlWJS6CF/nX76UKpflx8Uq29qZiwpI+mi4LjgYXk+KN4W4uIj9WhSwtXwFePYNDUIRTY
mX/ig3UVUSggix1DvKxEXJvWzYIyQVzPWZEMrmR6Tzj5hHPjgJnkSBz2qwg9w7ZEx/OIWx2WTU0d
kkl467Ylpk2SkhGwEf+8ps6NZiyOPY4QGQI+Q8rxvJF3eHHN2+Sj5rvdMqxk6EM1f4CMvMVA+tQe
uiRlMcmH6B7jG4PK/GJ5o990Q4sbsnt0IEIujBr3nZVPKYW1aGdSxdbrZ+k8p0SKJ/B/EiMT2qPc
ywfpZnLBvEPLDYvu4l/QcuvULPzz+hlhFXcisJ8uEjrQSCbKryeby0DGnrPP0JifNy/MwozHX7Tr
pSeKPLXTcKVtUi+DnTRZSgVu2C8aCWyBrURjy5TLUa1Qfc8JrafWNNfyIavhwFpzmt81fMBKVc41
Hr1Q1WUqZdxqMJl0nVcMvVC68DfWU3FIjoV7eFgkg2mZg4NBQVSko+lvOTo7C3Cbb/M4q8GqaDB5
54gGRZONn8UflU+8xzDyOPLQ2AnFfb7c5KozcRZ26A5sHw76S1ADBM5optFkAup5q02SsU/y2HBg
b9LpT29HFzBCw7Zpw3sLL+cf49tc/3ZbGEYOgqGUHmELqdf9oiXMsYaqqzTLwujvu0qLWSlr421s
iEXOKW8qWDrj+R4kC6qiRF6DLBhMEbpeUbO5Ak50LDGeXioDQzZ3w7PxzPutEjYGjBnl2Q8c4snZ
gvSjt9Zu7AkOQp0ujC8bpW2LIVHIL1MAV+GYy5ZaIKU5g79lwz2u2BcNjQbY9BpIgHErndYZ7jsR
jOtaLoIZ/A+WeKGxh/JXE3deLW4lsVBUDl6j3+deYbsrur4n4xUBQqh7wKHg1kbRHmX5uui5Xik/
6K9nojE/I6Dw+MEMiW0nsGJyCSVa697z5kTTs3y5YT2YO9g6gXottMm4gSwl14osMmlTLiKfgjbc
GmI6qRY1aB61p4GJ4uKc5xv/ciZF8Pzx6jYQqCMxDEQ+qvM3UpLBSM8AY05AUgqeMEwdQyvjufnV
pBOfeEnFEWGGfi/fzIy3A+Y4HTadZVrXHX2Ny657MiKl3DgJuQ+Xx8pH9mv7AkuWrkk7IeHnki+C
nqrgASUN88po5Pf1A1zJuu6k6GGxMWehRUIapFPkUMma271j2/tIJ3Ad4IF8K+76TeoBQCcu3VhM
Sr/n4KaBLvNYad3PHh7aeWehM7ima/+8ikNGnTtEqj/+V5XXou++ipY1Dz5A/Afs0Z/7hqaUO9uv
Ha2iSm/aA9ZRW9C9j80sbI8v3ELQ4RaWDbvb8aQcj3QJB0vb7DaxT/xJWk3OkSrLYTVcTPLft7vA
d0XLeCr47QdoxspVJ9KAhRj4fsW4bZ0PM+AZ9MuN91RlZ88FTDtMPK3WPyZ6w8hv755C4buJSyEk
ULtArj75q1GYCMjKAPb/Hdlm5tX6lQLdLoto95kgQ9T/C8gIsjJDZbzmpMEGB0fm8t06XxpVP4xi
9050AA9QWQOEBPIXAZlfx1iNhZSvwDes2juFrYZBlB7Z2+Cbu+OjjeZ1QNvf4Fl/ZP2Vgn9046+k
H3BH+nhi4Mj2qzTtCzQXaTgPtZebv37b+4d0bVRFbAJnd37N7ngasY4NVWnpMKiUW8lj7eXnWIlw
lBqTb3fdgiZnSsKTTH3XWVYgrrBUTSXjADvuNKmDs+GShKUHb9zeL6YAmiC8TCSEnaE+g5jzC06J
bwIR+hnuktkqcUc3b1PgEhZUiyhxLAihTH6/Nt5tFhNvZaNy70aESTmzzHsD37cDPMq7wpmuym64
GsLwJQPhME6rAwvr1WSgIi2iHfH17PeHvpV390TFII9pduwfy0q8VCkKUCVo8gUZ7H0g0IpoLTUV
75wAlxWsWnNJWYrvcIqQlXjiWwwBn8YP8EKEtECE4T/ub8Wop+EVvjYaqrxwB6H8h/YgkZP4CDV3
LJvRtfeMCtUu5f9HvWjMntRX+1KqVyC5EQjDkMa2Ww6L6bY724zCShFoSLLWuUjGXFu3WWcaQq50
t3dls6H2v/DzDWmaBeBtK9MEnvP6FHkDCRcaEDbMlZso2X/UaThM9bsH4dCOUqTOFhtTc209JOQ5
qPBudrn6bwR/reE4Ozo3RIPlpqn81vfHC5XFHGUacUbwgq5oeyKv8nunfX4bOu2K27glLqcipIZU
vdounUjGvER8O7Jja4E8BuMIEBzJmFGiURnt+ZFvcE9W4stYZx2m2zubXUap7CS+6XTk7cXe3cTq
I7zmTu683cFHPbU+Vt8C6j4Ai7in0X1NfXoCakEwA/bdCaAXS2wVS3Vc6KBPqYhRbBfgUkuJ7HJ3
hrP33CvcpAnjCzLj5pfg/VIGgHHfDT4isbSHrVYtojpu3CDHl374OJOgHsjMzPt9TeMpG697WRJd
1Ef5TueO3Arn4zl/a/+WQjwF2t8hEZLWRRDbiVwUemJDpEPFGnU1kz8N3gvr7dej47tAGoJO5IzB
WrOVxDPF1dVzQoiZnSnPRvnfU3aULaOi7SE/Uz6rqYv70SQhPSPlaAu/zjaInUuUDPoVjMiTln13
rrkSSvA8+YFEUmOQLq7P7YDoHMY8fAPZuOX5Vf0CuP5gGoalpYfg7vWod/JaJrKNWc5JVwxAeWmx
mpllhvc0wQv306OB1OqJS+sxQLyXPUmz4c0Dlnpql95qVaOG+a2o00qSnwlWygzJe5m7c/QV4o+8
fB0F7YumomACsPTnFf5yJ+HOiZNRLE5NRLJQumNc6/9VQySsmnhgknYUW20M6ItPZhRODH+jFUrG
rMpCNBNIezQuIappVkpMqDtA4pz43jxK7eDeu8PDlhcmzc1RicpFu0HmVNbJs789LcK0P/lOg/6H
v8MqmAU+7325fjgTNjBJh95dnWMdJGVRBUUTMw+IMDeGFQ4koA8Q03WTRUpmbKReHjyTRUsOsIBZ
W1Aa4AF0Q6Ea5Yozxg8osxGOnfVmnWWrhOCgibk+L3aJib+ZIw3wH43114rvRC690CxzQUU3iCtU
XH7TwHyiBUE6XNzTuJC42g3zToI3TTSztt0SIASNGibZHmn/UaBlf7aXlq45o6TtBH6KY5Yzkrgg
HBJdmnpZJNsJ06cckm1RUwbrnYMMEFSoqO7tnFd+KjT5FnxdnLQ7XcdzkZLTc3aOt88EB16ouU2R
ovNaF8roFaL8r3BZ4cR69Lis9CyD2ZFexPBiejjOqqmPc1OHuiZQr5CHjdLz5+8ZiFp3jXkbX7ma
cU1JU2arv/FAbjdqxhkvZZAoWfNyOMOdxeP3SmMN8CVqiRE+YlWVTv5+v9AsBt6DcdMrcSCTK1Ry
5Y73iQzK9Sshtms06dHXK897f3Xa5OlRzE6l88oJvV0+c8Ci5zkT/ZGV/FS2/9oCl/HDHyVBdUHQ
7HMspBcKkXtoaGwizZmZxmWL71aTzz4faA05GBd9OlqCacoAsBKBMkgJx3SqgugbFR/RFnvSmKl3
i75T+D47Qe/m3ey+mD/A9ER1XEl/4sfq0lfIxkgHh4q7h63f39kP9j6cjDBD8V1vLxK3F/QMKFdI
fYrCWB1Pa619uM7TdoiWIYUJtqNvbqgPih2dtbeuyelLs/jWFvl31ebjpcd1IX/vNNA7jY4s6ZQW
jxEHC10juqO6dMHdEJepZf9pyS+ye7xV7YodxsQ+hscvKk9GRFdwK0fNi2oCvKkubT0E9xUoZkE/
Y/KXVzyMTQbErK3mFHh8+BKnV1dsEEHI36AfTgrQszKwqawbsnARTs1xtg00rEt+GLOcZX16eQ81
RjEpGUIIp1Jbn7jCwTM5IxB4EFn/omZestkYR6IGAKqhpyhhOx4outFza7q+o2nhTMr+o+9jlA5Y
llpcHfwabgPb7MXeP8TVVCoPLoZM5L3DSOhot7IYWV+F99G6IyUgzcScXaPs+Xbq+ZSJCJ1znb6X
+6K7QF6oGv/7K2LbFpjslaJJ4wCW7fprA9897imcJytmXOYsgBTCfuE1NHANc80orvlU1Doeildg
oX6pxo/hjB2KpgAHbrKIUnydrylmjeP4R4pOGv43vkGpUc/ZoNtUgNCQQTa3UOkXK3f73Xh/x4bL
oEBbKJvDPTYSPhitDrIfVZp1ovYn0n/UTYTFGokkf5sad2+3BLsI9moIg7/Du+7zH81tUOxJS2+5
O2sDZoxnksaLZ92s7P3zDezkxivKN3cXpnrZQMMbytGn8CG6Yl5+X4pxRfePxHtSquFkUbFytxRE
KMBmplWhR7eREnj5bYxeoklo+dI58NuQtBwX3CSWKN7OFQnyvor0xl0rftBpllPhuPooEY2WWeUq
I44e1ujrvV6BySs4mbXUzm9BVuLZ2L/ZeuDO6X34V+SSNCGgAJwgO0uSgAms9UtikLGtAI7Ti36U
1c/jP7UeA5YwjymW6V+SwyE4swGq+67/80042f7cYA9AbaWlWVMHv2XFVGYw0DWxr05QtFXivD+q
t9wo7RgM5AXV/sCikygN7y2CN/A1UNmGVyJV4/xK0R70Dz8Ii6N7WKpQVfrWp09T6O/5i2HQMKdu
6Pxm5ngToAL0NVCF/WSNXTPMVaMN8BzgaweZca1ci6gaP3WGjz40SFY38B9eyj4DgHd2C1OLR0YL
hNsQPXay1fP5uieJ7HTtZbion4qf+dY+PD2AFooci1xsrQby9bNVFHTIEwzTW9LJ+M8Acxc/t5ao
Nnxco57H+8r5Shi0iZpWtt5FdzPv0Nz99BRGEA3UxQzzZk6NshrAx629AiXIjvSED2M2eZqLFy1+
GbdkiNZ5M7XeWDCe5+3t/5ZMCys+mnVNVI41zXRK5zMAiLaYJt0KGcigS0dzpHnD+4E1/P/q5SEt
eFVAD6XNhydrctHXUdenn8fsnCs5qfjBQQXcM9dS1rKr+dM82+Cpb+dH2PuRiiWa6gkMZ9pf7S6X
9h08c8IiA1QPWWj0lEcmie5g2mXcJo+CQDyjO9xO6fbdhq0NwmqZoyXYj6MXHCSkSxfUX4RtTRqX
99DRoeK5kP+KqPFxGTqN4KNKx9LvqWMG6rX44ye8+yIU4LrYgT8RunkEVqX3gZfUegzHmcUUiqmJ
IwiLrcCoIoM1OsCaLS5SuM70qRcHMgRCJkQtOx4sOuSrfLrSRTvhoouuuLy8/IiZ1/UEWeXF29xG
Q1YE0dkxZd1nsdJH3bU/iE3LHNLcGRbVJmxFxAt5JxFnOtiQeULO7WaEQuoL7KJQtW+9xRY9Mycw
WqpZ7Vnk1R77X0+JSMyotio7YfduC4ZLUrgc7HgSsUxUKpvIIfglQNax5BklY3GUAiJTOYB+qh5N
QCSbGxTbTfbrzOLn2Umtw3MuSzTc+CGRod9n9Hw5vFqw8w9W7dIsHo9aU7K4h8RnuxBHmKi0ZL5z
2DBWFJKHRpr2KGGvBQlNDi5x9KbmjYbK3oR68bZnIudYgFrOUvcmZmgboZKHxEap8bOza1iqw+QB
wQpIgk8dFsPAXOVnYcQdixFgpB0egs+ALeoe7TDpcCi4bt/LNMsA9na3LM7SOZbibzTAaUN2rfx7
ERAFHE5q6+XdoVogIuXa1nmARgzYHEsYAhKNMEYQlg50wRfwVpeN0cfDQyZqIE1frU0B7XM+BEDd
pnKFdJ8wqDnKI0e08oUKr4PLi1+ZzunLX/0wJZkWs+ZsDzDQLU/osESh8eoThPBluzEPfGKR3521
EkxyvVr7kmdrURgl+iHARzwaNlBT+CP1o/8N8B4bWXWPRyDLxVW0limUWkG18umRG8dhcJPHpvfQ
4kDe4lUzE0mZrfJlEILzOl/euD/pMignYaYPDw1iNO6IT0JC6uDEyWw8dAd01rjFENpz9P9p0dXw
FTd2iOwryMdtbvVkQmxJJqBg5pZcy6dnBlKUcCubqdHMmtyNagP1t+LvTXoAEKCY5EVpxAUfpyUE
r8aNgUE+8KxJydrM2dpgCUjqx8pFqkPZKT4+Egq+lXPS/gAhH2+nFHndrN0ZiO8Q90oFJf2iD8zE
363m1J2+vGTWbOlXIBkHghAh2Ksa4WIEyLPsbdktIPTlLk9g+eVz5KVBT2L1DH7EjKkjPc+ocuQ7
yNI/oKTClXhaEop7uTKgWaTGHBaBZnnpQEUAtcInAX49aXwbgAsKF869XSAGBwTvteJ+JDnNwv7A
Mk3q5/e+RfVDVXLofwGdtWa/CY+BtdxO6iUAwASXdR41acOXKUmCXwmkt9uJmCi8Y56hlCrSWFYx
nJu60EPfWSH9fuB2u6M5+D/FAxVv8pq4qnTPyEBRhcgNgmVFWJuvus7+SraNgscZ8oLkYDTa7+6u
SdTzMUcoJ2OGEBg0jXtMhiPs41dPYAj+zWsRp0bZ4U3Gv+Gw3KAShl4+klr3vd3Tyw92dl2KXtJd
ij6mP9s6/Gqgg2pNB4cAhJE2O9HCtS2xJJ1O4hUs8WEfo95K+iu5vTCOcExVvXs7fhH0rBBbDxS0
4+nwc3BFFnvhq/RxOzH2rmkE1SxQ1sk+Fif233azSLsZGqKbuckiwvxbrF974ARAvHjJ3QtRydeI
Jwl8imF8pEQ74zV4qwsaTmDPVGsNTAbqUeCl4c7WLbBoTlrLIFyc95tQSqfarXs6lc5KXivqst4K
aJjdU8KPtyJAVtOb7anrzVzG0ivMZbImUUJjMOvBcPjgcr4BhFDNhOPOdhwNXZtecdRVJGpa/7ZQ
X0btBjmgF5gQbBDRcvb8NXjlzdP+NTZBCsGvdI0zJKOKAb/oqxoAOHpN6QP5N//DRdz+igeVnbi4
pf7INmkyalGq+UGkQAiShWOYx8S4hf5wUHVO7RdDlboYbplFf/Hcyheb8kaP7o3WS8+fKoYzl1GF
uc2Wvy/gz4m9EktDaVUVPyYIcirqMJEFEpU9tWl05EnnrO1J5bNlzeFAkz6j474lq/fhRBM1Zp8f
RwcvpsjXaLlR023xMXqdEYaZ2z8zRx8qqZmH79EAqBTVK9Uv1WOlO8/RhAwup5D6Y7ZelCa136yq
hp7uxnfqE2GAbRkAC8n0CVrEnTpko0GQRBkpIchNs9MXuHoF86zzE1b5O59hpqei9ELA8bTQTaRA
G9ONuGfgn52AZGd67WrnpbER7Ch56kBBRWQgnt3X3OSFRyIC6bILVWzaVFggac7AcEJWbQFFC6XF
BdC5xj6MMZBiWCxJrTJhirygDKbhwp4eo1eTX6TkxkL4wP24GZdzeJa7VOfl+t3m6ZUMrlJB6+cv
Hbem+IOQI+DHVqvCbFUT8Mw/GiWtsKTCx7gwwnVXAA6bXZjZyTJiR0KcR9GMf6Lb1gviCb4jaric
Keb2u/p/+ape8KdRzQWwdyoWYrOpLCYEJ5ytgFoqTcrlJDdbEOVEwkAfkWlH9NMzWPApij3sXe2X
GeOIGdRPl8piGNkphKHEh3HXVqRTED4731+eg2HTy4gxBW26HSAJLsGqEFsnbtbaupGdjUQ4pjMi
kfi1tFHgycc+obu5V/FWJWukN1tYjo70PwAmccwN3BfjN/6MeMAs4TEux+2MBXR7JPhJ1KMKlh50
rr3Wn8j+5pE8WjIxNe0kFQiKNDDaijG3OMERWY5J99aTMpQJqzpdqub+/iQF1bzqBCSOw9HYTJBx
MAUAY9Ph8Pkd1FgGxlGWt51DdgEqF1KryH+UOaoSIPv3r5arXWuNKdDc7IkNTa1yuXV1aaX/RMM5
s0ppUpS7t4Cfv2PyqrpzEVuI+VMTwNPYWCe7nWQOE45kgAqgCQHZy6qnsaoAhhWQDIFizzlkGs6/
3KcXQhCSg7aqGqMJDU3C+Pv8WOSHcoSVZ1igU43EX8B/nXdivKLpn6lR49Q+n0ik7T69BSR9fR+a
ZUgba1+2plaKpQbfzkce7Kc0t8S8hvOI+9jdZdPGSTTefXp90/KtZf/O+HrvGTmueobh/1811W5P
Z5zQPxgx1PVOqDeUAQ7thsv+xHROn4gz2Ani+FM1yWeY5c1Nb72+dzFUH18q91DGALV9XZBsnW2W
GUiOs3qUbiC09Lku8Iry6yi4L4yCIx+K/DNr83FfA1wn6THjDh21Fr7GbYryWSxP56trexckxwEA
M07P0N1ib4ZFFmacvMzHGdmo5GGDznZsYFCqvYLCC0vnVzayMmBACHafWisVfbsbdG2dkBHAAa8I
tSQxKszbuYLN5+xeFsXlzl8ZNhQpjwsj1eJ2yn9PCRVf6cS+sOpXFmaKwM7ZpYJZsbynSN1u8iHw
jnyv/EJmRkD0tMHl/w1gbA1TcmkldtK7s/eAa0J06l14Jbfnet9EZ93XPCTn33fPPvW1cZn0q5Rw
pUGVyxuAMCi6uEcKs1kLG2K1PNAhITz5+9Sa/AVrAhVsupWF2Qcxx4afAcqZmpgcyOonYg0BqTeZ
3KmCk1EZnbsCSQqcQSA8tvkGFagUJZN5yK0MJ7RfVtYxvaW7Len/ZcpxL2ckg3mTiV96YrCdXur/
zqF1n+EPywcBJs0/UPDAdj3GS0efC3Y+XD0XYnJQskDXE3w1guKiTSCQYYZ4ZaIY4s922PzKLOEJ
unWNluRRTo1A0ZO4Ae1NSsfR9pZLMRpw7wk05XC2nO040t2NcWEq0FmaPUM3rhCMNGqo6yVI30UH
dcTKC0Iho8HAP6HwQA6kpGs3PpLrQaG59qnJnN0Uz8GwQSfR+6iNQNUEE/4sBNT3+prGHpP0ROBw
Tp3R3cExfx9IvTeMVANGGCmuGDoEVl2oGFSZrPvkrlKgfXWkM+87SW0QHfFZMxPBPh/zuCftm8mj
NL7+CsZrcikyNWtL0G+CeRpkwlep471JrYIXXIyFjZfLKW4yXepUXlYmd+ABFcGm0yCPV+sgcV0H
Xn9y0RLmS4UGuYFz3f/xOHzA2s3YM3oVY9lS6wSWeBESx5NPn5YjwZTqBKWES7IoG2XwHZendMxL
KNN659j7iUWyCTT1t1X7tvFRjbKl9Z4n6zg2FL70TliO4TNibzhf4WCst2ejS4kKLDpnuHzrD8fN
ypHwQ50b/Kk1sEU3pw93oCXZbrymCMba49DOQkwBamayXhgtK9SurCi6y59jJweq9lzglD+kLBQB
lWlBpCL9+df54pftRopRtyxpo42nm08JtNfNJqZRq3ItjCchjPQgpM28Rh12TQcET1veFtjweIcj
PCb2gRkiSLyhnMtshcAxOy/+J9j4m/1RNLIKe33UfIGk9bdKQnA47LmMMfgVcx/eaADrYmWQ0ZdL
ByyTW2r4cdBARMOZz0CuHTpIz8rVSeiCP8h5KZugugXSnR+rcvFkSZy4ZwdRaEV0fSdsB44el+4w
s37iHaySzhVBcP6k7kcULQPbnokYqpXjUJDV4gUuRbYuLDCOtO1w3o50DqtVZxbaebuTlsPfkUiK
Dvv5sexczoISAgES62tCNWcZGkt54tJsnvZGpUw8uEKr/v55sWlpJPmvldWg7p4UOr18f+5d7B/f
g9P6HWwrg3QZewRaHA9tWgFN5zZZ+5ZkzKI3uNjqvbfPTLudgieQeEgjgh527GCeq2s1ezfYHZm4
KMyZqed7GdkaXUDTMtGGANJOqNwiBGrc8IGVmql/S0kYR311+6nAklJ+tpjwSL5YMLsthj7SDQxP
rlyCPuc2+KAAYkdugcq1BpqljYfsIeMcTshia/ZkqBUOBrB+kf+wKg9XyDp8XhhKJJ+IZO8vzNfz
r8+ogbHDeX7LbaF/18lj18m2EDcjbZu2GPbLfO/iGWysrZpKuRvdWi07MDYoSL53qiV61lvuTy2o
hNTmpGshSVkP7uYMqT6VoSCWt/og+nwkOiVoZtUu2JWF4e9uqiI9Ub7g3YeTCwwhR1NAA6eYnBIX
W9kEbyGXG9ugnkzap9O1ahfxdq2JLJZ1P7VH3xeX8Hz9/p/cYHxrsZCsmjM4xNclmVvj/D6oEMQm
UmjVYzZgQMWMiLPToUVgPgafA6yzbWtfNud/z+qKxWAu03oQQlEhHK98K/JP/EFPzdQG2Tlq0f70
8k5NOH6X63yxMirGBickhRTlKaXj50aqn2aWW9koSbLlbxXzFYO9Vv1zUI4J9I2krxcGwVxQPWz4
neBrZ+U6lsJhcyDfETDIggSZSCCrEB6hEd4zIzhyRCBVpvFJFC8g6BaGH2YvyzMzeTRPEx7IvIT0
EeC/n8Whzq1PBl2UaaG1PZ0+cIGWFrPNiWzBci7giaha3XDfVYLun0yALR6OFkCH8EJP9qwtTcnR
pwMPCF2oq72fuhaY3H1R/NsVxkZMWlxULhzZkOJ4JK4FdpEusPBC+iF4quLcS7dyB/mls4oECUSM
GTocnNiSFz1657gNbXdNuNHcloWnk+SHNUOFxj5sVoYWKGav5W+IPgJ2T6Pij7pGgKheSaXelxQW
+VPOjTZn/y1rwbAwE20KfzacYxFjv876rZnmOkT9GKLTuKL9pnHj2pFfF3X4Jv+e4FIM85s4/Dwu
EyjBiBzq14l/CC0vjPxkd8bjBxOCl9+Q+umAvOSTMSbVsTE/pkuKQUOro1wIeWmNE0QMkZuDBjns
3Ar+GPXU8AnS8QRTWWOSkjFFY3KN/a5joPpWxEE8g6kwmsWSuCDcYQRJ8wGJNe2FBKIloxqSv1eW
0T8JAH1VXzHrh1qCPjDvzBf77XcrI6++SoBqNqYP+Fdd7koybIl5fOiOF1g6XwlTaQ3MqyfV8/mA
xrhSz7IVwh9CYajrTOvk4vVhw6shdCjBTzN8mT9BxxvwMCrft2on6Pw18PPlbLsHFqU6U2OG/lYv
m5yT2AzGwX4n6adlZRmhj0s/XsnOXeN3TzuqaLfejAhi8LqOn5TRI6YDC3j+SPVck/8undmmdQQl
dLlOzUmhTYLREEEktTpi5JAhLYRaLlVRKNoo1UtumuEWpVIRzmoI/DpwDGIXaFUUTX0/9HV1ZRNG
lF9jXjOx2cvBrB9kse7ZEejWINrF0JPr4np2fHYlQsIr7YxHPN8+ekcRuxEH8PKmeatf85U1i1oo
qWR+wYBV9odATvQRIeEFELkBuaxMUA8gxdA7DuXkzxy9SFwobwAr6PXwL8ot6KQa2KCTpFvB2tSZ
bInS0DcgjJKQTY2lBO+bfDdjoIxsRpQRExHBsfJb0P5Qs0iqBQwz03h/OMyDLNRERaliHfEuukdq
vyD71cn7iD6A8jt/dd0Y2srl1AarXdbFDMsb8fP9Gi/5t0zhKkGGX9OE93V/vmwGO72xTLSIqkNN
G/TRoSoxOjZHEDRi0e4cvZ5G5kpa3gS+qIHrYeE0UDMIA4vstDXrHFebGb6FsovKlJg29NTOep+Q
ir1DVqaLUPa7wm/qFvxjrhAxoQXMlyfKF7t0lnY9ihc3a3tPPH0Y45EfJG1/mBBM5XltsaQn9Md0
36U46kq8fayQ33SMumURobaVyi9hqLQt3toV7KrocuuAZSDBcDofXIvoOEE8uy0PRD5zGEzL88EI
QIGvSzP3ZLw0KNV07YSYsNqDwLxRzmYrJrDr7Xl0Vmg2TYkGRpqoyqX2pzGx3sFHB8YkgRUe2qf1
dIS4X1hwyZmTeRzMlju9GShZr6lJUhaQ/TenlcV+ur1RcmylC1Gw6OeghtwHVLfHg/thHaLh9Onw
eHkT7sVMNfLRTQX4UrmBI9xVDUgQlh8g8mwLK5MAY2ECGEuxuT0t2PZcf8me1e0DKJoaq5Z3TvGa
+XK0n5PEW1FRaFUoAcVU+HsXrnFJBf3+RU5gOZi88VEemUmubEzD7tGqI7voHcYNEbEztYbn0/OE
Djp9S44U8RLW0NinfYMlalzOyBq5W05FDqBJc5uKSUpTsAwE8eIVbBd9j10BKOM8B15RvDqI/L72
kLdXyvRgIJSvqFD1Kh9HmI3i2juOuLmlhWVpcxJVM7hWIa8UDqtNGcO2YTomKkuPOeRJZ8yJS+uW
52DZzxl+zHuDQvN4UFxsPqDz6Vv1ax3/BKivkCTRhpI3/OCOGG02uqqhzFm11Z8fbaVEw33qglBZ
JSlC6l3lV9maSPP4ig7Z1iVZxrrcJyc8Bg1+jcjPeXl5Vn7bi/uaJ0chc4Pg9cs0EVfPtV5EdmjO
PAu4OcaMaWxWzlLABz/7FrLu2U0/wmoViEcZVuS2VWtw/9pTPvnM/EHzLVw7xkGzMriH0wqgtEYr
5pliRed+YE/+Om08HUtIeF+JDAY3oAUiVkzFTT8/K/c7D5SG1wCEZnEGhKrAfDugoCVlHgrVyUjW
t1jPoikZaL2kEeMnSaycMbZ93W0mB6fkEQObjmIJMjrmdko/7+4Z6SC7ZCToXiTAUbfaOhtxYwDd
CTQRKibrCoB7+BNPYmLeGRNorC4CQOVm7tP8AJmFnKxOaMJf5qDIfj0QzxeDmjqsmtnMJgbh5B7q
aTwxiavVqSytWxvvrFc4eCU+F9h9FA3bAnYDbm8nQ8H7vHm5PMwVfq+6WjQjvnALab08VxzqQNRc
T4SgRz0vBpfWNkwQgJm/frTezDaJ1yJ6PW0YCaUrX4OtfxsyiwTYcoi5Fx/VqYfvit//EqB867Zq
3HaFsccAl58tNMTOM/dfEHiYUUQqIxhbDYTs+JyPy7XOdLG++bVTOwXbMh+DMVzTd+SZevrfeKhO
gFJF0guhkQX+6LOOWWF8sGNegovISZkRTWbGouTcbFPIBlf1IELbPVsJkQ7QFCxbAZFdkL7VmXvh
eOmlBWSkksrRNz5yc6tkxX7wSQk3JcUpg/dXjuNCZGGwIm+pCM6/jaYihgtMYInsinWPe+qKYwfq
Vl7wXF5fbROGG5kdhbD8hUY+Pup1x7rgQhe+AG6R60hKZI4rzSeehSnsXFSpUnHTgVy8bIyd7stR
ZK+TZuEmmNnVyJKJStMtfza+wzAtXLURLx+vHm+IuTMLC3x+FWuL3FOlWohSqWVzASluB8TyUTEG
7yBG3QTvG5drfRbFn8wI9/KASJh86jeOJ+Vz7hWP/GcTicsf9GN/hvjo6RXqHmsaOjCDBJ4Ehmck
Ir80LW3rvKw8PxpcBGOOpNdc4mAx5EkBk+H+oi66KL2k7bPmv6xWXMIbsFoHcu6JIO9F8kqZ0dtw
NlF7lIdzFus6xsZyYqcUAwSlS78p35MliIYB34wV8CndqNEtLgCKskCXnmuryKcDkZLuKbIRetHS
Ss1C495a+/AHe7j9ubHNM/SIu1NDZRcCcahUqumZRAJv12ay7QxAa8NCJW0WbLN8a2l1Af4gZsUr
vqro9+HWk5wKlRfy4zm9TdFogbAMq6TCY62FFUxmY3ZCxen116JwSaK7zIlCCXJVwXwx9Y0vQD2K
6jB1TDVQHFnlK/z7O6phdMZoHfwu5JQB3eArWsXdZaO3cvjvCr2IRqeJIgKvGUHA7GpfwZyF/z0k
JGJL5XZhfmGZiD4zA2QXv9BC5vU4v08oWXticNQgORJYf3NbCTO6c0tqO3awk8my0hupzYnmZNNZ
MuYFf71TMg3QSOtdvCrk0C/Cw7BQU1wNTetWSSku+26MAWd+8conFQzXNpZMFVUpH9FoOf/Cs+1c
puPuCF8H20+/ep0mKfT1f5rZq5ZIkMEIaO8VdFqEymiehyir23+kgF30TVZN+WjZITGF5aEizgwn
E6M/UR9IHpd/Ds9Y7oV6CdA181OT/d0qkQmzmkG+/SzJ6ziySUAeyieUBSG8O3IFtNMF8/Zm79lP
ElGwPD7152dvAGSEErVvHJVlHsGhOCkZLKeFDWUdqV083dsmzTAmOlTa3UpO5umdoaMIc/NkRg92
DA64TzMsgciJO2QtO+MGZxO+miLjF2rRh6LKM6V8W6rS4+jvK6NQr1lkd3haoaKTGuRIMl5Q1vfe
qtguE5ppAfUReSHwbm5ofR9Thpo+EXEwgs0ctdqj5c+R7r5PV1sGpQrlL7Po/fj5Ld3KlYkZl2uw
32xdVQMAjYMcvWOPfTE6vsTG2VlDTucnyHuNy7LIS3AtorYnHE/Wj0qsmj4AVWubwDgbqE4CimHc
lQz5OzXGqbY7sB1lIthaHB55OCGBo661Aw+t6rnWmL5+vQgi4Ckag6Ij/Nze+FqmYGfkzt4VvVCT
NKZ+ZYss3G7ykPYOZXxvwIRB+ujj/gdL2T4Ps8YthpvmwaitE3BH0nCk/IZm1JPWR/9Qem+MHyWa
/ZWP4/aj0DNPyxDuXpfq8PHITDACMubUdwc9KdjjHKEg3wfsmBF2NUCK+LryXksCd1pgrl4wZVmX
8myVk0G+o1LjxLZaTXd/i9atrO9qkoamxA9ImMtZzLarv38TOEcdQc7gRh9BKoRIEUncRifwIdzf
LKydcjKPOX41e/nRW/D9giwiqVhSYwz1u5GUIa986TsTi8AzoBrRMtXNqe5lcCJxmLPzxULxUS9H
bffO2Q9MrGoj/XUqnJ0ERDVgUi9NtTgxNwVnL1IGZ0K2L6n+vRYbptiLeGR/MSEJ7GT41HeZ1dGI
pxGoXyQMh2JJLbZek1eW2dkHFOa9jIWVrcsIoxEekMB9IGr0yVGGUO0VdtKLZioWre/UqOx4QGJf
FKSW+s9s66yDDQ62PDs0zB9Wtko+o4kDcSQd0KyUR2Pnrs+vnYqs2EIgyP3yiIeNZ9O5ksHLAIgU
4kTtuI+McCyM5C+Sp2RsrJI3BgfMPEc0FzTL9SfnWmWZVJEbWt5oeW83xCZkF9yJvnFJk64D9czZ
3/nFor5ac07vyknt7miKhzzE+1RORiN4Omd+RKlO3dfPodtVF5INKE5KoMpJaZFSkhDWf9GClVlF
AvS4MYhj1utPqgGQGablBT1iCUl2Ch0y95Aphl7gA3X4gIdcwVCd4E+0J4WjhEpkwG6EaJWgxW5Q
uxMnhKzKMwWQ+LNxzGuSM0pdzSa8Jem/TIVyvzAX8/zZziwjEmmvNBw6Fz0CqD5AFDV7Pn2Xfo/S
v+LdlPa5Jk2PDIMWH4LmO6j8yNSn+f2rx8n83HM++U1D1PsGvJFXX5tVo1mThcuBWGGLOm56bif1
cjpfYXqYIDxmzIGFK0hUasBtlDwYbPz7ZPFkp0VtRtvxv+oyZ9g6MmmKdTi7O7MKtnxywMT8yd5R
EX/UlZ0LfGe/YWEi7+M9oSW/Fk0H4sLCRkJfliwLFULUIw2CgGT4HTNn2SRtaToC2L0Zb4z4CkpV
9Ynaqmrz4Po3aHxjxVQ9uFLCO3qzkSDmlPy8SyeSamguIOAXquF+2hE17MWSaK33TlMMpn3T2g7J
HabUcEfNLfAb4ReTfsxGXCu7xkTsZkg04PsNtPRnEE+9EUsNks4w6C/FYqMFdQu4Ex5l/pj835Bb
H2h3HV3+IUkp3PwuNDA8txRAdJRIwkG0jqIIWAVYFEYkmNdPSGuWAtkLqWbaXH8sOGRo9NpBccV/
TqWUaEmH8ybmMhhHsrYoyzEWW64I09nxOiMcKR9gIOZ2ECT3dryeQPvVz2tv+4VPLgKLrWZWNx0K
p+ekDsv7WHcVpts+GlGLhvJsfXtS96FSvZyFU9IEUoelusPoUhdIrbegVT9gNAmUT0X7+57+IJ0+
x5vrc1NrzZLGXWALGXzAzvXFSq8jEuw2OaA4dMS+m5Cxk79dVpN6PZrHA7CD+R6F8cBvqJ7mCDK6
NImmP041H/ugGZpW6O0nAeubO/k2IBNJEvYHqJ+Jl+H8vHIjzP43unHDBcs7FsPKb1mhx/6w8j7z
9VjIirkZPIapWkYVTHoKzJ1G5bOea+UDEatE//hmiQLJTmDqXyYDwMvjRAtsoNP9n5eCgMcItkrU
2PAimZL0H087h1BW+Ssk7rv6hWB1bMkUtRlY/LbYmwsOVTeIyZhOoPwLJf9UmYup20FctxjVEOeg
cXDL7X9/AM8jKtaBvZGgef5tetchNyUE831dhyzIMdkQPz0XeNqETt0VU8MJY9b+e7Zg/q3f+g6c
71ErgztpYlDSOnEIqVVOlchsIGPG5ZzglDt+hSVr4NLo7NFA8eUP0gCgvNVGlE8nTB6Qt1I3yV50
ehza3/Qw7SAZyfLeAurkW0X9QgQgfriAbJe4KonjF4YoK6l+OIblTDjmVIezzRF0MhaQAbumFxqG
hYH4Lwm1LWbzPVPbVZRTw4+WmxViRpQ3AA/fyZCwqJr+kjSPHgEXSG4pHGro98ArGSLZmKeDGMni
khcwyT8UcshSq6q8PxgIl7xh+v3t+8EwL00IaQYByR7qja9kxdLbDzLaCeABvEZt6rtXSZwEUhDM
PT5REvrxLOrP3gSNsfqeFCoWweXR9oweex5NcN+NKjHaogoiEelqBCWN84h5uD9NHQdq2GhcUTvW
Kj2rzmjKk7KMa5U/xWEgordeWPnLsLtP+EkmsSUE8OAlQbrqb+T7F6VLBjYndyk8V2m8fFzpVFIg
otHEmJUa8jh7TfLTm30w9o/d0IMJxKSZEqE+Va4rKM4rBwm9XYhoRZYB/PDcpjiiaon3vm9aTHLX
t2boTB1N81i16V5yNroy9Wyhpak7BNlbCtP2FT0w4QG9k0Q+NtQrhS5Qa5Qj3v82fM+pVTvoAG/E
vdeUnLpDAQMS2K+6+lEIbs+HeqEc0FB6WZtjRbku8Dv00569c7TgUYtDLIhk5Dl230b7Zl2Bryfq
sNPx9dy8Wz/0jdO1AmDd/XRDB0bQNSczgl6ZYcqLdP2Q9kkAuJFkqjxSkm5vHHhkAnf9I+3KBO5g
Z+Wmi1UNek9hYtrroDKwY1+O1yiLtX5EQxaI1mEfIV9nDw1hlg7P4Eq5HrmbSCnl7zQnVoqULGsI
VSJrzzc2EF9JTTshSUBvK2tu3TWGm6IJHHhtLMYPUVkhH1XhE5Q8veK6KlzXiAwkNqMmGdNpVCHZ
niQ7Y9MQ6sg0P2V1ql40oJz0AvXeurIAcnF3/vSihfSNOEaIT/9JrKCsgY36LQpyT7Xc9Wk3X5o7
Ho8ODqZhT2dG9UY89eGIUp6mrIuHfkMq77flWU35Sj0+ShLQnj9QZQzswuaj+4xPafbJgWuHsLYT
XeF7Z7kf+SbHgOCZLAGGsirNNhQPxRg8IyP9tjsHolxlh7dBkLLeFoEhDWV0hMxtAE7Fe5MO+oht
OHhky1H4aYE3qeLr/vn0rsRQ62ciAiFEDyfgW6qNE6m1AAwhfB1qy8d+I+CZYZ2shODUKws/4uxr
G633rXCnprWHIb6+UQ8feE3iPB6umFzU4VR8uqkItDBW7hEmSYq32kcSQrc3YgwrO48PtGzpGAzB
XTBMK9vfM0yJIl9DLzIqFEfp9mkPXslnlptRbZ7w5+3zxtWk/Hm1E/OTq8/fg4aWpqsSQFY4WCM7
VZ6zhJ7bcOiJ5NB3YN8i6TYvKdr0Heq+Q9Son0fn4EOv6vPIxDhJVxoHcJ+QOiSb+WOop7LdyMaJ
oXbEGQzIq2ta1p3Z0SNJKS8rLBmw6lfllHPrY6LR5xbCmkrzxM+/KSiWKzsCUuT+vyoUS3NulZ3/
pKLeig2Pjv1twPDaD2fA2Nh/Ua5diUIoN2/JkFCzxg0ajnTkm4TjYorZBAGr/mqqHlMFSLFwnsBk
XOfBZAmpTapml0r1j7NlQ/96+OYD6a+vsbempPdjt/G7Z+VxlGF/Ls+Eae00IJ4ye04gB4kvVh4u
LxZBNLNJInjQaen90tu8sigfIH4FZYGDgoeRM4wl9RlQ9LzAOhRbR7UHPYsS2hKBGHVTCZW8d8mB
VwHvxENDFf6jcBlMSXYcJdHk/ABLemu5yPsmloNvgM2ANVobjs5J8OFJNquzVfNZLkxudT/RBt7w
wgdK69qkqNXSuf6R/ZCC4s6GdV+fZ9lMLeT17lXBZdOFuRfz5KILMx6i1qzc6WJ9HCXyBlB3QzNe
jsmLUI3xINlVg2P/qv/mA4wSR1P3mjkqA47ix5l6Z16F6M5pEi8TNmAsP96wVlLfyxq5cxztt6UG
1MYuc46n4ZX7BnX7VTI+W2WzWgGYg5yWYQfoeyjqBI6rplaNVgwevqxi4Ipqrvk9jAF68llGwjQU
Erm9t6m5uJ52ixASDP3B9xfPMC/27bxv6EpGpXOMm3+nu/96af+6YlDAM966AlDZz5t8ru8hnGs4
Vx9lTOkNpJs1sdXIbz73/fmxAFlFHgCmk3Qcu1g7BoInaV2vj/JqOqkoB9/buGxJzedyEdAvm3Td
foGhc85ffBeDvCDcb1JDWiId2YN4ixpeC4YAcAjvQRwpEnjUv+S2MvsQw5WkohYX/CXyIvCFl/Tg
Tfjj8jhKA7ByDX/cYhtFMXtn3HWoTurv9rSR8aG3r8rKtnXu3yJleVJxiwhWW9iCzL5xadbWwkzj
cMPOMvwvRWioJ4jHM7904AJ8HVVZBqNKoqnJEAP8lUReEj8YhAyiTe5gXjdpHkthaA4PXwnix7VQ
qYJhJ+y/PC12g5DU2dc60V+ijJq8w4kK4aWyIZy925GUBTYkrquS3CJMVvuIMFEv4+rqOCqYPiN8
rgnh9MTu4rrgsuM1kiUdYrrIv6uhs7Ao8m5bH9QFAKX15wB0quj74w63uGe5hMycMESyV8U4glUp
5YqNCT9+er0v7189GFf9L9pRbkCvgsqZbj4tstzyuEMzj74xQtykqyhiSlWb2bGmJrkn4Sd70wA8
UVd8A4iJpmEHZtC0G4YGgx/g9BPIHLacfdr/U8LHNKAO9huGdzH12UQ3JxZZWe7pdAE/9Z4EFcrx
fWERx9RsJVJoHBTgRH/J3Y3U+saCs3iFo/1FyU9Y9WSgH7gHYhEVNKOsGrF7LHeJDC9ledHTcveP
SQrOIDHMrlmrJjwWrTBcI0fCLjOv+FBEG6HFvsz8MjJNU9OpzhFA6dhNz26IPbryOGqnkzs0pKi/
MgzMsczCuxoHty7XFBPmnf6Rh19z5ACOxejxlcMeD/3LCF7uDzpjBkj5/Lj6pwDgSkjcrP9voIpr
zFirQkuzCocMlYA4wOMq6my6leZovMAErJW4RTdFRuPJuSei+GTaVhmaI5yvrOTETHUUZUm5v6S/
60AmkZZLSxRrOccvIONPdaNA7mN5qIsuPwrHu9dy+eVxBM9ZtTXTTjly+04/lXmLnDfQIDmWkjDV
DjTU7k7jSQdU2AvIn4xXNcwQ0QxOIybU2CO7KdBMgnZyR7QYRPQhZkPcVDLlT8f7ReY/5lGU+FFw
DFBh2Fjg+tl+kwGxBjmPG9vfuR4n/wT7eSSCAh9x+yqbW/j50+2euUzQjRCIO2/IKGORX5pJMLNg
UyMI14ebqoAnhajvjqf5AWIERoCKjvhfrR9/0W2CnARwIJSsKfQsCPyYsDvpu5g8zUSgf3hrQsQT
IOxxKPhaALTWldF7z0xfs2fwpXh6X5ph1QxoxFNbq8oLyMUTpG6czo+tcT3Wam5tkHsDXbmV9J7K
Sl1SIPOGLvKHth9NNNhWaCZHmYbBeyltLSEpFDwccNp5YBQPV6eIJH5xPSaKcW4pr/TrTtT/k9y6
LABMLZ9fs8bbaWGHcNGpAlpZxieQ9S4cBliBIJ+U3hbpDijymxyR3quydLfDGCG86OH8Mj3n1K7f
kXwDCsF8uQTMinmXc/9Lw87qNQMdbbTEYddHNCnpc1hCDBdrrn6uydUOx8Fcvk0igzBjvunZfqvN
OWOP5/1ASW8i/stXD+hhx6ZU6T78TgRst13olbjc5PyjylvCHCqoKyHfG+XD7JJRq2zjxPDW4Mf5
AX62xxzQfLsw3AmYx3CuLVx5RJ4243cyCni3C7E2837RQGxY0Kv3Bw3V+ofW2C4EyzrBUyCZgvzA
QqBWAJvlq9xulBfTy6AL4OZrFSHI9WLM8NkmPUNITcvOliQ+fepf89WpPutSvcM7RPbxJHWlE/Gk
sf70+RPKQUfRazKV128g1c/B04c6/DFdiV3ZgkBFT1bP1TxVJ6dXSpFAqoVXjgA/m9EX/AxRQLFs
zj8AutBT86rkJSvGnUFLGYbL+lXZFaULmBL+/jQXiSB9RC7YDSP2fdidrzFcsQFuliI6Tg2efpn9
7fVn6A9lghxxGqIlU70nDySxNRTKufB1MXPfj7fTsUNXDR576yxosR3yu9QjVHuUDguMT23MdvXz
aZfrd/duZG8/DrMTfvecWSUeYVLZrX9+mgM6rPdLhu8nPjfUbENADRfXG1IR8VWhb/el1tuGq7hw
7YCIZypfuYmA+MxNBDDkZIzhrGIIZF/s8ZAd07P7kbPkwW6OUsz/xgqNqYJBy9C1cYAAcgjo1Bp0
5SIS+Pb0ADJa51LsgAFZUvViu+esMJR+++oPRqu09Z+meCEJJDaxXZy4Qktg0fd8H/kqjdXr5k6U
gdACnkJnEmXLld7tRMY3kj4wc9TV5zzakM0lrRDsfv6sXLYgri+b2g3XfZAB6vAKV2DUwI2C7cGE
qCKxBg8qCCfH23XKuEUcKFKEPITpY46o3Q0dTWj+QTYBIhcwUczooxLgmVJCO1t2TNQvDMyRUl0r
N8/gkTZRNlHuW/RAO0BZ1SivE5UWai8QG1T5YagEn5nlcjU9ASWMKQ9x6hYcZyqM6i8J8FjWlgBw
15rwd76V5d2XmgA2cfNUUN4fAsa71YHCwk0/XEiYJfo0fGGkDX1V8rxuVBWMyb4QR+Ay/JN6H9MX
aNmCYSlhB9LMC/ZybkWSnzFcZ9zIXPtwyEST0mFW79eJiyGEOmnq/rTvdA6LanzlCQ2aN+ygdQ5u
4z0qMFEsFm0s58aev8lPbDdiikV3LgfU58rqSd7TIM6YHc/SgHDnsKbzMOK7ANjmGMEuWJn6ld62
kvAmfX2uW7WZGfZB0aWRt7nkSAH3hOVG2nzo4s59sniIebYGLyXRqg5Ear1IzYaYMFnuP8RZ7uF9
Ikg17fogs3ZVF+igDmFMZ63eiEy1d3WOJmpNhkBZveWHZyzauJSgmDu3Tb1+2a9DlkkvY0yc7ENK
XngaksiZi5AvsfoNW9E6Q2Q/e/Xd1UU9w+1g7v4dgBYIoiAyLoLubFcZ2+VgM0F/Z6IYe2O72Fbp
6bmOWhvw5PIk64QFfZTt5sNsubcLjY8oNXa1NKGdVCjyxTQU5zBNTZ+sKjAcqhKrqiy9/S/lGk+T
DlrZfLX3gyvYgxoMilUPJa42eMhTj1Rmgal9AnA+45f1YsDxMMSU1tZUfzcs+zZeA/xtgKu+CCIR
riYqeQteMEyATEeFUSfuw4kGyzCdjrvrhGKD6XbuEH1ZeQMdeEUuDw9/sxynCOrqdLyHZa6xixUn
vRE5vae9kVmReDMhRg0yEAgt7jjQtOgRpL3z6LbuACkkOUjfqIuspz+MsSIXqoWzsPvZQjAtaIM+
MF3zVHygJezqU6v/bU/4IKHy/5XOCcxpGv0+C5k3gfibJijqglSl91eSLUND/IO1TrXX3ODpXdO8
g0DG+f4czNPNE1zz+9n1jx/0bMorw5oFzn4byt9sgsBXnsC/kqT5xa3Ncdx7wXKo4JLqHCzCH2Nx
8XK5RyEdtIEO6pR4rhDA9q3lnZU1eEgXol0RV+4kyHQmz2wXvYlsAxFQoGY7rVnZkW8OnezY7bVI
AglG6EusYNrREPsatKqrg0ixMSCK+3OFDvbhZEnn+/3ToW7oJmYrdSX27Hu67Bh5+PLB28P2wcXy
hPOP1jkn0O4tQ5wzt+1lfvRKiozINR2oFzUg7jq4Z9pMTfrxkQKXrqatFJhiDpdb9zP3JexnPrdd
zF4iUAnoPcX45vrCE9kS7fMcjuGjBF7/BsLsLtGD3/LhOByfnX3rcigub/2fN+o7uzdL7E3lJ7Yx
aj/pKy63KdlLrISnt8pkyevIkvUpajWSui/s0c0MQRDQNNzfkvetwLeTL5KmU12Sabw7iGlyNS8R
NT3eYvRZK/87ZAHEVJ7r+O2CkoBJ3Ph5JM1FhPdJbWKEpb01Xjmx/IuRPpEwkKW9T071ker0ZHtJ
hyX+acjcHHA25ayl6YFQT77HujXVjoja+v/rSAN5RuC6RL3fPNw37dPvqLiWVoPxBYRnFNpCcBqd
DX9rZpBq8W3q3y0Rwxw4Ff/Po8hodH+s+Qac00bxBG2DLoU0486IIT29ylUhhMjazhkoo23YSYIm
21CpMoS+KR/53HRdBtxqXnjjA2jv7QyjZKSwneoH98AqLSHs/R2q4qqImQrdkIEJ8hZBloOMxXPF
t3v98AvHHsfethTUnIUbXxuFvMdzHShtECFgF3W7O8eKzwxTayns0hYYkxp7WbXDRLMx5W5Acwtr
8tSUNmGAXyzC4PM33jD7hqpmIlnC880nBSgRWYF0LfYCabXaozm8oCpGKL9nWoBuAB+QedCQ312y
qgrCi990JkTtRoqDrZB9T/J1J30++lMWcoJzfFzAGu13vO8CwBgtjbOv2vWtmi9CSl7UmaUN/EiZ
qSNSzNYR9qbXHPi0A06Ey1sZoUIcRFRjiJCKPT19U1aq6akNPUi7ID7f9RQNQnbDYpKy7cm3ukGZ
ion6B9dxLdsK6q52qllw6kuDIQYVQJCCmsmSoM8mh1JNQXesEBD5s5Dq0Mt7wy5xLYsKum7qK1yj
WF35iD8Iu9u4G8EVQtn7CM+X4N3gGfZRP96FF447elB5/xdtNtIfbRMU+fw0skNqa4YUGwqHlV7m
32kchEuMHs2mlOkhf9WNmnnUb3lpClxWPDs/6N6HnYukBtUBQXXarbKiMthkgsfQy701b4Y/ZIOo
TQu2ZmC2VScuZ9Ie+bxWOohdjkyjsVaPcpWKaO4YyyvPfj/g0DfU7Eq6Cov1n8UqojpkKAZNQP6q
heUBZqpH1pqm/V8C2gzMmCkFxEw/Sq8P7u+s5nmroI9EdFumiYLYQHflQe9k+0zHrur7eKQw+EwK
HUs6HsCt5+/PKJvXb4I35XpyM1l2/ZFfqvM4I8+7K/OIdYF6ATdwAnWGE4AjO9kEXTols/qeaP/3
avxLkYbpj0IYCOGgV43HclBrhjZ2bjv2pXIlSY4X2Xr3WpviB7QgnFXfP1oUWE5zjh4p0x4IGRhN
dfJtLeGTYB/WbRffOqS3KQilfVGST96YcDHvtoTYTmwQRPp+/lfg3ResiZrDynwFSaALtS6vMUc9
L6ZkumGLTdYAoiQXMuIZk6m87klsHrlPVc3C507RsKgWviZDbDhJCisKCC4e9mONQthDqzuKUltg
PUYxlDT6xY5ggQBW7UGZw477z4U62YUqnqMO6EgnlauYEX2r6WUvZN5230PMWhzJr7XLWByL1trw
mI0CtngpszhbAU9L2bpRl5Mn3AOsJoZ3GvYcT39Bflly7nrS5KjnwA1MH9AkTBU0CAw+aSTUzVeP
QMpPA8AtP86WV3dLfFA7u7G3L7sEc/QIVbZ9WEZPXHaQ1IRhmvfBqjUDeLB1TZlgGJOv3wMRSPQv
jeNCe28nuwNjKH+8Zsh/0GYs8K6OetcySNGXKQpa9kSQ3zVN1I7e0RyjYvW14c5g2useUsWLpcIA
bG4rQK0k93YhS9WVcIseD4badw7R5+iiLXd5ywBi0P4I6UvKqU2abX8WtUEMLRCURnoscQ12Fo+r
J8Py1iaZFlfGDf24usw5GGli/3lDPVekCf/vlWyix62FPy5iaZKlIDQy9P63o11MfEpKcUB9ZY3h
SDtkHcJR45j7ssEovDaoJGUqfDovkxy2HvkTrWYKdq41wtcLW6zcUcvE+LxafbiMSukJk7n5zurH
pAqFShpb+YRSwJL5npgUbqxjg6mnL6f2YTTM1ZvU0/GdN4K+ni4d2818H8pYbx5MTXeglaavQlv9
kHD7pC7N3DuoAgx8HwAizNDRr4JNYqIGyH25VPQ3iPcwZF+Xx7sGjBIRqjoLJY8Q8/SEj5NqtQNB
mbDfgu9MK4jvhhdX3ySjHRN4bMj59GI09ixhgLIjG34f6zDC+vAC7SRN3jnYlyp8FgeKfK4Q+r+O
7xzxHzv8bAXXPjjwGUcoJnMcTF3LnZMr7OZ42Oyy4GgX5qulee5K7Qfm3xzKQZqP8ig537bI1gqs
+bdfCWyo6eXGF+3a/J76csVDlQZRrYAdwPxvDqc3R7EcM9y2C6eK3J2qaDt5rAh5BcKKkPdbFaP8
QKyrXQjA+7IgUhWS8cEaLGlK6EDMpGq2mnqq3L3wUZc06JanvFsUf0HiiXO0ZhaUCloXwQA5WQeV
Y5vrw2EXi1hH6jr5hi2155H0+SQ1ZWka+3ikS7nQfBwwOLeAGiE0fW8xkelVIgIygfxb8NV/30yD
FYahTJYGAWMsBxA/vHlrP3x6jHfLv+SinoPKI771v1a8adgUHZhjCPxcNyGie0Xfj5X8Mb58OzSA
jqGMnlkoRCkXaJFMH7WSFNBg89uoEzOS8QJm009Q1X4LSbP+VVNOikJCPRx6y8fL9+ztKiVboY4/
6qOZQhGm4wdl2kCNJqBSrOsIqfaJVfeVNZsuKPBxb0kJoN76EVCu8GIImMrERjcBxwxAXMjYN7Vh
ElVPxSHoNh3KCpUH9OBXfrf4m9sRbja/svOjA//jEkUJOfc9m4IpXWD+Bh66z8QY5png3pjGW9HF
q0TZwTby4BHqqEpljs3iQzdLPxYSRW3pKN2LVwbNAsfXEAri5zOowZ7bHlgyx7IrlEdsY7TSfvF/
VYUuKID23My/rTqC+Hi81j7wsi75AZkOUGZVTbgEj6S7ev3gAXyYSmPNKxUX6QgGkgTfpYO9OHdf
n2CCMU9hPWKUWc7BMjXCZ7EY5npk//cCsiSIphKAYLRSEwVqdYmLkfLM3MfMsOREG7UM1Uyy9BRu
tJ3xpjbBzmLrVh8YvGBeRCJ02ivi+8xl3/C8DsyjF9btF7VnLmBj3n0+Xbo9GK/YAyTl4exoHOOr
+wEldLY7VgxiWe1N4g9zc5JOKWcybctnNHrctEm1lOvNBRVegxuVffuEf2RYc7N2YzQ8msJvAiKr
og4DfJK+cSpkLXHfI04KZeEo241KJvF3qRIHZA65uoh0M6O5lIdyqlxjvrNeozgmyVsT2jIO5VYu
k2xT9oHlPu/VH+DJfTyDxQ2jrKyCqa9t/xx4fMHO/8TuEQkq1sfrobTwTgsALkTsgEIDG8SidGnj
Dgwr4EzGKDH7LTv1Lw/hC7ndeDnD4oM8F95dGGo3V6UqZlHPbSSEOj7oKjbgAxV+UzEnSUDDRdht
YMboBSDtRzu5ClWjfW3biyJmTYsuQlddTw/wD23jT7K/QrJTOjC9J06SiIvW2bePVeuFRGAe5d8x
bN7WOIlQF6JZbuOFZGFaiOJud8JfqOy/zbYLiOfmib8McVrb3V5nONZ6kgFiinql6w5J03LFBrBv
SPsJusGrMkLOQa5Juja9quBNU1m+bMuA5TjVeSDR6ZuNhRupMwWPKroRdJkt/ecYStqW1b97yaKE
4SpiQ9Z6+/qV5e4hLupycIPCjLCljJ+VijzTIoZiSGjiyDGM6VV0UZVLm3DiohbNyXN0UhHD3Fs1
dD7BRPO0EjAcqixH0QLpf3xF3/rIz1JTORfkfP+cCWKZ8MPc5jBtrgL/chnbddbTz03dX5DdUjH6
3vjq/cyL8lX2/vRjrDxhKMRBRdCNcVW9IOqAvWykoKD+V86cbDXcVLgfNZFGFGVOTy4C++GkbFK1
ZjuPOAQBvRHV8LzoIsv2l3cjFhmxCUXgr/vzR9f7jaFwG0WWA40haGBWh7gIzGJr9SNTloslRTWE
HTKzw4VGkKvwB9nqZx5iWI+dC4zEkKzqlm3n0D7a1VhYBvVs8F8s5BmvHxihAxiXNhG3N3z7rzzO
UmTvFJBwKU3GWmEtTcyXNj6qBsf+5L6t43wRNLfqj1+Z+098ORm/I45t2hSIaY40r+dzuxCLUiYk
omS0juBYaUdwmmR1+nJ7mUEXknZtgFizwqZ8OgHXMA8trPO69+HH+NTi8oJ+ezxxM3Jk5RNNNZ28
IcPz7Tz4LdJCVOOpJh5Fcq1X9F9HleQ/pgNu8BcpqO4TbBEiz3cv4acWGB93jR3UsB+AuF5HsMhL
6KQ34bDjU2EI2+ztSagwuSGc7N62qeJ3N4dRj4BZnozrRE7bYi2a0ELZbmzdhaOviUaRCgxwunS1
oN9lQ5+ZPfnUvYEqElfNZwwzpKSZno4uYNPL16RJctQYPKx5uu2tepPl2dt22suvBuT0nfTyQVcA
mHop3/CxHIOe3PCPQq2J/gcJrNfCJ5np70iWHcLgcHIlz6po7CH/coY8FCBt3gw9qyqTxjG1nYwm
A9PLMMYHTCUI9S+PnJDOeThvbfl80vc0y82AYRjPzQ7ak+vkS4MA/4JF4OvljnmyiyOkxadoA3KZ
jyioLGG7O8KX6PDR1Phrxj1bN00r8t22Nasy+r6QH51GchTrBysFYWIB/hJhvGB8Lso0/srtbcLY
bBaE86cyQIa6gcnurdBqrJ21n97JltG7Qb/QJXjZ2tqcG9OCCd6DnjG5+tGM4kCfbVqMyTL/aVMf
mMbHrnADvGyVbJfcjK6qBLDvKFu+2SjlxE2BZEWHBBRtM+OYGkqEK6onub1JFRsAO5LUaRDzkXGg
N4+mKbQVJJI83Bx5iGCb1K7EwGpLtLyDws63UgLtxt+RUYIfdtTe5FUBmSR1SK+Q9BBjByWCpSgr
kXBWXm4DRo//+LoDgELIszv6XDVq5eILUNRczRxZznSAhW/plp2q/YTVjwObIu5ovmOVUU+2V9Yn
FFhcwn7fmD6EHWn1x7OpizM4dK0QwUX2kqksSDtqmVT3gAUOwVTjFISfJc3DcjSiBZQMTumK/7Vk
RoT8Q9TvQFtiRj16Pw9EL5ci1A70dUMXIhWGsMzn0Be7LZqR5G3cLR7esxaq/Rb6YztWsch4bkPd
AlOG/pV2yixrxnmIO8nugw91rJsTnCTR1uSnzclYJvSZgDZUzort7tr60X8HER7fUSHLggadij+1
TruS0Ciqg8ukgwKOXnKbHGL8ZtiWdL9/9SOeISZy97eJ5B1cG5OOM0A9/HwX6G7OJ+BMQZyIzQEs
yUZ2bkMlLNn4N/2uWKfipI2oUV/TODbZTy3G3WsgxB70WFwcUcuZmFDEwsajrgJWqEx8DPlgR+wO
RHKbsTE5vz/MYAsF4gngfShVuVPYUkthnGYed76TungkjtYPNqPhpjvG9l8KAk1nfFro0MjKxWRO
WLsr9FfspfuI9O9kMNJJ0tnCCm6NmcXmCjwAtZTar59oZVBn5Z09HFlON28FJ3qzcRT+Dxjlk8ta
eBW8ptHYjxKrZMYPFLnHv13tQeJ14bwQxUT3rug/BZbIS3ESk5ALC9DsBa9SAs9MNcUob2cYgOIw
2+kzmD8UHIQFyH5Pu3/eIECz5pvDkQXBYeBl1B3lq1Im15z5sYwvJOe9hnKb+poYI31alDjBI5Sb
PJV/dImlIMLg4+X17lKveUVkX8s3qI6SWJ8cfjm9lxYmiJOe6iNkzUSVs+1hgwaM5RjmuUM1AHV0
MjrCnvHrDkOvVz0+AKtWn0eDsRxwK3WwdSRf4HO0gMFkDY3BiEFOb7yE1dn6H0ouu7PSjR+E3QVS
me9C5wnNCEfncS8ZbnJVtMMALQW2bXPSviECHpAVfx6QDLSJ5CUGiTICrdGuA9i8g/o8YsOoRLuj
PzyvJ6IsKNFq2YG1lcc1blhEDg6xDHrlOkksxTPTeGcaA7henxKnT8VAOOQlTO4jlrhUkY5rSJE2
BDf4WRes8tEUFzZjGYSmCC0DxjSL/PhyZdMpM6zNgbIXINdW0UXa0ggfGdIJ3DI2bsEV9eWBQd2G
lLf9hw0GxzMNakZvwjD6puxGQHpEH44LS3n3GdqBNwGFb5YcU6cQ52PM50WJaEnaq9MaS2uAaCIU
DAh5BUdnMQucR6B932RbY+j86E0hDLKtWA0lg1QlJYPQ+K/EJu4KtBdVfM8IXtGUjyyLS8JfBt6c
WzNkqgEYjKdWANd3KLyUBEGDjZvHezdb3/JNUSpiL0oDlRM4n9HZ0+eCYy+YwZ733giBubuZV4Nn
/rh+w+tGwnI9CMe5x4eBbkozsaNLzuEqppjn9MFpXEvxSl4IzYP7273hawH3JLpn9BHVpiaKsmYV
annNzkXHyOcaKIAO1SJRtpohhpp4VEwVpuh+IbIah1zalRxwbxTgWidDccxG+2zpoG48HGJ9l3Ti
xNr/jW6o1UfBRDapu4VyqG6gVlXA5SditP1kD/Rk8YybxsvYwdo6OEwXmOvAbvUMUvJi05IWS3ri
Lr0HPM7VLn7KtcfMlkLLWRuYbUReIUHG4e51eb5RBrruz/QNc9Gf9nM+xGzknGUh+GI9zUlIDbmx
9P/ImRAsH0fMZ5xM//VJU0MpuVn+AzgCcJx6rb2RuPaWXOpsPSwuDEModx9/W3JRDELlajFes9hA
kcZC6ox9MhrEQWAoM6Hz9NBGb/kqMyTq2D9kG5wBN315kOnU26aBn0SUamlB8MF7CDmBLSOMckLz
0MeVHjVTqoqFuXfx85opBn6+MHkqrYhb6ZC377VIjiJb4ICUYkwo1ysPnwBSrw2gKkDZrU2EsWEK
iRVJuUrASkycY//tPSdso5fgm9jJBko1xVIdwGjtW6Y1/U//1cFbBMpCPG8t6Qnc3rh/v68aFeG7
heoEIH6Eu0gnVVKPqnDvaCzYaQ/qi+rboeS20KestD5EMHDOgYnABwzXKTc+M14ytoNefkuVNP9e
xhs4jbhTWhjDikVkG/06ZbOmN/3AvXCGHJvrli5u5M+nQJj4yMdUufU9ObgpOnV3BBCKNW/2qC4c
f/IFzFNCZP63SAOmutPN6ZoYrG9AI/oWi3Tzda8NIJBn4pv7LfV9ogO+45+WvvYkFOVdmeiQ/6QR
CmjON06+dfESDnkDY/gOgEfH2xzca/bymRst7XXkB4zfGgYQIEZKvZOuYNvl7PnL3fOUqTPCAZ/P
7DD+j1RvQUeDk93H93HbUZYY+ag1KUadypOf1tE1nKRWs7ernD48PByet7ZGIW1a8jeHxdzQZvVt
qO2atTaPu8Pgg0OMk2kY7GVoUv1AgNsFhB85VKrjYhXtUUAs4+IAyM69TyFi/fu0JiZWMdO0H7fm
+Gx1jQYwk/SVcQSOoiDGA3wWYY/fN9OJUtJ3e5MaG3k3Dq42Wv4eMjT1Dcy/jFX63giNm1ytAlKs
ViyBgM1DNHwm6bhJGHWUGULGwCkN7ROlHRWDlUjmmaDSloZl2gLEtBjvqLBpfK+L8YNZI2hbz4rS
HmVb8Z6xLyAthQiKqFy3selIc2QUC8Hf2sg67pE9KYyx0ZGVBcM2F+I9Id/01YnmHsharmxK7Zlz
9W1BDJoPZ5dqWf/W6PMbbYd4k8nDxUJcVm7umvhYqJcoSM4sI+O/SrJJ8XPIDYvNtP0kp2n4Pgml
yiWzztuVc/oe/hFjcscpB4JPOTcqrjwFaclGD+skRSOKhqSJb0bLEYeSOLtVPp0/0QMmvBx+vq+Y
NvlATjwrL4bTuGFxD7QtTzMdfb/S3Va+IRrLnNcrQOqq1E6gYzxW0ngY3egjqhSEazYiGjeKeiik
wsuA55CfKa+HB9GPYAEfLrKyPQ4lIL52Muc4Lu7fpgRf1GQ1zZ2w3uqdbcDfN25rV3UlUQyuSPIA
OifVlecyIjV0LirdNa0SwhpAqBdhDXA5AV2DcMYAIyIyUwaVWwGAEDhH7AHoJ/q8yjkt7FZWZfDQ
x33n8EcLAYTkCBP/vsJUL3tp+noc52aIR3ykBibCBS0A+b2bhq5vHqUvXjlRbH68tz8OKU3ybRpH
BwJh+FvH3zonxC8Agy6ii/hDWVjPDISDOn/N6Fb14G5gFAarUnxl35MWhEJ9aqaQWQ5RPCuGkXi5
r+a6kxJCqnT+E8JO6rb1vnb8eyMB0UUMrfOiMNe8zJlw/GpzOi7A1EBCQnrZQ6Lr+e4iAASZhQVI
tLA96McQbH3DhAB1+usJKxpZSyKaN8XEpQ4kAcaqjhUpxw7H3BvhWQM8fy0XjZ9FIelO8CuS7/V/
cMD9L+ixilm0oKxw2tRWbAEJyHkBmfpbh7wpAxSSKcN6kxYhZkY1mOYL0KIvBqr0YU3CueowXnbH
AAu3FV+KkAJdmLjzXepwFO4po1ghxEFC0oiqTrvKMG6z7jPlHLFyFjixgnEXjrQzjQ0jr3kDsOQB
xDP2YsZ+rgLF0/3IvWfporHmY8qHALBYlXC2+6oQmXKJ/xGbAvQn1wxQhW3ywdBfZh4596qJ5I3Q
au+D0+ilxMLJqAHfKlgRiracwRkNCpJ4OmIwzimv3O8Ytr84onOxSNEUyWgb+P7l+nKS4R2fYUED
csAwM5pCU4lr5l+Kji7PnvR4cFu98uPQO+HVvqlaDFmJoYu3E7on3JHlWj1PXUF5Wkym+t3J1IuF
5h97IdFhMQp0wo8Rf0eX5O4pJbIN9FNUPDrj3eXWerBFFa7A6fM7tQleMnKxfnqbhU2mxylxyyhW
z6A4UrF5iPc5B+3bqCdl03CZcCH7BWhjRpmemUTKYh2UMpJQyWaX+3fpCLMN+RB0B0tZY/2Q5cBh
gswTbcK+bIYI9QTObNFyVnuRJI4Ww+WS2zYz1Bjsk/cqDQtycUbaoRyBYMkJmuvVFgveoJHSPW7i
GoKE4/M8XM6qiPCyRNMP8SOSpm30xVd8wokzRdu4KvW+zfLwCB95yz453hT2ezkXXS0deR/mw74z
JfHDa5yYv7hal/sdyo7wh8tre0UHgFy4VoZhX/KNWMl8Ot6FMzMzR8+HJ4vgakOkfm78IjRFOwEs
SRe2jznutMCrzkMJoxDi/S6ym2Qa/qNL9TUFKNBBh1nQ460Zo6VuekqcZTwMTMkutrm7cXl9D/T2
rCf2XrlvX8iISEi2h9WI5oRyYX2hSyf/HoWVTnxDEjjNDogg71DYdciJ7apneZl5RnQfv/8E664k
VlWvaI0KU8xxhCx1vlQl2Nxr5si+n4n/F7cBuDe+P4xUW64omVOcylw2HNkEpMlba8KJ0Dmm5h3b
bKt+SqF9fxLP8ohnfS9xtAaxycBiW74B0epzAtWnA2OdbafhH4pJ81Jpr0av6vfHkCjSDzJtq69u
rP7vP48jygByrW7uzEQMcRO9z2YT7cE+LntenpzPCod7Srk0nTFQ99/glJMh4ygSA1fSY7yb5AsJ
wFlYqdzlYEjHj3F2w9FVNB/R2qJr8FAE2p76fdPtcHyzCtW0IBD1kjfQ7yDEzyCyfnZGJGqEs3dt
dPQM8wjO12LyGoI3+ExIXXeaRqf1tHsRaxaKyO9tzQBK3WSlk98FKNKlBtcuk6aPa2mmJhM8nkT5
siaF0X+ReG+WWnGQ54v/4mNTXhAIQcT0A8jjepkycb0cLPQcf7CiNyzsZdEIXBGvr9Zr13FIw2yc
7yLbWgM1GVX88ISKBCRLs0phnA5wdi5mXoiFL5xJ6ZYvpsUJCGrRM0x537bSsxAx17PJP8uiF5Ja
FfJ3fHkygSNpHQg3j9qw6diI1yZgJQo05Ash7T6J0iICtxnVFZSttbzMThYhMtQvOh2YW3Rifesx
nsErSXYiQ15LYBntAcXKEYm0CIe1VYFYdPdwre6M8roIv9Z3vHlIlbOFLkjgX5wlWLxxjP/mBKkD
xpjyaCLAOxMa2nPjIJo7n9oDXs6VWgGNfBlwrrzAl37bhm/gks+4mC9KpCNuEzqtjTQ+AVdnalsV
Fp+ERTv+2HVhWxA8XmdaprnKEWF3f5XfYCnKcE2Zrbf/KDiFesTQnZl9R/Tcank1VkvnFr6Deyij
/ke09cdF+dZ780sVhvTpoZq0/Yzdb6KOHcrsjiSOGDzUQdQiGLPwyMxPolx8Xj1o7/2ik8t+n1S0
966sm1bnx2/7XN8bp0+6RqFVJ/ShsiO9FuxNneupLEKsKVY4meqNULmBuw7OIRL3zFG0qCUyy9fk
O+zZmHZKxmbhCyu4dAXFrjrxjA15xfcWgwjXilUDCtaHE1yQbQx3r07LYbsE17KuV+oUM3EVx76L
dDD/kWEc7DtVUG2sfglXkLZ7Jfmm1Q/JjAR7HmOt1YRaN422htD3iuKOwtRx0nGnVVFTVTlnJ6Gv
U0Ch8llMzzE0shb+NcXP7JtOEQJPRPr6rI+4RqLZOK2jdalow8PhKKEW4hmaDAFAYmG6Glm+bLOy
QEhm1W2otaa1nBCQMt8w9RpHqTI1UMdm60Vr0cmbx5MVu3SkHRTgBXvbwopTJk0T7lESKb7i0kIK
Y7Vtptr6wgKLG8M5NfIDBQd8wNt3kaK2fGXeKCs50tNBeJVPA92qvWsdIz9+aJ64HOjRQ8VXsDpU
1V1gIKd7SCKUtbqKgaEqzcWHH97duI84jyldbBg0qIoodBZ/7F/Kd6dr1xT/6y2TCZ2j+Bbvcum2
PEF8WNKU6uVHH6I4/NufqtfpQX+WqNHbRqtsAoWR45BfWMJt/m9W+Qko3kNEz994Pk+Dp6axWTaR
qippe8DJ6pqO2hy3Ec4DXi3L248aXTyTjLXbSL3nwWyMD2mAeJYjW51fpfgJszR4r6AUZMyZw6Za
atC5bSS1IbopMpAuxGcAXEpeoNC11dqrhRYr8tsm40pjyMJ4N/wAHpl+2oMHLkH2q8qRmVWeNzFy
Bi3gceyUz51US7okNXQo9BMjbOdUgU2MszxT4ZYL5eabHnFPdVjkmiJBdzY29G4NupfIL8m+Dn6B
P6LTDmAyii9AQsuoxr38nG6AMENZcEDeOTu3BEz8Zr1ndCmXqZqBuRkycgdMX9511fqlw0dqSbe+
YIwCxk41FAXnoWPpGfnN1sZP4TbNhxdBGd3CDmkdu8fSfM57ruuZGOWb/6Jv5MdgxopMjFeTJzgD
M1ujsW4lzon5POyosvBV7Vlje7KHmtriXRHMDfkUDviPtngtyGC73ZUVjfo+BwH7tsXOuGPvPKDO
X7BRl4IEXrBYnpY4Bj1CluRcq2xnwnkUHkghc/XWbbTpBznsdjKMdICDhR2Ln3guCo8+euSpJKym
6mEqDNDJAfiRiMzCtqRRgeNE1DTmEmGP6vY3dM3Mh7z6XMWhJsn0xWtiN2+2cmv5K5zAGcrXeDhw
qxx+GUhEm2SBk4kEvAlmvFVBkkSzNouUBpL0i02GTdSnc73TkK5aXEdoO5WOJdB0fGYx9f3Q3Dir
uGOFzq8PZgUDLPHeqSB6OjKRPBoqA+nDjh1urXSvuqaUf3bFQPQRjJOs9bPba3E9nKKSt7qSHSVx
dFgm3ZPCeKUodnuprgvG5gSy2EkhG5MfKmU2JE0rJrrK4WvNiqkbLTA3eNgxxONANRScJ8WJ2ppK
9g+njpMZWgqggQAtTbJ52l3YGS0vTDNki0Od2WM7UoPWQoUzjGg0un3tyaQwL8HLtE2I1AOtWgG1
maslcTejgrN1udxCX02XnSSQnGCykq+iupPuulayDM3wCzg+oCiAfPCrHEnU/5OOl0hxg8domLE4
yjYMMySJut4irDPS+Ffe1lxKjpdBKtR3DsITqlL3NGgm7X9fVKYeaYVcncZWjXJRAmQdSrY3PTBs
yQ/yQ9MRldpJ5cnxg8RkzTkP9lFYfqVetnz1tJjhXCjUJdBMZ6zVnaXmoxbLo8VMaGPsvD4CDQ54
0NMMAHPsjAeFKvhQNG5/2sz+x2UzhuwsGCEvP6HV+k8QTFZxvircVX6yI3pa2BUQFKEPy3VYUljO
UkGCqf2qTq5FJ5RN4gQg0RfGbiiGmdI1tqicFjGG43C7uj5S5GQtD/ovh32KXP9k7L5pOw6jTv+Y
ghIuiB3hD/4pY3IMZcKrNy/1NgyC7KjElTP6FC5mn58K+iYU4IKzlz5HrZbK2irwZYwDJMnweqtF
8SeGKwNRE//Yd9UX27c4uuWRXX2QOfB/BLMNTjqnm7D12wKYAwKQnPhfoyp48HAVzVbz6I1sTuay
wMRMkiRsTM+LOIorRGvbHx1wdNTagMFJ6YIuauP4RjOOF83fKxBdho3twH0qFiulv5ArCsG7JiGo
Xw4CMi8I3cITewUlhet9nu6lxcVwuIis1nnMDZ6tXhoc28j+s4sXWprW5CqrZ3wMaCKHV7GF9cVO
sPPyTZb+tcDvCDD4hCJ5BWaUvRRFNPkgOxlci4M9/Fq+zQ8Suh7ZbKSfu3va6ctrQj/J9VU1aBp7
tPeRejk7Ca3uQsvHCOtTrXjpOT1gAaKGtDKQqsjOyJXOY/QXBGVLkq947JWtUL9x5ZLdxoTtVR57
Tb0+YIw4XoBuE6rrNv0pz6vZ0KWhxcarWCzd0x8PxH/QUCF9RhEWfd8RGfIMSy+iZ5JHWF6y4Rgv
dorS8iUiU7Ki26F/Z4I0Uhz9QdU0pXX/cGFyVkxrCWuUCTdjE0giztzedcDgMHkBHSxh+IlHJQ9w
+/NZujPdj0AGXPJK+tgVONDxCaJYjLPyh5agGTEgSrzliHOIdY4m3ZB51XU+hbH0SFTX6vQhhVBG
fXApWIrzsmSuJnePVCzt2bB1Qz4ZZ/Z8aHqZUqD6mVfkvcjWGOPLl062iHpOa0zWGT0DxDy0aO0Q
cZgpAAhQ1fxvalUlFi5hUeUcsd5REGfs1Dsfa/2FNPcQ06nN/SwQgtcjtKo0iM9h86EBBUc20PJx
pDUIs1mlj8Drd1ZMk11VGINPFYlzURT1H3ObhVGKXJViHQ2Zv7ucSGqJ4epBU0IRu6OFxE6aM+xK
OS0+mZD8BB8FX41ow6e2HtqT2tTBozOHU3QbLchiXBAjc1bYj4LO/1+1OcUGZQApKg4KraLy1Vdt
Zq27M1sLXyc74dVapu8S1TF6nhTggcNre/YlLWsuE9ro068O3Vp/ZnPy5HFbl/H2hjlLDhEW4dx6
41XzqXBAN2xvZE9yUZ3i51gY79fW6jEinvpbWyAQHkeqita0wijvK3pe98/MjfajniH3tjxq7Ib7
1U/ZeDX6T5/bs9Rk7yf+axWjGfwI0zqTYr9P3Hxw9ygeDcqzzDgn6ipAVzDJzyWMmb+QCxKvflBz
o03mUG1eNT/NnKM0OHBZJOlmVrB6QN5lX/EMxfC6wr5HU1kQ1ZzJRCfTL7d4xD8PbVupOcCKTOlH
vUsRCwJKeU7ri3dSd7aroQHkCmPgxCBeECj37W4cURzMbCe5rqmcukxn6KRr93y1MXVH9AwmL2a+
quiOaFiWRw8UXPp1iqpHvVA8BUTmp8XUUyK5jCo+FRIijwaQk2BskagK3FiKICFpba6MjrphA2/D
OwMqR6zUEN+uAgnTX7sKk/0bx80JHNj3KzKEDDqEF2VQDDtwZ2+I1luOKiA7wXYbc22N/Ard4VC/
FA3wZ7OcmHwY38x8tE8MnRJFG1VZAsTbzgJkn3JbjHknZCbysilgOnSs74yveBa99JbVjH8dpotf
E75yqro8LhTR1TvOWk7Rwx68Q5nxt1oWjBJhcJMk13tDoppoplaeuogTk4fFbjO0+O7HnmtbBmaW
ELiRxlWlUnjhgUFerpiAsKkgWSRHF60TS5kKTbFqjpfAAByQL/am2b6aGIm33GIAJJ2Qak4D5FCV
Ac9+ipZyyp2NGwwCyMghAO5U5SOJTCJG2iyrjAvK5s2yD8qxqbAsvGBkexMVAM45f9nHitRbAWGR
d4WjpLtHTxHkFVhZJy90M+k3El2EzE2GcwoPcrx1R9eDVq06QpK+52sCYGrX031UMFe1hF1GRbCU
AQAgzHijSLfW5FflAr0s7NS/BAsTHklGKs1pjKhIsffp+J1e89crq306HjBkTl7vKWuBRCs5DQxk
JPbJEVPzgJFfOi6eJ4S1Oah+Dg6HwY3LS+Jg4XdpjE9LTyExuZw7MSQ0JStIzDG28xsjLHpBlX3N
KNrEGkE42FUeWii0bVFZWfFR2VYLpzxUwpVndRYfDhib0pQCuxji3yRqaK8oooht2wA+4D6xNGWy
vyM0jsbjdsZzigztpFAaRyZlilbfCO7T1MmNNd0ywpIlBZ+5Qih/coWiSQCzNj2fTEGBnYus4EpM
VvVzvVY6f2yYru3LrtJhu9S5oxizPhLjG/DQJZBk30o410yb8oD1EtJsnGYq6HM2H7jJ/dEVXNhE
xd8F8IqVCoMAi7jE7b3nmbSIptpbVwS/Nt2/ucq/maZiTZgmRUrT9hHI804EEuWEz5kzVTqH72ye
mlVSjUyHrdE/VM4Z+gIpBZuU1H9WLbAOWk/LGYn8XRIjyV5CCo03ip3Y48lZ+6e+EL/fJ4IX8HK/
YNne8SW+ph5pxOBIRxJYB0UQaGOXa4rNnPgRdE7VrnGNq4CPIuWS0x0A2tfqqF9gc1S9Th3/z54w
9/L+V4GKzweQoxsRPY8sVqKOB8AUGxGU+P+xrnSSIzNik5jXN7JbcxMZMKXa30li5KuqmA6gW99S
E4Kvf/Zo9DhxHYizMZ6Ln9tb1POpaowKPRKIM0a14+crtDFXjvtT5r/kvLPi1Ooy9eLBYIxPwX2K
V2IXvKgQ6ELWiN40BKmXRZzNijwgzeGBTDzEvA2sEZuCkJyn8HDus/C4kV2Xz8G1hIbHSpuLd9Fg
+dJzNbee0197iki+NDPDFbU9TPVYhhuqtTBGq65rgAsiPq9fBhdwrEjfjOje7/gNz0PlECDZs//Z
ULbFwALKXOiypUtQJ+r/aVJJUsk20jmPq0kKKM3vqMHtOsn/aJYFtjsD6bowkZiftb8QMAA5+IRx
cOmeyTPmOx/IyPnIHDW7UN1vsyKxc7mZj9b/TCzIhFNvQ7Yzgg2Ux+ffQpxZN5i+IxisfJWsS0v2
EorxjWMwOIXJyje8BLGX1rZN32/yLYXYesOY5EKtUKlP277T6AnaTGvSMJFCjRH3tWC0fS3DPvE8
tG/irsgQQhN1le9nczGwjYHf107GriUy3anowqsdicy6VPTxvPIudrF4HRE2EZC1HMVYmxnVI4vu
7eYB2ZANUOSIcAycKYxSURQMNkz4LyLjuWJPJ9+98OvPhX44dFiVsH9UDfd7QzrLWcEGPgwyDnEB
8QeKTTusMuBK45o/N+fcMzrr7suoMkVe17BxvbkT2DwnEhFhIx3aUERZmKFtVgwEWrmHl2v6fkLR
4wNP5Te+0XAHEUOmsRJhBLPwci8Sia14tqY2cO91mPoazzuox/hdEPt+5bS+pTqjz63NfoWdaVWs
qq8H/cQAOLcVIBM0PDCuykG5SCluU8yl0KB5uJyc1wVtyWZTwk/4MhdvDTrt3w7NfKi84tlHPcYl
ea9xML+l88NkaYxHmIzm90aoTu6OtoCiMu+r9N4GRJGaJMk3oetzdSIDqPZ766HaT1CiKTpn4lww
4sYLXyjkn8H/EkEL05PoWDUv+sTaPNPuaMf7O8rk8XnyR2SvO9l7QTzOvrB5vgK8vE/HPV4wCI7W
FBbHoog5OD8vneJUnghEpRhMW3whiBLLOXWd7AAk+LPiYcw5AOBJHU9EiNPRW9POXXaM4jLcb/Gm
XSaXSA/S3t3Tin87pIzTsk3HnmR127Sxl0TdggcOFMn1fVt4tIhXPGhTl23hQJzaI8xnG60yj14f
l/RFiAKHvBWc4kWf7GQL+fJdOmeftFGU5Wo4dPvXImrXStNjeTQohUxopaButpa7hhHopNxyKb42
1oH2GC3aInZOwB3nFsJCz85foLKG9r+ooXDZ0r0ISLl8pFg8OT9mPsU0NU02ZKpvZZgFJ5+ZBMwk
amUGYosf+MxIaunmXOdX5zOH+B9hUG9k+DKHfKgNi/7tWOaZv9NXDZGktuxEz4PQYihvtTv6EaPp
nGv2mjjAI/cTPRsYZ4U+g0ZImBbqAzrvKXzXaQrxkyVDeYKJgg+L3LHo7jIZF9bCRhPf49rfZ0dE
fF2kb2KYu+ZtJge7OBgdq4akpWaUidI0+6vj0hyN8jNr4oQMWFtkX7mq9P60jWA4AYCFBfcbC3Aj
u8sFf4z5/K3mmGVxHZZC5fOxcamlb8Vv5OcdX2nNWdH8vnu+gLGvhp079C34tWnQv+MKrlGNgbUH
63pTXakjFGyNRxdwrB2uhHioeofAg0KBOi+kTy+qx7VDb8VRagsIBwP5eixCoZEtEb95FhWCe5AU
u5m49vx0A/Ua7y0Ypvlr5mNobLzOLZnPp2dhXAeUzYJDgLHqXluJjyXwTmidqxiT47279IBIvKSo
82Sv3HT9RlOfYKndZZ8hAq9GFWxVBGwJ/emp3hgcdL/BgexJiPPnVVnyvJJ2Rb+c8GJtnVTNnMUS
HFagyUgdkAXUWCSqSpzwzEPkww27Ay4ibfXvs9OOEx4E8ECt7WziMuSBa95jGkINGW18C0vf0oFD
3+Zws3gNPy5VGuGtbnYFP8063Gkc5zAvXI+RbnmwxIdXacyuwmpI8pwrJOw4cb6x3W5D6mN11eLd
/s+YGhwgTsN7l2Wc3TN3WXaJYob2Tn3sHepRPVTCEGC7Bq9VZJp1wkLSBBTygU7J4kLWRKbiRSfY
tglZoWLHfo02DCMBYqqIQFi8mlymMrhE1TClLh2AZgPlQKCCJfHFiM/a4AQPwmwi0j4ImbaKcD4a
VU5QO6ntnm9UrLAPYtspeH9fN8AzqosMqjtecGa6s5q0dIN/2pd5vM2Fr8Mc9qakcQTsz2LidYXx
jTNQdZaiWovq4v9MHWwL4Dx056qHhwl4Wgv5EjvbZZS8gSfRqQBRHOK6NvD1aBFAafGgsitJqo7b
WvQ8pdS0s1BBHqlSkCWtan7puPD8LTm55y9ies0dhAxw0FMsQBtDXuki1BSDxdCxz0n5DfUNtCN5
7U0vx97+iZqXam97WQ+Z76DEiJwELuVIl/qcaY5S+3FY91dbxt9CQPzuRHQ/dy98raqebmoOy1qI
l7Mk68RXtdz2ECfsOGC/FZH95z12YarOgXCI6gtUCatWnceqD8FVvCsQrvUAUeEsx2qaR43UGU/b
4N2CpRTyoxBZYYgHh86ESHcRQhXBIW72RosKEp4bWWEzpgjpKWkPySsgAWYBb8nUMYoG07NNgwCS
ujD3LIfvHkFXIq0FbyeihC4EP2a2im6LXxGdPcGpdWfBBY8ZASxI6g+pZ4accAejJqTgfvaynfIT
y7aM2d58z8VK0ANNPSBugHhPnHczKsZEI4Mpol1ghZ8EsQRcG0Y7Fk1p8InWvvM7o7JtQ2mD2xU8
2/8zyjR126Ury4PU4NMtzIm7vDTdTvI5O5yNNCi6deXtaGBCUaAhETweHYEusUnGQgu2t+vMXi0d
NgxKyPmJN/Mpt8FBLDl7nOoIE1StZZLgxGkZOJns5w1C4Y4q+2I+JPp4hvnp8jZq3beXcbPYOVt8
ofRQWYjZGJB0itBiTEPQQlAfiLHCkzXgO4bHfTKmAJvncSzWmq1isON9WZ7hGgKYbOcjxIzzzxk6
iMTJ8KhAN8FKXijy802rRbpMoLaf123xhdyXvkrqv7u3kOei8COEFPl5MQrfJHg6NuRQJn6brsyu
jSlxyGjEiMHvPl2HBnwlDRfvYiuG3X53P5JK1Hqw0ZcRhZmTLBgz9rAFjA4G48WT7IXZjQLNdXqI
7rS4gyHkjWVN6CMbH7bs2w+rpE4lIzuGO4qU+psYinMLWSaSwXTf8wx8ARfl5vzhhhVnbjocOQK3
EAl1BDc9bgYnL/9ajzMBmDNvzTN5aFErJ4asGCBLhFGLIBLGonJW/thjYjfTzJTgmUy68+6cjc5R
Vm5DupAa5zx/IbCY9UL6eqw2KG7FQ0ddnmtzffmZW+eiZ5yXroiQQqFZGIGWkzgkfXzL6OZsO548
bcoVKTimDvclCUt6dGvzc0MSFV7rQ6MK+BSaQifNyUqtECyS9WH31ACq/vqQzXCR3o2PGe7TmEYQ
HLq7kFSZzO9F1XEasOA3cQ9PxRf4KZl+kmEHt3QGg5pyOEQuFuyayF12nU1KCaSSWafjgTgn0CFd
qJwApgTA178TawY/kXzZUbJQazr97THesaMql/lhx/tmDEARZ9GUWpDU20RSmPH04opLkttGWRQk
uKjNk4q32GpkEKzyCxXEFTu5tQHf2Q3WVP6vUhU8ruNLBha3tGHtCZQO4wXag7jRqxMyI/WVxyXR
j2MqGPdViiNON/YiArHaqARfPVbpsCI8nlpPrSdiN5SGtJ2RyZITUowYY23nC3f8l0EL7nuwNSAS
egRPF7Yrr+/oXIf9WLITgiHe03la2leokW7lVSLl5sfDmsL/J+TArEG5gr4hEAHTdCyyuB2/jQ6F
PeCJf9l2LoUD/GhfUksql+l3IdQc38PyJ8O+zWEFWTDpSddFeFUn0N8Ygp4OnikXA7AG9A1E0aLw
QNu8vuEWML0a/AxN+FTyItdGvcCMeB2LMnYMYF4C7kgZjBAOe90sp3y4p3xai8JQ7ZJ2C9rqrd9p
8Yl8N0KVibWEvFIeq8XS9IBjvzmUt4l4TgtF33PugNenXE+txHuYtIH3zei73wMFCJGe7gXw1NFG
AIPtcNwSl+qM7rYBOu9sD9P4YvLW1mNHKPXrY3KYBrDq/DzVH8nUQc3YyzAC/K0qtUA152UCyzm2
IX6x79arxkGx212raFUlUydjnVCdyuc87oqW+aMg4VsuJGFBmtsqvy2DQNUZiJJyPgbmrtjflq+g
fPhSsxyQYX9iaPTbomc4qghzlNhz9ycYCo4VHh7U0tKOWP72DUBNSrm7PfJxQ+rGpkwBDgMhVA+7
gvjoYKcZqGpBhVXQ7S5kkJYcSgQ1HYiEsCyATTeolwVbdWslmGmA9g71vV0UJeNkddqcwlhRfZOR
BySaVSGS5NtsQ0uKjYI66v4Pws/Rxu4LZL7MRC6sCVUky6PAGcBS4aWoIWUkc++oSvsiHvDH84r7
vlSDLrwanCSV21Sj74AJllp+16tBiVco1Lpzz7nJUN6OSHYk/Th0zkDg38MxohcuNno4wj7AHsGV
Zw0l87US5sLK1Sm+5U+S/3JrWj7QfmN+66iVQDvgGQRtPoIItRb8xnFH2PkpeU3TcXIWkIY51h6J
MwVH/giU5qLl6wEDE++kZP50cYzRL4JJiDK9tNyDjpeftBfXWPTdYRmp6TU2cZBC+ZOGKPOV6xQ6
XndurrVOkOUzH5kXLxEyEu5OuPxFgcebr3F4ucDhzM6RIPZYuh5uyneYkuepmrz4hurYNNueH+zj
lTL1bCjHXRYqypQjTOKfL03LHtJMWT7OAMhVtbfDM63mvXguiF3539V882u6F8AkYeJ94XmcYuA0
tX1qyXQxF/9SwmAgf6cFcSCTBLwgSGZ2YT4NHGP55M6auWn3wEN16wlvJSfdFz2kOKyqifX+5p8U
PGCyuWW2GBYvZfiL+DCk9hUUQ9IuuoGGv8UM8hoBUFiH3PmigY0nPCaZdgdQmO/Fb5p5zpY+Wp/E
NHVxUTKFNgTL1MnEL+tOfVI1GuB/mp0fOUR/nYdOPrTQc86XYai8tl26OmkZP9qoA7ezUBNcp0jA
mTDT5+IxMwijrNUYF1+1WrcX3qW866q3Htg/DXtH14D4i4Cg/TwpZj4AnjZ8jq9YcSw3yMmEqOxQ
vEffSQ5LzWjBDcPYI4OcZeK9c+uh2iM98E+GLPwBEyJlaFuPnzE6NAJJErvELMfbiA4dCZrY6zKL
W2Ivw6UoXCzUdwAZ6G17Pwi04gcMtWLVElt2roAyXUImQbanyJWvBxQ8pGwaA22o08DpAr8hWDyO
aEj6+qvcHW/Jth4x61zPq3Mhj2RcHPD43W6NWhsYumkTFX8SmxIP92iPc/G5uCArkiyHb8L5w+UX
Bdp3yjs0pW8VsfQPxKEU/QSUgjLLjgau9m5a1BWiD/MauC4wZjFOtLyOJwDhBrsEDbGIhYtdQvEZ
O+QDItHpDsUkOwCHXAT9EbI+OyU2+O6E1Z9ne1DojGcPXItIS2Z/H/1od3/gO1lEQarzcURpw+E7
au4v5ieIo7SVFrSKjjyWnSc/59HwWLQtP21818BACwnNVAcU3uqdSO3m56CALV1odLe8ZtNtYqv9
CQO1vNP+MbVwksg1htQBwD5uiKozr7pcKMezh+KkQr8vjLTuQMzgQCxLk+TXrfcHCLGGosAWqE66
hK6i/VWqcBIv7KDjcETqC+Xd/NEyG1yb7cDytUUrsCKBoM3YApzS74I2wWO7AAGsc2fPSUuv/247
QrczMON9BgLBRld/83wu22CtcSBzylLWwafnEtKH4qNHGOy9Pv5xvvyO4ZA7abWdTo6CQlelmIUh
96L6EoxE0tWNeRpdXlhCDFkxyNF+jAT4A+/J7cg0p2u+k5OriFXzPIvjZupPehTTEn7jl8+F7rpY
atW65Z8PCiZCeoi3njWEDdUBqUqXkD9B3X79S3rs/SVMuYndMDsNjD5iPKNGF7M7lxgPE7TakSGG
1Y5j6nQOy+J5dNifRuw5faXJY/AWw248Ml3yJ6GhcvtaCVQtu7lEAwuPlxTJpWjWco68ja50hHIb
8HaeXbIIH1sOodrwRu6j3VZIE8qmM3ahJvf3oVQLBii7QnXVCoiQKa1YqtAup1FHhreF0UINN9x1
qdo+RSMoxlqDVZDQgTUdPVUpiEUcxzf/lpEZq1eMlshJz2SmA9evHodhg85u6XUkrJrx46+RNS3d
3vHSibapA9JlvZylGUpbGyo6UQAhTYdh9RpdhcyFnI6xG0WFB2cp7WjrQCm4Q0d/acDEF2zRI3By
PEzgTri7hddFcUZZSnkMDn1a9b+w4mHZSnL1GPesljrptC61LSpryM61AZRh/b3K4o3Rq/fFpQYC
6304B8UJyAXEtLFhngR3AxccsqEQGiafYvpkEb1BXyfkeHTptEHwJPM/cKbSwiGWuCAJ8OMOuw4y
eElHFVCRpZVUsvFIDFCgd8nK2Uwx/U7gzMVh4SlYcIQGxrTF/xgMKiBKGgAazmlWcBZEZ0RxVJ/8
+xhISm7VY/ixLVGs5S3jLVNSedFMXG1EVmuLCW/PPN2rHLsDxS3ckL2pKTB2Z8AKkVrRwrYimQz9
NdeCJlvpynxrJB2LmNCX6eprsS+FmkW1MGAqJnTqkqUCZF3O28Dk7ranoFSdiX7geoX2kXG3ZTcO
gPMjOMb88Eie3vZHasaPqkOHR55EJqFUrUzqR3Q+gzniDR40jFN98zTC2RuWUV0BdrysbMNIpxgV
6px2c65YfgmxfAO3koNSVvPbrtuKRepUBtbRvF5cQUIckiCLEs/MCX0922uIm9QX3KbeMTxA/KMO
Ep9ler8g+09jvtqxKTw1gQdFy03gMcJaJ2qVpHhXpyh9F9pUHm1tye8lxrCJXNRQ2Dq9GADNzJtB
kmxNO7F+N3CnLVZE4gJgsoDO/3lVRpuKkd7M7BICfMYH/rg7k/vur6G2RaQxofLk1Ybnrj6ZMhe+
kqUlfWhvuHrtbs0tFEqRdZGgY8hcFL9PRW3vKGI0aIWA1Z5Zp5idxb5hvWkK1q+DYPhgGqFz/XUe
rCCVhOB+oNDSj/FOURwVPvLzMW4BEH36NWXZTT+YoAo2kXLWcDy4BNKuHCdID+tcuyyxHDb0PENB
k0lTcV6xj45ryQGmEeHyFinPl8ro6QabcH5TqnPE/fLdZ7c0MDwXcF3z8lguewkMwatErP/2PbV9
jlB2caULNhRjhhmOa4vBW+TAQ+pNAAXMUh20+mbAweQQeTJp0XhlC/EAtC4cgfmRGDr+YqeYQqfV
aLdoO5BmPvtKtGBQGs8qYSVlky6BH83RR0OiEk7A2DD/XjEg+By8GLNBV6I1lUP+BhpZOBogxHh+
trB9aQgmT9+kYTBU1WV00N8Dkb38dVezT+NF4QFo/K6Euzz3qbrScJVu1OS/vAJpjwzNIrJl/sDE
9o9Sfcw6JfxtuC7QdV1QQlZIxsBNO0LaVETisv4v+OXNyB1ijrOIQRUh0/v2nmS6WAcoB9KTfBZ5
sGzWxcuJgoxOaaBEAq8D4+sacZyS4H6Ae+9QUaOQi/xmN8vroZjePU7tR3ySqW75EiruCVWIzAbw
0zdljjFzJ0U59MYiSBWRhoKDGJDRH/wVhWZ1PmNd9HPRVsTELMaF4VfRGuqeMXilw39lU/93I12B
p7gI55R84EjbXDJwH5QObyCP6za30P5QcDvNbRrMkf+aBjsCzRZccpVNY34L/ttkwCgDsM+/CC2m
yqjjnCC4/JWtGY8wr6D+SKycYjdy7J9sWANWy+AO7m14CEoc9eDgmHXmBflHWmJFSJpQNTFjHYY/
ZezyOr2s/Ddj0yCq+JNSgUhpwhKa4ssbY9OD3xRC4690qD81AaMX17jDTozNR5kfh7ZU6jwpDx54
Exy0pfPuPWmmLv3XdmLYXwU6EBtbVSKu7PWkUT75zVcXZey62mbTMs7fr9wFqBvOH4o70uR3v1bh
1w4wd/XLZegwW3MfN1ZNBvJFG88OM5u12S1PHKRxftzLW0LLt9ZYL8voUyWjlYkv+SApvOpjqtax
IPeyLHf5HrtocBu5Dr8G84Lob2tFD21fM4aUnIZRpvym6kqT61oQmGEBnhBxQWgFxZrfE2JCr4Pr
PfwCFAwrNVSWY5YjzouoiVUXBLBBKVMO/XPsRg6DlDyJPgDmLaEjJbzcPJnI5tHIxMQeRrcXYDgR
5fPJ49Yd/KtLduB94Ikm2rL5tjRyOgEXvE9q3KABEDhGGBQgPtOUKBOVyFP5L7v3gOWuJd8qXojF
nV9YtsCh/xKCiVhl2qZLsi8egjIsFkUBgoALalEK5jC8kFL3uNhdCaWkEuPcy04vJz6EEuJFGWqa
SJmGR47oakSnFfkFzcqcI859dQQFmLmhqdftnszLzPp+qXt+2Bbi8KXDS5Ge7+dI0yJoqso9n9oC
IOT9R/SiicEuqmJPGU/C5Fpf5UEbzpRKfi1M1QjdSEg9n/ETZf0QuTXflPjFXM1juIV4azTyRPSW
xZJwCz+avpg8pYvwR490iYP1O8a5Ua3tJHvfGKf3rTbo6Jx8dVEMkbcXxueAhsBUEUrFWMkfNDRt
wsaazHE4b50Vpms/CX9ogsZqmvXAYoz8uhROaTvhdYiv32+KuIkpPGxVePcTmKAeZezpfOp4bn2r
70RruMXuXoTZ2I0gr1fET37dwY+b4uY2JvrBvsKygpuwW8MLBYg1H8XnlFpBri1hEJfX8Zy7jCbe
Ai8HM3GBx/CSIUALRnyKcgrlTvLUrBat30MIxLpZNFDmWhDLFov/3Nl0z1HjHny49Sv8A150JfMA
+jZ9LMdaWWJWyohBJTDiFRgCAzbk7rMKHAZuH+3WXpRBanKjBiyvLfx+ie7w62mPDgadB3pAjviK
yjYJTAxP92dUHN+2URoQYKoTlo7tPyATFTqQ0v99W+MyU0gypa8HeE49qZq6GdSzBaeNAq4Gy1Pu
StE6kobcV3jhgfO5YoFYK5X6fwjngp8uQd40HiN61vgja6+qr3gnZk0F83wlzABv14zKR2e/uIxw
Bp9ejstQ5RQmo3DC+1z0rxtdGrRZU9x28op0LtmxzIgRBg+14rOldxyADsC9xdNhWeE2sdG6dtZZ
P9oJ3Ir3MbcpfoByoSM2DJs/Z48MLjXQSdiRsOIqhc44tE6uZ4MfkLqsFyM9CzO/gPRJIuWf9Ab3
urHJ5/16NI8S2knn6yR8sMiqvdYWZPBTFMmHBr4fF1VP/vl6VN/h4rVRCDAM97TNZvbjQ2g38/vE
5u2zO1QMZ6WNlljJEbm2ygU7KTyVwV8RvzCNOhCU7/BldFAlWOMWA+vqZHxcl7qFJZh/3GyFRsiM
APD/aNq+MNCC4Q8zvlUoBLKBxKSp5d81LNMGk+/fNfcbMsIoDnH6YiKNoEm5wIN/1vbzSVPmhWV9
TsJ1T17aZKxsF3Or4B7xhsCoGNjB3OFbF24yzTcpUIRqNi8reoJ9q6PS/DZYD8aWrpPiN4lX3aQp
2eIl5BmbdATYqS1VnSbM6GaX2WNKQHfmiGWT93Wbzr95mqPUgbjwE8UbfNuUqFRL6qX6Rk7YXyLI
XoiyOz6ZMJ+57F/cakOrYZ+hZfTidI+TxeqT0CTx1qWD3VaFF43majLfTh6/EKe53ybzImz20bhS
/uMhaHJpwHRQ4BOnLXy3nLjbqq8VWQu3MG6+sIXINCQDxP526ymf121hPGFr2Thvvd/16KoTWAvm
eXL8G6yoyYPoRmyUtqCg+RWXxss94uQjfzHqXPTxzQg1jOW3GKWIzmvhaRwbCMz9j/GliNRrwOnD
u2c1uPkgy3iBYm52JzsAfKbFfSK2YnVWQjeVJxHGErxLcw74BGklRke+Rvi+lUW3X4nqnVdeRUvj
j3RErqRI1wio7h3gR4cZCpeWeZygSPUXxw3KIX/w+VqHSTc7+bjml+acuVLAvVGNWx38ScLOr+hC
FONh2LBueOgtkjzly+Efj/yxd7xOpnjRY3guBrjONCFoTaaQxX0+KHF8s2GDYAZBfRqvS66MOoZS
3CrBKOlZMhmhX4QnwqE0WJsZgK8UKYFT95S4l9aAEUhMShiJVpytXdt0NULTScji404w8wjhVLgN
tTx8r1sIeXEOIjTr6IkRF7ZfP4/O9+2IYv8jG4kvxOOgHRwSHaeWZHDYBl6ksCKvYzFKSsftTF+q
KdgURL5HkBJXLghK819/GLhhSGg/lguTEymzQUYeGl+bL51ZsXIOBVNtxYy0F/yvBmKlNSWbH7VS
lW7AGRtiRv69PvjJ+Is21LctejFQF7GVdliBHFSosFJ0MZNE58SQsrUp2iYdUuhLa4EXka/bIK8X
TSswRkljImDAHIZN8yCyuVTKVC3cBvggESy5fmJOX8YYlmqumTSEFwX3gtzgfyBVLP+BROX6sNYz
GEirCvb6JXPogDvBeynU5czAPhjLhk+ug9AW+S7GmCJeFRxaM+vyPhjOvEmQ+2Dw/NOPrNVHFnkC
Lx+/E2GOJ9Yzg5LgR4GoVAbfHlylX1RbNyrd2oaedZbLBXtmjIewrBc4Kg/YOl8kr3anYTclhU1Y
muojjzXg5VuJPVOTfM3z5BVGSanJtlXOdcJ+YllFdEZCql9sX8DBylL2qscvWpzHFI4/6eODSVD3
H/lObNGIeUci6oGXOySN8DJlzKvNPmrz+H4MwGsotnQpKKlrdv4ZbHXK/OzhEIKrKyc/xoXXjHl3
XsfmtSN2pg47EkEIP3s6kOhFAzH4EIz7VCOkEzNPncRhyJFU2g6iZDW5FnkfzKNH+thgduXQy2Kg
gI672rF2j0si0AK3jxtA/kyP9L7EYsigXhRCHJoJqwGLfuxfS2YOcBaSOC12sGB+UVylFXAYcd5e
BUeJMGbQYuijSoAHhV6/75MoldrDtnWnZ1ldbrjN9SYYj5npRPb5qtNEmI3c3gCGK12ftQ7xpdcy
UYQzNzjDtI3cEyFRWWZrhmYWi0PmVC5I+tIG78M14IjpBGwC3leb6g94VtugG2Kq5+HUylgn3TGi
f+X1G4h7471a1DYhbBI50Wqa0qD/EbQqjA/npib9m2YkNMO3Xzy1fl4gjYFk0TmYdoIcG64IjBod
OCr/9bhWf5wh41b1ogGb0aPOU0cajxj5abHpvEJFQlTwYIvxe2wc89/O00zhbtadAyOT4Cqd0uh9
WY6g4y3D6HM43Q2WPYh8+Msp03xZtBVZyJfq19p7laqAjl/kMqXShLD4CXneNDDZ9Ggg1KHM3GAq
n72xm2FdA99TE37/kQ9Tw22Fkd4jC3SsVUdaLqPTzI7qxD8AdRt2yLb4ebHIGaPbhvb+W1p/S9gv
MzNWdCtvzrDbYwFbIhD9sgftQpiPsXbTLvhJHyXCupuQcHEXjGnUX3cabuQPrOvCFyfrCj1Veq9U
xOadF88JKCb89m8wvYs+1ydOcRvXQYi7DmiD1Ue+p4JpPXBGxicjL5gWcvcksgqMwd81GcjnGy9C
sgLqBOLtggvDeK5ZTyI4+h8g6cOTEy8VcmRrK581G6PVMwaVz28smT+BfC7qjLjHYm3BhN++WwYB
8pk6Og9ZpvBGdt+dbgT7kjsJ3+FEU0t8g8B6mR25hBUfLfRd5MW9QZH9D3W0JLqx0mqB4kGHzdQS
ViF8UFvU3RbRoY+6QsMiLP3LOtHeyesfHLLO3i4BLxkdnvD28qG/zrbNOk+ably2uB34e8oKLh6w
rR80ez+pxMtOyO8Ap1oCiWPdlNXBGQ1GGZEVdTEUE+HFkrhf7H0m/3MxFYxJGorHG2HTS5zPtN6m
OWyqoDTrJsiuQ4goRjuwM9VBlZzShkmcQxKiw5XPeJHPD/m31vvSK9UEHZsg6R41Shulcc4zt2aY
ogGibvaG7nHG9VOG9lGpUr52ycAWM5lAEM04Bdo1cj2r6jvnm94uKhi+F0K3gQOpT6lx7NGbqFg4
x7MgeIPcPfmVBgRkvCTAxMmbDMw5qR39HYWjTn4gVP9FLfxwlKbrawR2gBeEXmRtkWMQ4Ni0nKRL
cd2D4zhDCdqFq7NN38CkjiewXWDov9JkouN+k4I7FhzUeKpPyueDu3D1O/RYCWZVhKjnSNSlYQAc
XZWCIv/aCiB9SFVNinZQNlrWNJaHzmjYp70zW3VORYOy646i8E1/XhWIt6CcBSKS2mBEdXfET6ZC
k8tRd9jdRgljqTAUZpnFGfsRNyT2I8Dj/kvGtWCTciwoJ0g1H/fEqIS7w9Yqt5AsRuxhxT/o29WJ
hNCEgsx0vp8YBngCjMd8WhAB1IpNkxtlLkoWsSJ7Ws/oL1391FAfTSv+UtF68knkaqq+F8Nzo/Vu
NblxWg366BWG4Z+ZxVzVdI1RnrCDl1p26IcY9gZhLeCHdMlaf+UTdqomEeDeB33Mt93nkNwVGylZ
uACLYpum/QaVN5NDDfkLSEkcj3+XpPL4wka6SQQV/SHdzY6Sl8RhHy8R4xLRL1dhxsSFLS2LqZUV
iQU7oE6/GWG6PKIvTUHcvBPdvoFlN9MJ+5Zy+oqxhuDVKGIvt1CnPQVtq6VqoEVD9S4woQbUYL2C
Yb+kuBrTYpHbAP5bs8aTCBaSCw8RHYL5B+JU/Ksb4mNPTq4IYiY/a6SACdSAJ0kiRUv0PqOrjFop
ylSlbukexy1yoU4xD76ljyZrMNGD8TuksPnhepwLWpYlJfoZlIX5riYmRhAT69rBdlWF3XUAYrZV
8+So9FpmSohMT4YoiX4EZkeBJB4KjG1qfDT3tBzNmcSaNjV0Jz1pL2Af7tWVlbXICeGZxUpJZ8LS
u0CgnOD1IG0jMkV03eJkPpowcD8IgRfyMKtQ2KGOMX8jCpHGt8fFSqxloIPd98aNauS6c9xwh3bs
pisgaHvpx4VNLgH+qCzU0PRN5EGGhu+AgRpsn+tfD4PZZMn5aQEmrk5n3DROUHUa940nW4LsE2a4
5wJfRKlciFBonQJ+3hRnv36MC6XwNYzqDgYFg0VhvDCCh26nreCMBMzD5TsATj4bmc6fBoR285BS
8ajtu/N2c5TowQZwVvJAlnCstzc6flmq1e3gQ5DjDsn2mSZ6nbuT2epS3ig5Zk7edBuZpbsJeC3/
tlcMs3s9ZaPoGlMa5nsQsBOZAfZzUQbCD/PsqvDtO4WzFKo26cTtZVgkyYTmi8UiZv7S1qJCZto5
cNDN/6tjPf9euDFz5TVoDddTCFpdHHUjVwJj40KuEe5Jj8noz+qrfoowz0fzYmRuMDXfAuwgzCBT
pbLo1F/tFd8Iq7GltuLDc3cLXgGEmlCUa26Fvhawx3qHhI5UJyg5N07PfXF0QfdL9/BH7YLx1st4
jKF8EoqgJ25FWg/AiHDq00gONJ4787sNAvi/VIl/tItOeLCk/v++J/oqUoyd/w4a3M++uxfCRDwM
/XLgu/9+PYxwcjZwUyXLRKSRpkiioHG63n6tJM13F9OPZ06sgYfRDx3yRs/v85Kk710OCeTgXeH7
GLLr98kEtwLKJD38cIvlxG6kFOIMQz0InlmMWxAkksh5vY35/4ZnUIJYT/rQ26Wud2gEKEJK/R3d
c8NOjDuC/M2sz3Pc8Y/SgdqHJwLHh2Kglp9OZb4Qm+Y8aC9VBeFlUSPRQki/sJ62nx9b4OYDpR6f
2PGoauClT4JuKfbBH3TixL+0BcnWcYK9EvRF87f7VMJJhtvI8CnnoCEdndjsH90Rza7FsAfUu4Lq
iyicvdKnEQFBIYDzX55djGIYwesNKTFDO2JV5jqBIbF2Ulkf8TB2pJw6/3Z//T5hYx9GVf6MMoaF
KE/lXo/+FS4MVRa8gvVb212yFQnv0paNT/BJljug7FVpedg0w8M5JKcTDnGsLf3x9+VE7atCwkAf
CzdMBNYJ4lIaz+vKeq2cLjdf/9vaX5Za539ghbxeT66QTlaTJjdiT/4vPbtnHOj0baiy/tq3HYjG
nchL1xD4R1gs5Q2Wcerljs0FG6WUOyAwWrGbermGOrEpK17SRFZN4u0fvMiPNQ7oqdNm/QUuHh9Q
34ctGpSTCHcbggPtzLQ6wLyIcsQ6t+4lmmLkEdNXO3ka/D+IhiLXbpAXO7XDzzrtiENMh+jYkFDr
G8NMA8jz+YQHdvohnk1Sm4MSePupynkQzH9tNor0CNpzIDNloybBKuGP27PVv3R2KsyfROa3Mbwc
ASQR948Z3Vw9cjxZmBlcCrjHHZvUWR68Y1uihFTryhuhmunAhU38IVZudGqwsjWb/SOLQLPKblyk
MC+O80wqDo3q8zPWlNv6bcZbKaR54xZOFWCAz/Sx63iOsOvTzVxzikX82gjVgflniUhaemdy4V65
vZJn6ReQ1SPvZkOTMiOekUfy9oMIyx+Xwrzcrkv0papm/IOCGTwt2EGuSGq+kpou7dD9qAcctBfv
i4SQ8RixryJE/yYMKNlKy1LplgWi3S1KjYTKExwuHaYcQg9YgSH5EZehLyu6o3xaaYaVhwyFtG4D
mlympkxy0p+icwme9qehArQ18ikMg6VJwjSGJy43hy+DRMFXPcQOKknVK57bNpDwF818c3lxIABU
5MRX+BM4QpTiFlUvpiXMUEb7VYFx5BTQoDqIVXXl52XO3EUOJRso0ZemC2ABwcGgFlNsbkvvxfK7
UglMBTFGBHjoMqYj4OZDaQiHH6WsvtXTzJtQVGTvyDy4chrlQ6PgN87B2y9cn0PS6Qx7JTyZ8c2s
MBIyw6AHJ8nVVZBk40w9Ttq9oNYHu2UoJrBKKZyHHVaaAi5R0/9GiQlcGCjDmelu0misGNih+ae+
OIZVT2T8ILLfq3cTqPAmxqCKHW8UGeK1kw5uKQ0fYMLnoEZO70BOPAJve3pJG8JhEMDcNNXSp+oc
u2Yab4baXnbrIh3J8dVDjeMJls3lU++2Bw3MZxims1yCnVZRGmtyJxkCzy2h7dW64Emt1liygrTd
7e61AHMWBb0U5B6Muks830fM9LPJULP+0wHja1+3Kb0l1qcKF74H1VmHpLI/G6L4nRAw68rndfQ+
pRku/SifBMdbKk/6DijZVM2TS7CiogbbbdKGLs5w+pycum0VjvexId1xdR2WRhGrZrDf/EeHO5Ci
9BnJdCOWxESdHkUZAUMQ2bPEKnhuI+C3HehcdEbHWJ6UYEkXn/lak1xxBism9+phqWPtOJopqzCz
Z/J1gzUtspSD/tSIc+2axtpUcXAynEpVxlYcsHTgQDAUXhXAEyIjCX/oSlTZhnSkeEhsLgADibX8
zneWTVC04n4kXqhWMntbaVuBzovDJHv3w44cgecIaNLMv7PHFdU1xz4LpRXlxfn4l3aHm/02wvwL
LqjyGdsN2GPOBwjk0G/5Oc0tOgBr0Eml8U8o7OTR3BCAm0JW3DNAOun6GY8fwYzdJRtvS6ZlXPEv
aSICXxBfXVxBkC/q2fFo3mSDrKtEYgbuvKWDKRNbjoq57u6JC3ehOAfeoULdVxFLFnyEXvj3ZeIn
egBApAQzCcAGNEE3oY7YvglYfUlod+ra+Fxy1GubeaZKl3EFISCfg2c6P3dFWJ0N7T2k4Yj4fSqC
nI9EcCk62hxeCSRYvqOuz9CSu7IihCPrl4g8f5rcWyzCOEbfhSUIAlHdcGJppwSiXcoy1cBBhSJ9
eezkD6tGGD8VctmEAp9AQmftFTEIyucdsaE+3uwZKtMXUNSn8ZgKuQ4Geyn8giQmeIaxl3ETLbCX
sXG7r3ImEzlKxOAmHi4I7J6WAnnuZEoQZKyYziuuaUf9JeG+VCl2Kn6B6qhlhWsgcH4mx1xP7pC1
qxgDawT4o36yrLwhpgLWfjjvB6TZTMX7WyjP8ZW7M1/vgx/jYrw90z9ShtBriqM3Mz7B3IaQuigc
OKF3ubNj5sFPSXd+Zy6lJ6Ux3cK//+yxRPCglt/fwW8yASUa3WGkNuR7ji2TvEsrQwTk9NfTb5iL
FrzLR7UWIMWCYyebafdvjSNsw4N0Pq9dhxAvIJfs91lGWrqnntvUylyCoFAu4J+cKnEkeeV29aCA
C+6wzSW4P/6RYQ/Gwdwt/lbxa+V8nY5yZWeIsCUlRwdejHExnuI7tCHZdw1xMdkw1M79ovHZwPAx
7kBrJ7HUDO+dSasFDoNXRDHpbRjVMRGuulPlcq8BvbK+rovWiifIFWcpU+wHS9IjEMwROyro9Mtr
wRXQ2NORhQrBUWPauQV9epm+xM1YohZQLvw2J3UVG3lybO3wSS0Llusn4HpHDvBkrJ/I82Ib07oi
1NXnI+A1efcUfKSHFq99RhXMCfwndTjqS0iPnQ/graUfFp+gZQfhN//LSxgElcTTSAJR1rPs6gqj
Rn7qB+Q+rRLSOGnp7MVXslD38MkUtIh8NQDiG4QaMhz5qgnZ5hzeh3JTr0B+/25YUw4DxPr1n3bz
FG5KwIUDMaydIYl5P78j120XjGsgqb0O6jwhFTBMJG4EHkaEe/Jr9GhFcz7T1PBsvmDpa6JdjFbG
+KR3aKpOco+pQ7c7ATjijDZxdgPk3gCqlXyW66Uuwfgz4HqVXOzUmzNu1w3qy+/hcV8nKzFm6OsJ
PeC7+8QumKWpHEEuUOSrLoCHwvFc/L5zB2esiik49wZpiw7+OS0WcHFjA4kP/92f83ZxS+rW448V
jK3SJVTcc94IbHWGNBZGj0NH3KhXsfbPjarSEzteZfGU6cJHZWzFacdYOuZ4jM0JUETT94w9CjH9
dC4baeKpPKaLlLwi04lez1LrlFAvaqD2Pu+zEE6fDgAQ+cMHqFNYhx9SlQAM9jrbf5TvsdFnd7nv
xXO0zAWAO1Vvj6i86p8PAzjNI9dHg+KVVWGs11wWIgs4q0bC69tiiVfs49fS512g736ie64l5O6r
u13YYzdNEoiLJtsODyF7cELayFS1ef6m4OG8TfNaYAWYSD9FMyI2QFF9/f0yvEPuy/NTaJNtubuj
p9WGHs2iaJ8t40n411mRZyl+kD7zSXIW7Siz2BNHHIuYd7nAX/n3sWRuM+ULHOdsf/rXGC+Mcc40
GnucT0elQ1xkSwPmXniyM59yJPDc0sWKel61LYqs6qtDeTAF7F0EbSSrUS/GII1bJHzatWDb7oa5
FyfME/AHBbAh/36RSN0PC2jRDxzl7rHxXEEMnmOgC1vKuM/bwpm1FMkGBx9k4Yk3nMxGgQrXALTY
9niWAR0oOg5ajTM5bDxZKB5iJYmlumGFcdzlIfH5hRrx4wOK5ug0tlMG0H5xOx6HSrU8J6V60/qV
zWQCpBUOPNU5cvTip1alLrZfvgevTm8Pje4F92WIGNfvdH/UuktNc3tF/BjocXmMYqyvdS4zxU6r
E+KULiEb2yeQLtnG4cpZjG5um8qj3Qb8h21oYXghbDGbEUCJPuKDtnTmiwKDRqANvC16UnkNiLi3
N2a1RUgQs/1g/b3FM73BqA9XhFP6nu4RIogjvXOQtyA+4gFO/+D05DzsNHbCgFzk2hFe5TwZ/3ZV
8KFNGbvEYYfVi7Lyp36qh9HQydQw17fSvs7CWRAevjMKp8M1xlMbjo4jO9WlWlraDNTh3GlQ+0p4
FffQlJp6gPFao/7Ev2r0kAHgkv1wx+9Yargqnc1SrK+zzz2V+lAtUj8Dh/j5YkwukbcPzM1UfkgB
sRfegHP4KekB3dSMYUNpia7Rb7OciQIjLG+i3hPmRnvC9u0NNt2MgVmO7c1IvOtpMgBRUD7IqklZ
P7b+jEAi+1+XGeG6gMHGplB+4N4b2UaH2e+TwfCbvwG6wfUXStwmkDKYYm2DSGiyS1MCYbJq/YgT
RutMjf5ZaA7A8V02VZaKC7QC3e3shBQ+NDryvOy5yjzRHx6p92kdI5AkQFwLyPunwTyoDRFxMgVu
JvNl6EsoOrUH7dz74KauiE8RES3ssjJeM45uwygmkKWujyX5R/ZclX4LIi1ZTjXKv/nGChKKerUB
1cCKgNs9KchtBKK9oQ0oO6r+uT8d+ajEqZviFjcIW/aKa3DroH9tiX98H7NgM22k7qqI5MuTAe6U
Wh14IBOd5c22BGW2uoS4zIQvhpuRHj5ldzkL7U5I1HAc+OogzG1PDSdcI3xKtAfnr3RUhnWbq9LA
lk1KFtQ1WV+Abx0v4ef6yZSX53LRaPFAgtSa6uNvk6fK4UcVdNcvLBafgs1UcplQvqIBGgygMIQ4
qdJ8Tew+QlW+L6K+Y1ACxIzDAnREFsAnbXJ2YM6ITWDGNovrDwEWqsfB7NlL5oTIVXIvXkNwGyiW
9aGXjHuJhd3+E0cTqi6PHPzvYkJZq7yZkQYtXk8Pi0Ox0gZn7uchNjjcCIeeH082Q6Uy816NO4f9
WfbuM7vDJ/ubE9LshzbBd28pQyQ3IOIxEd7QM0zQQNrY4G2/78KaHGHmWIQHbXxIm/C6M1inN5ZK
Lz1elFgDGNUncSMRFt4z7DIz10n8dxjP6/m0BHk9EtbRzzrB1C4OAccIqF6aszeQlyAovBDJp2X5
XUjyDLfhXddOUXPeBhEn6+WOi/C6Gh9kz2JfJDmwxcoPlsOEix/M+FTa8kv2JikhSV7A5DPkb44g
micBTyKE+WjQvCPo5IP4/LScxtXHSTdTdG0lBtO9J3jmwhFKoPVNeu9b6UrXAoeE4KfGPD98h5pp
gO18NI/P81LSJEU5yPI2I4/oR04ld/snq36by8wT18Ouka0Yn3QMWzbLuoYwEDMNG1XAxBiTMo0/
Z3dbfC+KVixD/IxMXwvLRrLM/0t66DZ11WAIepLRX9EFwJlIfZ/fRZjVrO9VaqJKpAgeQGa4poFc
dV/ntVt1F5MlEY8COLFVuATPXFCDFdrHYtkInLZvLVUbixVWGcdngcHjYpkr7HsEtQDM1Tw/EGRw
9JAvEKycwIv3y9C5UrRiAS4v474UmTgHqTlSVAePxHv1AMRmjrncHdr9qOwXS0AzIK8w6jMSPvSr
VqAEs/bOpvl4daSmef96MenqgcvOUS97qP6CcHoal1Hgk2mzzfiX+Xham5d7KVtkwcHh1OqTGJYX
yTBvEmJYXUsiGxPAhAnjUOu4DWiE5ce1Em1MFjEovMU7BNTBBdUGv+ODAEq7MuM2atENRmopp1+X
4ffskblvBby0JeLqf3eLFmhe9qnOz3mOZrPQBfpagaogBnwuytvGj7SiuGUXY/voa1LUh/t94nyb
pp51k/rOIgBl0ie+eKAUdK77LQU/BL88k3HolL0QTE3NrKiR23u4oPl0EObLKjURrraAfMQCqI2O
SPHHCDQjOvdU37zSnKF61p8cM6YHftSz2sEYoWHcG4jZVjKxejEgjDXmFtYfdWBXmOdZTO233Jxo
v3oQkKl5+691xOIHcOEs3oepIB1Ad1NHAtjcPkJWQ6z5+41pYASnwiZp4LmT3rybnkgmBpCUDUTC
PBmU7fhOhXwsla4OQDIodPQAsHJxh6v/7EIxHOcyLCCeJJmAiYYSxX0QpdwRlsZ9ultGLna3y0gW
2Kp8ncfMuKx2tUQF4uTOxSSMUowA4P6eiU4KXe8U/+W6qCorfeNQnDUdohSPkE77dU485tVS+MZ6
AOKXkblJyS51FQCqsbvkr4vRXArk6GUlyagge7mjoHxkRC2LyDo/hMCzk6FxVGmGyQkHsyzQHh0/
LdXoseIMRcAvxhmF8HbqZR5hCH9UClBJO/3K7KlJb/bdJxOdFsoWyO/0+X39FIlMvWMnNWt759bZ
yuhG4KJLatVk0gnX5bdnZPsu7nMftdg2Lbz2BYRDxn/w1njcp8dlln8OwSxculr7eMRt0jVCYF93
xpiOZNbcGs2ijPh4V9XveLIOR8gi5SjQzmbNok+RQxlmoV2CPA+Ho/zmN/qz7/1+ZlUfeftYsV6/
D9UwdLoDxVFNTP6qpG9xMoh4121o9v9opJU2xMzTa7485mXpAUoeqTccE7+CAEwu5bjJwVSN9ADX
Ooa2Iaip6J3oPDJDT+xrqpvuW3TQr4a8HYtWJDbp0C17r2j739IudPrZ+q6jf0IL5siD4AFPnZ4Y
0qIs8LChY00DtNFdII8Joj70Zq3CTmFuFe3192sAEozdHFuoKU6oVPMjr6KxTA+6g0T7ikSMXaKE
UIhmsB6vupAo4BJ+StdIV1BkE331w8hQbFA8BjOsUWBjipY7/0j0uqKlo9fnUkdjJp9F158QVo+p
VxXLwSwNpXLjio2gLarj86W/e9GnJSKivdJRLWQSL+E20RzFVkeQryqZE5eNo7RGKOql8J5Lu3j1
h0edW4zVX7NarDDYGFHre/aXWX3p9yOBXnOfaN6Wa7ZtzJZCXgKeYueVHAFjMkSS1XZL59V7cJes
2ArXwbCN4RV8r0uaew4RqZxh2ESXbeekBS2U4X6aeCtIrpWvX51gJ4fLTqPx6lWuBOTiCfpxkomO
//A+FGPYPJoDdnYSkh0NdcHABryQ6ZQX8P6uKBrSpvkF+9RF+2fheUs9reWf3+C3pVotS3EgyGoD
dI6VBZmpb/k+Q2WvFyUKSU1+7uIEKjciZDiaxFSOTmzHHYomJd4Xh9wh9049S50ZuobV45t9FRmI
CAPh65RSxnT0xTWCHIhKDKpq9oowKxyIv+DDuKPc7igJHboBECWFxDM7Ojev662IgEc1gonRbnX0
A1K3/XKdxqrGfQocLmQZIVEAdT7glA6v66Lkel6P6YcOd287qkVwKd536XaO+V8ySZOkhXYgXd4V
8cb637ItQtSoxfqsj+4rEOcpdPgfmluF9auPNn2NGCPhjoSV0l41truDqGBaBa31XV3qM2MRibS+
1n+V9j3Y4Ozpx5HzaeoFZX9pC3WtnQnlsCbRhZtobKzVnRO85aUjDReumXOJs4pEaUXyXC61GVio
77fAV+zPciCizyVg5BTAFERlPvOTjbk+9XuvzY4ED6E8HNFpR8gnfglRkELGlqrFwfXVUHpVnThx
u8STARGqDlhb6RUtGOteizdySE/X0mLsF5//WtEK42Dc53SaDMcovp4cwiY6kSo5h7VJj906h01Y
TgSxE1vGBUdAOYK7qc8Jkh5fVQN+dzZyfq9lw9dUkVBpugoDhgLGIkmIMKjaVBwfnjQVKb+kKqjN
yu+b3hLpWsrZbXPus+bDZa+SKf/hFDqSqDJURce1noDxlUgVmbXcjesS36s4M14HRhLrmUfydPi8
EBz8Z8UgDFSWLA3H+fSz1sPuTV9Sow+6tX/B4g6a6t161W6WieYd51g4G5OGwNlYJzjlGghoY7B/
gRpvI4pjHIlx93dyCzQXZXLl1C0Mpq9uWZoEWdOlQoLOCBR3MyZ/gaB3x5HuTwH7+LjmnGTB/ZlI
hYndeKHArpP5y/gy0yODCOXtxcMcXLbhuyBA0oLoslR5wlUClRTapvgSHc3Zt3NLcFjhJI10cqNg
BOm1dmhqCg5GQ7x9QhZdTofrripseWsjJI/E6HVN63lrbM35jzTeBKWCHhwj2gxNSx45lTf2j/f+
YHrtOdWNRcj+mI/bmu1RlRy2wCltFqTfRaZ4Y7L4sL+bhP+RP17/tRJAlahboSv/QcXGTWEADwDX
yf78SQhUiBme994u9xrFPReV2wIsljYT51DMpGpvai6WoTBxD2mDkiMI1XXYekYcrcTFnBHkggh2
RcwrDsGHGFZZMip+aEya8SKBJaCQ5/DDfIlnN3fqnbderYd28crnO4jnoEq7DeoxBFxLwwH8XGET
9MrqazhHyP2UfVdM9GsIBqZJnH0A6ofUOYjKqOqFztNISUlH//p+jRmtNLhGvcAy8JMhyCkfTdJY
0j/zN1ZrCzKAc/HsE8rsK+ihuOs2U8kz2VdFqE9PLVWjdicQjD4anO9QdnBzJM+Ti4pIGajt21JV
l+AEPoyGFJ4K+vDL08A1wHNgoKlHiz4xDBSHi3p+vOZ74Uanr8tSCcBjVyEHyL96vNo6ptyvzRPE
ImkjSHkgNdZ7Vb2Jffgzk9EgEhejIrDC58pVw+5sTzJ6vO8mnNC6RDfNFmxUd09u0l4182facytF
6hQ4bJoDyXNuCvZG4OWNvmT1HF6SKQi1izFS2utBchmUrDdUK18HBkP0Jrj1HOT/OxH2yPnRP7gD
wv/8gEPNFHOt1vqMZ+j/YW/Qt1p5E1m1bhHVt6WptlL5asTNwBnMw13I0nGXnVdLPv5RXifDrlbL
GSRM9xvPe5CGvQ1DrlZCf3vlSuYinx/nZGxBOwrNU1rfaHrlkHrJJz5MTWp5pU6Gou11u8TGjKtT
U87WIquX1HQidH+rf20ikXCnBQL4JxyBe8aVL0pdBPDiRTsVlmeLF11ATAPui1AytqVsoxuAvwdD
HSu6LEVihaRtS5BVGETW942NIfY0RdhhQRKOMSH2YXjkInm+U9xyD5jLoaxijUhiDrlaHCBdNEcg
iYp87Dp6lMk8m/DJwHotYa91zIYwXUvTNZonfkzfuGWUEaCYMYrVHl99ueOaNaC0RuMZhriXdqVN
20Balq+GvYGDJGci0qAJv3lk/gPXTSpo7WxuhPBhFvVdDoyjZZ2OJaRwkIOAHE5eZMRKtbcRrUpZ
HRqEkZp0Uh80qBJ/ENcmwsiiUdmAjF658M3UvtZybSqXgFVSxrPmWYz/X2kfH+mVL56MNYtKe/m5
NBIjBzEL2AMl4YJ4ahyYqvTKIvHhUrtTthbc8hJlissu1h9cV1pNOpqehVU9XL7F2kqUORERzGl+
qLgHJ/2kw18NkM+kbj0YSUVzQyiXL9Jv6CWxHNsFIiD9vDBcwoW9Mt1pXtv2cn3alx/2+YrFElqz
JLqAkwl1nZW2OZ92yzrjeVkDtSo1QupZGViNp/+BwH07OtLflN/PB8SMQuvP+8CFTHeOhVon36am
GrhQMn2MXTjviKJ90GDHTF5qoRjgXOnsPuLx+y36DqsDYMFSOZksTcM3Rd8EvuE3MMvfcB25gU3Z
mLY+ZjWbOr7Q5NS0el64rfDKj07lTBJjXKFMF6LJ+OTCrGG9Rab9yR8H3zf+Fst2Yw3fDnLHJC6d
4znsxWoGf5CwKTjrSEPsmoVgZlc7fg7wPXKgc40wrJ031N31/iTO43ojhP65J+h2GxrPVmOLRVYc
D8U2atE4lf9f6QCj0Chmjwny0/aPQ53IzfRQs2BUq2x/Z3GbUcemwtUWqZD1YI2Qc7gChoPG76Pt
qDtraTZ9pC81xjxFyF2xUBmbxIJnM0rXlW2Hggebwb2mExA41zJkSwIQ0RATRquANQPOoAmqVhzT
0IWSCCI19HgHdjp8GZ6ensJwIQIzZvFgCJeIFQxjd08/htJNZidgT90ZffATh0Wihy3FDJ0EHZrx
Y5w35lr/Qhkb+9TBfUQeIp0pMPzUdP/7Xe1JtTkPn73L7sEMnyGvvzFeAxIFX4ANNl3r547IBDyr
EmbBtamZd8qJtaUg2nhb7phqZhiiZC2zXzAghQ7ednIlTQzreKHA73rlOY9IV0ZlKicnW45j+Vkw
u5ZNxf0+hCNohR5tvgFNkuGE7uJIInru+Lci/nCZ9h2G3LKNA3rGbIdLsNnG8JCijKbGDebkRGKw
fVcaMgRb4q/gNF3KQZg2J0Uay2ZW6CFXfURQsmL705LYpR9pH24U9A3nmBAtYH6d4E2Gx+rN1+39
S1aymAzHzDhUZtDWVW/kUpdF5Qf9J7vE5gfSLSuyakxah9KY/Yb+tWOmkyi7JpYgh+CAz71L8ufL
ntksoJIzwjRvfSCpD3563+jz0JXZiDp0E9L/YPDCqTZhrTph+eNvuVrhAm1SI6/FwsRtM5Vqc7jm
xGMPodQETa3OpYvA6zatNSjgsiqg21/g2EKFAXsTCPHgPsTv/zATppy8ODFhzxcF9MQnbxHIozYD
Vv7EtYtmx4goHmVTxfTbN60uvaYEGPXetQf8JDeu74dINVqKSJa3T5DqPpbLrC+HcigVzftqI5Gb
gmKGN8zzSZrxlkTA5tSKUZKNQ3VAgdtx1MmlUOarpCCbxJLjS3ZLJXumXxJViN8rz+eJ7eHE/frn
qyX5tW7AMJoYFcsiDkgaCqbHrRRuR5O+eo5evE3rvvcl5lpa9Eg8vRwHe/KOYTd0cogYjzu2C4hO
JeiQmk5zweGlWjec4PTXhQq+A8vohXuHWrYAq3niUwgeFwYqRW6j3Um9MvNUYWEIguBp7HqfmG3z
jS3rD0Z7BQulVZe7RBwmjzFVVcp+qbWV/zP2IIdmBVwTK3V0mpmYE2vYRbn7hFb2C5lE3rLwIDvX
y2XhD0l9gNr2RiFVQOp3GZ5aJ1KEmz4WQJNze0BktIGLQQrxA0J9P5cbbk9/X7SP6IKAkQQ7StBI
hjLzx/rlDxuEJd+YJTEfjgNX3rKG7XjFaPw6s9VNV7P3XPfdCXO1qV2XpYsNw8Ecc2OIy2AZFA7N
pnUBFo0eqQvuy+/Y1oKPwpRxYkMZZPLSVD1r0CNjNqp6GhDU7UgJa7q4Il2KtTOqNcK7wbRIO5L4
3ePNWozt1KvKgTesAc1iB3fw1KTczs36o0v+su2GXK08bZLJZ4cN9RsI7B8x6eBI/bBwd2gkenvo
Y1goHRicgBkIl87EZ929/6/SYIQG8SAYxf9nTKOJUw0d2WpJOgjSAaeFCPvG3FH5IkZdDCb8CpVQ
1jWXqRJy2npU2wDb7E8yAY8mSuB5nOyeuX656C01tND7xksQO+H3PeY5ROFqawIjNd6Nh1Fb/fY/
O6PyosbhAQ6QkCp1DOO9h2d4gsQN0oP8HQSaPK/EVrI73cl1ux8Od6qzsyAmBHTN7M/Jdlhi+rUQ
conBbqzEWcg0GXaFYGr9CUKBIitNeRUJzWIPrKMUU5fBBWcqUYK8jatspg4k/pagqVYMXS/w0vK4
MscziSuf574e7Cse5jl4H5k86byNI0F9NPA/tpmjaMqcKH6nZKQ4OeuQCyudbHQe+IE33ZucSWMJ
847wID7roXBFdwcKdmskDgEiAosFVseoKiYkofqhccQhhJxg24cdvcOPf8BiaSZWQXtMhFCddfOu
tGNlJSOEunR6VfbSPDGRNGcFAR8wRfvc30RFlbvmCm1C8BReHpeILahEKT9HbWraQcuJGsY8jiWE
GUZ7jpsxVxfPx13PP0Xu6eXeqNOAkME7DfkTWefxiX9lBumUZRU2vcpOxRz/DoC58aXLXIx31WPt
qOVA+ijbRdwcimN6ft0OPmMMtHfbzGrviOh90EkY7RaUEPMWCQ9d2/9yPHDK656Lpucb1T1m1Spr
rnO8jYrPUJJknzLm70rxL4qAC17mamTN1NTCvM3MfW434+cKi0VkZI6EBnh5lbqsqeclbyxvvaUH
X0UvfptLc/pjySGaCOWFQ+IZ/GwQjTiWKhgOAtMt8mXRxY9BORU4EsPt7L6DueFAv9TQrgXp8yr3
bv1zvrGYhueraJf98fliHxv+gXniecbzYOq5OBjtIThIQA+KXLXiayUCw7NYp3FeL1F6ag/zWTab
WZ8IvcocPzt/osd6epyAeuNuHeLHWCrg5FHa4Xo364yPyxwZXN6TWaOhFufBdBGa+kHkdaGLW5qU
jBkTp05BHTffW/zTqABtnObRyDlfD+oi+Kc9IQPCGG+Xfgc4Iwto76XHAn9CRL8gnOcmxeDjGnHG
OtA+kkhrkerbNc32lgPWV+RV/vL7dalA7vuACRybn13672MAcL+OISBNCwqSF+T4JVYiiU+PZb6f
nO52FQa0s8EEzeiumaXncwQgRXGuJ9nkQw8dV1j6JkthW3dTo0C7tw3XUP1EY6916i9bJSKrYwcJ
cICnlKp0UCodU4TXPuo53nIsGLNzuRN3XjuJeTYhVKXc4H2BmTAdyH/lAAwjxarS9UIzy2UxNFcB
VKWAdWNHiZQ4JX+WljWUS9oMWtzxWuequBEvDtldtbC4hYpXcJCYuBxH1+TjrXji6hDdB1g26QYz
3qHnAY8PUeYecm4IBk9WPfKHYgmimpfxZ6tcG1Xh6OxOarvXjKIBBNO9ShxgsiJzygxuE8BrTvGJ
UCyXLTEvk6GkP/qbmpz7qKgwxkRYH9ZLaH206cTXGcaNQnJjrQd3z80nYtnJVJJrLP36HeaCjKJZ
xJLg/Rg5kptePdFF5S0Z2WuD1ZOqeYOVT39XzcTLxTGjFq+miMk8DvPR402Yv5BvW5b7K0un390N
Tl0t9uCubbO/LKan2X+CWZkN8ySyEO7wcdXYrrJkD0yme1Mw0cAo8n8GkyO+7wga839SAR1EqXLX
4c3uMkXJzNdAwUFu6eWLwYxTWz0UImzJhhv0Xg8AiT0cMdVwLFQXKMwOyf+EqJe2mA7x6QnDfNRv
/WRWq3F8Rb7LYioIztBMT2FRert4BcnFj81z0h6F/UnhIMv2U7eveF8opqDBwsQNzg0ubvZWjfze
Q+uf7HJ1dCroZbZP5FOmZHynX5co0qdAkmwClt9CkXgXuU4yQ5RQaVCYlwBDlSepl486aI9aBsf7
RMXBp9TaFH79QDxP61IkMzQ/k5FepRrd6D28pefCVrJVWfzmPcvDjstZRND0lfxFGpkyns/7LNbC
OYJEehapdqJtOV0bw+7u4/9KS2zGCmEHCnsiqwBr2RAvnv+EU7xPRHrXDv5exmjPJAbFyUb5aZmQ
pL5P+0cXkDg8+TYwuqyhzcQJgPXXBcXSweEsMa3ruZRplt2lpMWGKneNr/Hw4P51S1MKKtE5+uix
stAFr+Hq/loF204Yq/KyrhmkxN9sRXj4/UXVERdTAZJ9fNjX9tPVs7Qu/XsAStAoiYIE/BKcKHsQ
ZXYM/52QX0sm9bk8xZy4viaQYIP+6iZRWyYa3UaXobsrHHWi4laxqR7PfBpw+LZAdCFKcVDEZRKi
v874gU1AoTyra61X0uBbIFm1PHUR63NmPqSbQOwz0+kr59GWr5MMHrGaVEgTL38A18Fdtxxd2TAv
6Jjfytt9o1u/LKjBjjqDLktOTHw48kE/mUBV26WI+TbXvhRk0XwUeZIqt79xbORP1rhfcGU5Sjzk
H39Iedj2B4af92x0aTlknx3drx78fv8bMuwYb5pCoeRvzodq1BRZmcQBUfvmeuCQ3AN7yLQflmmn
ppWZ/ExfK4W2cZi5VCCZfX6C7VIxI58XiKaIXzsfHJg32M9QU2SVEhFQ/HJ/IEhRWcAMP9osmbGb
KLESYEneesLSIm7KvT0Zko7mmKl5KnZRtA3ZCHFoQc9ruLJ14KBvo81iexpbOh+AfxjmUsH4P1ir
+/cy1nt4yuMq+ivp8X9zje9aRYYAQDW/0u7jrVB5KGvDLPeV7VpLk5Rq+vCDoJ8+FfoDna8JwZio
xCedAryF6GcZCX0tKitD+Duc9jDjCniV7aZmDV7dGOtwle8BfROsREE2ePZBSeNhvThjH/YArvZ5
L4MYaBuYy4ZSsB1vQUWrzDIAL08JE9xxtZmi2HxrCpRVMwpiOLMS9GggbbTGQOkB/nlBtS/3omLd
wycMCY0cKWvNhev6CXgYMp1uQDjtaJGcJCSflBz38uIbGlacNOrDrGMsAhx10NCFgvqDZ6GPY6T/
Gb7oN2HWVk1KRZRMl/2XNKMuqjUG3Fe4Lz7yXneSGq45bhc2j6XWjOBpogep+uORv2tC30k76Wd4
vKxQQTQDSe0AiAWzoRrVkkexmllP4UjaV23Zudqadi3LASl/gaRl3UMklSn7ZwO2Ps+vLsQ/GR1x
0pMLBMtXnFpiqGAdTlIAQWl29hfrim6GpUW+NCyJegpNHXM+0bqveO3jOl/3BjUFQa9aL2fGQRnV
ZFvvjZyi3mop0+jmuFmmmUAJDx3NqLZ67D8iBGDyrCUwKms9du7zc2DSPBdqnyDxmqce8+uVQFwp
sl0te9d67qI/qdLOBh7KaI6mJWcc2gSwbdixjlH1KWQWIMYMSP4/6bza2ZmbCCsrTxxwoXH2glpl
pv11GcOWyBkIb1hiqOI7rlSNi8Y/CjBiGGtSFONIn1zsHTGamRdzjI5xFmna9pgEkVCIp48F+H3X
Tbl5WVCsHBQDIuVRJWngxAJ2Lfr3pFdu08pvwNg6//bvsorqXlNVK26Xw0AivXm+xvyMqGMCbO/d
9YozQE8ib1JeUCopndilg2wm1U1XZxxHQLuFhjeGOFoBKcDMNclzFvL7N3/cGWOeOqNWUw0hYAir
sp97cZyRsos2+yvpQF9RabNmTOQbKLi7sGe++GJQmtmXudYRIfQy0QhTEUzjFTESwNyKe8+hGw0t
EPqpEBF7I3JbTmAwPJXZB6fD9mn7KSZZ/VLLI7TuV1UACPg0yIPJ3XYr56TmaDxM2ur7dOwVKPD+
R1IPUpnq9ewNzYvC3xc9TnE1bwuiIPQJv6mmhBXlisHeynsXYRhfDJpIfu52tZETXYrzrkzpswBz
pRdTMiCTxT165kQiEIA4+y9rF2+lThfPKA71VYGKjaAvnzDRa12UIRWvCOyJcn6Z1b2v3Up9tGTc
U/cVYEfx/qn/zSZLlkFuthhRmKLAuMRA+0aWDlYRf0Zp1CbySzm/+pbjMi/VJUvSRVz3DoeXpa0i
XLq3z8TL+GpSAhOQh6VRaQzjYRP4AzQWirXygm+VMtRXppbu0Vo+cdH6cD7QKNPwC1CzVqSG8DB2
HyNwPbEYEs85CjUzzEtpQFndCQDJE6MNiVHjyBDlOlAQYF3popP7dtYiqa9RkQVAVTe07H0QQbv2
+DUh8tcOEvx9+KXWu73LqZKpO7RCesRxhZ6azS+UY5+QZ+HZFj/f+g5GtevLkAF1KdbbZgYDqHq1
DeJonNzOF+DRcc0KxcJACueqgQLdmUDHM7JC2eBPPIgz2NKPBaqnUH4NO+bUw/TDXb5c0pEhZwaa
5zsL/TeX/cK1TIXYv6NVqe4VPHToWGZK19A4scZPIIVQNBirEV56QAZqNOx3FgCyoP96g9vm8o0c
tGd+Hzyph8B1lRSnr9OKttMIoKdQXMgz+aqJr3RAT2kkaVIcPkQmEKJnmuq9MH8q3Le8+EcfMe/8
effdbdVfDDrqB2B11XZV1aiw5cegvbnyICM99AQVTqej94mB56M6n4pGFxVLSvbuGF6qaiIGVobH
JUfVocCGrtzKjBHkEyAeyS9aEXn9TfJRbsk3+6O8LmcKVlco4aqa9YXoCj//t7Mh2JaFwCnnNC67
Pxf5iEoKrI+MDiRSh4MMv4HpZV0tcrj+zxXxi680ao1etxTWuksV4XgPws+LgT4wtm2GrSu2cJgz
2wiA+BYFX4uwk8lWqb3DbzmLbPbhiB+pXM+gullNMxY9fD2vJHvIYilC6bgkB9Z5NJkUnWoeAqgZ
RKl3aEM70W/QWtDpPYYvzpGm9nKzBYK89H/qzaTMnGRv+Vq3+lIKr00e2QHZfMzm9E4DAbjSni71
O1fK0UqJlS59f1T51lbTxOyEKYNq86HoLFL+hBUpibS0gau040IUeq5jzX2ZS5MjR3US6Yk/fTym
j+2MG47SyNqj7aIgh2W1EnuFiQrVA8kg66kbhr9+ewDHCse+JI3p2OSPnDtAl6u2Pbl+p0AXwjsC
HtTEX5wDBQQajn48yw4afiRaRLNTQ+7XGCd9lCUhVFgcPlWC4uG8GgZjmk/Sb+THI65Z+D2GOtx4
6pioVFrUh97Ku2XGykdzn4ld7LNqxtngsYvoG/CoQgKqNIydbbE3UkZMuHnbgUeYtDFy5GmVkjWa
34GJutePmOln2+smjqPD+a7JpFa4K3Cbo3x8Zmqg3XrAYNx1wnZA66oXxXpY/Yny1M1ItpQ+ji1I
8csTZpS8xByp1OVNxur9RY5UO+s6qbB0Hmp4f0P2luo/fRVIJGqWzrru3S3JlAzaSLhh+N4yjqqh
5xbydp8briOxMvkx28SUD+S+JKlAtmuhlxoG6mmtxygsV2Se9zCL/l5AO0VMPcWJSboj7zza8jn+
79amym1VpE7tBr6DLQ5cGt7iyDuY6CGSE44Bk9Ntz1tZ50hlO107D7a/r0DOn0qJS/+tV+Uf+iVD
ReSXftRb9c3bk+F6kZRmn3w/iL4wObGgkPOh2wGoisMiJGyTYO2f1hRpT+rmpR31YkiIXqCvisGh
RMNHJwqV88HYxeJVjd5ec9+bbftNXW2evvbqLM4+kHxK+4748S0ZiIkVh5uhaoJMh5ip3cyzsu2Q
32RxUpdkVDd31N6mSyEbUuu1QPs1riC7m0A+LlOh5B/pZJPMlYYt8STRCfsfsoMUdrrJ3mYbekOR
UqqNxAYkHgJrVb/aKBtaT5nFzhZx+Tke2Q5usWqQOEGaBXUwZGNfdbWCwtTlh59tbJ5SjXxGrPKc
TyksTMH6pcrKAHETcnaGFaId/T6XgdTNLlvaKvdaQ7/BjB3FkH6WVzGLaRdkbAbOaI744zMfYU+I
Gc2oH+73B9IkgGEXX/UZBJFJ/cJQSW49BCaDqjdgYp+uca2Zi9v4WPeRy8eDVRrGNHCm4YEwEqJV
1JjXXJDwrM5CMUDjgSxHzPvlQo1bdgN6MDBZHV6069D5NsqkCUzDMA7dwIkfVeF8qMtR6JymEUZM
HKaa4JAP3ifDvGcue9GXVBVmlwFqIjH284WBM6TLKZCOXy2O3jMoFjTKTRwFHixzqpr0dkfDQQt2
TYN9Ul+TFVqQo07fgUayIwhwMY/80XdrNXt7E1f2oLikBo1P6QTkfhY+DL/9jaqAsIn8EEnNIBEy
4etfOxp0wOfzaoUqza+E1iLm5jXp1ok7TWtvtcKO7m2+Ix0EMeiKOZjaAvW2AlKlbpDEREKvUX03
dG2lLEuLPWiix5BflyWXxT5mafrhsNiqpOCm7VlDweLA9kky88Kfop4WZcEzWcZkbOic1bNEpQnZ
KYYH0eAL3u9H/u4aNANnFNCMBf26zliE52wE2vCYcFR1p8bz00wtPunXku7oXP1Zfd99pZ9rRs0r
Qfq7CdPd1n6Zavjk0x2cGP1eEOIZbB9Q4uBIxHsfYEd8CVFjrIIw35xPTepJIDnoFSEsjbI+QQZp
tcWjyoUmGEHQOD2sU8e9NmbKIEZhbl4/7QaSUNmE+ixRcMbszmmYOHl+FYI9ZECM+3gWg8xY7vgw
NCmpZ9FyxR3396f7fjFTeg7DvDvt9q+ahOQQOJL7/KbvH8H+L0SewPQz42Ck/k5FoChkLp6RSRM/
Ul04KAtdAtSgs6ogil3vrZEXgYfjHxvXiI2iBPxfwjRTqKGr9CFACUz4IFOHp61glmKUMzjOSJQA
Rli4OQOTTVvvyh2ShtyuwjRsamjUdRcd8osvmo38iLX6iYGoWO1sEpZ+AwWxvB0Ru0hdBSMFpnKE
C6Bm7TdSAA//O3vWcKWtofl0lNt9hM32R+2iGORzMSA+SDfvxQiJDyzpJLLyaDQ9uU8o9zSGaenV
4nurnD695aEzlLFMghDykl2Uf9ip8mi7bz/XJZiFbqB28VbVXdNnVZMlf6Q64kyPxo7ahDdrjN8L
rCp8bSehfuCPNK50bKk4stv3bgQG9cB4QTjJXsBA9ANs8FwYx/dwSpaNajqDqXtFGDBmSKXSLwQQ
EVPMnVcE/im5Cs7o0kIvzKWY33k91HBdSfVlFbuj6AkncOcoU3/dGhPY3uUzGeVGYZ0ircQKxcr+
b0RFMoIwaPwnARkzRStSBW7y9b/oBM41soDri1y7GOa4jw6AvO/cBZ1ysIkK+Sko0HSX6/3Ws7Fy
lVEZtbymHOIH19UUQy0YzmY4e1AED6LF51x6JEllNqCqN1KB1PCqcltbsvnRXvuRZGv4hwyyOLYm
yPAASDWaMzMM6iBh2pRkPyMR/dPih8wcUCjdYdxW9MMKCVOnqRE2h8AA47JSQjSeG5rXuJ31WEOE
GWMHd/vQRrmogNJrHYHVLGXiyZRO4oIuBSIZD4GejZWlETIlybpP1HG/EsHMllpJ2dGVZ1wbWAY7
tgLg6LGp7t6zlMpjzJ0A37EdE2Ny/+1pAvbQRdGmKVZGlyShod7TwDcvFa6nE8wztkDSkSTfyPdL
YNwCzXCokWrRm4i6MQumcpQ0rjNekcMtIyr56Z5NjutGPnYKsbuIFgVezbE5eaE3OlqD6zBRulvX
tsYe89HA5WZqFLb0dItU1w6ETOZ2L4/jSa+eeuYi+Rq2eDuGp6gzh5d/NyyO7i1WMzgtiGYcohPL
h68fQiX6OTJuV2FTwJKTs+B+y+a09mTMqjp5X1TtVP6KIo4I+EPWZJqakvmPVcpJpSH+C7ou12Ll
jLnrz525xXJzsMiORHhPvYUXFfYMF3KgfUBDIwODBnZ/gN3cU+vdT6r+Fn8Z1pdrXUu2R+nHVW9g
Au3Upr4V35Bmyjqgt6W6N3w8590U5rL2yieidRxoUAv4qR1uwr31yxl4Rb9ITNGz13bTb57fmEY9
FK4ppzheHwNj64F9RyUFMLDxmwR4bxvFNWs6gP9jvl0kVZSBrnwtweQ6pUcWHtSYjrYE/u9q9Yke
L7s1zEU2khqWtaLr89vkmmuQ+QQyBDS/dB/fwmTyZXkmqIm+Tl5j67mCQ4drQ/HN+NEpA88x7gdU
jaBFuXhGcIMJxQ322Bq0ax6CpGEXBkJoQu1Nbhq92plkjAcqySQnL08WWbRMm/0Z8GNtPNhWySxt
8mouPbv3lnx6qoITYeCPH7n5EfRhdnxJNjq45Tjn9WpdTgV11/VQ5xHpPtZUalCzCnzKzY8FVMtJ
Ct5ihtdSAs8FrEz4/nqQnl1cACibjaQBDP7Ws9DRth/Lw9fuSMCRK6/lqCGz9X5aCVPh35/9G/01
b/Bee+JRMB0IrA/YH9BlSrj/KWsU1fO1n20vGEMsgYrCn7D7m0hB/xkjEbcR17L8IGNshNpYLOUT
cQRFAaR+6PRTZzyGekcUaiCM689Q6Wgv1S99jVyO0Qrk/xY6ltR4+BEreBZIELaBHIYgYZDH3QQd
Hi4TlX6QGR+wiosX3zcU8iU63lytFQz/BoIUn0iy/cm+iLJtBoOAhjBUNAPikWFUiARSDOpCUhll
m/2F6mVQxuWG3MFJTZPjJm7iQgR8f07rbzd+6WkXlq5BjT8+QeQ8Sj0m6UKFo8ABKtyT+J/GXp6D
uG2PMUJzDezK4znxgK5jWiP+W5PzQBa1Vx/nmMJ1eioR6soJ2+dYi1wYCfqF7L2hdfRz0hZ8QA2a
FKu401JmMzXqD9nNuPJmy0eBQkOPZlAuG6x9g3czvJv9fsB5+2v+b20eHoSIllMZPCEbaakqHbFu
UkR3yjJPI6+oZE4jqIuNybCHMdNGOhbOQBSpnRII+trqYrb9o/YFjYsiEeulfYJCE5IUgW+37OgH
4+S2Z/pVUli0Fu2WRX138jPBngGu0HDC13NY+FH/re3lYvgUUgLEAEw0dfswmCwF0TZH4pJVN4KL
U53FwqbmYeF8EVlwGE68CyZ/dR/Fzd/biMD+Y2hHPnen5vlh9zeYpIGweQnKlmpSbxaYNrW6Bkyf
S7v9PMpTGWcUUu821qls/6jP+DVFFzLoi4JNAfsvcHAOCEkmJrEQPWszOiVRtvnhZMw16M6uOG6F
sQwxaCaoIbDFzaxI4OImIdgPC/6TOsFwVbvjeZ5v2XMS0uCZ+R0QUdTdBYy3yVBt8gIPCX3QVbK4
n54VPGGMcZvamQ63qJw7wpWjrmmRiF+a9rTeQxbsoDVuqcETgC0aTPKu+Ho+YH6q1pSzq8gEQPMO
DeLqixMRcYNZD/TC6UYi/Ll06Q+btXtgK9tzrym6bOfJbYjtp8nPyun3I5NIU6hLlS5skMvu9HSU
SeaZQkQ7xB04Z4WH3od0ZLAzqQgQVpbuu1TBL9QV3vK0jS8tJQ1NUjt7lSJOHzibYiaDdBqDHBWU
kKMnK45AkE+LmRG9gIvH/phm6D/UnKZFuOSUhSsZK/c6gVU7MrTMDlK7WqtnGwpKu8BYf1CEC62v
BWd2fSrV1dScAgC9A4THs/GNuUnhmd1eJGqrUZxP9oiw7CpfXMXsCnWK3KLxmv5Ho/fMLc6eVgEt
949IkUL4jkVkntMYzsuBJeVQoLpTwmyMFxvinNrWKflSEBhsDBvcid5Xzmkz8kAweITwZH9l3YP1
KjegOCqg28Ki5Kyrv4T49s3GqM9HbuU+lFxHO9DVPTE73qXJBdHT+P1mjQdlSa8mrpvLiAeEXtJ1
hqKJL64yIn2T6BGwiCvySwoRLWmJ7/ds9Kn90e9QjWNKkdcPTlO1pdg+vDeYLByz/1oCv/3YcThI
dTFFjLxNooBWqPw1VlOHV2LK7CXT9BgtGupuo4u/U6XjXi2ENnTFnIpJq2mpyWmx7JN+1nH843Ew
E8O/Zo6GYKFDsRI2cLiLZowyZQd/aEoXhqtaSbadIEIfwN9+MFFVaCAQHBfTT4DYb5G7pwPYE4Vw
kJ1Ey2FXcEXQBenFL525iBjU/PmR1NqdHdDxpN0WJKHRcy1myqP5ozOmklTAZJaGusL6+28kGwao
dTaIymGnb2R0paSam2RTj+WrnOvDsOXjg7QymVD7DWHCF/L6zVaFy/q1iQENO6A3/vtU1qwaBMH2
PHZ5o5wn0wKXR/rV44S3rNKqBV9S+r9Y5dIlb6VYenLfpcARtJ01/eVpqlGI46oKTujRLz8JnhiS
tjJt53KYmEOvlfrxlSGD8dklK7wvhUzE/hqADDMs7diPgvmosedTZ65WKYEqiHD+6AdO0Rw5I8VQ
52rhf4KFze+/DWDDSTXNENCmDyyZrmTDKroeqfXoO3yvYCHJZWDaCbS481x7sqlvAiAKqAkkeD0C
xUP7XFVtxEiMhPJwNRAeQR4eE4N93pnpy866oxO827Var3viTpiYA62j+Kw/gU5tZhCMuL+YHFAO
peCi87kEEyRD0hzHa/y89aus6ToTOc/IW2jx4a5b2VjaM2aiDWgVNVcOXKNPo5VfCTdI2LUs3ZKM
6Qu/6416C7iTJa02eq58SOY+dhQKrdhga4VRbE460gjERWptTQAT01CuYY2TVZTXvO5XjsEpOq0n
SjHZ34hwXvg3UycU1VpXWXUD1JxsI/9qFxRKW2v9GNIBq2fQKVICc+5GOlgbj8LmaJNQvfZZHo6i
JsFHYEVpVAPoIONgTWWZZU+/maIFkk/dJR+0zjOqBWcge3dVhzr0NQB1oMPpciq9DdHDuUiKKZkV
AWdgFRw6z1UjAX0PWFPXamE+GVsiJybs++ljdiRzbyV31YGBeAAa+WfxUD89Ly1eBMJS9daS2jbq
Nf0FogbpT459sZqmBNHqaLXZu5szNaxpg41e3ntqF+PqkG7Mzb01vniGmOset1yKLA2B1h8mn9yC
7NukKIon0cUIin9pHHGI2MDbQwAWIOajKORhUT6wYAJie0JX1ES6QFwJXk/aHNeDqyaJK0JXn+4Z
FVDsgKtb4HC9TIcik8cnOLNgYahwKQHfJEUlTsE+46ziY8R/Z6Qz4HizCDIPhENnBkrEKz3Cisu7
Ab7wLrg/wdOD7SfQmEsUYgpd+w63guUpIOENcHS2CKZfSs4Xrx9PxUIuNA3Lf2lGVniY7ybQZ9iQ
MwzL2X7QYDVPtXnhJH1lyYe/V2kGgbu/qQaQB9AwKaeFkRj3j4+H8Hg1Ie4/r0eqHbhBwVDhOanN
oaLL7eKeqR8G8B4/ZVVKq1gP3MQYRGT8egXJKAb/aB1HEyaY59gf1mKVxXcIr/0wr7I8tHV3ecd5
uyYAvwdc323K78nn0hhHJFuqYopvI2nCWmr4OPFcE9Rj75/DSBVxF1GnIly2fBqY0GAjAYil1FeR
LpkZGwC/slpkKb1VMwPdxIsz8h5SZ94enEyCOZrnFxg0noTUEMPu5Gk8WlDIyK/aj+sbFQ7fIodC
bH/7z7bIJT/bjozQL+gqJ2Y6+seXC7BMFSCVWA85NRNgl5CZcvvPzwxyLNSQH3+yJUn9XHtKH36V
+d3Y/7v6ITnkG8TWKTZT1Kd2hkmT6Z+wCeSHgff7rfDJ/DHI7dL7xyjxfLKjQyNTsljN4aj0n15f
6gQUFG3+XWfDgTXdRWBr0A9cEJgdkLefzfoynUi8TRvz+1GrPL1Idei9rRzk3hsI67FU3QnWT8Xe
AeakH77ruAr7fxxp3sR0SjMaYtmd9dW35Ol2lBD69GMtw/JwKk6QbmEmcgTmervyzjkfZ76rKXzr
gOJgHget+Yt4UmLBS8F+CEb+Rr2lYt5HlR12oKahZhGH6xgtB/IOHFQxwYZ3Kv/o80kIA0eXKh0L
NDgcb8QZ4Dxu8qAALO/BlBbgAlI5wjbROs+HcdDlOFhqQYlNfIPrQ7icqA0gA3u1SWIhvIjFMKKc
djYJlwiEBJHXenVOqFNHPkRKlZEof2BF4yn4QozFY9rZw22pqwkL20+LyHBLUV9MHDOb0z9ISlvn
45Cj3W4aZ2O5mft/0KZ6HT8JJ0XVKw8NElRfzw+YI05CKO6C9XLB7EBoqYaCa7Hbf27jz+R266Is
xyDHGVzne9SqKGil/T+fHjInxjOQMr9x5cQlZFnhhHYkNJXNdrjFnPFdTV8SG22clA0UCUDnhWve
9nE+Rxs6o0CVl6zm77mFucSDTGV/nICkdjIOYSXsE5djAENn7vbvAKgAAQWH/IL4RFSovsUSnOu0
j1+4g+61orDNArj0aa9itKHojFvKlooSd+8qgW02zmLeqE05/5zm/oJKCL/bjYabOjJCu56LTlH3
qFx9N5e42ahuT+M3MIteghRbfL4FwS1Hj3fUO5ojci5iDC+Q9+oxLNdfbDfvQ2S/F3R4/BHLABwl
ays5CBkjCpHdbbKkwJsMF34+5mPLOt4M4jNvNpQzhfn/aTduuXFkogBfvzVqE0E3R1yqOGqYD6CF
Q1OMhf7G6qHTq1Ld4A1L8qnknX6EF/7JRxHVntVNLPMJJxvX3lMEJiHRpNdnwsq4dKRDcoGm86yi
HhAaDSmPPrGkkSwHuY/HaKMtNd/iQT9joKVE
`protect end_protected
