`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4176)
`protect data_block
yFTKr3qn864qomTWOK3YJbF3KpGSMjOUd4MJGfJIsWoACwc/FhXYysggjs6064dxNcMw9w6pvL5p
pj3T+1E3hx2JV4tLr0wfn1y00jIiub3Ml3bdruPx8FVVWgN20MI025Ox8aOIP9/hLeJlgSDy/RCj
btfAsXW+Z7UB2ozEubXNHeEXchoBR7mC31kD2HkLGtn7QOGiedV+yZ9cb8zLKBpkNMa5/9nKv/Mk
0dQsKJRw7UsifPs5tOOshIeN1ZbXf8m1y5Wid6XL1Nwy+o+b5w0mm0tkCISa6VPbHLxExcHtp/3O
dt79SJuE3uuNuAiUu/kVanPbxlvNLDNLOmu8493qgmpvHinxAK/mMwPdHJV3A1+9Ap118H4FFqRx
I1pXzz43dFhHR/dC37cHErjyzOYdctw9Me2CEFHDDJjXZ9MvnXnCCrlYoNfKEkG9L5Wd2i94Iupc
ENI4+OY0j7oD809sV3Ui/TUHfWY6AEddkFLuW3UPe/n2uszs/WsTNWAsJMu97pleL2k3ylc82tR0
DR/d1X7pQ6TLlFmf2WEdNG1nz6Z2oHlNvapHPqoaulX7aQ7HdLpdja4VZVvP9yzVr+uFiDl4R2YB
QU8TuDrdBf7R9jZAxB8bf/8MwywcgaJBAu7fqZrRZpjLId9VKXrA9kjg9rb/72vy2Lt+A/UA+xrw
/Y1l+bW7bgIKaLOZ0lVPMtKa1cbHfS1FEAa3SY+irETiVZtxt4lm7VfJxFD7Hm7nrAA0Qinu49vw
ATC3gsWPGefDq6QP1n9yzeMwagVQswcBr5MAre21tTIiNdj5RjaHqfBBeRRWCGv9XfvfqLmCWiJc
CEgAaIy4K3A8w6DdomdcMG71sZVOAOHv/LOInGUyjaZe5MLJU7shW3fNEKIUmALu3jMQ114P3Oyc
zFSYDK32geFoCofFBrdEDDTtOcssUPRK0RlywwuXS2y5fem9h7vPvizScOYp/wbTIB0FerNIXxqE
Qh2SaIOUFSB/KGnkdFaSX4QRpVksSK2ViCSq7MwychPsA8rN1vT4ixypAihDIAyMEwXMZUtkEv+h
56kUZK2PEVBLgBVJADcVGXWdwO57Xh2J9qE+KeTP4cg3I8uzZW1Ey8GzJN95lfS0Nxcl0+xdofkw
7SZEtXrk6Y20oQvoMvdmcOvgCypkcKcla0gS2zZ8Hbr+OuoTsWTkA/8iT052HjI8B/vTaQjumEMw
LHSOEuHDwDrEad/tIBTh5/hD2WtlCFbTPsYY5YTyrPsWiaKhKJziSpcvGlR88jLRROd5BJPmmBAC
uroaJJ1IRfDZ+Kd3X70BRM2JFTdctW+IJhm+nENcBusNg4fwS/bCRWVXudFzLWNv5xTxeRoLiWdh
iRmGKLx0ty0V90NLSE9zm77fiW0arQpjSx8mMOtaPI26fhDZMCFvx6EWI2BlyusEHzC87g9wtYd9
4jPoSP2XCSWf5KpvAV5rebD1OhED17FyZmY5kcJaR1406Uf/1EIumiHKAJxgB3YlaeGx52LdhAeN
nKkCKcff5rbs5IXIYG9LyQwB5PVjkvhMFYN+ttguBNcM17WRCa+rfZKreAv6loi5i7MOwO11YaYM
wFehF6mY3PqUqxduNAc/I+GmRSpiRfzaBMpuv3F+XMI9z3riO8dzRD+1oScddwhRRVGEYWCpZ90Q
6i5us9dQkCNjw4V5Yaj4bm7INczSZwR0Jv5C8t6I2JOSPhcR9RBHQd+kwz5RaGscevZI1PW6MwEN
Okt0jS9G5fvsHs2mWrZmhE0Fi+o05yF5bLdq8WLyAJja+IfttxU3HW0MQTpefcuh4qoCO0yPb5pd
A5BgVqLR1UNFCKJbvWB11xBDySE2+MgjffRla/mwnrmIqBucINNYO2lkD4HPPNnJ7PRl8KarP8vz
a7kCa6BUnK0bUyEbusRHL1HDnlhMcaZuhaJTgcn+2ZMAk4Vqt7EfxNg/OAc0jSYSttAi4XRrHfNb
Rfm5CkDjXx7n0+YEJIfsaC92pdGtTfJbCfQVWjzi2tjVgnPzYUFf/Z3OfigjpKz8+5gMXMokU9II
gqaorv0Md8XyvB25oJ30gJZWeLkb8OdOmgaueQSP+JasURPTRltvjPXjRJWO4ZsxFAhTKqmvGPLb
+e8+OWonOasvb/aL5D5KI1qOGzrt8migSlISCfZvKAui27GgFp1QCP8aSabM8uiG4mcPgqkSoFRa
+Ehe8Yc1eVHDW/WWpkyDTe7USKtWTgQHZXZ0ttfYbSvIYa1SbHhGsZA3xl8wTm3pQOFP2yHdTbZH
Tedip27XA5sHNlUSd1JCaP73bYREWf7XPDRNqTtoteWiGcBUBV/YVl5/xac4uZMbsnGncl3JNN/d
0I1xe06tg3TLa2nq45hvaVbX3qJN9l1iOBzy99hue8nqKWnL42LRDeNVeIKMENarh5EGc77FVGrf
vhqnFkvv9qYziu4qml0rJjOs1yq5UmQezusRmXl45gSf6YAh5RAxAOdp3wQjWa49mnEwG5CRwGVD
5qqunLNq05j/elw5aATuQFua00kdqDL5IqrhAb3y1qErU/mYwDTGOc+TBKsJv/AWLWAC/DsMaNsZ
A6uKVM6IVl4MlIKjQPISPSh/+sFuZQPcjoHImkPg39tsMNE6sRz3A0ISq4IxL3VXX//R/tySY3/k
ZlF4NxpZmyW1ZWm4hg+11htGigP0YZF/9QGGX0d56FquJQMtOxk84BLGJelWovk6SG/x1TqwnGhu
qP0Anfqs3oUFtig8xfnCJHqXaX7p+XFY6Z15ZaLQNGIsQufJcQQS2TnFQUAkpJCYISaXQLsiDbQ6
oNihJwXcepDer9jENVueQVqz+TOwRfcnW0U5S2b6m8+UZicmC5sJp4dKthUn+jDPd6u5HKDvqExb
EmybmXzv13d9f2ZC8lpUGLE5Ele6jPXLb9gPnB+BQJe3bsn/7FnabjsU0L2gl+VhziogKeZece7F
qIRldtmRBLhAhJwecDK2nORin4f74Own6iZQkihj4dEtRltXYPJct910QQckhtBWfnD3ZQTmzYGX
4UI4bemw61VfsjXOz8AgK5nRTesLxA3kqV1OIEqiexCAbUKqTdBeXBbjK+KQYiWzcq7obwIhg/FM
V7gOYLQni3W7of8tQBdhhecxUW5xT6I7fYf0/ChZMYimAtlITmvlM3RiD0QI6PXLtHBj3Dsyy5xh
cm5DuKPNym/UaPRKskWUnHTzkgvOOEMjw+t9oYS3ZzpQFpC5mQxUr1cblGupiq3i1DksYAL1xyY7
ChembxwGCwV2aBpwqFjQObl3fEJ+qutTixwU3alG4U5EFgoK7+X7Yn/OzmVpHsP+l0y8jw5dDK7q
u726llMQ69nPAjziv3IWZbBssvxA57ed43SBXz6OqxJ4ixWEk1PoHmy/6LQQ58YNdaW5foGJ4k/H
EmJ/6XImGKFNPw8fo/eh4hrYLcTcNbpjYGbxrJtYpCNfp/eg3LB5OOgI66xqVJjZykvNtBybqOjj
uw3YZW/WY57e/6H4QU5fWZ1Yw7A+WZ5jqTm0idUZlKjrLFPTgKQlw6nacFY0SJhyJexn/jyr+Acz
2mNm4scb5cae1MF1q23q3+LE1Za4mEPcXnjBqlP3UA6oig6z/Elt+9CRzfj6tHB+rxMrpAAeDVZX
2139XdOCt8nc6tKnkMtDbS+8pc2VOJB5fMqcKt2oV09mpZUvQwzhlmd/ivt5+xKPB1UrtpB/CQlk
KbWywbg8ONK8v8K4TZ7rBwHbo+Hg96FgFXSo/zX8JWHMf5GDLSWaySq5CKjEbUFZVgCVmzZcXBWw
S9OQH8FKotXg8DGIVpWT2rACwMe5ic26smcLUlryhyr3zykgR05vb2xHjWNmVDbSAbC2sa/+5TkL
HI+yjl8sOQGYEzVQgAa7b4N8jqFUy1zdQ6R3rcphJPRkAQsShveOmK+LQkFC8+RT/Jh6qwBg1UtB
uK1UJNpDB+eOT7XoXTReorZcKaA1bcbFoRSlgOdWWQlXyhiGJhFAZN/GazJzLQGQZdqA7KbPAIjd
2Fvh1DkGk4pjAJyLO/mWCtHRvVrQ8acVzQ9bYEWy+eiBW7HMhizDRQBPyZZp4ZBD7tLXg39GvcLN
9a7TGdkeSvDFwHsPRogYjZTzQHsEYa0V5qgNYMjptR0XhIIw0Ke8iU8iTr7UA6JcLLaJqJwfLMTD
60JMl7E9B0nDMrsFOQJs2288z/899z94BQZe12vZP7S0rgTz3Q8WZnCdk1EVczT84x/YmOp4Rluo
Nfh4g3JC3q12R/WweBT++QL618It4IQXoFDSOeBxLUaeXZXT2qoNs0sAgybZ59mY8jGnzu5r+jD5
91b8I74Hy5PUE/FO4QwtHMM8FlAHGgXAiaWopRIZmrMOnVnf0I04t/Eal4/sqTv2j978ivLNscJb
vHvECPT5khMjzkSLO163MXLl2HalAjYCoLC4DepqqEZ8oPCCWjgQp/W6zBRcJr8WN4iqqoEKDqWe
sVuLI3DpbOAKC9N9JxfCjFgRSDnYqTQWe16dQYd5Clw0LZFoE9ngDUvuwYENdpye3HJ7RVAog7lm
8aAH+xV+tI9XW9xxKQ3XNbBHEQiSrK/Q9r+MBTAdHMWd4EgNYK9UrShths/Da7cpPwvX5mj4RBWv
MI1jAAhuzZ/MQ6ogoJXBqoDfI7wV6WeqfcsXscR3zJKOCjLF7FZC9VXFp3j51da3kDkC2zXRVy++
wLdg8XXJxGbI4crysdvRAOSKl1yet/S2CoB4b3D0ExVOBy8KQqN6m22Tck+kyYNBcvSblsOUsSq6
MA/LoWxSYVbcTmL4XYiJj7r/3V6GdNavMNmr0KUmondCdu1qkGm6HXge1Byli9Ezf/9veLVOw+o2
lURKpqQG+8h47y1QIvIPaaFxywoAgzkZXvwg8DE94eX9cq+F5qTqlDAN8wQjvbs+Lb7H1d/hieBt
Z8GoROB+CoCgsYa26Gra6M7QjexQrxHRXajHXpfRDNtR2UeMZ3y38ayGWoMT6xwJrHaCTPqNQaOc
t8wLstL/moi2qbfjKMjbD9hFbiGLKVkLxvoP54C/FVPqB5Imklbt+LknB0JdI+9mKSOHzxKDgCs9
QJe/3YZlrqblnP35+clTJOlDW/D5WQ0gJxvBZ7cVLfe/dCecoGRCcmu3csC3xmwB9ARZJ7sZuccX
xe88m+vtjlgH6d7He61RlubtooVUW5KH0sM3UXBZ0Ge47TatehYX9eR7NENlMZnxv26JaW6fzyE7
P5RxzauTh2dby9N6Blz4hJaeZL3Lnd3dgis+fooSCREEobwtZJtyN644x8Bx7Q82TKtNDWf36Wah
kB38cYMfnFWPc0/g/0+J4AtUBG0Jxnk4f63kevmgzvfraln2JOkF9wh17VIdqK4vvExKTYhU3neB
1X6P7NuTGjJsfO0u0mJ99NN30UKE280Fw+l4dCL67QqwVyXgu8+bCpEmNu6dAelwfNTQUFXEz3E8
TCuMsPM2pGFp5lJTwaXeAyAblri4AIQIiDNQrN7AU/FnARt4MYQ53u4phUiLGRD9JcAuCNQmiGlU
inZcmQUnWndIBeKphbaf
`protect end_protected
