`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
/yWpInKArsVq/Nno+CLiS/f/eV+RPe/YY5VZMgUUlpL4967auqOV1PS6wW8MrPYBm8vdYb6JbGe5
eveuSUnrPHhl3vNu5ZXjZe07Z5spxRUEWiu1+uMTqs8rPfFuER6Sn9ZNqaJaS6gCYn/daTSiak5S
ye0T1PCP5MfcweBA3NkzmpO8wx7TEI2EyUMV1pQcF3oX0VfDY7ZqbI2JIlTuV4v7G5TbDVmyh5Nw
S2wWxqDUvd++VFViLXbmC/uW2IOJCegLkm13KxSQcqUBErXwGvdZFfvW9aYM5gDjNWMWMr+QdH0L
Vj7JgVmuNZ3D/b6B3xEEPgqsCVA3Y06NqVREdl7+qojyLaijOirjw7h1mX5Ci+Yq7sinD7FUMgwQ
MNeoCfa6FF8sVdogf7qEE64KJD53wQn9yN7EVpWDciwmruFS1Maogq0Ba49l1v73RM5nz3toHjFk
nWAYo5RTFMPlLU0+k7qq5f804O4bhqJN79lIZQgZvF0oS7aEsmjrNOIB5P3CzIKNxu8V0FWK4X3b
mxxenlQC3haJ3Cofxy1QONJ3f1Pn9xD21f3ouDMx/O1ArbIXFLXdioMWQ/nu1mj2K95BXVJjFjsu
Qs32ZBZgkf5mBMmtedu3QpOXJJ5yN9P1/gMKJopX+17qCEntRsst1WJ0JrdSesAnb8PxUjctizCs
pqcNkDNr/3CUabUPBvQXhBvn7PsYilIALzfL4QldS9sUFbE8hTtZVOEliwKznWZEE68xqA+ON2ON
fv3vdPN9wgZ6VUffU3YY6qNgKHPVRxBgR1iuY45X8sGo8fIDRNn26MzKMXZDWDSatDUk5dBHHfwL
XoKOmquhh+OCJJt7F2nv7BURGGW8YGDXbrj6FR/hoO3qD0fQhNYk6kL2ViAS1wSGfn/oFCfkhxKw
Qh45jOS1LDW45lmc6uYs17SVKxZRAbbhbz6jdJkA/rncHbGJ4DBudhtsFuStZ0JlFTigoXpmG7/+
JftJmRWiVbef2msmIZgPCQLR2s80Z+GlZl6eNPbEfAwc9F9CrOLkokWaC/dWpELTcn6sXqGO7hsX
V8zlnc5akRWisaRwLbKA8QFw77SBNYftTzo6VLMqaiYK2spW4GoyYzBR3ksiP9W69Q5Cy3gzLDEg
2/LAH2yjBilYLNvd/ehwsgstV2yGzlwmxUDeAKXxhsU6ZawffylR7uh9a2x8Haoy5plLQoymc13I
Ba2di/TcS12DaDmVmytjitYIQiJc7+EK7SJOJEdpS8F49ggNCFkptx0c6WRZxaGndQGI8sXZzfcr
VD11MD7+hsgNWglAWnfIMYuqCHEr6keVctlstnoub5x3ULkdiDJjBV8n0vzTqSLQd8NgNT+Xuiw9
KF5chPpE3s8NS4mVE5rVwOVyKr/eEHcH4ogdE+wdhBAPFxsGiiT5ToLHvlsWMB7JvjMt02ISzY0l
cCcpt7FjUvCQQyPNqAUmXWle6YPKCMErEXzjeSxTW5DLH/fRtQ3Rjkcw0qBSUu46EY+qUCcgTKGW
SILpYwYU9JxqoLC6YW96kL5mLfz61OQZmd50PlmeCQdjOmHMEXDlzh33qoOqAWo9Km552mD1Kl3U
HFvxHU/Yiz7YDyyeAJ3RvIcrVmOCfFTzAU47VVlf/ntg+q8Vyf85qDlU47XXBeqQ4oPR/F+w2Auo
m0AYHDj6w/OgT3Jtt03fx7mIRAhTplx/rN/qq6csBFhrF0zEOeYEZOfizc9at55NndRjtiZBD48g
rMTZAttH96nHmmwzFnBn19wOcHmoPXHEVZ/fdw2WKayHOSgpmCRcxBCd0vPSfgbY+CskXlVSRdDs
kulkYruJxeZkdKZBehiIh1XO+B5VyIa9l6HIdjO5ykqCH7FoLXbu4MNsF6LyvRyiswcidzq0EeGj
V1/L/yfM5KChdiT9iNeIC3IFw9+VIR+wFU+FcJKl6pDmODrNUFQ2UMJd0cHvMDFmRBfR+sxVYk/r
ctuY99QOOWUVY5nqjxlV+mb9Hl4W6v/idQVDLLv7kLENQ3N7XqKdaT4OdapGh1NW9//5aa683Tyx
6QiCwvdPfMCLsRbEtwsQ9zyH0WiIunrzfhqKqPIxZsc3dlmpTkZwKSpu3C/7CWWxGOfUWtBJU+hn
sZzoYJqhi2y6nQ928e3o8oUsV2AF94SfvvLzhGARsrxWI4X5DF+C0irc13dWAHLWg+LTxZtVDIB2
wFL3J21PumQr5hmRn28r8Zt7YRpioEDzcWAFXdA/4utI8G/zXWBZAEeodteqhY9zt+lpKm6EmrY8
7iDt+KO1STp/i55JeDCT903ZuE+BttRO9EACaNMYWnAICWrBmIMPbrTnoc+5qAHbHN9qKp8Xti62
JU2GS/FYYt+/CkpM9Mr0U7qL4zy5N0BI8yZiuC8e/kJUiDka6r/A59SATbO38ax/hARXqwL1P9J+
w7+fQpkBUTD2Md7tKvDlaQEw6sVBsEGp3G1FhYn6KwEyB3FXTxQlu9PmlEwJX+slp4EQIBfOFn1a
v+jVIcdLh+0aFjyop72g2S/pFSdj1YoxMrFROu34n08Vk30YazIz+OweUzRqq40OVEWJryqgJEwe
vGVbl3nJnRXcEX6huMInU8Ho/lBfGnCFx3FrppW8XEr0f0lfSoaJ3RyNhQr7pbKcGfZXyF5G0FyO
JshwFAU3O2/MgN0IIL+gz8SvYGKihhjuWVdiLinI6maA4fCS6OKZPOYMT+Hg2V3qobEbO43pVcP/
hpDBYnYZ5QjU4Stwu+24WXQ7TE8RyYpCQfnCwqDdtE7Yx0fvN6L6Be7hREERpFNly2durULKlJ2w
YGfzsDd2Meq0Ln5Ox/eeuG4CCMBlz2DDJeIbBnbBTYUfuVp/xqLGlHTKc9Gzd/uXkwsjBDkne2gr
dTcH+lyYABGSFqn2ZM6NEX52w1tyWJgpeY0pGe4qRUHnvb/6pPgzJs7T6qVQ01HY/VNGMV0WW4W6
eNYViZPxZ94eHBtM2Bt8kZAuY3OuU9qhoaqKYOxqPT4895Nney9oVfswdg8IraOuzfyRZ0f1zh2Y
NhaeV8EdiwiYLMVVysQz5UtAFsk0yNagvdM21BIc27ioaj7oX+DP3Mp2dNLdp7vfzqJ571RA0Djn
1heKYqfMVnwtEHVmhglAWUosdEqLN1juktCDr030knJxzIxzEL5gCU2qQmADrkcdDvh0NYa18JmA
R2Cl3GekmaGbdAIv2v1eG+zdJPxJHseQwTdn0ZMlQf9nAQoMJLG85M7nJKuKU6bWbzgbS2bIYw6G
anBCotHZTlG6ntWdmPXjnL8ac2/mw2E/IVh6Dr+9hvDTUFJyYB6WEbXoPfJ2H5DyvDZStyfuFLx6
E49oUmGclHwhECxlXKQCX3rMN8I0hZtsDz6PRujQPmRbQaBL+PkwIrvaX27UUH8ru6HCeNj2Im23
lAm/dbdphfXynHPuFbptNxent+AFjyLY2g5fIUQe7IwbtQCMTR2LQGYLBARvNHQC5ESzo6jrYZZk
joXrt3JE/GGUUVkGNwwQh9n7Rk1tYGJ7Aqpn00MbftR2bguhOYs92qdJausigkq7+DCHbng/kcZL
EuchTRDCGeEadOgsSmBFlfhOiTZCM6hh1wzSfoNCSxB2SeWAnNLREt/qWazzBQhBmimAWMGGkIR5
+VKg/wFXhqZyaDjmTJ1Trjf1lBwp68bgWc2GT8IlkRx1VAKbx83w9DOS7QBZqwJ423JJouWfbDNC
FEC4OVc1AXpAYxrEYRTORz/7j6Tv01NTISCpfliKBbVj/7OlcGWdfDpPX7bDsuk8y0EQyFWJ2+SI
+adOHPCekMLa+lT4sLoAZKD8ZEnVbT39qKo6FMY/Y1CG0/gZwjDeWl6vsCYJvizT+rS8/5G4NPWB
tqHkJ/yFZMWVq50FjNlRDt+DEm5SzVOouJ6SWCAM053KtrU4q2Jn5Usk6I2L5dB0ndIgzMACQkL4
c2x11Ju8zI5JsoL39Tpx28RD2T5hjRTdezB7m/LTcuim6cdJ6QT8NFpjTOolXEVri7bkfILc6mbs
TteXCsUT/t6VHGfv5j6BuMP4lUIF8dCqN2K2Nsa3Nzcuy0zn0y9EZ5eRsRILD8c+Y3Wao9IB26nF
M8BLDSMhrXz5U/ifLKH2nTdQOU7E9sRwzodcKKKCNyaReT6TiGA2hrjEVrHR83BGtVF8S5mJPNys
teupyN+Ec54aNiaJmyisJlzLtwfwB7GwhxpkR9q4OmY+2zlGURXGel7Y2C74ggzkqLy9+bH4egOa
bQTRGVtyR/kHTBt8czy3dsZJw6YKoaxaDqGaw3KijrMbW2629mVXXtB37EghPb8s1B/8Fvuy9AQY
17Ffy2ixhFSFzW87pX0dG+GPuaTFV+dwXddb7kwjgTdF17uqN6QHrx7Rq7d82IMw3kWKAMdkmaZV
ezW4gK5dpRDNSwY64n+0V9HxmJi0T4ZGqQH5HTkhxjA1KCRqzyoAQ5PPILWwhIYwj3Z1+VjyCMlB
maZ5pvnfHxgAFbWW7a6SK3NECn6729poZJWZGP/f0rPaAt6sMtxWU7iI+KRC0gka09W0UZB6R6BT
A9ohvQ0NCm4x0hKBlOqcTiY4Ug0YyD6t/srdUHnaWA+OmsKz65GtVWkSJuRNWRyE4zQtjRLVMbmA
/A9pjiy0ra3hCijN9aGNDr0ZcIy9M38bpnaeRGKpnZyx/k2JSHcpNoPDqnDO5h3wuDCedUtwtRil
M+CkdEaN88q/K/qDTiD71+wZQnUJuM3G6Q7FnF9jvRISIkv/w6+kkKSh4NgG1pibv5BOGDXQfV0m
FoVlnid9ErJzzg+xu1HUoJHlJnM+qd6oLS19nuiFjgS6zaQejc4/ngPo/2H6vgxk4YvlT0dd4wvi
vLLu3b0peAGeVlvCituAyMxvSawiwNBfuqJYebP/I7gIomoLogQIwLTF2kU7xx9bihqMzX12seph
+4kniYorYqblky9l3G9Rt97ZDCXA13qeM+Lrvt0YYWXEx2XlyaPPNvCIwxz4nVb3snHEOsjttWbp
9v/iVV+GJGIT8TOmM85bP6o8BJoeVqbNR8z9qsgjACEQgN42PT5HyeqwqkkRakQ5HYlHaIUDrPF4
4oFI84afFf8UV/ALD7E4ux83LgHfRW5k2Yu0F4a45YnhqBdqLF8yKRCNE1PHPVnY9j875pFwX+LD
s8muOOu4te/pKEpgDMsyKSON3qgh8C4oWODFIpT0kkqgy8tzYnuZx8egRe+mcDWSOD/pFzOK9nts
wIAv9RZqtnUefrz3QfExdTQh9vPeNp1s3R57Qm2Sf6DpfPgfdxMq/nFLZrcrxOuV1FgftK1vTQTI
GcfMBKjDbgDoUt5GXsN1oS3mhame0w5cCK+S3+1nTZMX/BiTh3Tr8R7g3bVzVbDcfiBz8IAtCPOE
N95XHI5ANmB+kCMBl6BtPJzt/xN4ZfJFvpuH3zG1nywLOMmWbGaLraKuXCl8UYsD/YiT8L9U1ROI
wj7cong4lczxj6Dps97oJmLj8W2psnKJk/0qPecDVDECfx5N0wdhhLmL7IWqLoXbxKA1+l1IoBOH
4G3MlJwPMOPSyc9VDwaIh6/5HLKszwAY7V9eSPyiCdfzhFpgvnIdiyTfwXt9iq+rrLFVUhnyUJpz
URs6g+wv8D8lHgdXw2WyHlvOBGW13tY0HEEKTP9KCqnYj0BtOSOAzdT5xxvZubpZobvDcYpMKb/r
pFM22l7rNt6fXXIGKHqEcS04yO5jST326tXRjCEeR7os35UAwv8dw5iU56E7U1AmcnmVOpATn0sM
q7soXZ0LuLtUBPuNcccH+dfvJf0kg34kZ/tpsf6mObJNCPH+7+Iwi2opTwUXHPoem9PyGNLDZMfG
ELKDxfba1eSVVmg26eyUopoZDf5xtNR7WnwkYV7XwmC9AZ00kHcTkdgdhckwt2LPhSzEuLEjIPkd
E7AgcpSAxUhUhXh+7PCF+mV+qN2evBiPZmy+hh6VkmCPfUjqBaUmD3an5foV49mAlGclDFh+cvx5
U+HKz8dYhZCBRmeNTjsSCOBTjmr0+vQOdqUwNtcJ7z5lmrh0JKxF7MYNAD3w0DF1HJ9jmElQSXQR
poxXOMBuivvct5Nq5VTzBfILY+Cgty6YLafDvOlXDABOqgo0FIwvloCpmAKCojJ+53CUudKuCHbt
K+uoJ1NCp6jP4D7H3KQKCpPucs9EkQWiKOEwrrWrlljSpj771J/h4xuc+zrN/EGA6i5BEvv55AlE
CaTZZSppZ3w43B/FibtF8UITz07rHXdFZPl9j1yUdvPIOrsw9IyDLc+I1Ii2H/MHvxWkPNz8o1Ke
+loVAhuPDD2ZaI2sI3Nf0BEJdLDCQjCSK5J8/4EovKjfWRICopFbg83lXwT6vTQOEzflkLCFe6pt
xglK2PoDJNLc6NTZhLHcwToyA2Hzhx22MtC9jmykqVkoUVaLc9qF4XBAfFEfsn8IIDnu4Ap+oZvz
K8KjzlqlPTvoeGnk3YhlP1rxgzeQJnElO9FjiRo8H1jBBbK45coa0z/CfyYfAo1NcZorlKUZlfEq
hjRLTgcn7IhtlbUXQ6f/Ga+UiXEpw2hEIc7oKvOwaSy46AeX/qcWmEwTy3XeTnQeBVX9hthZy2qf
NFZKiWM+QAA3X4I55T0JJ7JaM+d8FnCnFr/pJngFi/BtxLVkK8wvXZmDTu3ujOZkk9Njh7uEE/yt
8G0PFAEF/iNIZ7iEIhw3txV16Ih5PCiu26k9byNTzx78FNG9i43CmzyU35ONftIrjq4FDALYQGgp
UNb8aPgbxe0Fiq9Py4oT2GQGF0pPveB9d0hF06Osacwy4sm3SrM2aj8rcEhvGX9AdAMVo09yG/S7
xvTlxfGNfqyEBcjksUbzeY/US9ccH9u3ExbitfIhMufF+JuGZwQerZyuBa4KjN4s0V9lcDU84h5T
FXvyaewblTJJnxZsb9PUudtvgh+11Hndg8xacz7uItWOJQczhuvFcESOU5nm/jfy23C2RPbpYjEm
GzfWPJvnMBWShqwh+VG0JyAJ9sQJEyzs9BeIPmBL+0ExnAtGhENv/LXRCxKbcGt+eNpLV0ilXjQ4
WeadCi23KjB3i5+3vgCOe2EfXn2V2pkGpor0edHAX1sw0TfCcJqrzJDQeOoQQWWm+DDdeCLR9XSj
iiB4afJMU1C7UBq1fissIXO9AuLeCFHEIP1ZCLaMI0OoeRa5+iSqmXq88G1UUk33WzzbI+y1qHw0
Rkg1N+q2cXQdFJGI3gNOyOQ7AOVxWgDhsVOTI1Y3NfGMJlH5BpbCeoIS0OddaU+X9KHKEvaF/xOB
8uTzk2teIk/2PQqdoRglaPuZpC9jpv1/F3ZWL4bGrkn8okfqfXDs+u3J1TVvd5Rq77ot06XdVDpO
H2EtpDhQrf2iD0OjyLAUZ8sG/NybLDUBc3ww60x2Q0i0sLrEyLvlKEtz6icV9MBcEHEhooIjlhwd
CSE2M4v4v61nCy2AGcXJMHdfev5dfdc3oBFYeEHDWh5H/EzvQvRw4PyvlGAAbfbaHlmUp6oSbw2+
uMEOwPWzh8t6LrsULQLts4EN4gEEbdNTTDOPSDodewdnAUrLtLFksuaTASJRCLqTNDsnwdke6UNn
nQdCHI/Ll4zQUWcU5BzX6nmyQ9KJ0Hqm4snYozRWS43CsED9u4cOSMOv31JV7mZP5+1ZW134Ri5a
tROY8usbjy6S37XJerlIf85xUQQ6Je9YaAW7heEzsGmOd/4QCHVvZGU1t0F1LfsueoWmCJrYim3H
U9EmBZdV3psqvFXY4CKrQXviJQ4Aa8pljBaKU20RIfDymFXrhOOVuVJV6CzRUXJdKbWNfygRb3kq
D7g1CjGUm8cALUA/8OMJdBtkemAwiZAIwjlVhyDv+c9huGmaIax4HTIztYNoAXhRMUdo3jYpTy+Q
Hyu8FhQf/q07aG2qDOXC2Ot0SiKdzD82LwNWf8xo+buOeYhHOtPbbg6CsVeyHU1OXGm5HbVxEi+u
QNJuuKR7ym5bSHVxvB0fVBLdGT9DSyFxHfwvxjwwNDSg89xn5XR+TzWLmrkTS7AX5CddJBtsfkRL
xqbEMaJA37tPcgEkDLRkUrE+m+8FejbdZx7+2paTpHNu1tlyTxmcpNtcMhODSQnHj+eu5rKZpAZZ
9dq9PRDQ0IS48hqApRLLPPmRPDWzS+kocSwWz0o+ntybLqOS9hG0vgwJrx2Xqz/WgFq6SFSXH8Fj
ItTXpJr+WIkdtXbdiZPzxj/jXIV11zNpFOkIfw/bmA7cDYuQ25klZ7ZhAWzqj3J6XEk/8xBnQ719
cirSKidL//97nfdwJxmxpJiv/HVEthVEHxePGr11ggQSsN+7mydF5fcHlw==
`protect end_protected
