XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ˉ}>H:������I=9�Fh�A��Q�m�y�8M�^���Gp�BS��k	��ty)����W��p�,����
A�\耨"�HzGvdvi	ɪ��e��ͪ&�)��`J|;�C�����	<hd]�a?\���%mF�k�~��YB"�B{�p�g�{_2��8� ?��������p�fk��+�>4%=���Xp�^��s\<�@���633S�P��*&<�B�hĽ�h���Œ���3|�*����f8F{u�g���݀Q��"'��L�m�����E���Q2ϗ>?��d���� ̓��c�Qw{1X�屸�*�)G͊�k���� �RHV(�����=[7zvb���W�Y�C�<z����]���T+�U�ş'������9�ǚt�ж���}�p����^�tF�b<CEU�"AG��>������v�`���'F�b����фSH�۞���9�����	��$��8/فL�}���	�A�\M������+S��'q�KH�T�T�~R�7dØ�t���J�oB����t�!���g7Rmp9o�q�f.@��L�k�ǘ����m�]+Kl$v����
�y�粿A��	Z2��" 8���/����Z��˦$�3H'��S��A����p����3�o���߯("��/��`��q$������|����۸&����?�}.e/�����X� ��|�G<?5Ʃ0n��d����7�vf����:"Iʟ�X9�'ѐ��5��%tXlxVHYEB     400     1c0�d^#�쮣W�
U�o����ϩ�XZ���Sn�f�%�5u��ᇦ��+�L�����e������R��ѩE� "� ����WY��-�u�3OW��� �ߢ֖J��o�����=BQol������K˞wn�'6�"�Cod �Y���C[�
������S�.�<�$�G>��r.��m(�#v��?����Bn��k �(�i(P���POB4��q��Z�"bL���"tu3�X��w�l@�y��$ݷ�3�H9����o�B�O߄3�b4�����ɱ�	t|5�,��[΍���p�__@�}���\��r�'��5�=�)�0�����6�ܔl���VG7E��&�x���!��@���0�\�$�h=k<�)�q�>dvӚ?�iu�3x�z٦�g��k�7����a�_�-���5��u�k��XlxVHYEB     400     180zd�E�������A�����N#��E�8��T	,Bu��o�UW6$��4���  `�_��D~'#O�o�+�m(�t(�w�Wv%�z���kA4{|�iM�Vh���o#����V�z�=����p�U�G�ud�|(�;uE#7������葚���3�<�w�$�S��s�-!d�W�,(y�;"�4�*�Ka�����BsŴ���� ԧ����B�_Y۔l�A:�ِ�o���>�Gr�	[`�q.ZD3���
��j������_,m�
��a��+���<���d��ȁa ��@beY���q�s;�Ūw� �u�F��P���dV���8���
�����y5o*�"��'B�~�v/����H����o��\�XlxVHYEB     400     1504�;���s��{���8\���|o���(Tr���<�NR:��z4E�b����G�	��	U�"�W���ol�,�Tg���I�I%I5�	Kqm�	d��c��WzX`�wa�c5c�wB|�H�=7�}(1129Ɖ'��ʆ�;�a����<��l��_�#W�S#D�+e{*�:7;xʍ�O��E���'�~�71F��e����_������t�F�����}۾<��Y�.2;+^�-`�Q�|� N5&.����Ќ[KuSG�Ћ�9�&�n|���;�L�ȕ����~��?�CL:�ēRN
�� 3��7�ͥF�I��Y'�f��
�Yrˣ"��i_��)�XlxVHYEB     400     1b0~��c]0]r�s�~ǉ2�G���e��e���w�+,�K^D��kR�n|!@��)_�&G4]�含T���a�J[��]��x�˯'="l��%�(kFM�)���?NKQ�v�07�JOǑ1�Կ�_B5b�n-����j{F��ٝ��-(>�`��⡙�?�ڐ1��V��HX��K4��f�ZƣF���p.?R��C�n8u!u"8A�����/�z>,�\�����"�"��N�ՍF�!u�i/af���2��x���a׿�M����,�(�F�FfK#�#1~[�����I�E;�3��1ʏb�������R�<�l�q>�:R߷gU�1br@В�c���9Q�3����X��� _�M����
��4s�U(�uXG<�bC�;����\_�J�q <y��:�&�2;Aqo�~�XlxVHYEB     400     100�=��<f�ѡ���/"�!d��E�R��U�T�Bi���b��u�ݜb	�=�Y�־tq}[K�>�Q��S<A��j�%ej����ҒBZ$ |u�9k��n3X�ep����V��0�����W����	�q��&x�6(	��l�[��4��X[W������DL|��髼?`4������j�\��[U���	���� �E��.&�� ��8�U�k���)mxë�J�&諼]s��h;��l�dL�@��?�h� �XlxVHYEB     400     120e�F�0W�C�$�/�m��*�?X�Ů��'!�V3�ul��w����T�������)�JPP��O5	�{��4��M������6�%ۃM�fZ�YƹQ�1!ʮ5Cj4۟2�ֆԄB�(D|��YPn�YR˱�R(�r!�>\�ԝS &����wq�_���^E/f�HV-�9k�k��3H��Y�(�S��a�y^M� CI��ݫV�D��;}�=id`��j�4�E���Wv�����wf0;�S�y*A�����C�6r�55�%I�Kf��똠�ncn,XlxVHYEB     400     160��)�����I=�$��������a�s�w3���H��s M��ގ�`���t���G�����NIU�_v����-/��=�E|��0�'�kv��Z)W�ɒ`�",3�RiX��(��x��\o7K���쫢Ɋb��E(��Ǜx�O���釟W���	�p�����w-�_SI细z6�L��1�j�pI�r����G��A:5���QlԆy�5^B�i
�����s�¶W_�8C�-_"d����t�Wyۍ ^�Л��3��'o��g��&�s�(]H�0�T]d9ke�?,��rl����힁8�5�2�ұf(�1]�&D<�}���C�{[�s�W�>��z���XlxVHYEB     400     110�3b�c}�k�=�`�,�27��pd��9�������q���qˊ37��0����!�����q���*N�ܠqB��q'O��2����Hi�s_�!Cv���/�5J��-��y��E��D���]#�+��r�#���x�v���Ψ��HzbT����o��3B��/"mPH�w���X��<� ��-��H��`?|�ۈá�[_P�+è��ˉ�er�ڭ/�:{�n1�����=4�k��0y4!�l��&�a�����F�[;U�?XlxVHYEB     400     100�SP-���א����ܼ�B[�Y�?=���X3��o|n?«C(�Ǽm.��V���2�a0�9�>gY�={<�@���iq�(
�[��uwBs�j�'?e���<�r�U%��K�T�/�2�,��V������6$����.��'d1�2M����������&o�#s~ܺyoۗ����(�qg7���])Hu��гB��
`?�b ����,��Lք�ɾjs̅��m.m�]�M�ެ���JV��[cdaZ�QS=�.XlxVHYEB     400      d0�dxZ���������w���C��>`�2�P���J'������\���_0^B���H=�T�R���W�6O������!���jg��|2-~�
�3���q+g0.\�ı��H��7�-PS���E�S���y��,��i�7���%�aVA7`X-�w�Lӧ���
� ��6�d��M:���U_=��e�b��ԴyXlxVHYEB     400      d0�=��$�OF�(�h� ������ ѕo*U}�E�O��NQ��E�}m������E��L�\�si��v9��I�_��=��j���&��^Z}�U%�C�(�aLĞ(�8LQ�K���<F$E�͜B'&m~��D�C$�3�iL^���_�5�`Q�k`�hGc��]��}d��E���<�ª����v���`���&j��V��XlxVHYEB     400     130f��C��c���i����)�,@�V���@��,*���dG\�k.[��׈��R\*T�܍���EFI����U��t��{�'�,�}2M=�7������6�zm,�j%Q4h5j��Z�Ю�ΕI�8�xXo�ﭪ��sO��՛��|v4;�����E��#�	 w�X�̹r���O��C
�ȷ����[`�ޘ�U��ѷ ��Y9:�v�ɖ��Xߒ���G�l=؅�k���!��ؽ-�
�f��$�pS����i�Y�˝�LZۚBPU��<�����oQhť�C����}�����XlxVHYEB     400     150��UY�|����ѧq>�0�[c)Q�;��2�)��Th�J&�T��]�.�L��]�y��Mk��mBI1�
N�gA���h�jOm*�
� �կV���B����$!��m3937�F���q�9{���cr|w2P�,��Vq�G���(�(��i���������d?��^�-E�g��QI?@֌)�ru��(�&�����G��:�d��{(hX�#���3�E�9,��Z	%���o��أ�=�yP-Ν窓�nA�dl]���>��]�J��b�$��m��̄34ғ+�E�Tr�]�zw�x�Պ��أ��QVh]�XlxVHYEB     400     170�C<Y���a�JY���rZ/�U���0< ��nS�#�M��<;�-��������K�P��zL2�5��4�fr`�ͺ���qZ�P�E=-7��3�Z�Y��0^pݨaM!�}^j���+�q���c�oM��O�"�Xٯ��2����]���^V��ֆ7�K�ܬNޜ��؜�Ȣ�O��!4�Ʉg�@3����+m��a�B9U��(�o��P�{o�KJ� �l�a�ԓe�-��|��KB�s�?��nO��X!n�03�B0�T�-:%j_&7-`�M)M��jM�U��H0'�#��08�F9���*�S9����W'46g�ӄ��S�bu�������/�K����a��E�XlxVHYEB     400     190�\�_3���h���"�&����.sOfzTjT��E�f�
0M�{����7�G-X@b��k�Q�M2��M{ �u���G�n�,������7m��� �uQ/%�@|#��U!_�]�� 3��K��4�����'ʰ��;��:m� ���z�Q��ٲ���n��Q�rz�e�p��g�|Y7\���ʽҲ��s�����Nq���f���`��z#r(-�u�jK��F 󵊩^�l?|ц��Ko֭�<�� �b��a�8�>�b�I���b��L3�'��a㇨�h�8p����E0�Ƿ29����P�C��ۭ�-�qm���ؙn����U�%�ꔘ���3_���ُK��j�Y����R�Tn�=�+��VȏK$͚�q��R��E������_�v&D�NXlxVHYEB     400     180�?�����r�OX����Z�Z \Y�v�w��S_���~p��Sc	����NNu=Z�"��W4��4p���#s��k_������ڰ�������&��Ӿ��V� ʹ�ؚs�4�f<�� Ec]U�t�̏	h�j#���{\)�2Z� R5�����A)�GW�Z�Z��]��I��i:�J�zк8cW��v&�"�s%�,�=��3��t�ſ5������4����Zz�͸���sY�=ѡ�mT,��i2͛l��������f��x��#�Q�)����������Qw���Its�=`��[V�n30�UKϸ�c�R�XVЩf{g����:�b�
[�+4d����e�_.�I� �kX�?���[��t
XlxVHYEB     400     140ن�'M��:>�+L|>���������w�/nY::f��^�ݍ=k�G�[Y�8�ǃ�@��O}z]YG�Υ�+V��H�@�����*�
�R�yM=x��!��tn�l@4��"!DW����F��/]�Rnaۖ�~�*D� R�Mxx��>tlN�"�vDg|��s��P��XW��0��]۲��-%�Dz��(�!�6ȩ�+X:��l{.��2z�ؽ���U��Ā�#�;����h}��}�}�Q/��\^�z6�^�'�d.d���pP��41��s���PSt����ڊ'1�I�r�S�,Y�lmrs	d��vU�n�XlxVHYEB     400     130�Ra$�{�*_1�s(rC�A��`�J<E�\>���T��^n&���=�f�&�݋��E���9s�?Y^�3�U��p�|6�KF77kпF�G���v��U�"����{bâ�ag+W�\��^@��a6!�Ȃ�ׄ����vC���?��2�|sJ�&�U�Ơ�te��&��!�L7��d1�T�����"�cdj���&��j"@B���OeU}���Vҽ4$Ǳg�i�`�Sc��'����z��	#��Jk{��� �6Rװ?�Z��!\T<�ʚ�����b ab�@��(�`	��~	��XlxVHYEB     400     170�ė�X��)e�+�,
�~�r�9��3)�j�h��?��Ǖ�v�3����tO�Qn�6{gW[y�N#��G6tÀEK���UC-_���g}�s��ka�2l�����/R�����1��:��G��B���q秫����Tlz>�#��u��󸾀��sH=�8����9�l3�R�9�����Y�B3����U���?y�?җp����)�=�B{r���Q�s�? �;�@���#�F�8,���,2�8Y�ua�YPz��G։I���3��:�����]�RB+�20eĲ"�k��S@����g� �\�m��ɤ� e����p�{.��V���&��W;��e�;$�2��Y�XlxVHYEB     400     1204�QÖuq��R0�㯘gۼ���xs6(/?��neH�k�z�����,��f�M �,R����Bf���=���w�.L�x��I9P�-qq8n�V4�e�E�@�@�f�QC��2����T���A$*|IWS���� ��Ugi�T�Fe3���^ �\�#�x�^�M.;QR�����%�}W�`$�O*;8z�;��+S(#�6ǉC�Gw"b�'�!%�mv����ua'�<ޅwhZ�niL(�~l�vS=q\!0��:��7s6��H�˖p�ʕ6�v��h�K)XlxVHYEB     400     130��NJ��q���S�?D��+mD>��2$��f�BQ��X�d�z�A<^&�I�8V�PF,�]b)wn���t�`�k���}wx ��g	@�>�M� a{��8l1㟉�0�Z�2�`]%��J���[��r����\���Q�F�D�b~���7�h��6-��U1�5?ɤ�I��c%�� �d�+��1Żw��}�Y#�9��`��x�]7l��,�K��2x|M�!~��w�f���#y�,�IOm�,�'�����QP�p�p�h�l;�������0/D�zc����-F�+�z�6XlxVHYEB     400     140���+`��ڶ�cj/����D����p:~+3�����͠׌@է$�Y�Y�Gp2S#pQ��o&��ԣF���� ^P�}Y�C�{ɷ��Ѷ�Z�p.�LeÂՀ��$��w�O���֜���ti-Y�yA"���BDp���P�&Z��1�fg��.ڰ�x�6r !&P�����z��0�3��h���!�:Ma.��6��|6c��]u�=|u�#Ϻ���(��W��/e�G9XĹRW�:�k��D�e/l��������*�諰pn�E��S��uǼ7�T0�ǖ�Ҷ�Hg�B���|!�I:���ݐ7	OXk�酾XlxVHYEB     400     1a0�/�n�"2�*7�"���^�5Fe�<o����w������׎%'��yj��l��Zs嘅G�J���#p$)ٓ���?J��yD.�P6?MgXT��*�\�/��M|w�꠹Yj�'�&��2���a�}W��h���)(H��8Nޘ�r(�:�����H#�o��pZ+� @�@ =&AK3���*���e�����s4 �>��C��S��Ëo�7K����$�.��5+��@'ѣ�EZ�-��O��pd�1�4�1�]s%|@�����ō Q����m��*DOxm�?����M֘��YF.|��K@竮�qo'��fN@�	�/��XJ@JR| ��_��2������9��Gt��|�|LS��z��͈��j��+L&��b$���a��,<gl/e����XlxVHYEB     400     180|�8s�Ē�\>P�]���	{Q;�|��8��������TF����zN]�z�Zt�V���pX_�o�z�Jk��u6/�~���W.�A�C��ֵ��ka����m j��c2w(�׌.�gj1���qo��w��i��U�Y+,G6��Y���3N������%ede�����۶A9	P�C���n*�l�˟����7���{���q�8ϸS��8N ��H̢A�8�2�5�GE��<��C"+�u��K[�ǘ`" �m�(�l�|�B��6�ý@4��zP���zg)��1����}�H\��$Q��S��:�+$2a�\By5���"����!����;�Ź^c����z�৙VE��]��m���i�KO�XlxVHYEB     400     170�0�$���H�}&+�g�6����Wo¾��x���*�߁3z��j���alѣ�2`�z+��P�N0�5�,X��d��0�M������4Ui����*�=1�3{6�g<~"�t���6[�>8+Oo�B�RW�;�ןP�qpNE-�钭��(�Gܠ�uBP`ύ�-�r��-Z�y7�#���3W�2�g�Lg�u���tp���*�tPȤ�J��"6]�1hr��ْ���{�sWd���S�k@椥�g��!�e�2��\�4߾��b,%�՟߬ܣ���n���Ш�Drc�5�uAb��afaپ:V���l��Ғ���۫5�:�؈��\�:���{5a&��9IV���BXlxVHYEB     400     1e0+�w5.\J�!�_�hǘe�g��[����i��2�������}�,�5�����#�聟���7W+�y7��#��g!I>�7 y9{�Y�?��'^���o᪶!�S/l��L?�)�=Y��������2�(���#�l�x�`X̎J3�5�yэ%{��kf���FAb��Ia�O[��������\Iz��I�����'�s���e}y��$� �scYQ�[�sp�?F�X���s;���(J�+�f&Feb�Tw��jGX�_y��Ub0wI��ʊ���zF�8����0HL9�|��s�V2����� ���Ӣ�s����tD��~)fVH�c��¸�y�e,��Ty�b|�S?�+=�N���{^�,���et���b/��$�U[����pf�i��Ǿ�u{^ݼ{�=�D����r�@��?�-i�y�����+0�#P���<�D� ��$��=��<����%�ƌ��i�w#��*$XlxVHYEB     400     1b0�Ճ�����0w����H>�ݗ���V�.�|]&i1��b��@��c`ta_N�a��Ί\��DCa��z�l7�L���P�:��W��:�I�҄-f���9��Ph���������c#�o妱9jr��U�u<��ש"�PW��^;~�q,����ݠj�d������{Y�wV�6�z?
G2� �mZ'��(��|�4JL�v��~͓�v�T����L�g��|����墝3��l�{m��&Oy�X���~�'P����`: ���r��?�xh��r��z���ɠW��|���%鐥�S�d9�-Y��J�1/v�d�3J��}lCYZ�\�
�'[R?��@�#Ӟ����U���:�_C0�Ѻg}"�21j3���B$�'���5y�"���u��l�)$u�:����!�XlxVHYEB     400     160�z�X~�ӎMT�ԍ�nh�]���Z+�m$�R�L��7�Wz� ���>����Q�: �O��p�*`֕����gs�݄��K����R�D�_^����9��������U�ƞ���Ƈ�H��{e�oB���dY'�1���J���=ǉ.�J��sa$��	��@�+���M~T��}�ۅV��J�Hvw�	 ~�ʾK��g>F�%Z)e�:�pޝ�y$1#DT��ѹ$Z��B��ϋ̐���!���4[��hA�k*�'��y��* ���L�S*�)Όme�/	�yL�� [�ѫ�WD����2]�a��L��m���JM�eWg�[�eX�G���2�0y�&`XlxVHYEB     400     150M�8��5gˈ)�����gJ�y=r�Z|i]�r�<�D��߶�� �����Ő�\��k�%bҦwM��n�^�̕��C{�E���"nו���Xm}���q£g`�n3�%M̬e�=�Hr*�P����|L�W,V��%!8���@t��I=^���M���<-#��1�*y��)�f3[��P����y��y��)K�2�ht+�#/��MFJ}aw�m����"w��B������)��L?Շqno(k��)�y1l�q�<���]5y�8Y�Lє9�F2�QAs9�J#h��)O���������՝��w�����Ӑh1��Qúc�\�/c��XlxVHYEB     400     1a0�ݺMq�/���0�-3���N�Y�Na��L�ܘ��4����00F�M����b��˰�Wk{>�X�!&)f�+�6���
iC$���8�_�9j�k���|^�fc�ô�s�wFzy����"�1X��u����MӮܑl9��²����x�|G�f���r��ej&az·\��<����hP�`��7$����1V5r��x!�.8�w���x��Sr��kެ:_L��Ɖ��	�=�_��� :���Q?�6��]qտR ���=t���%P0S1��~����	'����S�2v�g�fK�zZ�98%QQ���7�{�q�L=|Xt83�ǹ��0�C�ǜk�Fq�ꯟ`C���r���*r�_�m����?��J�qP��r��Ru���R6�%CV�E�/�XlxVHYEB     400     150�:DP��ll�|���������)Z>tp���3ۙ�]��f%;�k��:d�@����Cm6�l����V��,p���3fX��M��v����A���&��:����oD��Y ��w`L�M�>*=�� �[�T��쾟S����TQk��m&�+^7�h2M˥�#��
��D�)�ZQk��.uEѲC�	X8��P5��(�o�\�ƻ���s[��
��`DKE�𓮋�6�\B��TR$���C�P��7�b����1'u�4/h6:��P�����~"-s;w��(A��c(ͼ�i0��hѮ���5��^x�N�XlxVHYEB     400      e0aZ��^���|�u[�`�������ɉ�4k�=۸B��>$���̋<�))[�A��&ɦ�˒����>�ZAL4�߷����̝��{��ĭQ<&�߃q�� ݙZ��q��!��5�2����[b�8�Q[��G�SZi�e�J&�ÕJ
������<s_�l�q��R\�~E��T6J��3��c]l��S$��K���b���V�:�
[Mc:/͌I�F6��D��#�XlxVHYEB     400      e0`߸���(%y�7ډp?��l1�'m�Sx�q�%��R�w,k���!��f�prz��Т,�n0�R�mn{%Uv����MD�/�؆Txb2���d��ޮ�}�^B�����%�4����g������$��0�\��k�Pܛ؝���*-�.>��$ ��(�(*HF��_G;y�:�I#H�4�-`7�f�,�Ò'�{�2����5�_wu4���K���?�XlxVHYEB     400      f0����Oч,�,�^���
���~����	y��*+�/�w�m�$|A-�ю�n�nG��ɋ�7�S�@�M5�^�u�d�rt�;�5�S�q�	I��������st����[��fcՁu-H�9x�m2Ė~�� ��:��`@
�X�[�}� L~	[���v��+��F���B �LP�Ԏ�ل�ײyAhH�s�2x�2����81Iy@\v�
���{(��V�c`̩Dzu�`XlxVHYEB     400      f0�ɞ[�CN�̶IҭpFx3�C��$m�b���s�!��k�N�q��Fb��a�@m�aO��-'~��}�����)���eR�В���Bc2�E�D�bn����h!��hJ�A��^�i�y'N������^]��Fox W0�k�s�����EBVm>�MC�B) ��^��]����L�����W!�jle_�
�鵷�Lɿ~��g�6�T�Vx�ucW�7�!�����ż��5vs��"�XlxVHYEB     400     110C2��>�<3�!m�����%��!a
�k�xی���S~ª�k�</X�v%�bј����l�PG�+:�M�̼L�J����7h�*�灂�fEt2�Q�P��ң:�b����`����GĖ��VY�T����@(�0-���Qr�]\����3�l!�⥆������b*-輞�?2KG��()*��W�?�	�?)�|�Kq��1�����r0S]�*`#��Bњ��o��߿�C�l��fn}�3y\Jj�
[�!{��Ao�Y�S��XlxVHYEB     400     1b0�XQ�I�]�k��d�
O�E�S�!h�	��i"*�״1��/s�Gey�`�O�A�Ynm����c~]�R�S������"ue1M�ќ~���k�f�u�Ϥ# /C���̯��צ�1�F�p���	���a�6U������a�}#dh�s��
��R
�U���𺒆(�bN���ʄ���n�"4�h%��U	��a��6hbz�/< �T+�@����6SOJĞw��>���4@��n�0���
���|RA��\9�K�b2�㪣��I���vE%��'�A`��n���"����|Ñ`�eO��_x���0��#�;�c�L������I
�����[s�~O(FޭP!��{�C���8�N(�L}t��hXk��u� "�T�����iL�v{���j����=4��I��5حH��c����2XlxVHYEB     400     140_��%�˧��%�ٝZa����5�	fԌ�S��^Eo��b�w�M���>ȿ%>2x�]�7j��Ph�P �{�[܃��l�����]IX$�Bq�w� i�+�H��@,��)��=us��$���Qǝ6/�|j}�	��E�.�#o��>��������`_�Nb	L	ʔZn6��a"���uۑ���rjU���S=si�8�����N�W��`4��r����K����_���m�~�����ۇS�NW��َ�ɔ+Z����@�<Gl�;�Y���m����h��n@<�xd9rw/�qc�x����/S{�,U�d���!�XlxVHYEB     400     160t��}g0S��t�3�.�8��o�VӿlSt�"9�[0��	��nd�H�`�v��˿Hb��wnU�$�1|Jp$�o�e��ú����XkХ5�Ӟy�k�`G��y�Rַ=4h8�u96$;�������!�Z%»��B^�eMv0��~j��<�c�q�HJ4@WP��˷2i�-e�U��'�"���*MFe�U��W6̂�VO�t��H���7E���x��ɺ�
��/�qu������ڗb�0ZS�ｩ����
(L��6���qԵQ?ŝ�
����eMs_��6�B���L��������Hߓi	�}8�����|�ִ����.��R6���g��f�*n�l'�XlxVHYEB     400     140�.�r�U�[�=���
NBF���{de�U�
�D},�č{�x߷jN^ \du��{�������ͩ��P�:on~y1ԩ��7��z�g��A�?ُAa�$�G�ܘ��`ps'�=kE��nd����	P��"�#��m^��;b8[�h�X��hw\���&��ȣ"})UE�	�"6�k���.�7ɘ�t<������:�R��5:#q<�'�p��w*C�N_p���HZ���s����/}6�g]A�o�峩(#i�݅;(�=Q�yB�	̊��4�gZ����r�8VZ��I�dH4?�X�����z�ոZXlxVHYEB     400     180L�O,�%"|�tIv��|M��3�/��>�n�7UZ���K)�����B�,���5�Gs������rRq��G�k�I"����������0����^hS��սQ��<�@k��������Ӣ^�ٽ)�-ٻ ���~�mEq�bU�k���4m ��3Ci��5�X6 �m>����﷚4?���.]�Y�[��S�ZJV�
,Ŝ��ѐ��w���H��C �C�(��5��x�c��ڹ�,��a8WV �:W�x��5ܭ݉5]�*_Hc�3قu ���&ĝj�^���������g!L�][L�j�⣄H@wr�(�,�P�PT�� @>�O�|�Z��T�X�����o��s+7(��'ϲ$u��-���uXlxVHYEB     400     190�X�A�+���	Ιǰ�oR���۟7�?�ݳ��з��J�av`a�aZU��5AQJ������@�o��CkY��I�e�8�
��r�������ɛ$�����Q@4q�+�;�G;�>0m������]�>q��7"�~�@{��x��Ѣ}�)��\��qO�ZUm̐؅�KɅ����C�R�`��ԍ�Q�j�E�~�Xȭ��9j&༿�L9!����XUN����z�-{��q`e��n~`���V$�W�%�d�~ ���S�s/�@����/oZL�d�G�d���,���p��~�C
���.ܞ��==�~)�P3��xü�b=,ӷc������w���gSm�-{6{��_oc����:M�k��o�`i$�؅^%NXlxVHYEB     400     150�R�lU_��@ޑ��O��Sn�׽B�����
�i{v��t�e|�����-�4�c3���P�S�J��Zт�y��ʗi���U�w�1�R�}���Zkr�l���y��\2[w|m.�3N2k��k*�_��SړnG7���h{�f����)��R��6s,u�e:ɳb �J�A	6�M��V?��=2�?Q��L�BU��ïQ/�m�(���G�O���6��8!{%����?v,J�c��Rx�HV&���9�|�E6�,�>�͵x�s�g� �F�b�3y��oF_�_�O�����hiX� �5��,|#X{�1ސm��W4>U�X���.p��XlxVHYEB     400     1a0/!���ǵ�	��I��^0R*�4�������d(s�
���al�rx��]]Խ���|�J"�T��ז8��h�'��uO��Y�K���?iJ���������kx5��!+KL�Ǟ�B�`{K1'̙�M��O�S>�񽍗�C��W'OC��۔o�n����D$��c���ҁ� �~E�<0��UI����jN�g6;R�2ƫ�x��YS��Q�#
�3�֒����RH��6�B��q=
�*U�e؅L�X�T��+mk�G8A���p�2����&��Γlۃrq��wKr<R�$߸nϦ�c�B4�Qa�ʼ A��������7��B�΂1��g,el�lh9c���S���(b�<�!6��>mWΪ���)��C�[�J���QnXb���H�a/^��}�-1�����1XlxVHYEB     400      f0NR�ʡ���"��>��i�ᴚ���BDQ� @a�=$Otg̀��j�`�8\���̊[����%�sѢ��̱��W?2����M\k�	�Bu˘��U��G-O�,q��ѫ^���\�"�e�p*S��~i���,��a�V�ZJ��8	0����w"��F�L@���=�#��`�| Dc{H���"8N��,�;��-���'����u�1�� G����(��$�iv�Z/	ֱ�XlxVHYEB     400     100��mTs*:O���c�Uu�pYn.A�iߑ:�'D�o�.��H]M��*�]ߕ��������z
*fAF}7n�Q^/��֚� qSwYDZ�E\�������x�d*�cYߧ��/�`�����M�F:��w+�		L�_�D����k�'v�.�v1ӊ+5�9�cLRB��_!:^'w�nW�4����1t����>k��T'�qb\�l�1�8Z�7 �lOa!�$��&�I�++c �����@d����ED�VA�SXlxVHYEB     400      f0�O]�3]�0/7�LB^����B�����^�M�հ1�s����H��ȫt���-�
��ig�o/�)d�t�<MZ�O��UM�y��ǆ�G`��}�t��&�A��5�;q��}���6jܘlLq+qÔ*n���7��z��Yl�}n�5�)P�Bf$�{�Ⱥ}>pDp��`.v�n�q��P��������j��>S��	|Y�)��<8�'>{Ԑ�
���w���;�ws�F���E�� `�)XlxVHYEB     400     120O�f/�[t���"��񶿓C��	��}ܠWk`�5o����v�7��X��9�7�Ajm��4VS;)�Yق��c��1�U�9׆�s����zs������A�
�{�I��M�4�7k_�a�[�C	xg�Sj��c��6o����wQ0���+P-ҏ��������gZ�^�2�t�~�X���gA~�j}R�hg��p���HC�I<��D$�'C�X�J�z����'�]�y^�	eׄ�ђ�yd�e!P���ݴ��8,7��Z�r6R�W�QL87�Z֭XlxVHYEB     400      c0�����x"6��Z�agG�7�S=4��SЃ9�f~��'�S,r _SE��VD	p<�o������x��4}���]h�-f�j�����>cM��U�g���O��������3��FV'|���Z���FWYZ7�|?԰g���P:;)p}��Q꓾�r��v�����e[P����gc�������=AGXlxVHYEB     400     150��f���3T���w��s��[���Wr�A��x�噑rQ~yV�>�.	ធy�h_����l�dJz�Vy�ٚ��U�Һ/�CDJvr˧Q�o��ը�h�J	 g��D����H��T���Ay�����x&r�~�w��iPй�Wsjˤ�oU�w�3`ז~jQ��e$)���m����Ba�'T�z��,a?T��L�۹�5w�;�2�feQ*���ts�!<Hbڲ�&N-_%�M��Gb��8��o�׈�P7��B=�����ײ"8iB�2/4� �bw�ߒ|�����$Ķbq��:tÆ=h<��Sؿ5u�qښ4�5 �+ό>7�˝�XlxVHYEB     400     130�m���Wm ��ْ���`NC���%�˞F�T������vM�ס� �s}2�Y�Ѳ(j�H^����Q(��=����:(���
rinӕ[�P~@�}6��X����!(81&�:��)jAQH&ώ<����{�k�x��~���3	
o�vQH�`։R=��#��\��tם\ {��_}�ph������*`% ���6�u!Õ�z_©h<�.[�0�SK��R��G�Lu�4�^��6�k8�"Ҷ�g6�õf��̱d�\2upl8�Σl8�=��<�	#��`�*��8�XlxVHYEB     353     160��ĥ?��b%vr�-�,�1!��/�֌!i�_�8V5֛�߂*R9�}D�^����;�uh�4�3CLt�����>'��ڪ)�ȯC�T�
K~G�˅�ք.jsV�'�X�'��P%c#�e'�ĭZ}d%Z�b+���!�O1c0K����Ԏv��]�g�&ѱ}T�Gz��~���h8l�#����/P�~��N��1H)d�<剚K�id�e��4G��9�~��TM��K�,-���q���T�q&w����+(M�"�p)�5Tb�zo5��¶��b�	��f��/V����n�ա���$���W�����la��2Q�OAG��+��X��p���