��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��К�U����%5���&�X�ȩ�u�MhBc+1��;��Usj�9�s>�i��-���p|�w*����@�ٌ�n��Q5��2��i,�S^���bW�X*A��$b>*�����Y�ً幱�-�
G����&�w�٠q��n(`�;�6z�J �T#�s�r>Q*Wv�]L.U9�G�*Cr�} 8�^u/����f�����Aa�}��b1�f\�������n҄��ىQE�<yCZI�?;y�}�V�'`�&Z��踃��
�9)���X	u���sD*�#FЪ4�T� l��n�l=AC���^e��,���p�,:*�8*��"k�DLf.[��}�>@��k ��Sa��UUr4?��%D�aї����šB�=k��a��������y��IM�A-Yڶ[�q����ު�����pR眢 n����A��Ӂ��	2�!8-�TrܳJG, "��d�;�� t�@��e��&�r�p=��.`��:�U\Uk��H���.CP�'��3S���u��R(ʡaG�CX�=雰/�� ��^a�ka��w�n�4������SJ���Xzܻ4�����l�a]!��Sї�.�P��L�\B���z`Ǡ�y;�����1�^���=V��eh���d�h�/W����*���[�p��Q8?,u�[�x>��L�[�`X�2;��?�ߙ F�m DRO�8)F0&���]������ s��h��)h䨻+�!�c���'ڥ|���P ƪ��h���
�om�M��ճ�f��/l���^ˍD�D��BU]O��ϩO�bo�BF.������F._ZS�HG��B+�@e�A��D�:�޵Ƨ]/b`�FN\�gr(���q0��F1�t&��VTL�l�G�����6�%�~}	Sa�HT~�Oy�3=NY��a�0d�9������V������-��3[��#��k⛈�V�o6~J?f=�-`�|�Ie��������qX�)��"������At�e��S���jZ��ȉ^���J�p1Č�)Ƥw�,K7/^�m��h� {=�[z�S�ҭ�d�F6"vǙ��p����Ɋ�8Z�;�V����Ce!�GI2�fw��p��u��e>-�I��O���)NJ�|��*��7�[�*�C�p�e�#+�x����>�'���ki�&#>�2��x���4H��$�p��^���_]`;n��UMnCp�Z�kԬ�٘�ۄ=.3����1ܩZ�c��;�8x�� e�h39]���� ���4��QW-߼�_��w��g~������� �|L&:@n�h�Ox5M���mǯ��aV;�������W� ]�W�%��`�V��ݯy&v1��F"�
��C��>f]�y&�c�C��[@hޖ���E����5H��3͈�+��JIez�������e+�����Y�����b�����G�]�6���b��C�IY��z��X�ֽ�a��E�&����呢.�G�9G�K36��,��Du<�ӎ�s�6�_fVq���Fðֳi[�y�ɑ�KD7|��Ti�`Y��7�as�L��+A���b��N����*mh�
*n�W��2hz����T�7�*�^���l%1G-�T������^3 �+W�.�o�sDV�% v��x|3
ۑ���,���N���k	�j�E���G�)cM[�> �)�$$�Eh<�mV=�eAW:
���LsR4U�rc�s�����Xa��n{=�̮zIs��FW���ٲ��"mF�H��$k���ojИ�i}#9�&Ҿq���>x0�aJ� oʐ��tߑ䁄�E�OR������� *�'m�υ�UX�{E��Ke�(�G���C[(}��*�i ��Z��-�ȗN5�/�h���1�����:��OI�Sm�@�������Ů$9���7�5`�u�G��3j����c(q�zu_OR>����}��	� �ﾹD��TN�1*�������"'Gno���|��ED I�5��	y^ŸKN��z���C�<�۴`p&��)6�V;'�D܎�� _�,5KA,��7iʎU۹��i�k�����J�p%f܁8UMM��o�6�X�A�4�{�9k�z�^�X����d�5�O�v��Ee��]$��с��2�I�Ie����I%��|).M}�ɡ�C��Ѿ\����ޡ��*A��+gۖ�T�Z4C�����c���� CW.������AW��,���Z�Fi�},�Z5��R�0���L �"�XǢ�������	���R��D��R�i�����G`rg~��+G�� |�[do�V��_Mj�:h�5vEfix8�*�PO���V���/�t���3����Q?,����$"[B#����3�2�S�҄ǈ�R���ᢅ����{n�� ��3�T�k;����n�"DF7��:����M����:���
7� ����P
z�;�xQ=`G@�Ld�;���Oqe��*����j狂5=�Zw�L�`, D����WcH�3O�Nm�S�$��X=X�5�>����w���?ŊŀA'Ğ�zzb�r�<� ���_�Q�ě��XH�??��ha��8m��)�������W_1�$�w�A8�}؆��}�G��;:�~U����J>�P�5�.E<xi@f�E���\]
����D0��E,S0Ǯ[9�eo� ���Wd�ܯ�<���/�� ^��p�:�o*C�E��*�ꦅ��ZbF��J���HB�J]%���T�/�C΄�"˞u	���M����.-\�>_����rD#�a�L�Ќ���g�D�Á�&��p��7���6�0�����DK�u���3�x�Ef-w���@fԠ��F:���f��[�p�g��BLKl����/��1ZK�q�'�ES�v��B��UA����Y�������b	�^���V�.q	e��c_#?ԉ��3�KEJ2���]��m+qc�JۙS�q�셦�1�路͔7\G�lv��I\��y{鉠�W��_��l\0�F�� ���h������w�N����Z�|ה>��Y�;��NL�h�G�i�#�.&'���1��!�	l�b�#�Tf����dŎ�GM7�U�)�7<�?���}�Pf�%���v~t��bj:j��U��c��=l��������6<����!�b��8f�)5�L�R�	�T�W ��;I:/�L-T�z�ݧ36�B�__d��Zs���B�_���)���#tF���a�K�D��S�ਦ�Ÿ́���y�9˭;�j�d�!�1��ܹS4�|��͗V� ��%*p���'���lGza{k�ѰB��0���:<�{�p���$5+�x`���Z2�e [V�����ɲq$��34��C����S�8n°�c2����e�(\�S�I;�_A�2ÐĿ0��_?����N����o���w�I�c���n�)��d��m��]9�XC#b�3,�UH,n�n��� !܂�L;���� ,�8�������B�;��O�f��!��͝��%L{�۟��#h�F�����~L&yB�t����<���N6�	��EH= a��LL8�n6��	�g�5��H1d
*c�{΍�;�AO�2���ȅ�b�m`���*у��4�kxB��������ʐ��g7���IA����(��� ��{��v���V�w�*i���,\�/��"S�/߳d���g�7��YRt/`���i��]*`��l��V�|�]+6rG&���Ҥ����b�,} 5p9	�L���I�V�c� ���m1G�Aj;��Z��P����$ǈW9n��9�����c�e46�a�4�wl-O!�^����6%�Wg�4����M	g5�s��{���1����%�2&׎���t6������k�ӡ���2�?��@�~@��N�{g��@N��hn��8�@ӟg�]S��_-�J��9K��������i�o����e�*�2��r����F��O��/�-�E�.�O;�]��
��~$�dz<��ܳ	YYT�����$FrlV�m�a!�r.|E�����l�"p�����
��%J�m?�^��E
���&��V��	A{����ɳm-����ϲj��z�tя��i֥43Iu9��ܳ���O�6�2��-����o���o�X�m��x��<�_�P�����2����+������ѳ�K�͜��\9O�^��&X����6��׬"���#�@l4w�&_� `ت����f�ķQ�5V=���)ݏ���V��%%���zev�C�w�\��3NZ>����E�^A�p{�P�<��e�g�^F
 Ϳ��� 	�D���
+O@�"�6�
A�*����iw?���\��Tq�.��Ice^�g��x�3u�E'�����zK��v4�pvc^G@aVyj{�O$o� �/��_�>��Lb�J)>��.�%/��ȭQn!�x�&�%�E���U�y��H�l� ����P?"�(_dz�{��Q�$N�t-?��ڡ�r��w`-��@�\WW�Uh�3�t5�G]��e��&�
$��hZ.�W�N�+��Y�p��5�h��W�bEZ@���/y���@�=u3��o�i,c.Ѵ�#��3ĺ2w,���l�����#/`$K�P�`~����`���~5@[h&��Z�Vs�郉%���8�?}d6a#�k�_ݧ����i�4p��L�aG��D9)v���M�S�(�0��	����gT��:�v:[%��]ZI2�ͫ�L+��`����MC�U���]'���(?��grgq����1�g�5�վxv���ٻĚ~��$��M�$�>^�����]�������PD��{`4�����}}�� ��]�q2��_9���yۜ�q���cMH�-��u�K�>q��Y��q��ت��Q�뽦��-��A<�1ۣF��_�F3�V�����爈�?�ܶم��A���j����@fMq�	�x�k��<]�z���5vo���E��T�l[�K�����:�f�W��7��H�N��ʿ(�"vܼ."���8�^��M8*�i���ae磱�^v�'VAJ���6�����IF��ƍ��>DW]5�J$^�p]]�UDɝ�fܰ���3��o�s��7�i��&��p
�4�)(����*��*1)����g���9a���b��)6!�q�R�oZD�O?�lpE˅���^m�l�.�1n�ϙ���v���·,�U�X�+��TV,�-�Sф47$�IgI��0"n�4y?��b�]���Ml+*��(I)'¬��).Q�'D��NƓz��*��V���'��sՊ������8�~	���*�:X��
�5� (�&�z�����_C�S�"  b�C�v�^��j%j��kK'2��x��/�P!�y߇p���!�duq���9�g�Ps�z���"�{�`���ff��Ϋ����X&veO�в�n��[�9)�˒vHJ�+��I�[��L��[�O!��h+�h|M�V�Lx�)ܠ���kL�"��Qp�&��D��w���N~d5�<4��g8���j��B8�����o�����	�(�,���EGH��ml��s����&��L2�豂���q�b���;3�h�((n��'���`De�����cO�Dm	����;Z[0���{��:Cd!�DwN��1o-���a�X�$�_�r�%��9���7Z�=�e�}lh� [R��2�婢����@<h�}x^�2��uN���
$�QtE�J���kr�����Ca75��Oq�;ʷ�����"+
�v��^�2�7ۅH6r���"�]f����Hv��������G�m����o"����?��kQ�e��q{x� �&���-uqg�#d���h�
gKM/��,����pK��h$<^Ƒ����EJ��2|��>��7x�ul��F˘wMH]���3��hֲ�#�k�{.�Ȋ��7o#��]2�v���u�Y486f.�� �8-<��^��^|f���v. Δ���[yԢ� ��<�<\�t���Q��8��Y^,Gq �
���e0]q�J��;��۔7�h7��j�����.��e�}���6a�MsIjX$�Ʃ�������@&�����QHy�ñ�wҬ�apxFkZ4sH�d�0�5f"�9��>���}�(���}
�aua6�f�+��Fg��:7s�Q_
��W�l�{��@����{�a��q�S��E�_�.0R˦��xh�A��N���F��[�w��f:D=��gް��%آ1�S�P5k �� �'�U�&�8gF�
���g� ��y�_EB���k���ψ�C�TK �ot��5��/�Ճ���Zx�)b\�F�c�`��.k�$8��xіc�y
s3�L̍ t Z�������<�������*7��Z�xg` �\��ּ�`)�@�r+���Tw�b��r�hωhd�~�ǁNç̝Z��~��K���7�	���?Q��u�ɆL���3��:m�*3��#r0f��;������@����m�ԗ�;A��)�I<�����#��T�2z�U_�Qx<QI�N.u����f^���C�o��;]�ܩ^vL%���Lr��ć�02�s�|���횡�a�0�~2,�?���r���w��8>x.���ߘ(�^�~���uW
]j���H�H�������� 6j��#��	�����8}IY�Ml^�IG�B�}B?PTD���n ���"����Zk6`^��7��H�Tb�.��y7W% A��A`�~��@s��spw�E!���sKC��9U�P��qj$�]�H�U�^���h4��
G��|,�=]�or��[�σ�