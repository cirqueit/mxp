XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R���	�;�\#��; ��������3�)���y�3�(9Lz���u��z��-e�#r��?]Հ'c�ۆ��Sv�R(P�D��4Q*u1�8Q�zD���n�mJ�c�K�r��Q�w2�r�\�A�zˇ��{��>�?~���nJrn�6cni�<PD.A
�=�h4]��&A��t��x��k��Fxg�$�D����"��}Fl����S�u+��*g��1ْ��ꄇ�Mgҧb[�ɽe�ݡP�j����z�ɀ��P��G���q�J�]FR�,�4�z�J���>�g���ڔ�O���f�USƹ��.��d��O�f�	�w�v%��aa9�#ǩ�~�����Q�6)H�J�+ M�����S���zt@�f�t��X�,���>~!dX�
��6A/Q�}�n���D�`P��7aM�'ܖ���B�~��S��fw���Q8�Wq6(��0Ш�f}��-qd�n3�z ɂ��Y�G/��t҆9l, � eK��g����^X0	Grj�g��M{\w�/H�_��8><�:O`Ћ�Q�þ|�5����V��7l%�Zk
=��`���j%�@jj�XM���Œ��q���|R>������LZ�F��U��W;zw�|�i�%�Qah�j0��O��Ѹ)�TbGR���|ݎ��y�/!GXPt`ݵ
Mw:�Ƅ�	�Z� �g=��K)�[ �K��{\�#o�-�����f=�2o�m��ځ@��24���x���Uʦ4���g���sVӴ$)��XlxVHYEB     400     1e0�<V�Y�đ�U�~6XA8�`��~��>���9�]����=3mӀqe7�q74
*���v�'㙻ѝ� U:�R,��KCŦ��e=@]�נr�1د x��c!4w��X�S��?y�ŭ���tz]�d�_|ê��e}����dkC<�X}�膫Y"#�� $��,�ߩ�4�qW��*��d�&���"�!�
�������, �Y_��Ϥ�p�U�^������K,!E�"�n1n��������S�[-��]5���8I��T�UD�������k���O.�3��_�k#E����"�ͼ�uJ�UI�՞�k"�SK�냃��Y�������#��A�9�.����Ckӟ����\U�}��l��}d���$*,v���vR#E��*&�[e3ޞ}u�^�m��Dx.&�F~hah<����?V����{�j�$B�(��>��*�|LY���kk�(i��v6	tXlxVHYEB     400     130"���u�~.����ଙ�c�v0�̜��f�d�De���[�u��r^Q���*�Nf;�i�Ďi��;�H�����dOy�AG�bR��ڈ��0K��O���Xs�,�5.���'�Lt��{)3 k���v���V��(P�+�ys��ɦ
p�(șG��.`���8�}���Z�S�n��_���~��/K�eڱ�r[�9�2���/��~i$��n�����b(sZ�x����%;���ʛu�ҷ�{�� WA�r-�^(Jhs@-:�zN0j�;T�/�������`����ID=�\XlxVHYEB     400      e0��@ۀc�������{�➐�8�Ι=> 	BI�3�J����7�8H�dG�+��S�ե�'c_h�4|I��
��6 �_ו��0\���]�OƬ�Qٶ/"j����}��A��yj)������F}E*��ju�|�� ��69���;�B�=����x�N����ș���sڮ0C��r-��j����JV;X��:w #�d���w��Q�
�S��> XlxVHYEB     400      e0Cj09eG�+���9py�X�&9�"��E{%��->bP�egڌ���c	~�O���$�ȥhD�����f��ۑ����D=6s��0?Y�	6yMs\����Ȫ���h��|��1xvZ��I3�M������1��}j��DF�����W�:2'bm~=�����-����MUm��U,4�_*T�=�3�^��I�\�
�G�ٕ��9�>X@UZ@�nXlxVHYEB     400      e0�j�;��;4�S,:��)��1g# ��K*E�������.���gd=��#��>�"�%H���v�.uQ�ťx���\�~0�o�e�#�Y�O�%0[B@J���׽w��E�����ͧ5�/?kF��ߒ�������ZN�����26�xg+:�7-0���z���A�H��^R���|r�A���@$;�[eJp��#���<�����3Β����XlxVHYEB     400      e0�k�]�����&�B�FGR�Ʋy$%��*kћ�G��x�#}�w�M���(�������)%��@�qc�:����R�]0l[�J�
����8�iy�vpO��%��Z�5:W�LY�d�:��mR@����/0M�.����OunC]�};F��Ly�rM�i���aV���0��i�����a�`,H���)�aJD���Wl8���*�f���w�TXlxVHYEB     400      e0� Ӱ��a�N/����W�����<,^]3L�d�.*J��슍��p.@�/���zt�x^���>@�r��_�ɂ��հ�#j?ѿ-���b0�Ek�����#�
`*|K\�9�{����σ��}'���g�������'P`�jV&A ?H'���rD'��W��i�S"���br��e效O���o��>��d�ؘ�g�f8�R0�o���N���F�.���XlxVHYEB     400      e0%���z�Ğ��?U���_���+��f0��U~��[���
K�~�.b����*�GK�1YU�_>Σ��Z�C�Ϲ�Y0wHqX �.�3�7�!�6���+�jͫ����12#���gk"�c�b��[m�D�?�#��`�u���.�|:z�A����	� ��`���<��3_���	�K3��6�2x�s6�
��� �,����P׋��)������XlxVHYEB     400     1a0z6g���y�E��lB�,3��k.�0�m93���r��r$�<�7���wd��)��eȁmq�I*��Xp�Z�q�*����������ԏ�ݥ�ү?�t)�;�MP���v��pH�GK 	E<pUeo�װK*TFZE�:!I$a�{hT|���6NA�Hp*~�O��L~Х�Qs��('`�����q� �sK0���H$� �"׏�F�� �>ɉv���*3w��*��Y����ùbN��t+��>���N�������B�ر�X�͂�F�>��\ATWc� ��$�%�:�@��Sc)R�6q���S���(̤D�*n�Ұ����oH�6���'���·��F.��JK����]T���'�nT�da������s ~,'����2Y����� v�u���v'O�4��XlxVHYEB     400     110'M1�a|��*p	�Ӹt����3}<o�l�8yYX���zg��2�o�I�����=Ol�Z8���)߹J1Dc����2{��zQ��X�����yJ [:���*����^7D�K.�ۉ�Beh��b,�����bH�7?�	���Y��v7S�ϭЛ�� +�/��E���k��̢M��FC�9/w���Pz�����j����g��2� q.�	�*����S��ߞl�f�ͅW�D%�1Mq^�M%���,�g���[+XlxVHYEB     400     1804�-��r�z��
`���� ��E�����p�V?���i��Nq����ѾpH�f&��j�K��y J��� �.�'�ũ������!�;�����	�\��
%0��z�ѡu�O�;wc�A�+�h��-� M��tn���bQ�A��S�dho��x�A��������Ҟ`5)�=a�T���}���Α�;��%m�h)�B�c᱑���- v�z���@�	��j�=Z�Z��輞�k��Ѓ�6+˖,��Hs�O
���SQ�=�*��%�9W(��(�F#�ŗr�J3�\9�K^q�\nC�
~N���w���O�_�B�>�gW���a���2�qf�=a��Ҳ�p�3�!ib��E��	vn?��5t�7���G�XlxVHYEB     400     120��:-��YH������,�ƓR�z��R9�#����a$y��>
�s��F?a��dV�0�2wvy�m_=�&�e��*�/����r|*�V=io~�l��1��x��l�[���a������xS�\ﾯ)����iFi1�HV- oDF�Z�/D�3
����XkI��G�螘�1��M�z�?í����VL24&#z����s��nס�/���S�.w
�1H������]�"%:�pj��atO_F$0�c���g�
r�t��\>3�V-G����ڳjXlxVHYEB     400     130!i�ؿ.$3�K���.��7z��6wh���Pz��g{�bnuX�]
�T�Y��B���v~�X�
�8��"=`�D�O8'&d�Ć��b
�/c8�	�>�놌���-�3�55��Moމ�市1�I��c��_����Fl #H�;��eHh����#�`ż1u���n����%g�k7a��`t&Z6t�n��}�cL������l�?������Lq����n�f�6 ��b�9��=�3L*�V,���z��Y4��?�[�y�2����߇ �`�O����<,i��a��rXlxVHYEB     400     120�H��2iE�ٙ�:�ay��.7D,�_�lQۄ�e���u�+�5����aϭ�nZ��|�]��9���z��}��QpZO]�T�*O�4F�	]���F^ȩ�����1��0���>�T���^d�!_ԛ��;7� <8�s%��0�\5�%0'�+O�$HG�kˤP5�O��Tid���Nhd�ד�o�%��]�E�H���E6�Y��	�o58�Uo����j�E�_q��V�q ���V&ҏQ��lI��HM~$�Y7�RI�|�q#��q�K��HNaǛ#f����XlxVHYEB     400     140�]$>ez�{=$]*�Cf�5����Q�d���ni�M�v���]�ظe���c-L:�4�eDNjBr6�4[�u�	,�e�&�bj�,�ဗc�v�.�(�i��.~)(s��Zn�BBI���b�lUd����[/���$d���+/���v�4:,�U[Ӱu%��l�%_=.�������z`�<���P�䢫o�
9�/ĉ*-���/Q�A\�<��ς=���R�;�sjT;iˡ��	+;I��f��B�):-+1j�4��A��i�!�
o��,�$f��r�����B��#�S�nc� �]�ʫ�۝!�I�B�)GOB��u�XlxVHYEB     400     140��it�YjG9q$H-��!�����șOhܕ���M�R۴�\\�7c��U��m�@r���Ƿ�?�/��L%8Cg��ϴ �������f`��84��PÁ�Q)Y�=b��@L���� ������p/ޡ����G|f���|#e��R>��?+!���0��)b��~�����&�,��9�
��x���	d�Y'�,�6��n���"�u~!6�1���C��[���Ǘ��ήi���k��Β���O�l%M)$e��ɹ�$�ރ�a!�M;d"cv-:��zݫZ�w�f{���ȏ11B`���0cn��o/XlxVHYEB     400     120������|��HXEeDx=�9��+�������,6��v��u�ú�,�JYd��w����Z�'�����~��b[�l>Ȥ�8r�a�u�(ew�Ճ?$I�%`������qL���-������|�>La�a��oGX�O-re�_/;��jN��7CQ�E�7��ǌ���4��ܔr�r8������I;��H�X.xV�QgjO`)���6���nM���IMVTE�,�K�u+�Ǧ��_6ExoC��Q�j��C-��q﶐b�L+xVXlxVHYEB     400     140�{�O�I�DC����Q�^L����ǌ��|f�	D��FEB�<����3&N�J-�8.���nN�m��H$u����Wl⛫��l{Dc�Z\tb�	M��]�q�5�x�զ�z�v�|�2�D���ß�V_�R>j'�&C+�Ò^OF�O�5��^,���V��Hd�#-�]����B\�>cΕI���
±8H� ���!w�B<珶Xh��ť݋[��F��5Za�^�W���	|�r7��}�'��UX���5�3�#ӶzN�~`�|����[{\��4ɭoÛ	P����J�x�j̴��)w�F�To7o��섫XlxVHYEB     400     120"�~D�므�O�B��UͅX\���g#ι��?������6'Q�\�U,%�`	����+6��#Tm�GK?j4�|�p6~u^o �0��e��q���m��wY�8`i�+2��/�	]_/�[%`*'�D��4);����(d����P�$D��;���4��=	Dn��Q�.��j���9����"����Y�όT�0��;;9����캙0�[�`��]��7���g �1���	���%��u�򠃽�p;]�C�J9ѣ�4���:5�#�|F1iS�9��b�ϏXlxVHYEB     400     130�v-M[�e����˸t�\XW���ˑ� ��ER�CW�2h�D���B�9=��'1����y�`��6���0=3����$�\���i� 4Ԭ�*��я��q従K!�����ވ=�J����4mF�( F�r)�{֖�c����6��ٟ��	Nd��c��E���R��ǫQ�d$ة#�u"�!�s����bȂ���s"'��=px�zb��fm��L�<�6sJ�v��on�o�>�n1�&��*E`�� ԬD.P;�Ϛ1��)�~|ǌfK��>6# �C�dI+�0�.�љl��r�LXlxVHYEB     400     120�7X\�87u��2���E����J��X�����P����$|��a�&{_j ^�Ŧ�u�!�r�3���9-Nl����3u_q�rz��;�Ȯ�;�
���Gv���-|�%H����s��	3-:n�u�tx��Ӯ���?9w�co&�Eh|X��4�48�)F�v��V� ���aI�s��pHEJT���h�FA���r���w���@���4�\�+�n�C�}@�ݭKg>��e���Ď< �-�]Z�`xʗL,���A�z�χ�F�P#��We�����XlxVHYEB     400     140����u߶g\�٨�bϳ��V�a��K��^k��پ��rn@O]����tE�rځ4`�>���%�Di3�޶���l/�Np7����K�kZ�S�)��d@	���Z���)�K����p�������y�W��O�jE�Z��:
(�-��巿M_aU�~��.�[ܪ)2����T]�<����fB^L�xEf.[�D����I(�|W�;ˉX�\��rj����B�Z1�����c��&&�����ox.4<�R"��BS�0����p �D���Um���\-ʛs�;6�HG��驰�XlxVHYEB     400     140��it�YjG9q$H-���[X�]b������.���1�x��jT��R5_�]M�Vŝ���< P񽑠�_
U����i�]ԏ��1��$0����D��C��m7�#��w�;����P6�Z\��ΠD;��7����0]�n�ƶjo�h���M��=6$�ܾ9�����ďW����ۄ�]�G�lvj��6��ČD�>8:s�YM�-9��~�>�lx��e�g]&�b�/���� �-�j̀ds�Q.��`W�<|��������2�!�S+� R9���d��+@(�����ZA��i�|�%�r�zq8PI�WDZXlxVHYEB     400     120vZ����2
�h��w�u_^'�q'��.���Mo��KI�c>c(�ʵƓVu)�D�Z\�8v�3�&ʏ�1�P	ųq��Yu
v�*l�wӾi
���h�� X�KZ�������S�EMg��S� Eƭ��d���U���'�Hk�#�5��d]R��B���J�W���Y�F���K���^8S�q���<�H��7"h��M#<GVGJ��N���.�3_����f�V�kw�2FZ�j�칥�~#���ƫu�_�[�1��"�;=L��۩ڼNfe��R;b���XlxVHYEB     400     140a��`OaY[,��!p�b�P��\UL/�>z�9�\��J���� ko�V�/0$��,l���Q�vLV�����]���n��qv;��"h���","T5y.��ӛ�(\I���ڏ���S�z>������j�Gsi�8f�VJ��"H�N�k�(��_�l� ̩�Jـc_���J���+�7u�m�-��m$��w�j���'�h-�NN�Yz��giB/y5ĲT���Љ6�s�D�޻���I&�w���Y�ڻ�'~S��6��7=�@��M�׌��
U�r����<ﱂX3��Tu�#���XlxVHYEB     400     120"�~D�므�O�B�����D�>m�Y�z���V^Xh�t^�*�ct�� {֥��W�Ж��~��;gdF� Rd���b�uB4�7���ZS�>+vV&� r�b�?�?�v��eA��ʑ�` 蔝8�C�D�G�z��r��jbFi����u���G;NQ�c��{NEK���dw׫/�܋h�K	�锩؂,�/�4GFdO�ur�B:�m_����+k՞�3�)jo��%�^T�����V�~#�h���-a<cVݳEɬȟ 񙳨YN\B:��)��ڇ����XlxVHYEB     400     130�<�O�m������k�G��R�*xԔ �%�h6�����Նg�?�J���@��w��Ւx��i5�T��]��U4ԭ����۫�Хh
j1�֑3W��%�,)�?~㢒�4�;���J��B;'��)��U�D��y���<�ǿi�g����n�j2��LȊ��iV`���'��}Ca3nS��٢� ��i<2�FXr�I�<<���-�zu�6���2}ܡ���M[�&q�_��]�_���S9� m��}���X/����Q��+0ٴ�L���v�6%�B�3�7XlxVHYEB     400     130H$�t�Z�!T�[�K�<3̾<�yxE���Pa��/+3@٦� I�5� ��5hd`��種�+in�Q�bc���c\�ii��b�uf� )>�i�w���i�C��(�q�)� �s�
e�{WqC�ar��Z%1����oF��J����p�:�S�ٷ�Ü#s�8���-�3��'��T(���ˇ�.��6<o8^�cf�|����u�F|5S�C"]C�c����<"�ٝ�+�'2n��3u�t��,i���@����y�vT�'�mP��}B p51<�#^��.(PW��65��*���FXlxVHYEB     400     140��ͭ���R��,ԝyZ�˥R����Υ���kz���o��d�~�����x`��N�^�of�v�k֡���)pFD�A]����3\��݉�����]���9�(]��ޚ=� �?
�&���c�
h}(e�S�8�;��_��V#Kx%s��S�T�~=�g��9_��{���[��Vȱ�	V�e�Iǹ(���u��2ю����՚KQE'��?�3#t����B��[��i��
D�Lװ�_�w�K�M�	\�jUx>_cW�r嶷��~��'�o���� U�5}>ma0��qEN�<1ڿW�Z�2���XlxVHYEB     400     150��it�YjG9q$H-�����ԣ>L",B���C��pMd�|��1M�-����_��P��?�iQ��n:^�h�r�`=d�{�Z�]���~8�T4��H#�JP�B�s�m ��$خ�:�&X�o!�v�G�m�T1� �L@��L( !q���#�GmƩ����4���A<�SE���P�� �(�Y�:Np��v�pgіt���">�P���FL�,��-��J��(t
�U|��T���s��U��[z*ݡ>��6�%���s�gŻ�9B�+5��#ٍ����_؎>��\rJ�;Zj��O6z�%��C߇F��Y�N�?���XlxVHYEB     400     120���S�b�Դ6��.�Q#\�yM|/�t��K�������������=��e�#){��`��=#�\\�������8��#Kz��.�z3D��"b�}�}كʦ��_e���y�8(q慭�;!a4��+;^��e\O�,4A�f{�N�E��jDoS��V���V"���?�{�|�X~�����:����bI���.�Ñȓo�=�*ޭ��v,ۧª~�$y&�>���l�,08���gОq���I-`tS\�E�C�K ��P����\��M/���XlxVHYEB     400     140��bm���'v�JȷZ���2`ŦTp�t�(Y�� �d�+B�]�cb�XZk�[T���J��y����>�7�t��o�͍���bRo�$h��Cv�gqZ��$�����Z:+"�Dp���là�fQ�g�g	�>S�ټ��4׶,��0��.R=^8�3a�N�d�?g[�Q�o��5M�$ S[&E��I+M3.���2�P��=�.<��P�٠"��.t�K�昝�����E�*GoL��Ҭ�F9>�XZ�Ǘ�L���ns��߱:l2DL��3�1��I��V�8�t��4�En�b����
�>Cw�XlxVHYEB     400     120��y2��c9AS���2�}��%b�k#�z�B=�8ԟ��p���I�/�2���"����R%���^n�s(U�ʄ�Hj�Ti���?B�b����@�*Y[��9=��u(T��+�U���1�i9Q�"��+~��#f�_7����J�%
�K%)� G��w�BQ��ˑfhK?N#*��g���qG1h�R״�h s�N�Z��=_�Y��b$�R7��!3�����3?��i�o��\����{aSp=���y�aR��]=T��8�^酕��XlxVHYEB     400     130�v-M[�e����˸t�\g���	CH(�� r�O�_(��[��]m��sﺬĖ18�������m��W�ee�jF:��W��	hPr�)e�'�*�Ѱ(��}j��+&�O��J��9�s�1Վ�fȯj��M�0$��W�cT�-;�kʈ1�$����:l����tV(�ܩP}_�V�Y�'Q����	���R�5�4X�=�W�Ox����;��}�mcj����R����r:�����'m�ǣ�Uu�*G�&��R)�:�%oڧr2��8\�w����C{{��o8k�arcPXlxVHYEB     400     130H$�t�Z�!T�[�K�<AZ������G��|�cO��5��HR\m,�V(�1�{{�� Bː7���U�uRU?���� (|@^�=p�`��z��S~� �?���!�x4�*+6�~K,�l#Ї�bx��2�WK%�6C��!጖v7��0&خ$�='��z(�'t�7���k�hhѷ
%�C.���n��^>����6��I(NV@�s�N$u��b�mjv�v+�qe҉f4�96���=�ag�Kv]��Q���m��r�(��SǢ����Z�R��Zm[v�s�lHY��C!�\/XlxVHYEB     400     140T�,Z�i,}������p𽮴��=���#eO8;��OJ���k��^��nԙĎ)9��'½4��J�� �mj)sWZߡ�h8h����PM��jV�4"��*�Jl����pIU�.�Xו4�	pi1'{3�A�= !h���U}[>�DFN{��`���a9�35T���,���PZd9P�Cx�N�AZzdp�s��ނ��kOk^��
��� ���m��D��	���g,͗��쥽���}�&(ҙ:��Ӷ)a/wB6�C��C�'����j!'�M֒��х���,a�u>n+�ڪ�2��՗�XlxVHYEB     400     150��it�YjG9q$H-�ᰳ�a�⥥��ͣ��E -X�B���N�J��Fa�ez� �o��5\� 3����v=��n�>w����_"n����Z�%_��=7�����U��v�pJ�mq��]�=�Lr�kr���؊N��IW�R���6)<.����RR�c����,�]r�WΗ���$v�z�ނQ/�Ô>�v��j	���"rX~�$9�
7�]������kYr=×@ǒi�N������eZ���N}�dP6�]����vb��\�xDy��|�R�=��Z�q����E�0e���J�RW�[��+���M�C.��.�N8������Z�U�\\�yXlxVHYEB     400     110|���B�@@��xq�
q�E(�V��4�1	m����h���]�2>8	Rw'9}NNK6_���3��NJ��RO�#@�;xr��*N�Mv���CN*u��ԬY�-h` �z��E�J���3�OmM�R�W�LoNDM=n|Uɱ���p 	^��Ф^?�<�nD�&U��I� lG�Q�|��&� *�ɜYK"]��ȱ�az��3@��7�!D�S���x42�Fߐ,��Q�;�íӖ4�USIK��v��q�d��/�8m�OXlxVHYEB     400     140�����:jvy�C7}���׌Xf�y�b��ek���7�E�>r��SPG�~[yMV&Z�W��~/�`��8�NWo%��>ͥL�b��,Y�W}&�f����;=�yL�QI��8�<k�9eе�� ��u9�qn���3ė�5 �Z���([�zmH�B��"�յ����vjk���ރ�u#]>��
��s�_F�?;���P�Aw,c�(1�Wuȁ���'��4�;�h��VP~4R��ք0ȬF�7g���.�2lJ��'�s?����Y�	_a�����l���)3�ʻ�E�[]�ad�#E�n���|�r�XlxVHYEB     400     120"�~D�므�O�B���%-ͅ��k?�;A�R�Sn��N���X�0U;KPZT�O����ӺNE�S�{ uz���b:j2>��(�'U+����.���1p�>	> ���1��R�NK���H5K(8@t��6^6�04G�ŀ,�u�8����\І֑v�G]6E0L���В�[��˥�}�4U�>Q�9�˿=t_S�,M���1jȣQ��Pgk�SV��Nt!m0���.
�,�&T��I"�ֱ�����OBȩ�R`a<~������3&��XlxVHYEB     400     130����£"�R�ڪ�]��C�'*5�.���6,����
w���ދ~R����ΆE��钽t�FR` ���������>"�����jdx޷�����,ߐ&ܭ
��	��ñ�������E~T��{0�S(sz�8�??*E���4�;dk������_AOR��)� TS��d���l�?U/^�_�U8s�,"��j]�s�����wG��WΏ�9ɜw��G��zJ��d���L_�MK`1x�h�,(x=F}W��5Ԫ��Kl#���T���i����|")ʇ]KH%�^��þ,?���u�XlxVHYEB     400     130��Zl��SS�͹fYnv}+)��D������֩�Os�ؑc䝍GI�lt��T��_/t����5OLgJ��<rX��/}�b|�K������g^�v�	�C��%��*���e�1�p�2����)�^�o�M�%�5�dΞ������R������*�1�*�~k\� Q��oWH�A.�-r}c[k�ׁ�'R��~�н傯U��	�/�F	��!5��hnN:<}�q�w-��jgT�[Kbu���-_�MM�,��V�B�k��G�]l���ǟ�H	�܊���-��U1�"�p�XlxVHYEB     400     140�[d'�����j�E�u�$׭��e`
@_W.m�q��/��׸e��|����s�����t���J8)#-޽MX� /�"�#��h�T�z	�Йt.~*�'�T�X�@+��Ok��`�9Ow�T�5I���&��'��l2�H�?�0J�����g�>S�ā,L���yV�:�ɓS�$��(�S���yT }��6r���A�u�"�y�gh)�| 8��(�\1��.���]y�"~��~���������f"pMW@�@�R�G&q)�-� e9Y�q�E��e�k]2ǻ�[�x�h��(�P�����i��R���Y�P��gCNXlxVHYEB     400     1600 ��d��h��k�,���Ja8��p��<���+�Ԁ~����qbVe�_҉�\���We�t&$Nҏ��'"���5��A /�^�o������� ��Aj�c��:7��%�խ@��N���Ik E����q�A<�g#��#�
�_B��ћE�4
w�,�L�+K�Z��~6���@z��zH]�t�tN�6��Уp0��E�����Z<����A`���`�*��dT��#�AT;�\`��R����tȩ�3�녴�(`��g �Y�N�F��/�&�Hz��A)˨C<�%ݱ�c�j'r��,2����bP�	sW-�^L㿗��������%�u�ޚXlxVHYEB     400     100�D����L�hZ��U+4a�Q�i�`pS���v?�7ua�.s�7�}�� %;���7B��:���s�U��K~����+P�Ci������hhz�
��I�4Q�{ya]l%����dS_皲�Mx���_�)��	9���������_��'�s���Nj}{��Ҽ$0g����������4�ݕ����RB�<� �4��b�-Л�G�H�e��v���E�� V&� �pU(�{xpyC(�!�� Q��JOXlxVHYEB     400     150��|;@����g4m�ީ�O-�x�� Y�"DY�$u� ���0���R_ǖ�Ci.��C����U�N�ي�~�<;��@�5|Z.aab`ߙ�_�$i�����2Y��
!�_��7��vl~n8cK����i�M�	�݇�7R��,h�Dr,a٠��s�r[Ҩ����ı�
�����GB�h.�Y��1�j��l�=X��S�O��T��_����ٷ�=�����i���@�1HM�Y&/�BĊ\�
ŗr��Wp�q�C=m$}��x�8�TMf�w)'i��	�>K�Ű��ϐ�����q�W;-0p5{_��F�kVt�^�C~>�e���XlxVHYEB     400     120��a��)3~��g�x+�}�e��D���q@_�tw��2���O	_�2A˜�-�7����8ğ�0�ڪ�L�����L{b���3�6�)�,䔤��V)-�M3�K�@zY>�RJkE�XQ����h�l(+v0�N�(�m(t���H[;�&?É:1జ��9AV�UEe�=r�L�����LclZ.%,�?�I����.ZsMc�.N�f��}��W�@��
�R�qL��q��ގN��8�cM~R�� �J�fS��$W�^��&� ���^�ʁX����a��XlxVHYEB     400     130� �����L�u�y�*Lhh�W=��E��Bt.�c�$b��,XUB�{0qE���!j�:����=0��F��u|�ʆ��;c"~%l2�r=����_���T>l]n���bC�JB	�j���OU�/��q�肢�pj��QQ�b�Zl� d#�u���!o>8���a��
'�bh���4��MM]��y�Ux!!��wj��K _�C���3�Q(ZT��"��O{�oFH��G�	����R�whoA��#?�Uw�d:��e���5R��m��>�9R֧�%� ×CG�Y��pc#���%eAXlxVHYEB     400     120�¢�H��l�Q�1v���wI�?୧ј� {=�8ʥ<n��*�5��p��b���#ϡn����F�L:)���@��,�?�C���#[B��x'x�9�H9�FwB�7�X��f�v	<�@χ8/h$�
���%��m�nG��|�����W�;	�[Oi�U]�Ł�QQ��n��w�A�Y�P߭n��Q�Ć/*K&�f��Zd)�� z�9
I��o	{l]��7LH�bӶ`i���aV�@�������Oc��,��)��%/11���)Pٽ�o��v{�n�HXlxVHYEB     400     140��{AZe�gZF���t�xgV�V��ͦ*COj�-F���и�H�@0�ۧäg�F�ȟ+̶
�L���D��P	�[}y��x�C,�� M}d-R�d�V���"��ܚ��ZSƸc� ���T3��"o!퍿��	�>�W}�!�
�fU�ѻ�  ���wI<�Qc>��6&�?0s_�sU�Ɠ�<9��XCl���c���)C ���@��F���M��؈S��ݞg��b�ᬌZb�z�vȴX���ns���'��R�>��HƏ�#��y�eQLܭ̫�R)?��V(�����{V8��x�ԿN}��XlxVHYEB     400     1404j���7*���Z����w��O�0.-�<����pz��G��_)�_�s6����K0�5��`�g�������\[�
(�yc��{p��`'8��n��X�c���bO1�G�DB��S�t-"���q��˼���nVg�m��H�i��&�@�t0��pP2��� ~��,�o��&�{]O�0�o����0h�G5�qA $�k)�� �i��=����"~jn�g<#m��}>8�?ւCZ�{ ��X!�%A���rI G.5���8��nc�� {W�(�����i��F,R��v�f����Ծ�*�M�/�-�z�_��I!�XlxVHYEB     400     120m��9<�v�Ѕ��R}O��+�#-Ӵ8�H֕Ĵ�M{O�)!�.���F�dŷ}o��r�d�^��v�����Ԑ^�|�|�	���9��	ٱ=�W�2���-�G��'��58f�)��~Ykg"�`µP���on��F�漢nT��
��k ��<�G�ou:/?!m�I��<D��������h&�:��2l�#́fH�J������a�_�Ǹ%����7:x�N |�54���w	��wV�%���Ȣ|��X_�)��1T���o�u-b M��WQ9:Yf�XlxVHYEB     400     140����UMbZ�/�ܗ>=��/�s�e�����t0W�Ay�OZ�6{��:Z�漦طb��VB�</P��%°6���t��wb}̰l"�r�^3�y�j�[��.ß����*��a��a>V�����I���fK�B�0	��ot,9�a���V������:+�(mY/l�_����@'2�����pbV���:�.ݱTH���W`1��9H�J�u�D����EO���r�//��r᪡�$�cV+C�\P���>�o�����?���i�����5
QK0б��	c�1��m�N��E<$A��p-����l�<�q�лb�XlxVHYEB     400     130íz}��DH�6�U6��3b�!�/۬B#s2�ô�yE��t}}/P��ޝ	��1dXN��"�b[��b&��30:�C��xU���9�iܐ�yz�����e����g��ھ
�f�`�?dp�� Qӱ��z���,j��=@��܀~��Rh��]ƆA�2b �3CQ|/�y��#з=<E!����e�3>~�!W���.4���q�U� ME�t�}��	a�Z�}��R���܏Go�K���S��v1���O�0)7��:�s�z!{�[?�����g;�Qq|e/[6{8��ٖ3�XlxVHYEB     400     160�����V�l 2UEJw^<���$+'q�hŤ`��V�gHg[���K�ѻ�Q%���ݕ"�|<�.l�n6,����D}|�Ydr��O~9PV��'�T1D�]f��Qo�F�]���i�~�Pm8�4F��Btk�3$��t4���$��Z�*������	���h\?��� �����٠�'��Y\a4���m}�$����y%�3k�0P�i���"o ��T��u�'�9�,�J�T�WL���1'GFdfi���C�c��ܠG�@�҆�r�]��tv'�6|6���,�Y$���/�p���v��e�Hh�������"_�p��0<+)��}8�h�~�^XlxVHYEB     400      e0�6p�$)b�T�n��%[�Y�|�Ϥ�b߇�3�Nג��_n:�M��V*�[����ft�܃��3�Hv����2}r�>ؑ��#J�		�uk����H@�ȏ����&�p����,�R�O��@�����$$_��lG:~C���vˈ{�n��1^&��˙��T#F���� ������Q1�C�=�!�bm%W�mu��������E��jq����XlxVHYEB     400     150�	��]ˢ�M��S�?əI��VE�*�
�(*�������2�వ8lǫ4�i�C�4Ht����e��٫���������n]f<����ρUv��bU�����B(j;�@3iSkQ*�6j�=�-F?�<�k.	�4z�yz>��]�����j$�t�!nC����#��g�@��a����۩�ٵj)��|���xZB��cdN\���nII���0��i<:��#������c,��NuY��`���j�m�=|!*i:�l"��Z��8����b��΅��0x�J�*(��Uy�-��i�����=2���M����Z���C�<L�[��U�H�E�XlxVHYEB     400     160getEk�<kH5%vt���`	�I���<Ǫ7���4�>d��B+� �[R~��*��$ڷ���)��N��r^���׷EJ���m�e�� �0N��c�L���3�(�B�����1d�g�����^F�K�?N#�%��eg�?y��5�(4��{�Ɣ1ATՇ�!���7Ov�*�^�7R �a̅�*{ 13�ڴW$�B�Lz��#�(���}����z�</q���3�%�v�@�|��<�_��+��v���Y^�?c<�g���cU]S�jQd�_��O��2 Z'�N�J|�s2��T'��Ъ�8��hw�z�uA�ح$D雝t�X��C�m1���g옍�'MXlxVHYEB     400     120m��9<�v�Ѕ��R}O����#���	��0P�/!և�/>�
jx�v���^bc]�ˎ9��D�T�FJZ	8&�@��@�fo�AcpD�Mbx@�����Z��gGg�̕b����m��GATȌ�H��sS.P�$b����m=Q^�-ym�%[�s/��|:1�2��a?�%�!���`$�_j����g(͡�8�_�l�$k�0�+����%\V�:�R$�r�Q��T�G2|Rhs�H���ϻ�)B�acx���_^r&�ms������XlxVHYEB     400     130~y�r���hw�Z��h��ьY� �,;� +����Е��y��[X��\� �����.�����g�"�`�n(/ZA�=C��33QPY�=�v�ȩ�Ff�?Z��۾xV
�,#5������C���:��&:�/�R�O�Af��7|%�C��H醺��W�[�z ����Q��ϴT�>E�X?7<�NUX���O+���?Н7�v��海���~4M1A/�*�o�%[�+�$��]2@5�/��M\��#ʲ?ʥ��D�b;PbUv%��N�.����`�R�Yw�p/#	(�-Uc�ZF�|�1~��I�XlxVHYEB     400     140ɰ�i/r�����+��U6�=��S7���Xо��ogwDIGq�������8�V=[}���s��������>����K��n����Z�ژD={Dٔ%m��_���`~��9�5��U��ś��E#�2b��xwZKq�Dp=e�-�	���r�V��ʂ�ejP�/Fq�߀u��g��\���}*�6#����v���U�\8�&��'��Z^�$���tg��D�Q�H�v���3��#~��ñ1˾C��1<�>�q��u�Չ�"m�m�5}��RX��F���KR��65����m�h������R���UJ:��'�CߎXlxVHYEB     400     160����/��[��\eJ��Ҩ¥�Zu!6}D�ܟ���y�W�3�AN����R?Aa�ަ�ad�̝�_� b�����I�rY>�
z���L?�h�+�ڒY�N%����	�|+�o'H�����l��wt�vА&0�L����T˯Z~B�ȳ�VV(	�6� %i矄r[���"�'���8�gI�"�
Yb��g"�ڏ����߻����1��q\�FqgO��p��,�$��#D,E]P�!z�Ŏg�:�"'���T��S�^]�i��j��Y+Yf!pP� M��Ik&�D���Z��T�/"����N��߉�s��Z�`�r��qTc�J��ڋXlxVHYEB     400      e0M�1
҄�H1=<:�6�Ҭ��Q����ɂ�@�٪����/�i ���C��^P�	l,ZP��p�U�F}m[��*|e�;���g�!�E�!ԩ�����M��t$	0�П ��<bf!�(��N	����S��ڄƿ���N@��F���O���bxVF�α;G��Rwۡn����F�����]|�����b%��J%��
�F���
D��`XlxVHYEB     400     170N�����V���sM�Ʌ�B�&JZ��A"�j�ePJDG��O"y]k�]'5t��<?���W�l�;�<�z�7�h1?�ܒ��n|�2�̟��c�a�t�����y� �06�6�V��*H�#/as��\{T(E�-~bs�n���<Z �
���r
Y�Z_���t9?�a͋\���*;���/�)�y��ն 5i�;��$��֌��UȲ�{y���*r���}�a;5�3�w�"tӰN0�w��;��X�/F-��}(�#�S��ہ�`X�"��}��rQv�K��퐅���Y���XB��l��e�Vҫ�����Iz���=Lp���p�|�|i���A�!J3`d9&� 4H�Q����k���+pxXlxVHYEB     400     150A'�C��E�XCb�̶t��$~����.��2m��::t�cDl
�Q���o+���|up�|�pm7�����WZLƕX��4�1�F��h���}e�nlB�8m�g��^i������)�K+��۰$yD�r�s��l�J	H�w�WF0��B�츘J�7S!�)G�+��X�%��,�Q7o�Y;�,�U�Ҥ���t7v1dT�)S$y����I�Z�Uk\�*�I�����ݲH���
r^��'�6s���fx-��|��F�6��HAA~!�T�j�Tǝ���y���\�.�_�fO�4��s4.2�_�<���wR�(�`���:�Fx���]}��wXlxVHYEB     400     130zU�����AHNZ)Im�m�XSc�eYv�a쵲'$��j9gL��3�U?S7�7�*�&�q�� �O;��Y:Ct�Ԁ� ���G������F6bz�6��J�ʥQK�e�;���s�|�Ll Y�I�@���֯����[�����~2}��:5Bn��5#8VH�;s�>���5$��$)��̸D>]���ӜF0xq�WX�!�?Z��9Q�A&�FMAPV�[\�ޫ��֑�v�5�q�����2۶�98��F���mb��~̄@��j�m������"-a�o�������!9��H����-�FXlxVHYEB     400     130�䛠K�q)�
�a�eI�u�T��;��T�Ԣ�����I)c��8Y1������5x��/D�x�<F����/i߭5�B�,9������ %n��h04ɧ&YH�6������v���_T�_���l��������p���m��_=H֦��������W�P��2��/͸}Q�mG���6�o\}��u$<��難2R�`/
�aj�#����ej��^�K)�X���6ݓD@��ʘ�S�^��S���˰-���fzqKי�f A%|�p72�o�d�4~��XlxVHYEB     1b3      e0��$8J�����L��Zk� �ެ�(F�����F~�HP�!���� $-;.��p����jIs bk�&�|�.�l�EJ|�^��n9��;�x�:]�܃�h��tpp�?�$G�<�B�V1�&F�p{ ��e@�N���Vē���U?�٠�Y���, �����R/%����ז�}��!�x��~϶��~qD滣��#��C_]�|�g����)��Ԝ