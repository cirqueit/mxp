��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����2
�`��C����#]d��|fBk������F����)�̑�Iz��:K̠��h)�K��nhJ���TD���q���#��!*��@����Jγa�jbK��ј��M(1X/)�Vb(���)��ަo��fG�3�L`� �pFG"���<�+ތZ���OT�-��hҬ>�a��+6�\Fʠ���˓���^/�eה��P;%٦]�%Q��QN��T�U�P�kiP8�x�y߇Vz��.
���R%d��:�2��{ܿ_��������H r~P�<�#�跡pKg� #�Ls�y�P�����"Y��w$=ģo�K��Bs	�Rf^A2<g�E��߂�`:|�%�s��*y�@5]�s�p�V[�?lr2�\������L"nP�h�'m������{�(�g��9� ۶�MYut��yZ�`
���
�.��b�V�kቼvv���D��e��w�a��


O�j!�<�4��=5�2ʱ����|��#S3��|>�"%!��/�FS�4@j���^Ə�B���$�'�p[��%:��y�c@r�56}��mFx�u�N*-�:����A�����`s�T�*��ݺ5�B��R�VpnO�U��o[Sa�X6E�1�;���E0q����4�ce�Q���D�GF�ᨑ�-�Q�Kv�䟏�(�o=��S���b����k�E����"BH��ThjZ��r�3��@��{���81] �o���7�z�]lE�3E�������	|�EJ���$�q �H���K���Py7���΍F���%��VY�=��\��,.�DT\�$Q���i8Z�qV���ep��Nyuk�6�ě�
��T����=0?=�`��=	�(d��Dhc��g>��L��.9�n��N�$.)��΅LG�,僢���O��՘_�
��n�����G�x,$JnQG�W�0�گ-PC`��=RD��v��n����YZ%�ڶ�^�D�y�P!_'8*6�~ ��/�o! ��N���>�:OD��˫X	���OZye�N;��!��i/���j��lt�q����\+cAk'|;�gNϼ�<HL:��^�-��6{ɇ�g�M�- ���*|1��*T�[DŸ���_j��FU{��K+���1�r�2�/Z��w����%�N��hK�y�Q��j03>��홅�G<(�؀�'�/脏�E�8�D]��I�7lڶ���v:K��i	:۶��	L凃��F|Y���l�@����i%-_�x��IO�g�����Iz�U�� �}��=o+V�>�]>��`''h0B���'l�;�;���7������E�d��;j����'uG�=��$$}��P��F���X-i/�݁�;�ͪ��J6@���HW �M,�`v��t�m�<�4��tR:��!�	������|���"�d�EQ�����4���~8MG�d�7��p
Z��a;

���Q�D�)��[�F�lU�f��.�-H��b���� c{�2�H.77�9�3���&íׅ�2�3���89	�Dg��g��AqQ$R���O��E�څDDC�!�!��d/���k"V�H��L�Q�!\[����yLl"%�����sd�����QW�ioR��8��/��'$|�����޵þ�d�~��H��K���ȱ�_��@������Q5�is�b�d��N^���eM�(Zl
��u��ߘ+kd���,�wd*�b:�}${����[�vB�^�j���*��I��OV/�C��#ڭko@�E�AxV��p�o�o��� s�D̚�7ii�}	6��od������yq�S3�3m:~Wp�yҢ�Xpo�j�r?4+�`��:F0����� 5���e�ۍ���F���$���IiP�˗+�*�i�l�6M�b�ז�7ES���јi�ȥDe�._b�2��Se�y��ً�M?$Ήx�c�d�X��w(r�uA���UN�V�_�: ����q��Ҵ�#�Խ�+�r�g!9J��F�R� �W�N6�ʞ=ސ=e�3Xi���gֿ��T�F��T>�SsP�!���,��e}��K&���td�^u�`w�u�_�9�p�?�`���z��I)���;���d���G~M={�rAENldo��Δ݀�Υ�6��0s&X��'��˛=���m�H���:��3�-T���})��ߏ�������4/��"\m��� pk�8d�ʁ���,��w>|���l���@u
߬�UV.�I��{�3�O�D�5zܖCd�P�m*�s1�R?�0�Ԭ���Sa��Il��竆�m�X$*�D�QR�Dv����D�D��dy��� 7�8|2��D����a*�P���R��j4�+t�{�y��)�S�Q�G��6�ς����g`�A�;�8�D�u��ڷ��*%�z鍯wў��76�=i���*p���>��l��$����<�t�Bt�iV~���g淿	�i\ *�"�/��ȕ]�2lN���9����s��[t�~�	�c(rA�H�m9mf/ؕS@�e����XOb!U����;{���/�%6xr�Q�E䀭�@�yΡI"��J�����\�y���Q�{;D�Uy�Ѱ��h�w�0�F+�������(W���9�g��0�o{����GDS����,�/N�R����q�(��B��G���D��$�D��:��j�s<���XT�k��К��\��YSr���:>�9���ml��V��֎���7T�Q'�����%�$yiwi ��g�1ϳ5A�#A"�Gt���:�.��9���P�)P�������e���v���$tF��$Jvjo�:�z�g+{�9K�#q�ڮ�h%�0{��4���M�K;�BV6��T�����5j��Dt�'�%�1��y y��E���looF*,XC�Tf.�}�Ŧ�9Gs���l��U��7��OOkfѨݾL3�3C}穜C�$s�*&�(�����k+�9F��-Ce��/�����p���j����zC\nUd&��<�������3`bX�@:J������&���:��w��ʜ��I���Ru��|�1e�?G-p��2��]ۖ�"�on<Ŧ�d�QC�
�4�S��bX��x؁|�� �|�̒>k�N��D�!jf�N��G�^��q�aY��R$�R�-��tf{PRW����������L1�����u��O�"_/�܊�q:XV@St
E�~I� |��4��(.�e^�Y������&�&O��l���~:�L��K/i;�/����Y�����=ɓ7g�#�įy��t--�kۓ.cg�XTU�1ˈv�gB�$|I�f�*��#�7�/M�,^�e����Mv`�V��z�yDf�����+c������������g8?�:�&�xʏ©�
���.�ߊŋjՑ#����OkE8�Kl�:/����YFtur�?���OjӁl�3x+^��IP�1$:6 �p�!�����r��S�VM��(ːG����]�kE �ݢ�d�<Y�������!3׊
n���[,�$�c�rߙ=9���F=A��������F����9!�*�g1;��i�[����+5�|j��L�[�f�W���:�n��a�mzwt��ܦ��|����T�(���/���\��;u[	�$�j
`Q;����O)�G���������W���/5����+��%�!�S�mD���&2ћ��\Q�sHXqt~��5�3>T�-a'�,3�x-��Q�W��=OF�-���`�owC���s2����4�_rֻ��5}n�Y\KTg�P�ms:6��P��jӣ�5�.~�G�~���A}�X�l�!���Q���m�xY�S]E�>�����g�|�R:�E�3���zU���u0yI쨮G�~�q�ag�;g<��G�T;= ����U��^��Vָ�u��n*���mSݸs �n�z��;-/��;N����#zާӂ|L�m��pQ+VP.�0���±֊�t/[SCT6��M�v�H��wL~T#��Y�(��s���20��&\%U�VJ�_љ��#e
��P��-XK]^̥���. �y��"�w�eҷ�Z��}t�b	��>J#cz�5n=��cO^J䃀7f�3N�P�Y�)������_��{UԒoTY�M�G?��3��%)��{(����G�y���	�H����a��-���J�7_�:��]ϼZ�5�W��g�!/\\�3q�.̐��nA&%4�F� �Q��d�t�/~�R6,�"ffr�WXX���_�N��lxޭ�g��(0����&��;&�h,t���v�])�w?�2dk�O��<:zw�~�B����1;�=F^�����Z"�>�냈�a8�I�n�D�ATM�p��
oPG!G�D�!R�f.%,�h�w ^��p6G��e	q >���QLRܨ@����X$��V����	�N�߅��`2%إ,|Mt�n$p��x��PoqB)CSw)˼]]�'�9Ty�:2m�m�E$m�+���vT%E��C�z�k�> �D]d�g��d�{p�M�K��Mv<�ۮC~P�،�oT�s`*!��l�+�1�U�`K��D�I�^�n��M��7;F��"ܿDv�ߘzQ)G��?'����� {hYZ2/��QB?�ϕI�P�{���	�"�-�,�H92~{�kL|�����Ӄg/l�H�t@7�T��B��>>*7_�9|C;���;�R=*
�Lܯ]�L�Y���@S��\)>/*���5T	)�ga�a��o�0c�J��;Gm1\�:�?[��ә�r:\kw+M��iR��_W{~zWY����yCcJ�^�!C%�-qt�kn󚻷��
��|%��� Dx`@����;ǕD���-T��E�P1�1I�YA������C��$E,�0�F8G�S)���]N��m�m�_8 ��)d)VN0�Np�j�C+�u�xBJ�T����%9`v��ڪ)��,�A$Ėv�1����c�t��@7Ҡ�'oP�4��;�p@z�I?4�Y���C��yP��P3�q��a4R�<{X�k��݄ 9N���'� �=��͞��
��"�e\9k�gE���Ƣ�@���
`�S}�	�Wx��|���-���+��x4�OE"��^�0*�Z�3'����*m:�@�4��%:qZHy7�d�2x�V��-i�����D)���g����AL� �tx�>lL-����R�Y������]�`�$.�p���ҁm�]�:��`1��mDːr�ھ�c�$��#��^j�lW1��F��)e���*S&�4q���୑ay�;��zƊ�4�3�tr��o%K�,��P�!o,EW�"w<)`��Ձ��y�Tg���>-��1�:
������-�>5�����{�aQ��N�	��o}F�RcKҮ7�D6~#y�Rx'�#���n��r�RM[��AX����+יs����\�ǁ�ļغ�M?�h����s�'�	�*�t��F�l(c��1����f��g�!nM'��8ǿz�����\Ӝ�eb+��������
2�]����ʁ��~��G�YC�bR��� h�k<
�>�VH[�-�����#��z�9�m^c��*3����wp�oC�V�����:�) W��eJWt�U����(ɪ�4�:~g,�u��A{ؘ�:�g?jdh�4��쭷2��}�UA!����3� ��<��V]����*^9Z��>'Y�#S�iȤF�:�G��+O x�1��w]�/��W-#��աۚ��K��W�l�����Ry	����>�D[k��Y?c����b��m���{�24r�K��yk�.�u�,y���#(�v[��A��9��6�n�/`����/���Ui�ә-����+@ؑ1r��fg�����ٕM���{��\�>_���Ye��[���q\�J��#6PZAa�'�v�{c��ʗp����w،=O��\̺ćEEa=�ք�F6�X!�_��y3�|1;�#�aW�Bo��/�o��F�I�8�N��7q�TH�s��,���V�w��i�[٪;�.G�;��|�"��n΢n$��]E�u�S�F"���ҍ�"�=�
��{e�8s̱�d�|�O��ߡ��3Nm��l�)���]��h׸�@����x䮸ې1�L_�0z�Ww�ܪ�bH^g�� #��QU�ʍ�����s�gf�w�����	1݁��{s�x��-�Ӄ���ֶZ��*zd�Zݠ�x�c|§We;w
�8��u����Y���e�;�$���Z���L�Z�7��E��6���?�x���9�!,_����MeD��Q`*�	�1���hl���f^ M䱙!"PM~t��^bs,J�-��ay��R�Q7���cO��e��ǰ|�` �?G�%�8�ft���sr� �͠u�����E^X��F�,��I���1��G�;=t�e_��X^�ސ/�x"G:X�]�yt8�����YD��q_A�P\��IM���[b3#s����<����Qܐ��D `��Yj���2�zA�b�3^Y�aL�!�i�0��w$��ٔ<M���蕼�ۂWP(���]8E�ﱎ�X$�뤘�*Ϊ���ϓb\���&�LD�:�8����&vg%.w ͬ득�0��m:��(�5Ţ���!�5�rN�9��Z����,cs����f_�u�T��Nٰ+��U�c�rU0�p�:�E���%g�jc��47G��)�RVK��l��i��
�M/.�OR��	������x�զ�TYJ[���_�AA�iD��ZU���cmN�4wl�C;ɵڌx�I+A��+y;8䋰̩͵Z�\���I$�#:����|�d6��V��U��v9j�AL���.Â���p�Y���$������N�s��`�	�org�2`:����F�n�gL/��I�43N$�I%�@!"�����I�Ho�6wԵcf�c�?�)6*V���Q/�ƾ�4�JVD�]��<�,H�ʍ�uv2�ɸ�	�/:I���8�"�;�	)��~7ە�B��uʗF�v����K_�Z��1�"l~)1����p���$�c3�I�ϒ�¦*5��7��ۿ�����cl+'x�1�\+��.�����I���>ߗ2�`��5,�"���.��H��ǅ�PfR�[����#�B��.۪�sq;(D����3��+kC&��ϊ�`���q�
d����C�9�ƕ��b_�=�׉������[?����f��*��zY�h�Ϟ�ޤ����J)+�TxaX��xGh�|���.��Gҝ�2�����$�����8ƛ�0�V^z��?�6YQq�B����a��-b�M(��A�=7�o�Z{(亞%�T�
�r�`����]����$�-=����@�,#?�b��j�4{AN�3�/=�:����n@dwp�������Q��p*�?�M`�嘓�
)Q(e�7]���N�X���c��[�*-VH:/dW;2�[j]_)qaE)�-7�e����p
w\��K��'3OA���a��Ae�/Hb��J�� ����N����wW4�s�������G'va)oH� ��k�0�żWǥ���E����_���N�(�-œ�f�dw�^�{9�J��gL4w��}�G[��-m����e�8Gf�i��|��nrHc2
�����i�/�}�@:*�M������&?��}�z��y�Yq@u��%a�]w�9���8 ��� ��4�8�E��.��Ħv���0��X�>X&M�c��%������,��\�U�Gi�(40�����Œrj�/���.B�m��jR���^����gb�Ӵeg�9框Tb��9�����8�h��4&���#!=�}2��TV�5�P��(7��(eL�:�V��Z��9N��Č�,���medi��{�*���t��&��v5ix�1*�ֳ�P�5C������Ƣ�z�"�>m��V�x`����_j��6�T��5�r��!�B3���щ�VM�Y���L$ͷR)�ʻ��g��C�<k9h�M��s��a�|���k�q=�ht��}L翔���~	�>�;�g��%J�|����+��$�'������K��3���v9�R�����o�
��FJC? ;N��#{�l�:��ª{_��9�uhȦX��D����F�S����]+�%�+��e�>�%P�p�d��.&���}���3������@c�7�Wc3E	{%�ƚl�_��2��MFP_W�7�p�0���ě��y���#���'ػ������ᗞ���Q(2�=�ڷ�ւH�6��y���j�+8��%�������鎩�1+���g��g��-1 ���?p��^7���q��qS�j�?4b�Gd����j	�|��?��w@�Nw�=Z�B�3@tbn�a	cry�Tbd����h��^�քA~*8���Ǥ���%�_�w@�H��$�u�����!ؑ��Q���̢dߕ#�ԴUך��̙��ig��)#=l�C�E	u��{1W�l�d�N��EK���";�XU���ڄ°�����dxӼk&�B��ڏ�(q�k��x�
Izc�CO�$�T��jl�(O�O�D��Bg��S�h�ʌ$zm�� ��i!/x�����A���!�;Y�e�����>��+��J�kɃkX�?�%<'
��%5�~F�+���v��թגaG�Dgw�2\Q� ��@ʽ@:! M��b@���a\�8�<��#b�m�]��ь�2�̵z� ?�:�T�o���!��	7u����+�Ѣ*�gʺ�}��#���/�Eat�����:_W�<�L�iF��o��b#�,�wV�Z �`�-���(�R�'3��.X8�^ߊ����E"J׊�G�����ѩ�?`�Q��!I1e�7�j+]q�>���.��@�a�$�NW"Z[��������q�O_�J��qq��睻�i_����?�6�ۙ2v�,�ؾb����/rݘ�X���������[���kgZ(�C��H�,��Ν�A�"���F�2<�9��D���@VȱQJ/��T�4��o��5�/QN@H�n�%=P�sφ�s���������C�Kb�>Z�m� ���iB�3o
٬� 'tD��-���v��\Ң`�#7cX\�rћ�P�6{/����1ݗ�p�8yW�r���c|�� �d^�;|Kj���;�`׿��1�e���8N���g9��h���.#����$���D4� ͵��v��F\ �B�)����%�~Ø'�w�ܚ��N��k�H�D^l��խ��������H��R��Z��GmBak����jC�ۦ�
a�{Tt3˻(7��c��;��<�����!��!��4~�_y��[����!�X��|A��|5���o��F�M�4�V�3�Y���0(��},y��f�I{�ɤ�v�бZ |:����ܴEk��l�oQ�Q����G�JuJ���Uw8�{�[����D�u�L��E�3Ŏh���3@	K	\���<��>��	f�u���O�O8{ފ�� ����S�B����3WA6#[�A)Z�W��:+ޫkI���v!Y Ն_3k��a�حa���+O�1x�1dB5�BQp���9����(��Ͳ��'���-u�b�U`�|�ҝ�`I�nB�v��c�8(-�DI���C~Zq`�۝�ӵ�S������)>�|�g���Gο�պ�a"d�+��T�ȟ;o��=S/Y��.Yf_��Hc��_Qft.����|��YT~�à0��yh}�}�6��>�����W3��Z�+�V]�4L-�i�u�T�Lq�����ȡmFy��nP���s�!X��'dP����r!��"D�)ؼF�qJ�úZR����C�[<��mb��W]��T&���P�j,:1\e��?����pz�O���'Yv�������A��;T��o��U�n�߼Ka.�>;΄���6x'H�*S~X9c�h�?YV+��ܦ��3���a�!��&4D�+��x��ź"	y����_sΑ���=����il�[�@�8ɍp�d��������կ<s)6��Ȗ6>�/�@�R��Ngi��Viǅn��YQ�	+�A'�c�m�P4�[��#���q�/��c�`Csk�d|�s�.-2Z��sw�"lC-a�by��x� �,�ݫ	*ء>��Nmvo��?��H��Z�l�U-@\좄�VR�2�(�����ˡ��������׺�`�`,�{8�O���,t{�0̈h�d�m�T�e��'S�c�N v���ĉ�ߛ�9��c�Ji���;��hW)g��,���}@�G�-k���M֘��]��WgN'x6DYB"RXס���*Pb�]of��nG@z�͎C�����\�JK�1R�'�$�.��
�	�_��LL�pi%;�5��p�d⏁��Jw�������b#n_�6
�C~�̯Wq����v�W�`���S��
*Ͽ��JS�u���77a �xھ*�#��.������E�)�6꿽��n��(�C���gV&ǜ�����=�о�D�����`7D�c5�l%Y��ϭ�UmMU�����B��G�b���1N�Xё��
����cPUW��"�Ӓ���X�?�������� ף́��
1D���$��~$z�]5�m�Z���i	I�OD?ɗ�E_��Q͟��P��X�1�muY�V�n=�]���y�B2ޫ�!�#̄�OΖ�8k
 �������{:�/L���#/@��(lT�UI$�`{WxNݵšQb�����Hz']4�~��/ [�،;/���j���:�`O�^*���M�4P]OC�|�8'H�k�����6`D����4�r�[�O�����S�T,�z�&k�@<�bږ<��Y�8�� _�Q��:42`�s��˪��;SM�k�O�D�}�F��	x����v���{�1�=}�������ɧ��$S~RA�#��jd���j*XlL{wx�jN���-����U7� x�YG\�+ے��K�:���B/�8}������O+�="��PG�� ����gʫqs��M�'h��n5 ��iZ��<y�W���$�-��Q+/ܻdK#f'C�Y�{)��r"�E���G�#rˣx�Q���v�{>J�NV�E4�V�dQĳ�r�[��S�%u�x�(ۻ%�5g���8U]9�����o9��cD�Ae�	,�j�|��E<�B%�M����r�{��T>��䒰e�A�
]�6���:�`���f�}E�|!�	��;,f8Q5�u��>��x�u��$�5�XV�lN�y��M��YQf#8HԵUf���[��p�jX>gQ��_�p�&��.
N��lYZ�u*��o���+�z^9��qѷ���1})3�o=��89�R~_��%���A���J��5��{Y�OD���b��^�s/���i��Lɔ.�3*�n[,��Z��?˩O�3:�G$����4�xx�O˿��uay�w��
�W����{���/��	b-��:�Q����"U7�2�
�ᅢ�I���M�<3M�Ɯ__y,s*i�>R��u�bw]��'�iF���j'y
�Z�Iۤ���C��2hrM����bԲa�G��kD�_�|�l�Z�q���#]�В�j���d���lL�$>����D�Y��#R���ȝ0b�M�ɼ�,��çj\�2������_�X�,�Q���!a1�J[]a��$������)���� �_w�G:�������)ﴯ��~&��33�'oݼS�v���s�P;�iɮ^q��7u��}W�M~�Z�X"�S��"�#�p�B�����
�ͩt2h!�u�	���pg�p���'�%�o\�p�����iwi�y)o&��PǇ���L��%�[:���n
Xr��~Ԧ�Ҙ`ph��%�����F�Ç���Q���M���T�����ݚ�@Ǵu3��eT%��Y��9fVv�py�����ᚭ<tV3:� ^x����~#��(��:*q����L[.��D��۳�m߲����� й2����7��{1��t���y��͔liW�Q�ͼVe9����8�A1�?ٻ��l�͉�(c~A�� s
�n���>�Jbx�KS�-3�ڔ�����X�P��Vf�s>�M<q�)�Im@���Q�L���t4�7!�Z�&���:�8�%Z%�L��%�xm.�^�O��(�$��_�c�8��[��9Z!6�]G9��]��V���68���Q�T@8���O[�n���eZb����5:�
:#����kdΓ�N|c�5�v
��,�ʜ�Ɵ�i]����:����9�A���:n�1��x'��e�����T��H8�2t��I�ˤ'����˞S)�D2k�XX�S8�v��:��Vh3��uV��Y
�Y������a?����b
�b�`n���ȁ6����!�{'l���=�]��Tc����C�-��Im����G�<�d�hK�H)%T��z%|k�U!-��C	9�����q)=�5tפ�8ȸ#���x�W����|H��"nC���D,�z��.�a��?�����4K(�B k^*w���sW��(��N��N��q�0�\"v=%aԡOU�ױ>�(���a��<~zK`�_ M�bs���J�V�wum����p�D�I�o	�����:EB�F��,��6�\�'\N2�/�B|l:r"�B�����A�lp;D��{������_���Ǯ�q��!��]����'�H�:��W�����e�"�����rF~'if�1XtY�h��y;�,�y�0�K��[0�Ѥ�t?e��z��c���ޯ|a"X6?�+B����k�յv/���j��ÉtM�(hv���!����K�:���!���H22���#�;�h|�U��G^.��ۻ�H�E�;������Qа	����ud_���#��N�D�g���x?v�)�������Z�J_q�q�q#��V�b��{���U��o��h|
_/Q��<��Ҹ�OB�[>"��]w��a�rd���!��I��R�n�J����. ho�^�K���_'��r�� C	��@v^�����x	�v��f��]<xM���p	�.��,WbTO�qŀH�z�8=(��A�ퟠ_��^|���ٻ���),Q���g��ɍ}���B�q>�N�b�Odh�c(�@�>�T�Ծ�i�	�x�bd��G)VW۩3�(0���Ljyoi�+���H��S�`:,��w���P��2.;�|��3�Jn�s�D��!�O�ӚQ����P�˻-���ȡ�^O���i��L�U@e�\�	�4��&��!ґ���45	u�er�}�7T����ɏ�d{�ތ���������=Nt���B~���Jƍ�I[����i-=�}���¨���W��[�U�@����/D�[b��υ�}�x�����s�r�gsEJ%=w�*�M!n��)\����u�P:L���]�0em�-ŏ/.C)^$��m�9�u�q��Dޱ�>�9�J��r�-�@ƺ�
�C����Ђ�y7n;���j͠�\�g��wQ`�&h&��q����(L�b�lX��8�w,%�_>�nڀ�$
��&�\�l��j8���������9��U=�2�ũ�j�4f$�̂65�4%dK	�YU�4�<W��W���CXUjq�;,t����?�6��ZxfAy�O�SӺ�ۯx�Kg�n{2<�	E=)'α�K�˔^����<�.Px�Z*��ݯ$v8~�KU	�	���Y�K���Yn	�2���V��P�$zʎ�?���e�;Sє��6x�z���<M��n�V���UX��:3�JI�=�Az�̗=���\��������sN�m7���Л��)�j׷��A7B�b� I�vs���������3R| �lR��KWoY���=��$fDW��~
]�h3���(Rʖ�g�d�[�4����,�eMC)o|4�:���O��`t�+�kz�e�N�o4���O.*�e4$p�}*-̻���P�jK�3*#�b^(fH��9ن
���ҽ� P�i@�%�-�����p�w��xj�W�����1|���nL��ե_�CiN6.��p�h
g������S�&�,�zY�q˘C�ٌǗ.޼���1�X*�Ku?H�yw�r��G{^DsЭ��q=��������Sd���Z3_Xui"%���R���1��,?���rۿ)2qpip��Һt��A�%;��<��m���
1
QJ�V�ô�p)��{�����ϕ���{a�BjUSM��u��8)Ñ��dH���f�d���^�n���@Ld%i��z{��V;�\�oX����U="����#�euk2��4�g���ǻs4�7�#q`�q"�d2p\��g�ٌ��39҄�.B+��-t��f'�dP�cQ�\�L��`�����j^�IJ��*�4d=��D��t��1R�'<6m�V%I�� � ?B�7���Od8��F���3�CO���+Id}�\���<��M��R��[bw�l�E�2�I덏�S1�J�Fs{��-/�]c�S~���|>��l-������$|���mW�%F(�f@�J��D��A5 f�{�&�I����<�J���7����`�<�����|��¦ί��z}7;>�ՑQ�c�����<
�2��q��l����W*�u����BҎ���J�.9�dD��#���Ó^8
Nf0�hD��[C�>r�Z��ҙ��ꊥ�T�/��L|����¶�a��J�$����lxĎ"'O��j?��3�a���[�?��Ĕ��]"�%�޽5�S+H�șC��>������,u�"�3ʼ7�ja41��1���Ε�u{�X<a��y	�����C	��v�Z�nW�����QK�mZ�2�{ Fc��ێo��������M���`�K�����H.��jL( �N6�J�ag2|���+bmc�q��H��c=��c?sk�ޞ�꼣�+�nѲ��,�L���/{�@Q-nì�Oc�ʖ�9��j �p3�LLb�z�^�z'�ܥ�/@k�
!~He���ļ�
e?�s~��N�^G63�D��SO�8'���(s�J��4K���^�	 s4�J0��x�z�yۦ'c4�9���R$6�IY����5����'>K��!�(�O��
̀R$���#���<�^��(=��� ���X��h_p;�#.�uhT:��V���D	�m'��4�h�3�0}�9�>a�Ϳ:l^�YqA�:���z2����p����Y(S&I����e�#��BQg�o��<£�C�!�G�N����K�^D@���@~߱_�\/s&I�cE����KaL5m�
�L�n��`m�m������?�i��{aGW�꼈�Zɒ:0h�9�Z�I�w:>�{����i���<��>VC�~d毒A�U�Qd�}�����>t/��_N�o�4c?"K .������8'y�pDM��Q�@��\sVm����Q0:Y;�t���٨�_`i���D�J;+�[&J��g�L�є�t�l4���YV?L�̪B�ll	���b1��RA�|��-D7{I�9��h5��k�4~s��5�T�d4R�@Jƞ��w1/.ܿ���bzV82����h�=�QA�(CH\l�2��@�8�~��4d�ů������)�u�,��oD��Y='�O	�7��������w��,s���@&��y��=�0!-)��]��C�Xil��M��8��7F<nX�4�uȏ��TPc��u�OAU}�{)0[=v�w�#8��?(���ٹ^Y�
�Էj�&�(�h]^��tyڢi�/S�Br{�3�x��$~Txw�0���7Y���>�!�n��q|$��]H�q|�A�#�(� �� ��)� �����n�7r{���N�a4�K����Ө���#
���aN!��^VK��x��=Y�vl�J�~P|44��.�Ƙ#��Q"kZx^p�7�L���� |FJ�@ =N�7�}w�/�����P_y�������7�$9�j=R,�Į�ݢ�=j^L�.�|�{�ybG�#.���y!��Y��gk���m�� [z�z�iťN���!��^���׺��� �2����;
���������V�����~�p�	z]0��m�:�)"h@M >��g��5������7<�:�}�vh��ӯ2�5I}�)2]�Za e*�e�K�sn��;�h���̢7L�3x9w�너�◺���<HV��)����p�p\'�܅)e��4Y� s��C��|����r�"UR��R'����/�M$�%����Q����D��j��Oяm�E��=^��ϕ��!���0�3��YB����}?�:	���E}I��4��*����u��*)���P����M������G�\��*�:�Μ�p 5S�zeځ�W��<�5D��+N�no�=�PG.%�З"\,�J��~��$�n�(��s���T��Pd�y�*_���RrA[�-�����#
C+���na'u��6��QÝT�;Wh}��?+�е${�����D"��8ſ��c�(���D�����W�(mM�������
�������DT2C,ۖ�v@�܅O�Kn�a|�(���p���72� ��cT�ᑅ0[�lR�^���z	���b��7em)��D2�A���.X��!ѹ.�,��TCn����t���R�b�>)¸:DVV��U�N�་�
WC{T�aC%���N�аuG!ʞ�4�sQ!����K�+�ТV'�������ξG=t�W���?0ԡ�w��R��X+�mV�ѵB;���z�'���ǃ�&�RĵL���7���B�GHr �y6mJ��ޚN$Ψ`��
�ƥbIz�8;��{���ˋ�E�^,A۷����N�x�j���� ��o��ŗrZNJ4���,?�I����I�5��:�GUdu��EoDF|�?��i�4Ձ�]#2�$���S��VZ� �d�bv������m������F�D���Tp��`���R<pީ(�.qt;9���~���J��jRBt���;����Bx�nrk����P	�.:�P΍	�����F��ThO��G���?�1��$���]�e��h��!,`��m���#OW{�N�H#�)o������)��h�%Vt��cis�y�Ê��ֳ�>Ӑ�=�5������f�t�Y;�5�91�Z�wO��+tF��Cc��_	�	��ԕ�V�u�] \��Т�N����:�ħ%�q�w��"�q�d�e6V����:,�15;���b���Q��~�����^����q��с{���T�C�v���fRƦePD-�\�O�3��9~��~w���z��G��8�i��űd��0�	��僗�Ջj�L�*��<%�<$�6o�M�t��Ar��b�NB��2�� ��D�ݽ�[��8E�z�W���3��Z�ߋ��D�P3|k���WBR�\���C��e����>�z������ ��צ�Q��1�:�s�*y�B�M�p�F����	"f'�*��=9�p��k�ża��S�5�Z�pJ�[j���U�����Ns9Z|�,p.�sE���׺��IߌxuA]/���a]�e}z`����]��ht�A�Er!%z\��Հ�h�����j�\+,~r�QWsO��ۙA}�:�<	ҳj5+N>؇��3�F�}r�RƑ5<�"J���ǾӔ$-ēN�� &�F�"�=�K��}�t��š��݂�tr;���ZF8K?�xU|�R�J�?mPzŹO`q�5E3)�)�&�I��3?��X_2X��+�˵���9�r^�T�1|���ݾ	Pz��j�4Wd�#�vV#���Vz9j4Ϧ,&����O��wdΈ��ɤg\~2r��ƪ{bƈ��`�M 3C��X�xVw��W��������b9J��'�y�-%�+�,Ѿ��|�h���CH){����h�B�}�&��)�~����(�Ȱ�ڔ��R�!�-{A��ǿ� ����})�ҵ���%� P�(F{o�����~�h�;k(S MB�O����8�SN���+?-8.�ѶW\����LUQ��.�2`53;�)&�M�����8>$��15~��d:�u����1@T�H<�����p) ��i�QU�1�$�v�7�fi��jY���Dn��,XI�������:���c���u%{���(���xW�;����QV|S��'�v�B�sÕM\���2��h�7�kT���:��Q�I
���#T��Jζ��|������#P�QW�xd{��xޟb2b��U���뷔�(��V�*H=��S�C�p�*4���gY%�+�FA���\H�T���a���?�����B�ڰ�	�/���`{H&a��8�]��i�&�()qu
�����S�Ee�ӓ �G˟h�߳�m2�ф�U:^�&T���P)�<�O�e$�a?/��M03�O��� ?GzIO	�,�o����3�����[�ͪ.jY���OԶ�0�J����zS=h�`	���$%�5z+�3�
��O�jtx |�wWѩ�' �z}��t�!h��m�Q�fIُ%��5lZ��m;�^���x����P(x�U�r(Cϡx��Ǵ٬�X2��<�p����]/�f`¦�5�v����wY�3s�.ޖ�:��p-�qt�s�.q5����w��rm�<�ZB���G���Gͱ�$X9�~����P��b�!�x���)z�|�jv�E쨆Q��O�T{����(���Nd��S�˟�t�h�Rԫ8=�A0t�� �n5N��@�K�j�z���ИD���k�G��&f��D�����q�'�Fl��e�.�,I�t�HJ$�*u������2QW��=�+�D.�e��'v�G�/�C����=�3q�P&4c�O7(i���w�k@� �^��,�C�}u7n"�Em�L��N}zVH+�'	�J�cM:9e�X޾'����3�2���;%�l(gb�/�oh��m���p#������!��H���6w�P�݆}�9aS��}k���+P�>�9��1�XQ?Dw��yǟ7"�C�XLzb=�=(���N�7��/�0�0����9�N������
���$�U���#�f������w��s��)�����#��p���].)-̼B}%��a����g�P�6��G[{i\-�hu�P�?wq�x�Z^�NX����͉
H��0J~ss�Y��Ǆ_'�9Ѽi�gf	�=�Y���DKd��e�75�I�rD���澌��Nĭ���8����bG��i���U��7c	TiL�d���#Tx��(L�9ZD����*;ޞ�!�qB���1N�v\;
��S��W��@0÷GJ��Q�������Od����mJ�5��VR�-u��z�C���,Ӧ���y(M�p�����wN}��¼��cmW�����Jبe��N*��i�l�;��y�+J����a��X�t>�RcTd-��'+s��)��.(sC���i:�5���d��G���I�7�)�*��A�%��CՒo,���)�bd�N/=3_�6��� ��@Y�>���^(5�z�C`:��SD� �Zi�jljD��'Cp���8��"�����1���{RFD��[��a�c+���p��).��oY���,��`�7j����uf�ӒopO9�[w����8.^�B��m����-��/v��:7�	
��ɴ�(�L[�Z����ׇ�Cn��nG�� BE�ksAg-�̢w�w�!�c�E���y䃔m_/�V�|������*7D��p����D}����":v3���3�}:��� ��;B���f>
}�˥�k��)6qi��fؾ-�.xذ���_ʸ��L���`^�<��z��3_1�h�ܦ����-1���JC��!U��� ���§S�-���|3ڕS�Udئ�AV�Oār�+��Ǉ�]�~�Y��da���PSm���s���*8�j�^��HZO}�e��2�,�gdG�-���0�n�U�%YDg �$� #9���[I�/��v�_5H���	���Ûʨa�ct͞�?�3oB��c�]�'ס#Yf8�3U,~Oqy��$��?��w�}�
l�%��z\Z���,�As�Y��k���@����r����l��2G���Cu�d�97��b#��{����*� ��-�3ȴ]�@M�}��y�辙���; ́������eeq��hu~Q� ��
I�:b��@�h�:�vv5��e^�,2�b������M4�m���:��>��e�'�R�0.��+��;� R0z;ky"�2%5�s��"/-��n�L�ͷ����������O���  �N���|W��T �D}�iO�Զ޻uH�[��P���z�"*��p�jhi����-��P%���F2����E[��u�S��h=��G������2��۠5�Ĉ��dWEd��P'��?{]}���+֡�Nš ��FT�=]l492��Пx�~J��PZn�����]����8�L��U*ޤ�]q�:թ�l�r?�@J�y�?N�7��X`�KvX���7��)!��։��P����R���j��{�uC�h�K��D<�rk��}؛�Q�b��j�Ҭe��/,�t)dΥ��,&�XA�A�ϧ�9�5���t���K��K��)Q"�&+����F���&B����0�wȖ���zx�"k�u���!���q"BR� �?�V�e��~�T��������^��b�b/���|�e� B�Y���Bj�f��J�`_�%���|)7����+����F����)B[m-ʾx$ߒ2yHY�##����5ɮ�Q�������ٸ ���
S�D�L7m�ҝdr�6K���[-�A�ͼ�x�,��J �����Zm��c�M�=O�#Dx��̝MVʔr�3#f&�1n�Hެ��{�/�Ҕ9kܘ�T&����ӡ�܍Ŏ���"�ҟ�'�Dg�o�� a�n9Z�j~u1-��
sh	h��y�;�%�5Dl�[^�7)3�� <�nLt�`��_�f����YJʕ�n��ι���1m�۵�v���S����w.w��v.&y)/hh�-9��4D�h�����$Yi�p�ѫ��v�`���q��[��8f�1�І,�q���ì2�MeP�&����x[�f믋O��$���p��u|�מ1Ŏ?.Dw��3?-H��~1Zf�9Y�#���' �r©�7м�����m�ٻJ��ll�Q��(��%]ulV����}i�:�u��$�Σ��8քe��"^����_Q:1�C
o��{2�gη[Rv<���d���)����2�~�L��� ���*�׻����(�T&��dݗ�V�D/8$ť��+���>�wǎE��Og��oN�x"2B�H8�7�zx��d$j�e������!�_ý��u-�!k.\,���Ɉ�ą*E��{��ui;�ܒו~[��
��,�\���}\��|u]���
ʘ��,�M�!���"��Z���b7����Y�}wƈ9DQ+8�Ӎ&�܇Do$��+��O}B-���`��ܽR�@�u�u����{����Z3��A��Sgy��W��e�6~O=,�~���Y��k���w�ܖ�R�lR�r-�"j����"���K�A��-��O%-~xC�{�-�X'����\Y�Q�~޺�E|0��SwHU�t9|uej�|
�{�׹ �?��e"V���'�z"Hc�jY��f#�O9&TD���
~E�H�j@J� )s���T�k��}�u9քXo寋}���D
>��h�.��/�w(]����>�L\��$�fPJ����ӎ(+�x��؀1����s��?KE�a�3�#n�n��ǜ�&��4��Vm��y�Q�y$'O�\��⏸��Of��ŐI2`/2!sz�&��
��}�+���:��?�z6	[��e��n��du���<b,��iu�ٽp������W��<�ѭ(���l�X����P;����O3�?�"V;$����Fa\�+?*z����+T�;����erf�e�М�������T;*�h<
��P�FÜ-�HL)Ҽ0M����L�.�z��s:Xҝj��dPQ��B�7�ůh�2=�f���I(Jy��
�z=-��E��x6���5/$����n���=����u����v�>����3t"�I�=�$����SQ?�u�i+1r�Y][�.AT5׹vN��Y���Ɔ`^����;��y��� ���u�4X�7P�.�Y��N�ķ6�q�y�%麓U���'$Ʃ�S-k�G�y(gY���$ ���V�J�:�Y�Q�v&�����9x@@���a_mP�Z0X"�y'���9R�Z���j��y<��qx �c��l��oC�Yq�&�)��؟���uX��t����3S����z�[6��lq%��8�uM��>����5�`��$xIΟ[�{h{���P���5��E�\�$2�{�%%������$r���ӏ0�G5]��W���r]aw8��M��ʨ\��}��n��� �U�G8	���j���wp��U����~o�p�>�"0�c� i���(����9���\�V{ϴT������.x 2��P����ݏ��5!_�{y�}l�ףcl�ϊ�a�F$�������#�Ai�;�(���ѝwҬ���}'��쵋��:�˓``6�nP��ց�9#��C�m�e{^�"�گྚw�Xe�?B�����C_�$n{�}��NFt0�	u\����+�&pw�15/�.�G qx�|H?08�5&��"9�wq����@�]R�i�w�fV��D�5�' �s�N�q���kU�n9ΟkZ��!=j {S���������;l�����c���]��,pO��4-�p��3�,�7��赛xd|���?�h旛݄#��]=2���=�U:�[	=X;B+�=�����O�A8��W��gz xw�k�����23��q� �� UZ�ݡ���������UFj�걔��0؁�V��Oh����[����`I��:��{ɐ��HQ���i����@���;��5����)c�	C��}�4��#T���]�E���6���#y%@ڞ�wtX�0ը�!���?Tp�췭6�D�lb6b�u#�a~�-=k��X�y�b��N"ěp>:.}p��fly�;���'
�ğ��ۂ���G����qJV@&v���

�2��ڜ[�'gDYa��0���WO��Yub90b��a���%gz����h�V�=G���k8{��!���~oW4!1n۵t�j��C~�XCdD��B�<����
���y��ڥ��h����ZK�z�|
�<+�� �'YE��r�#�c���o7���ɮ�Geر]�h1��Qb��s �B7�6Ƿ��9��󌜏�����)^����~�"���mG���t����T����}�� �<=e��S�Ö����>���>��Q{��@�8Ϣx/c�b� �6T���b��؞�2��5�&��@��rNd��;0 =q���|$s��hB�ڵc+�=����
]�H�t��X�F����RDm�f͏lå�ܓ��8��5�(XY��)R:�=f�[Ql|Ff�;H"�jr�� h�wO���r_՛\���ۆ��ɻ�F�
Lf�,����`>t�O@���Puk�
������?U(�V���9��K���"��q&�^o�X�Z��$~�M��A��Z����d�/G`�~�"���8$r��:\bE�B�7>L��_�E�$d��_怅�'���('�X�r��w��0K��s\ ���+y�����(v���aק�i�J�t��;�(���X��I<{��5�@�	�L�ߒ�)��E�R�@p����R1��������D3����j��P�?;�-��V�"e��S`'2G�U>j$���������1�(�ph����M%�_PŶ�^�b׀[�}� �o�����mS��V�Xh0}��%�<�����Ŀ ;[�o7_p��cf�2gS�7��r�4pVg���{��Wj���N���V�ÒDu@Xg�y�.��B��,2,?Bȹr����e�$,��C�xG4�L���T��u�s~2��.3E��3R�9j
v�Ə�xf���uJ�jV-���FF	��?t��#��-�x+���:���	���黍�p��,���"����&�7	J��q�����؎)�����趤1��MN���PhnJ|�n�B�؛��y��$bJ��J�	�AfA��};�d]� 7ri��fz�	�XV�w��4� �2���s��������b��_����/�Ji�w�FND�ւ���cq<�%�_�|-4�,�x��]�%��5�K� u�zIp�U�c�{��HV�yqt~"�d����v��[E�/�"H�:5s�g���B�7��wgR�w�-ѱ�0�E+�����UD�7�X��v\`4
.G��GR��I[�,,#���X�,^h]�̸'�}m�P��PQ��蕺?�~�R�@���Y�!��1�'�����4�y��@@���Jͥ�<s�e%Hjw��pL�?*�TM�D~��QdO����]��2jR�1��.�w
�����ap\~�& ��c��D�t�8s�=&����Ri��b;��ޗq��UKa���xX��ʧ�f�����y9�?�
H�V��A��;���>��q�6d'I�\rD�F�6˭|�_�u���q�q�+ &��6WW^\����<�5]C��zɦk�F������=sH�{7!@I��#��0��wg�YߧY"�מ忈~x�<'�U�-����>-k<�ƃ��}��r�C�A��B���)`��EF*��@M��tX�E~7h���{#.�c�8uA~���Uws0����Z������JUV���Kf����8D�5�=����'�؍��3L�F�֜�f����5^�Cf�|���G�r��8JV���ט
LѦ�U)���(�����9O�f�5��v>J5Zy�<���I��{�]S����s3�\D#i[}���܁�oR Dv�q��5�u����]quA�m�07-2��H+)��%�¼�}n��g�m�࿮�����/��v��L��MZ�btT$}����w���A�|��&������m+��ޢT�`����=|��R�xԮ˘�x/͚<M}�[����6[�f#����dq��.!��_���^�Se7�Y9� �ҽ㉍ZsT�wu�z����.���k�9*��:�����<C�Ҹȳ�Y۬t/�<��%���ū��pE��J��[�=ȒE.H���h�+����I<p�"�v�p����L4��賈RTϕ�?Ӓ��oY��0:p�\����\���56���Fkl��ٚ`"�C53B�p���.��`J� �����vKф�e���r�����-g]k��q-�myk�9��4�\�f5ci��UnE�xw�CFhV�m��h��n�=�庝�v œ99e��0&ϲ�U�I�Ν'��d4Kq$G\V��YZ�2��@ũ�K�I�0�}a�N�NK�ulv��S��Bڥ����J���\��X��*�"���.�10 �x��⊇h� ;}®Q�H�a݃d��؈H�������aQ>���f�`���4i�����ɸ�����~�U�@��l6B�K���TG'�����#T�8\T�Z���br�KC�U��3D/��a5��H^��a��R�	�Z)�"������.�����R	��((�5[��\{8��%��;78��_�0%�!~��]�x���˷�[?,��yMS��jۂ��b!-E�+Dq�:6x\m��*��o}CK���O�p,�BK~E�?�(����r�J���T��MB�.K\���P''�6�{����Ցfy�����v]\ٓ�����fB��Ϛ��;�|i�j�����`X!��6���͐�G�h���s��B�I���O���_���&(^��L���Y�N��v"��m��o�f�h3r� �v���?NNt��)|~�&��&��BDH���������S°id]�wj�by
�y"(��'H�C�Z�v�IMFXj���L������B�_�A��ŝ���A!����������cp����l$��R�qy)D�JՈ�x��5�0l?BےBQ@��-@��i�L��{z���I���w��8<��jկ�d�x���]�ӧ
h&�m����Ҿ�F@^2���C�9����Z�v��a�D����B�tg/��ڟ�m�!��OQ���l�q|�""�hz�6���-�Y*��k0�	�q�%RܠP�A.��aɃ�ui!��v,��F���N@�߱�4���}�|@�B�sY�ZS�m��]$�E�u���0���J>r� ��k�����hi��R��ֺ�W7[�Ik������N^n?w	�S�o;��nY�ν��s����{����D[ga>�9�v��jw�v�n�9��j�L�%n�5�����a�@/���y������"�o0�M��7��`�P?��٥:84QAAx�Y7�^�Q�;L��7�.FsQXJ�P]6��`x۠N�Fsp<�!8��<�b����D������Q)XOS��N��Nu`P��h���ȑ��!S���Nʑ��m�4ǋt<!#)>��j��`��]wj��~ni�jѺ�)F�lz3`�	i��ϟ��tT]�_/eC�P��0��-1���Ӯ2�B�>�9v�3�C
�#uX�7YI`�/��@3)Gh�v��J�`mf ����G�SЦ���=���)>4��Ыl�ٗ�TPv������%��!��ӊ �ׁ��xں��d���� K�b����[��M�Jȁ�e�jF��%iE� '�r�Ҧ?�%]$����!�c�S?����N7��BiE�IsN�"�u��P�V�aXx���jcj>���Tᕿ�ӓK6��/���(�Ѐ(�1�٢������`���?P�7!�۴J�W���#Ӿ�2�!i *-��]��e���K˹#����3g���0�)��M,&��Jly����bqy��<e~���'�+��x1e�^�H���Bq�/L>(¡��9��懬�&~��{c���m�:_jsT�՘����)%�U�J�d�&��c�{d���S	��>J�X<g�o��n�tS��)�\r�L�����ͬ7L��t�����e��/�[�ɳ�Ҵ�Ֆ�Rsv��p�R?�oE�k�&v�*�$��;�� �����I)w)b�q��"�v"m}�FW�S�d-� O�䙖B�Ф�]ډ����ڻ�,X:�58�TT�Br �1��s+�h�w�O�Kڱ��+��T��<`�7��^d��?wq�w|���v�����@!���J~�5��г��;���� ������t'S��H�|�v��'�FVe���:1l�)$H����S�b�O=�f��vO��z���L�
����M@��{*��vj�g�o�:c�
�)S��)���¥��tH�-��Z �Y�s#O&��Ƞl�:i�![a�&֡K��0"^��6V��1!��-��Aj���|�Z򲵫s0~���F�E�s?%����	T��E|`�'5uCL㩜��`�p!��p��J�/2�7]z��v2���P^>{��i�r�AT�K3��kV��bӪc��2��r<�N���֪��ee�9C�5� �D2������f�w�B^�B�G��w	{�	�i��]q��Q ֠q�޾��&ku�Կ�tI�G2�w;����"�ߺ$��&##��/� /=+�	w�X/"�2֌#'�>�;�Ţ�8�x����x�S;�Ɋ k����5{�b����,6hcֺ:��UzG(�P��Qp�l1<��1/,6g��T�l׎��xOp�n?��,�e+"<�Qj\P�d������E I�Z	F�?Hs���Ԛ�+���`P�U3$H�s��Cp�n�W�d����ubكhW{�T����P�.��u%����hJ?�����A�?S�É�|����ꏠUcr�A���G�ӡ��[���r�v�����Y�_Y�R$Q�|�CQ��t����`�y�w�\�=�Fc��ȴR���!��&���ߟ�*�@T��o4��``վ���ѓ�;�sF<k� sm"4����\��9`S\}e��Z	=Q�t��V5�L��a7pʽͶ֙܌RnP\����?�6�)��{ɝ����z��1;Te���m��;z�������'�y�F�my�U�O�az�)����"Ă�Aϻ�i�'�h{�wx-�1�mBd�	
�n�!p�����ߧ��݃������>�>i��;F*;��hښ�����7PF\Lq�a:���G~�|K`�����ũ��]�,� $6�4��e5ǳBX����w�'Ć1m�-�����c�=��d��?&yU�D7`̞jX(\�L ߽S�F4a$�#�Y)R����--�5�c[<�'���r����[ Hsj~-~��hJ���EB�c�>�۵�
C냜�"���$�+J�J���ݱ�_��Z�3�F�-Z��S6�8ٰ�Lf.5�WlbF�ɵ�{��Yh�'� L[���I�%��~��9j�;�-p�j�J��_�Z�]�p �S9"�0�3���PC�#o��Ѿo�e"ڣ�`�g�ly�p�f̨䇫�l�r��1��Ed�M1�~)Q�VJ	U���	8R��wO�l+�	�t�ѬtF�5��4���_������䎾G+E<�xW$�&���b�Md6�g��+Ku���e���Ga���+x����E��5"���>H�Ɉ�+jHٿ�Z��o��0���2����_���[��\�7f�n��ɕ���]YO�n����G�ӣ��	��ƛ؜�7�]�<�cM曞�0i�esh��F�C�V�٠�",�l��`Dͼ�KR�Y�Q>�kf-oKl��S��5Axq�EX�ø!�)2
�Z++����B̥@�y�q���ivhU�����$��L(N?= ���r����c�(�����3u���}7�:H���@������%�K$�<lZh��-eP��(�`V�����?j��N��	fE*]&���/'�.N,f"���^�gb�/���eF�;}]�%���ì3X
ˡ"�^���l��kr��5lF�8ߤ��n���O-�X
`T��nɝ��bQ6њp�K�_�B2>QD֌�ܻC�,����}<�����m���^�tp�����*�8抯�$h�8`��GH����6�CR���S�@�O`TU�H��uPMd�{�ҭIo��/yz�ߡ��J�|GwF8y���&���(�r��h�� ��"��7�N����%��x=�S'�$ty���j�Hb�ZC��T^;�A]e��J����ڰ=�J���	hnO� `�:Fƽ�?�����B���QM��#�݌D�[��1�fC��.�����]�3����&�b�~4W{@�f�����cײRDC�Ŧ�vMI��7��'� �5~eh�>f�a�H����=�����0�j|�<��]���Hz���|�C���'D��0Ȥ���]�ÊUaPG,��������"�0�w�q��:T�m~bM6q����2oE�q^�"�r6��"�b~��NB	9���&@��+d	;9�Y��3���I�Gk�|��ƄQ��<��F�B�y8���L�GglT�*�2&O�t*Z�o�r���º�){��1��vɁ�ϡJ����,Z!�fG�Q:j�sg���f;s�G4v&�����I���VM��UnE�:7��5����؛�e|7�F8��ymGA;�wn�xK�_aw����ʶ8!��8��?����	r�C�����f�S%Ќ?�Hw�s�/_2���>a5���lz$�$J�B��U�c� �؆��@0�p�`Q,H8,[M�����эa�ŇBĳ/ƪ]ѕV;�Qk��	�h$K�#iM�e��se�uq9p��뢽ƾ)U����f�d����Q�S�S�����F�^ x36a�UР��B`4"���[����V�`1��`F
����k�㍺A�<�����Y����T�z�o	�mN�H��Y�w�X��9䓕�!�7��Ҧ�z})^Ay6�� !LG�U�rd����2߇N��`O%|�:�����Y���dՆ�zx��>�-^l-�8�W��[4o��Б�> X岁5�n}#BN��y�1��%t~��FG�T�JTy��Mi��5D�~w�?�T%�H�&�3.U塏��f��42y�2X�1�V�~#SP�,�j��K��ȇ�\�G�R.)ّ|�y0��Q�!����ڶa�z*��z�7;��f�=���h2o�[��&��4�Ώ��[�o��kRY�@��J��Q������w�c���WP��oCV���mJm�aj�'���D����b��8lf�!Q��J��g�� �Z�Uq@��}z�>��les+S��cʍ�v�| d��[-^A�5�����{.��F�w!4�(���YUS�H"���V���c!T �,��5�4��N��ڢ�#ݞC����ա��$�X_�p�!-t���ߧ
X6��s��>�U��`%|�c�[��M�t�v-�<n�Y������)��<�Se���Q?�=�.�T{s��Aڨ���W_���s�R���p��D�I8���]��ĉ��~��^k	Q���H��J=N�B����Q/�ߎ�	���ۊDC������oثX�	\���K��l�t��6 lゟ��a�K�͜E���WFP�C,Ƽ�4j,�� ~ ;C��C�����߶�G";��[����2��.rR;f{�վ�"1�ce7l�K����X0i�v�H�O�6�r�uY���i���c�;N�8��"!Q˨��0=s��Z���w�X�������LN/�-�n�28{��z?(w�>|����Sŕ�M�� K�J�~�r�;�?�S�#� �v��ސl�d�s���Y{A k���E-�}�
_~ tw]��㑅�<t'߿�m ��nlO����Mi�����-{0�.�	�Sd-��Do�/��W��h�|���`�K�T2����q�䊼�>�����j&��9ҵ`i��rh�}���d�n��4`9�S,<���;�nC��M{��9ATz����z� E;gh��f�/T��=գ"������uG�cv)�6��2�Ō��V���j7 ��;Lͥf��>��g��G���F���U7H�Ù����
pM\u�Lܿ4��W�l���O�B֑�3��R��D���Z�@TV�f�X
�s ɾ$��b�ZF�z@��y�shX�odVzM��#LN���k�����0_���˰��b)T����s������,$l(�/�* ��:NQ�"��=/��.��#�؁��Uy�b�c���I{��*-�q��ģ#��h0�ExUk��;��jA0���)m�W�2�@"����ϰ[���v����\�_�!N�I���C���/�5E�$	���NA�f����=�m�F�������fLn�K��;+�USmP�bJ�p��c|+�?�y�K
�x�Dr��8[��)Yp�n���_Dٹ'(�N���a􌪖Vd�c�)����<��5�d�����k��uD�w�Fi��$�o�\d�
��ȱ��.-�o��3_�� mhL	��鄿�OӜ�%��dб�;�^|u&$j��i������#�� m_�RTOv��nZQ�h-����	�`�b����ƈ�����ذs8;��������:��J���/|.;��Nd���ׯ�6m�8�iuM��jrqe�}��N_��Ju�Jn��6����uB�a�UPA]p��i��w�y�T�($p!��	.ŵUmRT��-󵖥sj�	W�T Gu&�������k3���3d-���ю��앬��Z�ȇ���(g���3����&D�#	�i8{�%�C�׃H�p�"�M=S��1����
�cw>�|�Gi[Ĥ- r'K�־F�!S��/���x��H@���!_9����c�+�a�e{M����x5:�C�6~����'P�|�a%�K��G�4������[����U(F3�J,W/{Ž$+�|ڞ�{�.O�  \[;NXCz�r/���V�g%jQcc������J�:���nE�tm�%R̼�'��\�5pL2���-'��H���q��ֆ��)9�tq��7=<�U�a䯇Gټ�#��7co~gv(xylB7kAfNy�MC�_��4DV��1���i{�$���bvR��O�1�qBq��C�些�[���{�Q���%x����F(%�`�������<}��H`��77���G����_a��(�$K1�zn8g�m\��)��dWv��k��e�F�5����O�R[�x\�@;R�t�,~(��݃���xM}�]՘_>?�Ey�;���VY%l�K�I�d�hL���h�5"�.��H�Ϻ��R�<o�5�z���M�˴Y�@�-K�����É�)�+�]���pL��4E˽9 �\��<�^<� �x
���r������cdb��	��U~��U^?v�#=sH�B���f��i�ُ�_��9~�0�ۺg��� 2�0OpN7b��0և|�:�>1��6(3
%>��0�Ly�$��;
=��7��cc1o���C�C��L˶�vA=ƦZDP[�Ӝ�(hPfY&A�֤�Q/U�4s �^��6J��� ԛc�#��b�Z�$P3^��i�5�P�E�Ʈ��d�jY��f�%�����L��@��I��>�A�%%Pb��X	fd�*��'fL\!�Y��LH�9��5b���oU���F|�̿�FS��_ʛ�s���5[�)��V�!<��O0ӻ`M�^�?^>#�z��(����ޤ�6w&�B�VǮG��*;�j��H���:��/�����t�z�L"��f͆TIظl�9rw�3�f�	L��N��`q]J��tW�Tq�~<��5�"tE�#sN�����i�������`�y4%¶������.E�܍Z�H�@��Y�d��� %��g�UN85�8Xx.y�[�kהT'R��r�����nY�`���!H|ro�B��PpDF�;�2c\y��t��C��T�Ĭ�)A�+����M��{�c���&�{��d'8[��k�� ^���M�(�pQ�#�U�U��1�걈�v�2�(��,�j��9���� �z-]L���Z�$'ھ��%���a�^���ك�>d`W���Ͻo9���,�d^e����";<γ�~L؎RW3"�
��`��Cةj�J_]�bi!���n2��!��Z����(x0�&���^cōNGgL>j�J��B���H���.O��gwUs�N9-�#� ����o�PH�0y_4`�ȗ߯����r���a��ݝ�]�X�ݠZA-�{�{k��a�G�X�/�k)r���n5��i���YS���(��,�����K���@8���4x!�Ϧi4A�c!�k[>�����zF�5�f�M���$��D�7U�!�0r��sCXI���i����;��
�'8y[�qU��s:4p��ڰ����S�
� ���gnY'����#tW�.oE����vxR�v�Oڵ�"Z�QM�~в0�8elӡ��-�Ѫ��u۞�#�Of��O��[��{32�⒄I�����it���7��{V�zÑ#��z�r��#=�v,��
�'���dڊYX� �Qh�'��
x�s�$a��.繫��m����8n�϶�I�	�^��M�!��L���G�[��(c�3��<��̷�}�n���a(G�������2�a[L$�~�S%�;H�j�(��(O��2sC֎B�0�H1�]��S�`zį��F���n�6�x12i{���RVa��6�����	C�7�E��4C��h�����,UY�,����a��O~	e	l�n���3������Aol}���ߑ��#�����hs]�Z���#Vj�Q�h��Bds��ڢ:��"���[=G�_w��_З���gt$!u�WBj��:kMܰc�1ID����3�Pvǎ���f�>YΓ�=m��z[TJ]�=���UGf+H�0����k�Ȳ��1-#@�(�b�j%G�bsq3��~��3O;�
�F͡�XH�ގuiZ=\Kr��8+g{�68O[hp��e%wa�15N8�b0/U�ۄ^$r�xM�s�}� N�,]��=���SzI ��gǿ!�[�a����26y��G�
M|:~�@U�������ػ�>�ۣk�E�����px�e$YcPVt;��V|ٝ�JY3:��.Y�����z9�j�v;c��TS4��Ƒƌ��@7���5�Q��lA���5_�����t���G
8��o5�9��!�Ԇ��T8�2^C��%�U2'�q�Z���N�D~�����]S�sE�iՊ��A���V:Pԟ%�����J�sTq�Ӓ��g�U��m�H��UQ���˓?<���Tm�&��pߪ�'H�5�p��ڇz����@z� �I&t?�_%1�s3[nF����Ȧ0f�hi^,����ņ�L�ƃyEk:C�C{������֘�ܷi�CTm�����Q5����V��w�����|�a3�oBi���^Y5B�H����/�����5��*�crYn�s<E�L�F�~�\RP�KsT�������{������s󲨽��4�c=���_��R�������z@���A����רB�~�y�Ba�"w`��I$��<!�w���-��b�}��{ɬ7)��A㨧���K6�u�^�n>n{�@a��
�+�(�%��S���3����,�FDt3��>1����3,�8^ΘrEċě�X���B�A��\nH���*YwcU�K���]$�4,4�~y�mp�:��2ڂI`������Z����͒Ez��{ʇ���1��!�2��)w*���~'���O������~��K� �f�^�F����g/֚���L�!A�܈��4X����rf�������\V3s�y�s����H����C�Ĵ�8�ok;�$��'ړ.�ӰK��-z���O�r�;�.urm�s�ٓ���4��dTW+j�jQ�Ğ��������#�nM���/�5sΌ��ӊc�K Ft�G
qN5���P���P�&�li�]�g�@p��v�є���K�v�Y1� A,iJ:*��GA��}�Z�,Z���=C���a�^��=R�I��hw��3M(Gm�R�*��57;�	m8>��Z.�����@�� ��WEl֧g��� �~~
`S`��(^f(�F�AB(�������dF C���6����l9P	��[���Ϊ_|vN~d0����"�D2�o�]|u��y��$�ϣҾ:b6��ں�_`A`��e��K`�jӽO}P�
�b;���#���R��UAT��73�Yі�����/�nuEJ��9|�_QS;S#᭠�Dӫ�qto��D&G����r���7�0!�%kŵOnĽ�m��҆+��wЀ��l�:�������V���2����3�x<��A��dنk�<Š0g�~E��]׎�3�ښ��o�J��>��ѯ)x���8�s�o�V�+[[�b���w$L� G��T�v�f�]E���M�%�2@��H�0�ڠ0���-<�5��� ���k^ $���RnԺIλ���<֠&�h�!f�H��7��A���#�#h{=)T�K�]y���qL��xe�\��vR��"'���nvZi��6A�A�P����V�␼?���5���x���#��S4�,	�$����/�F�����_ޘ@�S�s�	^� ];��A�Z^�=Ю7۷�ap5���D����Q53�����㊶Ѕ�r���3�s��,L�x���zܨ�Z�kw�I���h�IZX��o\u���+���jUP~�(,�$"����ǒ �~������u�ӎ<8��������}��޼�Sy�5�F�~�d+�Xm!�������[Mӈ��Q�r�ѐۙ&�I��iޠ�����������=F�+f�8��|��|�ʀ�W��%	,�y�0�/���@7_D�	�Sto$�o�vS�;�,���H':�Do��^T������=�(��>⹮�~�勉O�?�S�P�PK��+|<T-��S�.�F��]�%"���A���V�I�:����g&�լp��x�{ ���^����YZa/��d.�(8���o`��U��x;�j�p�`%Q�+�t��z��3�P�D���O��7cr�*P�`��H�����E*��j[���qVm�,[�r7J���m�ك�����ݏ?FQ}��✬b$̧߃q%7�ap������*�*K+�8���!���G���t
XQ�x���s�o�$���C}mfsu����3*=�-C�������Y������F� &C5�=�F�IQ�{�j�a�ɿ%����T!%��~�"�@O|
ܚ�5�%�x�FN.�KX�Ҹ��t�;2Y=yg�Gҩj�����x�=��GԶ��7����=�ۧ����F��$lǐ+W˝(�(]B�C1@s�R�]�>;��& k�zq��Wח�����t]߶����BN�l���y,��s��#	J��F����*YQ��o�MF�>-AI�.Jf�֢���88�#���p;d�Y<� w>�Ƨ����:ȲF�����=}�	�S��~m��y4�$�ҹQ�\�Yi��){4���wTƍ, ��Z�ևc�k$�.o[�:����k6_�徹�=���%Ek���6βt�$+��\�%b�`��F5������1�������*���8y���E��I�^���m�Ҙ��O�=>���<W>}���Qm�p�_��5�eUF�q6&ݳ��T��RKn_�e�� L9��U���FG�s� 
�����~#�j|�� �a��*��iH��!����_��9OMHO��σ�x:���ķ��k�͗���?��_1"d��-W;>@Ǣ3i��/�dy�p�.�F	�-95���r�o���|�d�����Oaɠ
q_�G!D<d�QT�b����C�![�By��j����w��BO���.A���ֵ��n+R�fʜ �A��L���S��_OV�{C}��I��7-U��U��ݏ�r>:�䚩�L���/�t���"�d2����(�[�I�xF2O[��&mʋ0D��pyD�o�q����ӕ�j��$cg-�-�-����c�0����K�ab���������O�a�W%�X(v��u��m���?����������O�t��R>�Uq�=�6�;=����' ;;l<H+Q��5ÊO�UΆ(�ӶD��]�o.���[l���t��1�h���p#$��u-9�X�XX�RhA7RZb���`�-"���;9�%�0�FzWj�bR�>�'�+o��%�O���p�}�mGQք����r<m��kl�}���#�CVn���E�A�����]xZ�c�ȡ7W� ����>��l��F�0�A� �l��%ˁu�Y*�W�,˾�' ��P��|H��۶Ս:?]��p��ە>��Y�?����>v�ʋ%�A�QC�]P+���YOɁfA���<��R1��Y�Y(�p�S��f��|C�]������[�z��6p�Z;�bӂ��j@�K7��G4t�}��ea`�ic��=d���%���Af� �F%�_	Uu>�܌����ǂnP�BT�m�{'|����&��b �V7w늡�z�R�I^� �����$ų�Ys?Z��'/^|�;��ƥ�Q�:5�R�e�6�O��bĉ����%�7�-�Wcb�4"�/|�	��ʗz��ӓk�p��L���b��P������3�����L�ǫ�+	�!ʶ�$����c�����޻TR+%s���Ir%��~��:> 5���p!�b�+��QP��7wP0��Yr�d?<=�d����G>sZP��|2�΂�{|r��?E���J
�1�W,;;V�V� g�\�<n��v� ���|�,ܘh�0�����N�Ȓ��,y�U�Ӑ��I�O�RĽNT2_oj\~F����l��#ٟ��qO����%/�l�i��_�!o��H�Q��z�m�ގ�����t�`9����Ӥ�	9�
UM���2H0��+J�:o������~����!�X��)GH
hFd��p�7?��Vv.���/)O��n<�p�Ӝ�����In�]�����$���5����|���6�����oL��k��D\CV��z񾗉��_���w���tzY^��ަ���I2��)=�L�|`�_`L���R"�w�?/+\-��Z�ok>B�OɡA�X̙��3�q4c��8Jx">u�k�@n�޲8��R�pd!�n�F-��4[h��O�A�ښ2~5�3s�W4H�s�=�a���l����3^��?�.ѯ�
�a��EcSʟk���IVm��9F�(Q��/�<K�V�,H�j*gONa�`c�B���'g</�eن��~�����-�\���+�č�y��;Y_
gUCޟ���|�^W{���PBX��dL��wu+�>�jz�q���q�m=�.�{���aX�K�]��R�M���6[�����TE�]yy���_A!�#Hg�yL��P�1&��& A�w]H���Y|�c��(K�]k8k2���pDpь�\�2�Dh��b@�i2N�5���~6@��l ���y?�s2x���H�jKou)��~��`�O��րЁ�Qw/@G����	)��P���Mx��|���.�~�b�ǺJ���vPz*���셓`�Z�y���O˥(qcq����'�v����=׉��՟9�|�Y^c��nP�~�ܵ~�O�,'}}��N��,7�e(լ�?�^����"}�|]�3���CQ�@���uY=����˱�C8R��U�a�6�=b�ȋ��#���Z��[BY�BBݹ˘e�,�;�O ��'�m��g#�<���6�d.+���������&��?�����Tz#�oie�$�]H��<`�m�G���S��-�]Ɣ���h�D0+Q���V�����s(���D���b�Dm���w���
�9�NR�Ǟ��p�Zw�yH��s)��[�~�(�iA�0���S_�]l��(��8L��܋����6�-񍿬����^[w�\�?�F�B	O@ y(�t�ĕ���_���^�x����8�zr�/�R�Ҕ���겮ZZ/��xpЛ�l\7�cX�Y���"g���[3b/�4�<r��,����hx%��E���4,���#��Eɲ/����}���-3�X���ʆ��`��+�,N;,
�L}�A��q��H#�<�"��~��Q��D��I��e�g�z]V���HC��j	k�T�٭:�j�	��v��H"N���4.m�OaF�uFju�ț�+�p��V�{�O�}Cp��I%v;�����ٻ���,���*z�6����<v�S�6J��1�PZl��ޕܧ>�^�dNB	LJ��ن0hR"k������d����cZ�ԝE�q�5�����+�g;�!л�.�ULg8U�/�k��F��9Q��\�?�����7ϻV@㏇�� �������;_������:Q���kx������+�Q��(O�V��D�Z�Y*O�:kc��hx��JH �[��t��h����6�P�L6���Rl�k�����?����'��!��q��Q�Jߗ$�t�R�3���j~e�T q�#���y�Ek��Ӽ�Z�~S�V��lܿ�c^9�gaI3^|*%�:�O���6�H!"��V85�rd�n���G|߾�p�o`Z+�#��~���ѕ%����ے�{��:��cUb��Me`B	��0Dm�O[���iYD�Kk �8��/��1���*4�[�R�:��a�#�V|�4��$��m��y�)��'ţ+%� ��Zhm-6@]� �^M����3]�\Ҏ�#t��_��U'\u�K9=���4Uebc\ k����$<ag�>���K
��i�ݻ��&��S����|r�&�a#y���́z�����Ef��E�/�u�)ӹh\��&���*��/��jV����"���u�N	��{m�ŜG#�\ћ�/{3�������f}߯��g7���^/��w��6����_[@GT�z���S��|i�F���QrQ@�_��n��B�%�>�BL�
s�O���r4�`�p���Sb�M"�%=��8��<zM�Ľ��$lq��?lU��Q�9�8��FBٖuťm��4���i���ճ��s�_���j��C��{�T�Ã�xtb�u�Jd�YFp-�P0��oףϹ�:�����trO�ឪŬ��~�W	�m"f��`��i���ȱ������N������Q�!��
AYZD�N�9��9��=p�8��	��L��{�x�v:���:���D��R���KSS�ʓ��&$S��V�.��{F�9�B&�j#.��`�`}`,M�xk�@���3 ��jZ02ٲ�Hrt>P��5�>�����-�,���II+
֓��	"v0+t�6Z��GFP1�5��,��D��sc���qE�+��$k�-�H�,̷E	�&G�[\lóP�����W�b��6?���
����u�[��w�֙ ���� �*�.#=� @���,�=jGj���� 2g���"���I�tF1��N����b�Z14��ˎ���Q��\�$<�H��S�0��'�Ӵ�iԗ���}H�����]Fq9?!��Fplj������"��$aN=�V����Z�߰��jP�J��1��Gva�p��!�p�Wx��)�̈́B0xȳ��B�*�!@;��X�"2�WG�h�@�~��ryאK�����d�+��S����#��D�	��,�N"77F���XT�ݦ�%f䔥��`��s�B�sT��ٺ締�ҽ��X-�틈f7N57d�5T����jܔ��3�ࣗTЗ�X)�����]�E'���š+�Tn!J`F����R���=����5ۙ/{`�
�� �v�Sa��`��O7i(���c�;Mӆi��)���"���8�uV�}!jq��V�U���
�ж]��s�R4u����!�[~���n�6����nGo˂����sIj+3����8 �w�,�ڧ�I� ߟi>
t�ˏ�b���KK��`��U����������j#�d�FG/^��"18�.�Tf����b��!�)~?�9I�,+E�%.�Օ�9%W2�7R4 *ݸe��aSW�~�a$F8��aE��2�J� ZE��!�;T����}����l�(
�Z�| uq7��s]��/��b]�Z
�a���y�@u�� ���$e�a�Q4oٍ� �����z����]�L�Nb3,��>��U 9�:>Oƥ�5	3u���A<�����Uw�,�fۑ�ך�'��Cz�R&��N��y�D� �YP��Ao�p�2�U4p�  �/���o�6�%x���7�� �S)��c�E�E����K�.�8t-���9��9@['��O���u��[R�K+�Y�x+�JפF)OD��Y��p�w�ֳ���	��ȏ�q��lhKq�������|<��];ڶR�δ*�bߗB�.�x�Z�D�^�G��~y" ��c��p���̑0�f\g�Z?��xS��5���A�b��:R�aM/`?�".$��Dٿ�I2)�-�n�LcM�6�Lr���R9�`�[���A�/�b���c:��|�'K�Z�}9v=1�LŶ*��A�֐���b˯�[��wH�W9�����;��ʅ�M� �`I̟�B�m�Y�P�iq�`ut"���&|.u���+�\$p.�
�n���)��[�[�JӂƝ�1�o�^u���,�,ڰB���׽�3�o�XS�;��v�[:alf9�r�y]�A�囫��v*�b��X�����$�*��&�"���zc�щ iG%���Q�.�Q��i�օX����s���X�w�}=U�$����8*P]�V��d҄p�Պj�"���W��fopVO}��Þ�����w�88B,q]��^���e�>M�Z�4	��^��d�lዾ;�y�_�P�m!u@6���U"�x�+� �Dn/D�~Цԃh3��(��p{��qp
}�h� ���C����N �⹆ʂb��d��U�Tq�~�^�����sʜ�ȕ�j�>��.��9F�B`�5�~�.f�=IHv/J�Iĝ�I���\���N{s��^��������Z�z0�c�#u�c�`Ҥ皗���N,����obh��P�?�G��F0��X��W�4i��v��7�Xe\h~��b�%D�)�(c�
?�]��(Z�tuAˬ�!��}�䏾.l?@��b���lM���4%lw����%K�9�=�!~qMS��8��^�X�5,�t~�M)��n�֋��Ac���w u�_�ݻ�I42���xj��Ý���Io ��l��wb\�z�Ҍ2�D�7�;��p��M��F}�?dFa��7���H�ʏ�.��-�/"+��&�YF'���Viڊ[Gs�p�@q䶹aI��.��������@��X}*7�UzqT"��;��ʼ�F<7��#D�cV/A<C>��m{����v{�s��@��H/���Ĝ�����?,
�J g�^��9�Ѱ�כ�eW=?%l��Mo����兊���UX��V��?�����7-l�y��ٗ)v�4�޲�F�l�aw%��'M��.��tXp�8��7�K�E����H)�\�-^+RB�$�^8�!O^����'���b���d���*XqD�ԫ����0�%�,�wǍߡm�AQ�+>�G��p2�am����	ğ0ȝf���nY�zL\�k�mRHS��H%&GE���M�_å���R�h�hlO�I<�$�����+9�x��)ʰ��c��_�<cS{{u��|>n�����#r-�캫�>AQ�,`mE���gZ�7���䚵�]7�R�ۼl��5���.2�+�\�sʩ��i�����.�� ���~=cb׃w"���L,��)��W��`� �DB�()��|w�������M�C�$�2|8б�����9��
9�����-)�MkSm�"�U�����Ț +D��eL6~2XI�e�V1E��)��+'��;, JJ��݅K�-L@��)�0AuS$����Q�Ho���6�'ј�.�*�zA�Ԉ�pU�X��y Y8�ƒϊ���]N�sy�ܖ a����{�;��m�1FtL�K����>пK���g[,��W�g� �, �����Q'�c'k�C�%(\��o�c�e�����ue(�=`Ce�l�("ǵ�J�ȡ�N+yýmn]������P)��dp�r�M�uz�t���O�ZS�?���H�.��{v 	�L����HWV3
e���YL��Ͱ�dU+�~R (�0�K^�����8� �u��.x��+���T2	+��թAJeԻ�ۆ���g�5�͘�_�/m�mn��	��v����R�Bn]�~�����X�z�a���|Tj.3�C�i�!��<ˈCJ�e ��H4�f�Z��[	3u�>�#0�:r�/Cb�u�f$�U���c�	�$|u�rs�Z���.p���p��68a��Ms�R<��Y$��x;c��?��ks��#
�\5���]����Ֆz�(U
�/ӆ�ḷ�z+UB����f����d=Ndh�#��z
������;wL(z_�k�\��\z��͛�XY|f�y�@�$�y@W��ar����4$� FM:�M�q�O�:�zz	�$:(����� Me(𠏏50m�%dhf�M�8❂Mw\Af�)����/s�82��V����8�ަ�#�K��+���B����y>�(`�;8�� ��s��a�J�G�D���8�*������`X�*�y�k�X�}9�p�|�+�=���4v�r�T$��P	�\�C�B��q��]c�R�}��(d^t�L��z�ثir�d�8G���5�7_!�J�h�n��<�$�+ۑ%�[fj�RF����7�j��[+��=VJSH|ks�q+Qֲr�����R���q��g���B4Y^3F���@���U�A��~�;[m^MC>�oFҾ��Z#�X"���_���C &�u"!Q�O���o~���Y�L��4ۭ�_}�]dV#��H�рFY!�5S�v��Ņ]}�&�Q��:�$��d+T�N�%H�k49�wMr7{��a���}.)��V��qҮd�w�b,�L�7Xx
 �t4���u����k(�{��FnlH���¨RO4�9(�ڪ��X=q�+���mhe�Q���~��%:�V��sQOk���&���g_"��ߗ��4^�x�O���,N�<�
��͝�G�� ϔ�[+{�,>*'�cq�e�fM�xm��g1b�Đ�D���A7�F_%��.~
�$�&��W��a�S��z
�L���q9�]�tH�4%��$H��I�3�� \]`�d��&a�# c��qx��_n�T��֜��^��ƺ���8���H��WG/����"�n�iۜcxMݴ���9!�1LJ�c��O!���Vo��
����%�fd4�����p&�_�%��]�>��x��0Q�����VɬeH#�٠�І��W�>�;O����6���Η���}0ݫ�R�{8h�Pod��)���R���_n�ľ��7����
��*�L$��і|FW�%F���/���c֎��KK=,�H�F.=��EY�JQ�J��r%���U�,R١���+*1R?���7��=���h)���t�d��Һ�
��,�R�,g�kx/�_^/�����C���Y��(|v���#�<�ӛS ���zZSz����@���fz��\��М_���)0ͭ4]�ǐ