`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74304)
`protect data_block
0QIbnBTqgEhxgFZYMqrVOM/S+i5HSCZAv/Oo2cOKQk1iiIir+OEBiklLQdu1oNYN0N/d9Bdt+qzc
JXmkwPIRAuaY+xIMvYt4p4aHSg0dU9/cfBGMu6hv6OxtE1Y0+tWqJDXRdBNkWcbEkKxLQHKci4qy
B7lEOR0+vAb6gXDccNqd17Tj0yIbbp8FnwlQJRTeNN07Fa1dW3/iveODwq/tSpsgMvo7AB99W+50
kbhQIEiECdns0fYXp9DVbiIlv1mWpjV7VSEbhJooFnKe4hrxIaYRqvsN6AxK0TaP7fHeQR8QLbjy
0ken7ZQ3ptwloeONhFvMVZK3bdP7vzEZXpZCkIwStabfViDtPcRCZD004YTJqXmYdxV+28FP9uZ+
pKqYy1bazyU2b7xw8dug6yt1CI7USlan9jMltCzDfGkHZPozMUvrIR3q+2Vx4vliSaTzAZp1tUsv
SDtV9jIxTmXg9emW0CxWfgtNt0SEGWN6hS/3i4ZB7rv5R28RsZov1QqMRCp5WIZV+ylz6PUnLLEv
zxhsF2uGzSEQhSVZ2NOqrUwKAtkGcrx99tjR4PCpcdGLyJcoNKESz3ScF0ZsyDQUKc4uvrkuE8wE
aQ1IBjzdCvW+f1XcPVIIDPWmIDdZQLJZtf2V+SWc5xVDzOjcJv+lgLeCdciYTdrr4bmro6jgSAHX
XJpkd/YAYuM8Pbn0mExurheoSxGIL5sGHG4t1GGWJ4UqeYCTOfCEbCZXLUxsbTvSn6hisk3+raPa
IUbYVwQBmH+tHG7yzG1WqMEcPOAtP+PFwHDdxqWg7vczYtMLG85DOvyw26n5hGVIHPPVNF0yPFJp
zRx1rmcQzX5/5dexliYk271iryD1njGjayb1qqNFx1UV+9F9gl9ihmdCbJvXhHboXsuhBq0XbKQz
VucZ1mVtm1bFSYH43JQTbe39E7QqNH0RiPeFPbJO0Fc3nn4Nz6vG204HjCx/GJ5aNfc24feyJldw
HkLtn0rsWt1c5phAlZr2qreWwIHwhkL1OArAJFW/JG4yk60eSirnp/nKirHZr2PAWzGadfNAZYEQ
hyRorwI00KX7tnTk883grl9Akvapx7RuHyX0DLJx6uJqB+lDnkSQFlV5zBIyTxItkAyQC9k1eqNh
mox1E7rcGXtE1a+QWA1KgMiKczSas25krnOcfd9+JbzCt9vpbChNaa4q7X5n+VTPD7yTZc05waQA
3DwkTO7mUiuAChk9d0ZTp2mgL1lc2j7PR9y9tDaXP/DnEpuuft7QgcdrAB0MYWtgP0QRnzu3a87K
gy8s1+2AvaVxkCCRql1dmMbxMwvQ6k34U3b3R8oK0oJHp7dpjfUDVG5N/fnGLhaLgDE20B1gNt/T
TPvccPQMbjD8/Bc0CcFBcflKlAUSJbUH8VB8YJQ3Tyzi7IUI1Zbqeptk8IRuHOW3mQY8GjnIYzEf
pRx9+/ehaJ0EPRvAdLxrkWEDWuTl6LGl3zy/N1V7dZ2qpOeu4OHvUfckRAw9uIQHSQHerlfo8K0z
4GbwNqte/7fvreJb4rtySUz2axlFRziEzclhBqC3aTlV0kZNcHpkA0lzRWjv4uK/mnoavi26AGcM
YJUXRwy50l7YSIkF+wz/QXJGlmARS24r0Pd+fjJ3CjOKDRXL26J2+Kyhp+BIE3MgXL3WVE7fweGY
juMA4iWJ2cc2QphEaH5bbS7vMX8ZvFu4jw4g6KYEuu3SduFMmkkXcbfIcETWLigB+7YZ3bzuvszf
qxakKAqdNR6YOkrGiWEPNndie9Q7CO7JkxYcL3V0XFIh1PKevaiOCRWju1qH/YPb+hrC9+rcpVFC
UooiOntx6X4i8UtnJDYRhejBK0RSdk+hbVie7PJV7YeRNnxWvircyRHIa5BnSbsIgdNLdNqdvTW1
0Aq18CRfEXrDYTYj3oGnHilGQWpzLgojxfBxelnbd14GDSJQiJsqtfESeE9XmtTu11DR/T2gYaiR
apt7sjeAIMjcP519mhr0FXHYnX/fo3D8Yd7SaVytrnCX7nbTbuCn4KF5iVCtZQYGfLcqQYEpMr/S
/nb/i2cJIET0xKE60KrwSO9Azo1vB38zWeJ/lzAT0QaTRGwtASRe2X6i3BRseDE4x/VHK7LOqqcc
vQd76eFBuWpc8mCXCayiSvixmd3eGpnd4m0LHBhjwbUT7MlBfu0JkddLkgUEa9IaqEv5OzFWOtCi
vr4gpPh8PgTIfHtXQ0tE9Apk8R3VgK9owmY9kwbyPPIWyf0ETyAbergM0ZQrcH4UMYmD2aIO7sde
7epZFSH3rEHdouI7CdmlfguhUv4Geq7iy3qwKk7ziDO2BF90wErrIlJRolvPeiKKZ2AQjFZuTmhZ
qLMS76NQneGXfa3+RSj+DgF/vGcJzXet1sa/xIEc92SoX2KQdUPx/di9RrCukYhB0TiDDobBER6t
TBatpxrgx7F9U5mnCzxsFZ64+8JZnnTk3uWivoESZlz7oWixw74RsasvVq4FlAik3o+paiwKNYxT
LQVr08/Ioxz8LoMmNDyK2raGRGQxuumLJuoCTVT1E89cvzJsnRDCS1cePI+jgfb0n7ePAs0wXzqu
5b6uKLZAnGEQs5YLTVPVIPHlCdAoqaGGN53n3pxrgCBjFMoObj0pp341It9TKFnN65HfaFtuihnU
YDmF+FE93bEJLTbs72uVyNpnGyFWRF9q7jHT93vCrRhCgQ0bNvREgj55Go2t/LcOF8sDXOkvPLGO
8A1plRodT52cliaXcvLSFwnVVIjEc2EoVlyuFf2BGgwR0ANX3DtA46G5EOYDHkEkYMQezT7TuVeC
jQ+zAM8kKi7xb5Gch31+acOobg62zbT/+pR7+ISqXgj+h9k0bagsdhoq4+uItz+wey41z2ziimcl
cYKiYRctLQF+PB3UyI8v4vD22VkZq3k4H6qxoJ209uYWpDK9nYZ1SbHOG9o/pqCJ5tqmv8nW22RA
hVIY06Ec4CDlafHbNUHZ6SAGDKzGKEZlJBQddYn2vIvoS0NIvYOBW5WaurweKo9sLbrxcWMEh8/U
7CTRexqbkRB+oeCich9yjt57i3XREky72xDb4+VcIJYxs24dBJ6Us0DuCWdISB/W8UgNRKWJzfvZ
Qp4m3yLNcXNE1tjEy6FtIHrLTASNyEkC1exImc50l0P7saqG5pjUmwMjTapDiqpbYIGR5L8mVTip
t2NUTPvxdd4YpZJowMDTwcvqba3CZgc/J7DA0zU/+LnCI+dwm+byD1tETxjJfXciEH7FnoGCcwsl
cwjHeZ+kA+X36efYvZ8QY9z2WtNWHC7/129H6o/53pCW6RH1ZMhXjLrLA0cLFk/iDTDI/IvgLWsv
yYcu1LNK5do/tkFv7UHOD6jFzO3XZRboGZ6/gJzTMfLHYsJ6hId2DKt6OciFdcHNAHudvH2uE2lw
CbteF5AoCEV7Uan1b3kWzrmYqM9VeZIf7CiLquoG+bJwknayfHXIdgB1ildtnIQd2tq181o4jNme
ooyeOOTKVCBcpE3lQc7wZUF7XbcH10Sr/urGOWZYYBTp4sMuH4TmTmdBpeRmQ+vCrPPK4/TwX7i4
bQJOjlDdlpnt+T6FsGXB4eEWw3rd9i6r7eFO/Pc0bbpCVHZxJgQCGy6BgSsneeF7dgu0N8LRxKDH
b2IdEpUj6LJ9pToQRxCpdp22Lv7nFeFnTJXZsC5MPMq7OtemKxRRlFU+iuXb2mYjLI7mXysoZSKh
xMpqxK3lNnonjMWRzxu/1K5ibRTGlZYAs95Q3CzIgNKaoaxczmHCgusH1nP3D7Y257vsJX2z4bdn
sdMwhAcbYEYjFOeduYfhiBKwoUMAGl7DArUzJYaIh8y+kq75uczLIalMJZ4rCyPE+h0ZDPE6GGgi
nF+XJ2jYTFJ9R1dlPaMs8WacKnzJu1Fgv96oymWc2fm8CA+lGFrmzed5KsuzESscwWmF4zR5BKKo
qaoEudY0uhs/Z1Qvy7QPuDW4Jei3MgruJ154ZpsOBducVEf2+9k68Vk/Ye2w8XlsrEu/kY/5XI95
9TBvRdBc2xz3Zw6aiNdo7a25nde7x2h7D7s2B9AIybnA3gDU9YebkcjTT7t11gbVtLUID3OxgkLX
JFFvaz3OtSvym3Ms4CTDXMY2SQvYQaOowWKvczAI7BHqfZHrMNZ/U7KyKbTtlroRNmGyO9QWBMDh
dEcIKP8w/SvTqwv84qpS2eJduxHKDXFAAr4dhckpJrFJSNi3Iu7UROJrbcOHwIo6Kmti1xE2rHHT
+Wh8uNnUVyrKzRT2UfDdBJxDgsYHrgGmLbR653hQgpXTCjRn3eKmI7MBM62mJjgyBH3nCdRPIqBT
S73zJGifFyiQY3SO8N+kwhw/kTpteKgHQbq47vchlLUZ6ejQKwcsCm++FMnaUKn2AZqnrWzjO+Y1
qwkuX33aRbIlQcwIm5AQMpkp7TvqleUV+8VB6urI17xF814EK6syvcDV40qxQB2zfKaeYlLT16vb
f/NFJEgaru57SdsgheOJ/nJZxwc0CgRgAzRfT/4+7JxNElRdTLfqtMyJkjAI5EqAfpChVUBecJoC
dqAceu0Uz2tWn41gtHo8/Sejkj/Rn4ZES6x8cAe43MwNcrbVsXHOyKWT5yCdaiWh7VVaZEtS/pTO
g5uEzJ6fbZ2UuEGjqCXGyszIHXh04dtKDAe7a5gCNQ8fay2J6XJmtemHM8AWs3xkpQyE/IAW8J67
RSLCTtIE0DSVP2ITqzGrnhKTc/D0hOdb2+oOonGYgmwiJq+uM7bFxn1+fZLB0s7KWXPzC2rJhr2p
H+hqQ0YlPGJ1TF+acjQjrULEalHIp8ITO+y+2rvDDHt7IK7DxAg3EvSIYjx1GaCiCBBvWjl3o9u3
KeFRE3h1f6rL9Lvw8MvV2KBBi8canDpz2T60fwZ4VGunNz9yYcf1Nyyy8VBqxms0VeQQhYTSRi+K
HV87MoIRQBnfWQm3aiirl7zJopZ+51iqC4FpaPCe3ulGXNDx4jJle6DQGVG7xz5Ju81DSzZvbapb
wKr6ysg4VpTHkYlKotfTO4WKC4bAMUO79uiKf458uQL/i3UHBGoiNX7TJEYT4qCefApo97IH9EjF
8DEFF+oh5r2JzNUzNra0Jdh5se0GTGpmrFsY8dblOpY3EYkExE6lr04xF7+X07KKUhbluMmAlxax
espWL4UwKNmM9CTwIKsxk3Y0ENMnfpY4QggnY2aarpQPpEmE67sjfJWurUtnSJV+BkCt725nPkc+
miIxDQRU2F4gLP99ld7XfjyigLTetj+Viwp6rrrY2J3IaxypVj8/2fCfVx7wOyyb9YcGMlmXdyal
dcgYEUk8svmkwTXAP5dxwZidvJNiuO9TRWQJm/pBiVDf/F6J9cynFlPcYTFhOhQNGW8ew1QrA1l3
Md+VTrkjkAozdeA6NCzp6qUzegNBMwzdr0NvrGcnddtA3EfiMWiR1e0zTcmT6QFNOE17gNgRkt/I
iQUsr9VwBvBeKxVOfvNYXymuD47YmswrlywC49JxA5L0sSKWvoixcxs6s7vgy8djW/fIUVYCn4tf
OGcoroQ6FeRCgP8zFTFBol62plHDCVmdlotPaZsCjp/HYJue+IouZixuV6EapKEVMOnhfySvXQBc
hv98vkuXw+2H9es0bRa0ay/aM3eO5VDoTWI0DGZG76gRL3Ymi8BtWZaV+kz5yUWXsm2fDACjsjfX
caFyS8vrgJYxDS/EdeoitLPpJqcRRvk+KdD6w+SGncTHYFp8/zS0AndovFv9YRZhRUvM+M8vORue
dGTWPLZP0YYogUcPL53X5WdveUNbnXF2TtMAXzfJ3xfCogs+EbppFINTnuWcHkpFg1VkXmpzWiUr
JsYvzPtR/Ou2GdeoD/nAmyLhi/VRRuNL3CNHkULa/E51okONsv9rvQh0wgvhTkHsUy7n0L1sAWWG
4wj5ArG1XauFq+LJHevx3fNeKGz1E4/ta4g71rWnXxz3+vEu7wDJP+J9+4aSMKOfbZMCQzHzBJSv
i8Zjk/KB86Vg4OZoXqbGtSWJdGd6elTg5OR9n6Zc8VvHKhL2Z7k+e7RggGb4pc+kxkxCbWoTP6Zb
9urg3YfKUijXfosHAAur5u2nMAbM21YPXrSe0QkN0+iASlH0B1kuV6TmtoScJGLgXumLzBjVXcfp
cPXVEGr64MtYViu/eY+Qoy1I6Nkb412FCZNNYkhNIf+rxZ0cJx2931ccW2Nf9lNILmFuhlHobjRF
vJbiVhVG4+gZLy0sMD6xshqJbAp8hb3EXrSXjfpwjchyyWMDs0xvawpF+dYGKR2bJsv8TAcyNx1U
Kpqe1Z7PFdg8foJDgFe/WsqBjQbdIbBbb/hi/UWS/SX+VIodT4NZZrvrpH6kbITPCNOPxYmErioO
bNVXBJ1z6rt4MWYe05kDCbHI+ES4ZkDXz7o4OZ5yH/SuKl045nkxdD+vrRDJ51jOZo9OwcttwrOI
thwnCg3pdIfPdPqJBmCUmnNm1Sm/kYhJ0YWai3gXHPOKPILUJvaK9B7woQeEzHNqBve7KFwlxOVh
ZS0EbswXHaNTLJk6AsojYg4MLhO7NIPkg6v8gAmDzZGp9SYm+/lDSvu9BxhI5myo6uB7K9VzV4r4
FfKSqLn/Pl3LPKbM8moqTbhgKn0s3iCJGYf+bj8nYBB/Wtceurplg3m8pPNLu4xbqyiNZgdUL+1J
aYrQnyzHs/G79lZduUs0Zl6EmrYxPWuswnJU4vthxZzzQRiL30xeTcgirZ6WhT9i7RgcnFFXCbMT
2SWJ2JIebAv2lGsL2sdn+/RGrfXTvrWJJRFIS1ku6+VzPUiQC1Y20Rf8cypDE4zbu2oVghQLJ365
PdPUcwAhdxRY8hPNis1jGP8hW0hVl98bJDMa1wzeKDTXSjcDTQw8VM6niBQ3VRiDPKouZkDZuAyn
Cn1Z9qxSpuGb5HSSD45dz9H4Zfqf7u2kx6jTMFjZeOBWWJ4Jp/xFLbNmMCK72fDdJPTvslSgQd6R
zYpj7DQqoFnTJY3AOkvuuCcI6KM3+njaaHEM5GFNek9nfcf+9dxPPCNKxEezpxPMaU2oKC4I7mgF
Z3yhwBHqtax6laPEatLX+altayLxeIc6VjKa/2HZJDU3A07SRjURmM37qg8FQWA0IjoZSbWUD1td
n+IUaKhNX8+abwesPmWKSwhCR7ENTbiLs+6KNrnJmMzY3eY/iJNtU94Ufg0p0MJ7XnotBbgYpVUW
3Kbk5huwA+jjvymAI8W3xqbf+WDET8bhf2V4LGzwKBWYxvWz7azSwZgJ4xTUczJ6OCEHXdgHHe/1
t4L79r1dgYEyitg1yKSHGctmZ6YOHnoriAGtZkKfsN8CcZMJxHHfCDdDWFCQ9G6L+vRL3L4arcLQ
FZNoF0+PeNhJm6OS3aAA8XWMmLt/+JjthDPflUcrryvRjQRTKDkMFreuVdDeUV+g7xudl69tAgCV
uNJJLN2RMVyFnkh0OKAbgCqWzF/slYNsqsBaWWeJhhfyg1yid2z0ZJpi3LY1JAhRhm2lZyEKfdKF
XXJ5wBHwQrRMYPh+sSx6APLoks6+OKsWXEwh6wJfbOL1OInZAoGh3YLY+gNl03uS0U7LXP+IpPWM
zZS268G8aATv6eZIECoMi1ccgOEjubJdD0oK6j6u6oH5y3ePkXi98qZ81gfROTFrPrHQopXnfERM
83DICXaP2mNO9y/tzn397dzg0lNkfPbDhXMeZL+cpLw5amfWdtiaCJ3g23FiIXUBNeqfQzdHVEDd
Om16+aqOKF2pb9YmtI+GrjEZHEJfVcQoXeLuykaRp/ZKoMSMRoOFr7oQPxT2P0CZdmGsCjzAXzg0
70lRSGCxM5c9NfHtN7IaYEw/NPTzf8ket7ua5kTnEI15ur06Wjo2njjeILt9NzUxguek8sj1BmQI
4tyckoEGW8ze1SaBQVmpPE+2lKTqSfFPnfY69tPM2UA6RZMO3XMgY6eHHBI0LNyZs3VVl1BZMeRY
Fr1plrlxD+WOpLPcAnNVRvL7ZFnFB5MTkBZx7uIEZDSFqscEemk5Fpq7U/5kK2hdTojSdUOUU8J3
JkLUeOnJTiYfMBebxH+1/6X6XYgS3oTsJXt1gBKMADU3VSyTF8YrEngpNvyDdYg8q9pXWsK0CQdB
KBy7EONWQzF3eNIbT0qJnFWBiSfT7LPAyIZlZyLjsRcY6/rGPyxrOCRjOkUqSM1AQammxG6AdeyG
ssNohJhxW5Xo0H9dzIAY7Iluy+CN+Vk9Clg5WADb8vzhSxmuYn0mu76GGBCXfpDGVqtgZk/4Izaz
G5TDYXeIhyujhnTzTbZimbe4ua6EK7OyB1OCf6Eg3PItceOaxt8UEQsBT78FFi/LYfT+fdmCXHsA
G4qi9Wlef7/eft2VPGTVq9stjH/QhD76CsajDKcB2KfJaeEQg8RCLqbriP2oItf4IFrhs8F4z1sT
dnRUPCGZgAIzacdRmEIaO2aQNjzzSw4qDCrJ+6CJYGb6PQuMxVjr5/HVsndOKFsePkK3/OhcTy8b
pCiDWxabO6Qp0Pl085mUQJR/mGV0AddThh29d9kClPt2iJQvHeT49qPVLi6brm9ys4WhzBwnHgOk
wdYahLj97KjvmSAr5ez1NLDkoHL7J6GwcZsSlUBjVP+beCr7oQ3P3fHxymorysYf85qbAT1pYKxe
8gbtgI4jekifileNGm/0iSPxGwVnMc4nJaQthvcgYgQS7Pp5nIJRqt7XSxlrFQvDECr6DAeqHWjS
DuyKDZEf8wZNzsVvJsBwcCgQi8toPcDC246cEQuRH+pG190YLXf4VQhkP+gD/frI6+x3n90vZy6M
ZWaUFgYUU1y+nWe50D+xkLgCKyuePHAOailh5S3iBSuMIaLwfD7Fx+LwmOccAQGRQa1VN/Jgh6uX
QZpZgWs75IfsSFQEUL0mLUiPPYPzp/ZoAfTFVTe5APFNZcl7iEJli60QEid59HyPPchiM8HeG/7P
8+GrzK2kvBNkNdzEtGbsvpWnLbSZsBbtC6lE5+dOUOgMuV0AY4sIzxLB7SFXPMd5Y1Lu/1AfKVdB
3aZJdbkima/mPwTLLn8YjgPaBRTWq01x8JRAk2GD1fKoL+GrfKKKDhXz8cbCE+D96C8evVpfSoPj
qT0sfGNv456YlUZW3r9ZpuPxK8+GRxr5BxF87emyE7PkCWWP5s4dipDK5TX7SyfvJajQfZ/Swf77
fRf4GwP5Y6ozHNJva+OFM40ZbT5nsJXxW/OI+BetQPSRENBM0/CrsQaYqASrYH2Im2Yu9dFHhVD4
wrYTInDDCoDveTS/m9IlOU2qUiIm3xXRKt/W8wZB1C1HLvoleKFgJM4a4KfHfJl3yPXfoxNxLT97
/6oLZX/5RhDBq101s95DSU5c6WxqwZdNfVbs7SNTexYmlrD/WFdPRV/R53Gun7ZHJnocjq7ERHLi
tAt4fH5ZP0t6HDV9onUhTrHe76dXjaUKzPlVNHfrVLboKa/XWMXQK8qS1P6LXQsCaLlujauuMmeE
uShfhXdkZxSQfGCcSBpD041+/G564CBvg3oXhIPzyDkLn/wtY246CcaNZ9XokHN5DH1v5NSAWF/o
EuiYBEiLnbWOwnR+4209Z9m6QpyOD4xZtWARWVpmCX3xhEzv+jAf042kQsLteO0+dD/fnpRIWeT7
hRmTtJTvQ3DqNfPrGHs1eIn7An1pqe3K7+jWfAB7T15ckM0ElytLwjbXB4FfrMVcyn8fkPUf7Li/
eq177ukIxRtEK4CGsLnvhssw3wQLqhVU/nWbsU8zYNRzFFfVWMUbi9SvmeQYTcZ08N/jNl0n6ZtQ
54ZdYQ0rMUB9A1ZqRSw4uf2pWdT2c9B31i6sYocJXbyV3+fhxzwijCp/ZtFV1sHCUaHZNdt4HFqK
FG7TPrP4jr1f9QmJrLHqr/sXHcV/K8drQtkA8XedeNDGZx6LPD6LOYTynwhDzaezjIinIC/AYkPQ
sS0J7rlvT5UGZznuGdKaPrRx3mBKPleCGQ0uBfw6GLprCAT2CDmFUCWQ8K+hcPZg2a/VeNodWm+L
iFY45LeDULtdEU0joLL8Dan0T+WWHoZ2LscOmqXazJVh9+f4eYAS/z5tvGTTyd6BibrG6DCJIege
nYcN0B+PdUfUQ5vFBp+0RvBwslLFg5fq8ZzHP738OUCiplwQvcYOkTdhGv3FKca6BUO8R+liqu8c
toTfxO8HO/PiLOs9+P217ncLNbiywKXcU4B8MA/mbQi7LYlEITTtLtK+91Enjp/FnmEeJpTN/rwP
5fG7Z/xqe0i1LusEii2a3lpSmq5d7kKSy/qr7VOoTV/l2hijK/FuPKVRJcViM2fQMskRnqghD5jg
tFUk/eLZsoXLltebOHfjtTFc0bwg+gEM+9TQgY75t/Cf5CcZEc4lpIa4BgQwWK2U8yBc5J4Y3dZy
mP13Uo9EJfyNK5hu6bft/qfyT5qfZwUn+ZN61fx4rRgX9qyRJEwCJ0ZowHtYr4vQ72/VBCTVbSVy
JA81v/ZF4vILb4phRlvlB4gNdbM35hqHm1gKfX9pD9jcQEnm1ty5b5nc1BwB87e0Cw0enUBCIv2j
oRYiwn74dtfMhZohxgVn3yK33en49EsFY8B53TX5glkuDN6x0oOJ/8zflB7KbRT6/i6T7Fk86ACi
ZdHtFaOinvh64RTkxYsi44YUgmPcODA9e//weicWTvlUalFxDZH4CbGSK7mDDsBAWcig6XLqrVZi
1ZPb+eyZ6O45T6SHssn8vEaPdArNY9XltRoJelBzp0ER77cwwffce5YTjHdgzvwUyFQq1fk8tyWs
MCMLNsJ0mIidT0072uc9JHiMV50pxrm96ywQEKzC9MrU/+NcssuQwcvjTQxteZ2LhdX/+UNFG3/l
Bao0P+wTloWWOZVub9NKGwWeAntIdX2bNn6U3oSjo/qMMIrjk7At3OKecgbM8FQoGy1gb7CkEbf2
vJHH+2KJrWlhRA13oynwvwQO387bUNhqQeFyp7grXie/yF3nL0qOujEZ9Yt9kqkEcy7wJlgvl9UJ
muhUf+pZGadUuUvYUexM5Gq4SpG3PtkGKRKb79p6Y9JXrL6Gszuc50FRNwvyLZUlTrMx9l7X9JVC
QkEjjUBPlrk+Ejhkfcw1SgIXrQOKl+k1y+P1NlnKSkikvjz2OtfaISGAK7fxU8wjkbkFzveCH+aU
SHqfjQSaNsJIInE2dquSafNZo8QtPYV5a1s6v6JwOMRffxweVUGS/H/fFpKGsNU0MBRVs266GGmI
tEo16vrQpQfN2aFaZH2qxBJG0zdUy/DBIDnBoZBTVI9+IMNrHCliunY8wMBnAhCDV5g6zmR9r6rp
opGO3qUMXzoiAEPJ6QpXe7bTFXXi3i4tTOSP/2ug8ITfYb+MYms7f9OjtW1HjTBU9o5FyZgj05zo
iLz5zK4GjooJZsMvBdMz1gJpNZZG4dJ9psMsCffQtzvf1fMn4cT74pQ2YVmcP+EoxWkOr67vM/CB
zMDW0CCCSC3J58EDTV8PKhgUMZShl9N1H/1PN+E1EenEGt3OXxePcyfpJ0Zh08ZwH0OEad/6mwvh
aVVQwFso7Y5vwgBV+tva3EgqPQG2YOzlRBsoYJzSzYNsSKSjp832x2zsxGjkDXxgBjOz948ydbon
yvw+fDNgOZ4u1Pph2eIEq0uu/tpKlL1E6P7IzhAU6HcW3vtf9Ccyi+c+/uAfcm3M6fkL+l4PKnLh
KMJihO8+LY05oy8K+GFFaqRKab7Eq5Xv2WmQLuQ6E/oSKM1ONn8U9UFkm1NaGh0a4OphlcvlVO+o
mMuMCkxGv851Q7zjaHDqy89qfVvUBDwmpuqA05t5iyETNeSwgLRA0qucXiQrjAIGLM2ruAOA+ERT
IAtXGCWVtWb9fGk48WcBvxsbmDSV3kwEcZA98RlxO3X1znBjpBCLDA6lNVDmJAQe7L5Yj84UWyNL
mNss8AWU+2a1mx7/wEwiYGetWjdopGWNEUvzXiA0tEeyX2g/scs/pk8ZWDf9WBN1ae5GOnyoASnN
XqqngYaTFVp8fNjJYUhXO/1txFK2mPW3Rsi4hBZ4lD57+pXvI0EENlmnnK6YPDW6HxW2QNy1QRpM
GYSSUoSpZ4Z455QAPw5m4Jj/R8NOHLNuJiGJXDjKtpP+9S7EWtGRRUdNpTM8kek3LzGaznF2EGQ7
pBHgQ8scm5ZnlBvrLIGFYYD0abWPs+TL2ZaH82DKXNiHcjgSdC1XtSQLA5ktWxFRPlU19iPd5jDl
i1QwE8JZ5nA/zx8SgteV9P5nqPo0OmwtfeLH7ZpDJfKu7mZXI10pJpz9GV2kiyop39tnSymyJFfZ
qD+Ue+89TnNEZdTy9t0gh/y8g1KqCVScmharfUWqfjcScaAz64Eni2SJXgpvAGgkhixmbZ/mXC45
QxYIqhzVpP4wdXQ7pNJeOdkxTI1KEcQxjtaxG6XFjFRPtht3J5z/ETXu6O72xQMLnt0vPovCynHD
/0efE8zoM5fOqF+rD61pDcaHTER98M13R5zBbseyu3mjWEm3koP3mYYnAqMYmuaJ08hKmqkxaFp5
ndpjAphZjXgmI+LcZO+HzDlbC7C0YU/Sq2ljiD6E/UAGamhRGfpK/5kT0QhvsqzCSQ2FYJvbD7n4
wqKCLoWNnMyBmlT0/Um6Tr5m4r9V8TyWoK8ePJKV3YBWerxGq5vMfComMjlL6OG/vGx/yWoQFgk/
pXw96NPYp9iYqwGZUIfMnM7NpDL7gBlcrzPhbIJL9e9lKLlh6KOdLhWnxCeVv7vY3cW+6EubVC/I
qUKx2byg0OzzA6o1hMd53H2b3Cc7/X2BY4XV8tuEVvon1pagSQflQxnmKemwMYhl14JYOzWZHc0m
UoQqvqTnnUNbZ9DOTc5UIuERZ/gn/YfR21Ge8OUBKruYCevlEbGMaWq1w1VDTIogyUbN5oQ2rsxF
iKIcqibNmApmk/ApnNWtIJbt3CWnWrUOrYxYuZMRkMARHFAN3MbvRNezrd6Aut1Vhk4/JrQ2JGNJ
gEMDPYhuyRucOqxuWXbfPMYG6mJoaxNgWKv/D5gyQG56y1mSG6q/qZUvK1bHfJrcpUsNRLsY67O2
gLH8EGrTDEZ3UAQ8V+lRlpP7YkKvJn1yFecCnK0/mO9uxVF2Ex2yBJy4iVKR+vvXTEcjVG9SUVRQ
6cYlMLkP/rIpB3z8Nz3yfYt65IhK4g+Ggr6NOirM5D4uLevijpgK5rSOo1GgF0VRNGXeR7RZknx9
k0rgi0uiNPv1ZxjX843xcz2vn6tlTBPjhoe/osX3fjpclUZhCZPuUFPVFnk8hX0o1OldfVK0oIMZ
JOBd7A55deLUyy7oE08DQovhRHOcz64LyPcf5S0bCuqAaMUqF/ymbbfrDcvIaIUxpe5M9tcR1In9
envLmr/Gv+mEzkGrt5SYQGs4OjJP61zCxtT+dIxztCMJWBumG+m0cTo8ExYk0iiIGZ9XO6TYZXMG
gz8nLXQ/11H05PWdqPdBi7wRIHc2JLedFPz2ErbfKXvFfGdZ5hqceeV03BjFEYH/kJ7y+eb++eLC
h46CPxGSWAMZzBxjaZG/YjbRs7SMq/jt2WsTa/eg4jO7tHjnUiygo1vHE8JhR17XrUs2kRwVeJNh
aaf8vCGXkkcO9uWmkKk1pbLK2urW3/vqPLuXqxa1l6Iki8c9yZTWurZN94pfVeet892aDDHw/KCH
jWkP6nivKHlnopIkA1Dtx9mGrs7DaD3PKekIrKUyFTIL9lo8M0SdZtvkHcJdqeUrpCQLKWSM1UB0
B6x9MOlO+coAXBJMR7mOxV66JGf4PORHwAo+VFOrjpChCTeUe8vcyHclEgEUG4guTNv5TRRepAwO
OBdkXzIMm8N/GIk/DOzPfgXwrfn9HoViRiF6aoZ65xVp64nn8RgBR28zSU/T6TsY7miq6G+Bo0wY
zNbMUn7mmipAyF8OaLX+oGrR4GL6j0RYsf2+Cjf/SqotZeK7xWsITo5flAz7n6HnqE5aXysS845c
rujMxHDMkI3m9kog3AVay9y89rTWvaqhBauLY4Agl7Fdgjlysp7SQzIYDsfu/K+vv88tpFQbWPcC
mGfQFVRnJcS2LozmTXeW/qrV3UcdUiZrwb57adhTo8phmQ2TXQUv7xMCLsZdKHl77eoE5eO5rGSs
PQpAHe4+wBlNi6/9Pue3b6Ci/t+JjQgy5ZCRWuCod5MPYaI58uJmPqr2rz3QfWxSpmgp9qF/EHRG
CSZItCvKTLKmxq+qBgymhE6/GAhXxann3yFYwT8uIX1bMgVBM08YUVzR+/59wX4PBLMkqRwgRCVH
BQNiCjPlDtBBqCnSYwx6puqi5k0bC2cXmsAPasv0bgeXv/hzuLNpADOYjuuE41IOEjF5apeJ2dBc
+aa8ntpklzsi+oZG0df8zt+9kFUNIuaCpvg2CbEzGm0bIjRHRfTVytnpfm5xwNAb5WWvWLaw1qmA
Cr4zvAj6EKzXcez3BQJfhcljIGR1qBmEw9GnP2OiUO7Htps2ffNKsfX9Kkcq0tl5OlGSJrKA9qAx
pU4b4JTjDSFzN5ibR7fxgBDodoBXD1iTz2GrNjvAogI3vO9vV2ZAIdzi0kJQC67q2Cv8DHdm9bHd
k0PbOhy7ZFJ1kkj+8zMS82/KB2U9sRRup8tp/XL6soLUqR8BEocbSrJPh1+qeljT4ivE7PV9Xc7Y
HPFeRC/fgWPT6omnM2EYiY27MUdpHPI0YX8UMQvlachSLNRmh2pICa9xZ6/EKalMAVDWQJ0xgDsS
UiV2l3zneUnh3T2kAk1CnHGFZPHTIxngL1lT5uM+5qP8bUUz1jPwTXRKRXxv1a6uznTfgQZ4Uo+V
m5Vf5/oUpzZdmL21GOB6pY1aVmeUzXUtbreGjqYDYA9e6o7/iGobrgw8t2L1L0T8dZ2j3INZ/p2F
uBCOT4UlW0g2ObjOTke4xsP1icn0WoSOLQVwYDhLhrx01sNrhzoZKlhZ1ADr6XgOhAGUQR4xdA73
BfzzPoMigelrB8i4/uDxY8VrFKM6XBlzxKb7WYYRLFMZaYudD6aKskUzPjijv8FoXqZdhnvJ6Jmx
rmbIOp2Q1Ilf02ttqWriuaEZJfHKkX0ZmXk9gePJbbzNxPrJKmU+EoSkKbfVt5Z6gQYoDsWhsNDg
aylHoo/dG05aF2a0l1s8b9GGqUIQp0qiXN+1VSIMyoyYCp6J6MHNKwRCCOa+Vts+CG30M8JmJDjU
CDV9NxCYw01MDJSMSowBmQ/3bbvFeSkLo6dHilu8h8Z3DhoSsSmdC2akd4ou//9KT+jsC+UPH2rh
gFl/EraIYx+2bggoAm5qvKJzP8b5xSJZANL5LTNf3GkLqQHXVXHyqUHD6kWMpF4ZS4XflwV5rliJ
HzPgbrkKdm0msOksAclxKU9AOU3tY9n5bARumT+8ui87mlL6ecxB2GFetg2MuFlTUelVv5AvrArB
+DlvCkMcNWNPWBRV3tv9HuPnjilyBaca9syBmags/pmqNHRMuKLaAm9tRCzGx/KZXNzNuLKyoWGe
5OWwLEJ9MKgf6+hDdF9x9x/CsZXt/jyQH7J49PaZ5owj+IZMV1FPE1rXamz5yc5Y826o2TA3GAzY
q56QU46nMklGPiQwjDps9hmyXqI961+t8P1kei/vMBDZN6pvPGoSn/2U96NpVxQ3zudfBmAhncic
qd3Gh4QjKC5UXh6FduoBk/1SBLge9xI4Q5Uw1kJJzU04NDulwf/GAObsYZQeCCa1oJz33xerJ3Qx
YLInltOuEzM+41MzgSxkxXmTvB6pLoZMidRbEkCPXw46eva+CqvyHQtfazAkJNJvMOTXnPT2T5wp
LsrTUNvcsHyPf7ctzbEui0+8eVIBJxKFMm8rHvFB3pDQSl6di4o3vabNHAGoC4/GhkITK+BHFdhi
za6qbDiXNY+GhvVQyrn2A45bEQrLyaKvfeYJoo9K07G0oUJessohFHm35maU6S5jlCXLVSZd7vqR
qdgoWFW9guga8LXWnYxztAarGzlxheisWcKuh6kK4wZ7ZI5NEW7AvB3G6kAiT9mjh34wntUsBgIE
fVw0uE1Pbf5hcTD27affskNbKl3EskDnpT4M4qapaCtvWSRVP7rX/FK66cEBxJQ20iePdO4ssXuj
YOPGPIH41SQmHnxWMKrJqYVl9ssylugSzvcHjKjyROhO50ZTYBmGaS9jC0UFpzI4zykOW1FvNGH4
XfPmfm0jl2QJSc8iC7a1axJJkNzgIsIyZTz6k/klQB98mKt7WThhQGiL742Aq161Q7lNMXt054Qp
15B06d29SMjEF5TksF49gqZFWfOPNy3GdRF6YvRMjPur+S1C0q+/l1UOIUCbXEO+F2D4LzpZ8Fel
gRDQOCK/c24gTBr01w9E+ONt4vZ5rE1MEPLZft3xJrPDgs/U7FmCDPPlv87My/wpBKgU5tX6kEGC
pgZstA7VI4WGOK0Zmu6Htv7DwO7/LiY7nrgHbeTYLXu5zQtKLMItYBCu1sSKw2a9mqkmgss+M/+q
oL5um5eLMk++jVRRweRsbavmkY87vwAlXxlZZrNYi6rjq37NPkxnZixbo68YAfEXyyEiCPxn1y9L
dn49yMMhfOdd9biwUKn9kzmbQamXH18hvxwSH5rKuCrtCCSCbpbir+HtxiPjANcDD7WZ6QadtFLn
ItiwfyRBZvv9yNAG3NjnH4sjKuoaX0PCT5WnTBkV7CrYCcM7RU4ux/ZEBo+HwjzTy2UK229WJNMI
tCWsexuN7Jj6jzWA8PSrBtVMhQ2bzgt4EiJaMicz74tCnz0MhvdWQnYi9kT4x3WZi4d90eh52iRy
2gIEJJf1OE5f7KRR5hIvxQC2B3GAdq/yTyZnXLLikxwbOAYjEABp6JXGtiUlRHopahtOeLGdBnSZ
T+EHxyhGO/D7aWp4SjSNu3k+qU2YqKcV1vdQS44Cibffy9fRfVXhGHfJ0uqo95xQxL+ISbC5neU6
L07fc0+6Z2hAPgBIuDxkfRrljkj8okS/tfFwtx2OZHZG194M1T4fZAjY7WVDGmcQu1GWtoCYZ54p
8OWNB9npwPqU7mkMaJ6ZnG0fj6vp/txnZ3wydslLqkFdW0Y09+JXhz4BUzw6oCm+LO1EHKWCEAzz
8bHzl7F9lsakiUhqJwJ8ukoAzOwsftnJkX3lOot17go1zXy/1T+IVaWzFj0+JD1uV8k6pG83+YAm
PksFfqU+TmjYQ90igwOJWsLp8BEmnn1wqaqSCz1LQSUwgRhNOk3Ii8T+nVXos1S3QoyM7wWpxb1O
ElRwMmU1T174yPpb8rD9GX1l/94OT7Gh4NSiL0Wsy3DROeCAd1GF7J2pDl/vakjTXxz2QM+Tg2P2
rrOb1/CJZxYD3C622taOBmL1r+PCoB9afZy80xEXcXkaALo/ce55IoVFJmKC6fenofPud7o8geCx
7sJ7ORrYB+OgNjr3QiIzUUfH4gMP6sAWy4RrqjbFRMFWKcNSNiOgDyA0uo7QijE4ismJsQjuaz36
89n7JhAuGoK2zXpJicSeA6YcQAxw3/OhkeryXjklAx/rR77IW0wfA6+tyWGJzERG1iVyhVFtkmiu
J2A88nRCKk9TDZm5YwJkkssymhSzyBmAntuFextTYidYoED6AEIbuwVO2wC5GjixrD0Tf75MGjRo
d1GKswHXEKUf403xtPEO1eYtez8HWXk45pB2dAl4mRCNdOkroIHXQCwRkGpSmwYSSw3X21mik6Fv
iNVwdyseUFaaAtydXEazPiDT4y0xI69SDl7rWl8z5SpiTYK97kKYRgBzyTI8wtjcDqhfvgLEwWXp
j1sMaPwWAKPSr/km0bJS0EXAnFV2iLEbiu7StXFe9w/ZKtWLtoNpEZJYXNtVUcY42CrUnDE2OJAF
50Kvra86BPwMcRxnC88d/KyjIjiiwfKVT59HWkxmss2fRic7zYFIfBxVxZHBqRdxZl/4owuOwyxR
xQeZMSnurgFn0mlx0Ga6lpOWmQ1dAeRPjx60te4sejGl0UtR1dt53oYyOERM8rbaOeyosjj0mwLk
OjSrpHPPdH+Ocr2uXsZMdRMYUt0YENEhe1u/RYLD29QYRtRSxCP0G9F+pVtCgwFOIFeWjtc8rN1O
NH4rc1Iz1EGUrE6hR7XY8EUATUnaFJnTtgmr0xqQVDK0D0FuA7G40gNEu/ZnYoHTsV5Y3aPJjQOz
dls2DTmzUx60+IcjlTkEjyO6Pg/JwsM/wfSJcrLt/A6Z1T9dpsjOnqEA4kT8u83wJzJ2I0A3exoV
J1MUxtF2wI5qLj60i4PcCRDfvEoNPL+dXBJyrjBs8QO4qRJKTNbextNjFANKhzDdG/BxL2PIRhEg
JffZ91ERFMdVnnM8bBhBIpAPcTrkRSyP8ttfJBU84bN/y4LrQ/uB31vW1fH2L08TyIWJGCaw6b7T
W+FEQFkTlgcjTV2g+oLGL3ZZAvUUGXWhMwF4FjHcDmCfPO0TvD8vdpU6kH6wnl6e1rpgQSDlu10P
NV1NcbxjKixbjEB/Q4c2FCXiBGY48HM8Ky7kMHjN5EApfQVzj871c+GZZBtoLoxF1D0gbjXX509E
ZwItyXR13loRB6BdtHsxa3M35e/suz79LHEsfI8zPKXa0rN1051I7I3MBDBi59wCRiqqhU/bXWR7
rjSPfJNq46xr4FwolsOh9dfgiVG2kYF/unPq2+5WFCXX3UJp/HAZNx711ai60tNqU2hZd9husQws
GeAb90JwevOHHAfCcqxh+2ZNl+Dv3vCnVwBuubXfCrz33piTB0bS39xK3DEKr7FIEQQOxHW+lg1X
yjxCamLYz4v5+0l/2mJmxqmVwvM3ush4DtI/+l07ZciVNllgCxl+UFMV4p1zsjoiGdKLkRIhqJr/
/f3UtLEy11JtVdYnzWr801mNWYka9etTgeNYd8g3XhQBpe4Bl8ftaBchR4DsENahIRp5tgWDVQIc
OUfvAN6dfVJSEFXoWD0EKDiVIAvz7r/cc751L/q19aP77j157DxQOSDB087ugeA7q5I0Qt06mI4+
NKKLzuf09RCCEV9lWYvmAU3StEOLSaVC8FhRCGdjfSoMpiSeOjLmf04sK0d5ece0oRzrbLNK1V/g
z245Kpe7x+M7ycWovimpQGOYtSLIeD4jxW2m7zl35gWRdoKMEDEq6EYT0coJvBdwooJMpTCH9jpd
RMztO0wHN07Bw6vAmTusqGpzmNrBBdCSWaAwR5BypsPmgRmI3+ND8SMy3CXwm+JWVzBfeR7jxFlW
WC7uPpgFcNWDDwMUixp/ztn4Diqje7E/3w76Z4iGLbHpnFhCLBsEi83nz8GfzglnJs2RPqd5oe0C
q/B9OI8hvycmD+0/HBb62B+MhLayOlAsrTChkcELBSf5Rybi2gGzdJYolxn8G+f9b6RpYVpQJCGi
xzVO5YSBU+XfPptDRLeanhaqHyIWobOgu2cPrcPycb76D/4Z9z59MLI4ipN5tiW5EnIYOFV2jDzn
6YFUsBeRAS8cwXWCcU3fEphvr9HiUlIRuZ6Wi14tfXTJBrsbaB1XV/TIp/zIKTWQrmebWH8OsgFI
esIdX6vlgWksa0B+A20JJWMEnsGMr0m9fc+k05jePA3sOMWgYOzjhbbllbkCuvpdNRwUBwuTpRbq
yOK71EXFVCD4L4EoiV8oWILqKIBObn9oWjQOVqh912CE3IStfyPsRnqDHUd8QZ5vbrryBB+SI49+
d7PSLVk/qCl7ehLgpZzODVufaNCgqvg3pTmd9+EK3D8rdSaodBxOGIdOT1+QJMZv1t/fS6FLzGpV
WHWBr8NzkWevbGBL3bZLpq+7M1SRpyvctDzEeONuLMSDLmd9PkpvgXHtw5LwoGYoH0JSGEcgiQAy
w2F/5okoiM86oMcY0HDwnaI1IcISC+7JD1m6cfAtg7wjSnBqTUVLUjAptRz0H3W8izu9sXCkphbt
6nbhviLFzH1BfGJ/QnR1UXcsoKhiBYKSGzP05pWHeGs/Dr1bfYe6HTDs4gwpnkfWDe5Fms3oipij
EgVnI4p92RLGLwr99Ow4DP3z7PB4oErG0Qq/Mu77oNjXHVJZnS0I+MlOS09jDJ6P/d9f+fp8m9aI
ekdWk8R2F+bO9GVBTqyD3U5LLJlKcYfORFsZZKYvbkNh88JmdKDR3Ne03RpWI25ZHg2WLb6Uid+O
r9PBXRHeX1NFzHAH/ETXH5/iSO8nP3eiCl9idcMQgb/+Sz6xc2OKP6mqvYyfsAHewSnNHet0go+W
Rfs/av3+dxvo0ntVyokamOu9UxzG4dmTI9aTAed2Y5pSQQyBDgHfBYKdlZcLu8FZ3UMWcZyZD7bb
ajpR8Z0rIvY+9vixeexkgq0l384aykf2KsZMQRluiXTk0yJIAFL7wXYkaur1XX8Po8u6hdOB8w7s
7P0qF4pJCHxZCCZ0I6BUCrLFpFmaWoiF9jDtkUKQ0EpOfZV/bQ8GRfDowXjeiGTGz9m11UXyE8LV
g44Fo6SEer5dv98cWbf+l5q+/q03am8oJkjIWjnYvikRf4nBWqkCeOn1D3uGWKqaGyYtJNeoWHa/
1oxHfFl56kn04BFgenwnqmBi0xY5IZWEgTVc9ka8Z/j+uQe17BQ9PnuV5LvqRZZvfvAkeZ8uMPZz
5t+qrJkYyStYFCce5BfoHL1HVVXCr36kr611VgzdpJ+FeivRhqvIHkJ1KaMwEgG+qgqWABVRHfBO
XITVKKrfGVKNmAdPzfkaR3k0JzzH7zIbPk0nU1mTrqgBIBTbE/VwiCr09G06burvSKse4XosDliD
xUW9jekcEhWvbH0UbFp/bnXRvcOl1Cfy1nGbg5WyS1UU1ZslWV46HRcJRZSEAqD4GOGzP9FLk/2Y
HGpeBABowJRhzEqqBklKz5iilOege3JSIjnKxu2nO5K1Fc9PsgEWYy6XUckrPYPdEUofpbnEQodq
33drqQ5w3WMozRtXtLl443ACfPEK9I+QUgKdHZRxlUBZmhGhP4vJj5ss1K+nnC74W8L+fe01jFlQ
rGSjxQKAy172lmdXKnvHVGtvRbE15yf+VjlDnY1Qll+1THczz6cr7KN6jiCcwUJXtJIu2iZaEbuK
+rPxwGGotUd6AEJVORavEdgPH1cetTK7JbLDc5/fuz2BSEnYhOwFTvqzq1Ca6N/rKlNNZxe8Ic/X
hhQWVXta+zcpDAt5dJv1ls4joew/V7fDhn+YsvvmrGkAXi7XxDizkseo5bJlhBr2jaMrOnnoAcZe
mk9U6JJyR67CmLcsey7sXmiqmd7+qu0k4MovvMFBCvcl0fm2jLUUG+18/mQnwuUEYdNlHw92eRjH
sjFkQ1jKw66ldyBRmpvJylvOPNz4CwQoI/lKTipRmn1lGS+NiHNTdyBOX/C5KwR508cS5hkdMc2s
VWT7JEXEI5tYmT/fVOIX7RNt29L4+BjEz3YGYEVDn/AHclZ7VrMeDEvmt9dA4/XuH7KRxSIGJWFD
zRz7HdulgTomM7wC1MNVHowZo7y1tSH0ACLzfrQNJguvdl/lM3WbywAp+KMORJkRIbVdTwVGsYAN
7VzXJ7y9bv4GSNCBipFwugdkikYgC+k7ScLTQhYyJ6a1QxUqwr4QIN0QF5rgmMXBmahXReDNXvYn
eqr9y5MKU4kLam2wE5eCWIKz6zMgR0xtXxNM/QnifYGj0SXPpg8XJsB3piBMeVtJCeJNzlHqnhNL
I5CJzONwLELC/hkDA/uC4Y2Gpa2MD+vhWOslIjO1A/tR7mO6PcLgBxy4Bkzfu1R/b61fEUtPDVgJ
ZI/mRZm9KhlLqrL4GjLoiYhw2PwNeegcvnYRPRyjSxFBTgKQfugQDj+vrgfMa5Co9ku8zq3CVyBo
LQmC1qLffsntUAzpT6kIYezxQ8mNXQydIcJDpO9AmNK6SVNvnssMi+xaTs7DHwbObML6crWjaPqc
JE792KtqoUxVoT/+IhWmbE1Yt5RrzHdK1TgoJXoLtYNW2tihYIbTfVXGzFg4k/zJ5ADkqruOeFrB
NuQZFk2+k8i8r0PGbm28PQ1rZ2NlS7KeFSXP8A7Wb5IIRzME37O1IsKnB6yUEnpHYlUaTfy7PKWF
Ts+lixWKvT9t5U/MLvCUmShWaE5fftzLScZG1q8UUSNmCyv18+cvBOJ6yfA+jsht5sMGscznlZBM
cKsT8Pos289+56fYO358qYemnMOyJ5jH5molGL/heiDZ8Vzv0gInUCA5E2ddmVOvaC7hF7o7zcat
kDY+M8Qm6M9OMx9uZeg6lVm82Vi+S/W61IrGI4hDetXGAVgluyfLmEagh6Rd8MIaO3RtFGTwNoRF
SRH95A0KYzAqBoccIHRnEFiedSRq78c//GsSkUysxfcZUOnVSCIw6O3xhyY/TGhgRJig1lozuV3A
hTRV94xTRpxh8l6H5GS6KMhs/tYYOvij6QmAJ31BsPmDJdQOr5rKee+I+F/WphX6ta4b9L2NmpDp
peg3jT0T5Yoq1sOzNmVtrqTUro+wOD26zU+Dl8akH4NM8fQ7TIKqMjPIugQc6rzbxt7IX8GVzwmW
JytfFN4ysNoqvm6/Va3pxURSGWqBYtNnl4JRMmR4IL9D1zO7wakmMzGwlZ/vxcvBevm93BGpefbm
1Ey4aNnMYMzYStZHJ9y3B3fz98yX40+rXhUjmoN0axCDdOuoD5nImdh5ysCsD9ZUEH/nCKkk3vIx
L3m/2UCArKQ0gyRrGB0annOK4qMgklZFWTo6V+i1uzFNZAgzPLz9EDpKmmMY1XWD5UWNyLm9xUjo
1XPRxfSIzm/ij1gza3D8eIKBfrYz75g5RhG31lK5Ua3koduH9qh70m4XiBhd0Tx2YsxpozTaMRkh
LTUF8wGMXDLPgXU8z5uOrP/RPx6crSEPde9Sdw+XWrQG6APYHeJCdaZlgDbDSWjAMOIYaTRn4Rt+
6RFTVbbuCktgkR3djQwP/anw8PjrS59EIjkZ1Am/5aRAJZe8/DAB0JLsdxX+F3/0rc/twsAapM3z
SWoOPz1n9uEY9aE55uOts+B01lyanSwezNUAK5D85g/TCy72/Tw3ntRcihTqsmgXJZcHBO0QtpAf
gYRqmMUzBOm5AOQvnEpW2r1kgrPcaGMArb8iBdkgKx5M5+GuSQZdVPurZZ18tN1ss2mA7RvFo5pk
EE3iv6F0WdYk3LsCYBk7KXKoILBDVqCU7+5CsLZAWiFuMqHnuXfKEymKkOmRleFzkqe8JQClezd6
V74Ij7Fk//TESTEL3XKuhRZLjYok1i6BzFfyzDC33RWd53dOqFO8OkiTLU3pyXqywNQriu98TaKZ
g8BgXFWuBp9ujzIvfsace3XCyb3XWPb5jcvfi3Sn74pj3kw5fKBqJZy/2DA18h68ibftN6gV72cK
kG3uicNL1A+rRa0EXlK0GS+ODg6cA6ZnZ0R4BKb7INKVL/lhbMGtwtVGD5KAleJSs2gLfTaoIYea
uEcmCKTAwecvbRow8rBndBvreDaCrLD5Qcb20iGHK6/7Swkfm/4BaVrqwol3GYq+g01gIBVWXVnG
QcUyp+pUZiJRcssdObNxQrtuguE23L1993qHX1eWE2RnZMZmdFIYJXh5MEjgY+/Mj6RH/mfeUefw
7juf8H4KgQcemgZE7O1JJ5Kk3LJT545TdrWUTvYnKHDhEH590x4zx4TKnH78lnutBit0TzjIQcHL
+EPTdi3aee60maZC65oJvvEUmgAIkvGbExdcWmjEHJHAGZ95PkHaTgSFXVp5TC09g8V0LCadb+FA
OrMpwZJxhBU7L9TADOulY0Ro0UIw4DArhEZ4keDIKlSDkd2Si5NFohvIH2bJz7Q4E37cRLCanNet
JsQe8kfkljGfp0ao9CioUnzPg8A5XqH4FFNnqPgT1k+LWyr6b6Q+SS6TSJKdHWj0miEKu6ybfsnm
E8cEHuRKDy24fZUF9iOAnlw+gDKiWBs1oBcRw9FSG0kJo4Lb+fCfPsD0fTBsGXitWyF3JLkTWLic
qPUeZJ/neG+qZpqniOH8MIfRs40YAokuE4/QDiceCE3/GnMPerbXi24A7chp1t9SXd9dvTK+ghes
OKey+gZsij9mv2cmqaEJprTIPzYiYEz8TnAtxtM0nZIkWKzhzITFMlkM5D9Z90ttHjALPS8k3Pee
g7RCeFSQaKvFBCXBtJcgUeuHT5qOa5HOW9dxzMnSOX8kRSJ5Q3LJxIG82JfAjNoISxXkslQjueJh
c87QyR8Vj7U+ehLVX0yvR+3+ioU5s188frTN2sE8IH7T8UOWeQle++hgsDp9qS/9ES0FGf64ggDl
Ta/Hmm+JpIsByuFnRrBFvsshHGL9jbnA9kan08O2Zv6Vg3IN6gBDAIdXwVFhW4EbMlGraoSQajw0
pjiE1BplydY1LduC5C+SoQE/BkrGa0Ir8RjH4hmSfzx2Tl3+DPsVPpGeyRYJNgaWvIraLEBV6kMu
+WJ9CEMptGCbdTiQBSaQfsCFEW4Lu3Nf5Zw0d2c+yPgR7oanFuv9bpAr9KyljRHFJHw3m73zD/2q
HSKUfEgPqj+oBlW+VT/Mnf6rsXWMoLYe8ak2DOjz1R6KrR3IJL+HY2xs7KZdZyhvRMNVihtJWgoZ
M4Q5cTviwo1BOKWP5LTpueG5WLOy25chj30BLVbxGszv8MaP9Q/yTx0rtlqc0saHx9oWJvSXFATC
fEGcmybiyjnrw5xdRYXiOkzFQI0sNtqs/ZUGeGYAcW8zaViSWco9oSGj+PQGYcBPW88jROuT8h4X
qOaReS7JiMDSPZM5+L6U6Z7II6Kq3MrOWcSFz5coJ/YRBR1EI9jcZk/VuBvS/Nynmu5HIhwntClv
vvcIs8iRv2/LGwS2NfEPVRrWfR6FlrNMbTG0n3A7LnT1xd+/f28bRzWCjGvE3261Dm12R/41/ZpS
7q+Z58Eq/kbI+iHG3baEn1j4AX67UYuiD5THODHOByWMu6/I2PvrP3twTrzFM325gJM6oawuuDci
VQRLHL95jJFcYTJDfVs6Y8lFg51EI5sBt9WjpbnRgarUL38fNCE3dFk6y+2/d6xCHmQQN9rgzJjw
V5ThCCeTXnlZHFNmt6gZmSJ6tqQprfIE30OExpBJta3S6M0BkAMVN1WKoYL0W0MGekasd9lq7l1Q
tc+N2OgY7bAvv049+1f5bIwzLGU4dL+prsdV1araTgSqwte4YKkmjj2rQsq4gczZDJOSguYsOa1r
E/i4+JYx7GUsn0urtULi1M0/7yFvLaND36bPMlFWC815DnowJVCAJPNZGU+vlPtzgYCt/iEIKl/d
+3J57qaQbcugDV/bfqSoSntcBchGsNP15kuSRl3blEhaKGBJS1c58/dhzS0NLvhlCrVMbrT1zxbQ
gEprAswNQq7YhetAAoqXTXYgHLmwU9gEQzUKfNOhx+rCPqhBX5S/G9Y6s4fOgsfWDOP3VwraZnQs
ctC4BtOv+1hwtW7/SWgDsn7EyDgp5dqCzk2aXBP4601PONnJKgNcq1u00Dvk/bgnt0HFNeC9Ou4r
8x8H32Fm6WomITXqw3a22hm6Cqd/uJhpTu4KDXHRdiZAGV3bMr9jpv+vKLCSFVp53Ph3zIQ2mUb7
1t097Pp/fmxS8U3WG3azGCD1hB95LzVy1a8ejrOEn8mgB0k+YSe0+Ft5cMVpKpfRf9GM5sBT451k
unUHwadQK19j7M9CeXrPPKHS8GvaHgGux7KdTxgLH+AJMJ7Wc0VNSjIHTqtS8NblrHkrr7g18gpz
knNeLqx+vEHLZ42Xl3NfzSKgwosaTE0Wq96BZ/7wMl84rdHSPXRZCMv5lDIW/P7x2e/ihIiAOwhG
93RlOjy/E2YwoNyG73BgmZcudonenxUggA/OPRSuNtpKs7eQwEFqVeu1MLYRK/ov1eWgl9XE/CU2
+hUwJx3ZoTuBGGGLcov6pKYQNNThpGrj4/FlVfrMw914CrJ181p5Ja7b02utVLjHvvWEY8YvUC1k
nYQIvwyiGr4Qeg5C6b7EDbOyk4aKb7vuYnxLzhSQXD4SAxLPUo1eHwfV5CzNpA4jYHn4ho9QK6Wy
hD6ayOJTCulukVqqdbn3dRNG8dxt7hpJVRMLGdsMYeBKHAxoN5elXlFxx1/FT0Nug4KIKiMfSs/Y
xNFq4u17kOAYM8aYLaQne3oq43hKqwHf+rqattLfOz/CoYCgDALwZd5Rlnvhm6dqvDW9VWWzneoX
fojigLfRpF+iceCGpcDNFaiXQhSL3Ryarc2Ewl3m/ta+Typ6hshZ78W1ABSXxJpUGsCVo+rCu2UB
U2Ptu36VrgW84otNAVhoypUbIGY9URf63f2pXiUKRMOxLQCaQYCgVEBPJDz5dnrmzfHzdKnxpAoH
AFuj8i+RCzT7C7yKR+BBYIBHYGuFQgj97xutDI9/JFz+bQNkaOCfCsHk6tI3nWt4+TPIGy8fGPoh
9wmjBt7NCbCQG7mbiYHPV5aaLvQYb9U26/6Oama2I4z55/vmejisU7gcDh3YxcoD1EOyYJLz3y8E
uYgTNAo+etN0aIHYD/GdHM2LOyGZsk3mHgUYM771fQp3zPet9Kxlvnkl42F8KXB0/B5hz9xgast0
LmKfXIla2BNGpQzMMSWjw7RtUqhativ34PRDNBgSd4rZPi/D4hWfqpI69SZ9U9yVOF2cJ+Ukif+j
9i+lA6WRmeYIwcJnUS7OXRg4pQ1XC6kA4SdCBySA1fAb1CgBTqHXcfjjfbs/oTBj6WyXLleW4jYf
dI0v85fF95LGbanC6QQ1ipl1pEkIkk7OXPc6SgiAMU7nXGNwBdwvMMuM+Dzj20XTFiK+oexkBO1I
pCitFBULiHaSmATJ05CHvpDT67W3KBhXaRShH0cFDD4KkSfwR4nIqzX8YzwwNTp4v6gQTtB9V0Jc
iwNX4psTwpZ8nyR6VT43VE9tWOA+TsVqp9cGtEHLsYncfmGwBXEvvChkvUhXKPB03yPIsMBe+YfF
CNjPi78W0vKgIdWvrtIXTNK8ToPnEBEJNlc+BSPaff/hCvvVf9VrsM+Zj+raJMLxQfFS1YAzgU8W
dFdIdPVmQpaYJ361n4w/2eMRelBkXIRm191G4VMNyA0nb/j3ECo3ssGaUrlm3wDjZNIhXV/f06z1
i94W9s6xj2nL9RPPWGT7gv418PuGClRipSNmyIZKu7TLBCTcb6scBIspZ+jlCyOsFD/GXqrG8Lbl
FA4FLqsdG5y395Q+pLGjX1dxioGdpOLUnnzUSKx36Zjg+Rg3QXowy7uUI23fMeNp+7wTalHFigbA
rFa4I3sj2HveS8722GPsC0Gn6M5jayh+ULLid3PCuEu50Pfc8OFqCzgLsccLDD2hF3EkBGqyaqJ/
jhAFs/Fx2UDHaIrojUwk47dA6oDqVrI0JEew4azrxhuAoL+EFioDD660SCqgq1nuhsWDDBRjFPDb
UHI076yhnA3DcdJn7FpyE6507T5Fu2jhas1kb/+DDur6B8p3A4cwoay0TM9Kb4LlFDxl2Kjy7pqY
U6F0BcBdDPV2K5nMkmt61Jbqk1QbSpMl4vm6CskIUoWfioRIlVw9UK7z0YkL8oOidzSvnHSRrVfY
eJDEGIIFDEADjQ1iuvn5kQFNAFnScTsulT2ej59/cdnvX5rGcGSBNnxqzMupv5a/qaVRq5iTMgK+
oJ4xcN2cLG3Xq7DMOijYgLGgUhxLOYvAfIyXWEPjCQcgoDQjSKHYGkdSe80S5gP+n/VZnXtB4s8U
JAdVtX4AFjnN29yoN82L0N5kZ2mCv2gDqZhMFutkZw56+/qmD/8u5gH/lyeO+C8BYxfMN66fFZ+t
rQeBC7ULYfU+vzHSoKsM2HGjDA6hJ1EaPm355AuwimcvGqWsfZdZ0PPf67tb2RgM+PcV773aBZNP
nYJ5J7SjJA1NRtCIc5cRMbRgt7n+EzdcbN4+JMEw5A9ugYKws6KQkWnqW/ukpPq8qBGhVMoTu+mO
NwX5se0c9FxlzKfv+rI34jm5TnviZHBVTti9w/IQyBjZVuRBlWYLKwbkwyQOO+nfuAsHr5vqGlGW
yISrJDNLSH9I4q0/3tOfaE0/lfsm36LyK584m3LqqJRagWl1Zp4Cru4OEZpQcsyKA+yMYIq+zr8p
caYUCQF1R/Kb1ektmhIDrC1RujynpzuWnJOZWXsHqhORZaUCM7IVE2H7ohIRxl9GLCUokdrAamPJ
hE8MrK1QfLz2IbYMglVGxzWcwe0fTtxuUA9wwFdZCOnMeB7gdsqBV/YCQ8/+Z9CV4GJFQRm9vjVO
1aiYmZNp4hh3SpFYhUaCwboMA0ttf65or4KL8xhJ2e6828AM8Kd/dc/DqKnRPQxNVcsplqQoIhMl
0KZIli1YDtO7LXXfL3r2a1eVl2AZRMN8TRQA9m6J/XCwZKMGFHzhwXY/Wz7n/CX6x5HumBnhAPvH
a+YzaRIkLgjTYekONP7rhlRHWisM3k9XAcAx+E1xZlA/CJSgqFVdYjzpvYg9oC2G3aYWVcoUWiM/
Nund6u8Y0ASO+n230pKX8wrdmYNO2Z7KJo0qBiHw5TCpM9FRUtD+3X7qWTjdCsrbHUByniCOHNK9
OP4qXXwokpx/a/x6wTXzOkGxpUg+D9S3FBltY8gBFJcZGX1/29+2QA30jWo3emGqplcs6y8npbLm
En3WlT27PI1sG41IFjhKw1idSLEnL61FKSd/mq0hMSuE7+TWGdSiC0RT9wDLGXvqmkwo+X4/w86p
CIljDaSnzVRdyRq6SC/Gkq8OjAHAMuOoLNhLv9yq19W96QaEmPfkDepkWpU6T0T0H8RAPIqilaJO
Y0gohub/R5TjbzNx3AOvsSzzflaHgaqsslzAdZkktXJxRGnKYxtDk8D+8Ksn23WM8k0yjKBVNJlE
ULc41vmoOQbpN0fyJA68d6SafDvCIre5W6bZwSz3y2gNK3LZNMrbu0BVZKQm1+ZZmFIz66MUgj1k
udS4RphDVZdRoH4sTkSZnjf6+ck2Ay8vH5ehNMP57WWMO+DrpwZCdkww+nuD77u+RqUqfByPo1r2
aZHwQ4Yk06VnKLCDfjQZUW/Cs3DGmewwsMdV7nivKgGb552LwwK+WFTMZO5lFce2zA7RizquAaD5
fw8aSpItGdk49HwvmUX74ADiV15K666fjO+1PIVeJ8OSdOI113JbdiPJ5xnJ0RQBFOPjSVuOhiYU
rO8u1KfOwX5CZ94GKpaW7xTUNLniq0anIgAz6yJiKa44SqVZKTUyldEnSw7y4Bv9kykrzl7eAylJ
Yn9vyi184XikuT0WBw97pAVHf7KCmK/RBG5wDM4lgnyf1MBsk1pqzHRnmXWtln3DRDHJfwtsOeMU
sBoMlStUT9L56JI5/sXmRs2WmdyijKLcSxQbXahHLxGNHTnbj8tByVa3+DFoAU368cJU0R7Qhdyy
5sCWWNLms+Ebz5nRdIkA79LjThALCeE319gwIaxfOXEbxhS3DZJ0DVUBmYYZTTAqsX+FWKxuIHzb
oZ8ugmtyhYj0HbjpEzXXr7XhVW6l6zwbkmoIQqDNDWEQjkQE9xyv4aMKQE39i4HNuRtLveBwlmOx
wPdKvBtMeiBCgZt8KDg4ZXy0W7iKUHwdRAovHX31YVG3nI9CQHD+15W0YAlnGdoRN6uncS5gY2D/
xYPMCaUseDoLr/nHrwWcpeJu+MTzjZiaJ1OGazCECmkQYkjFe8Fd5kiK4pocPrWL0qTcqXcD1XpT
IxlyCdZOcG0BiYebcIYsKCr5nhEWofbkNEu3Rfi3d718t0gZVtE4cweX3ghQLuHY/RrXg7UOtDM7
Sl4WrJdCFn0kBZ0G+Ve8zEjQKVlvnREFu74WATpey1cvI6jujBllijCr1uq3/NbZ7wnrBB9k+jr/
9hYLeaVjfMljJ7YdphL9pfb79lV0TBufJeg3ZjWWZSwSydOOTCL8Bawfo5Gc0F3gAatoVviyp92X
VzXi9EB62KpVAgAU3w2nKY8EGmJnamKTlo10PjaNKz6xVLNGVIw33rc7JI0SzdzzKo0neGO39WtP
BrVlXkRl8RTQ4OKxgEovsbPMieBeUR47EkH29DOCRV1e6JDDmdadZGrQgUeg8aXcrOIpM/xk6FDY
dzvdab4g6MBvn3DrOBXKQbqh46pFbEhTr+UVGUw85uT48QinJ9FvHqPLwbAMLKrOQnc8hYCO/l6w
3wUnoSuP4UXCATnqYCH2n55wKDqPtljDYimOBc1y0YbBPBbg0gcUgRgs7tVkzklXMdOvUcCq7FQT
mw8pzIPu3Yg3d/Xleaa4/D6noCyByuq5SRvjiVh/uVh9DJyXEou63ox3xvQwlqCaZaLKiaujrGX1
yBLG7BF+KWlKNdRovIVoPMKl8loI/ij0AJvZP5HwDlLC5alSIHHeBuN2iZ9EqyBGqcoKCMTTnXJ9
ZiGX3x5ias4tq43xu/0q1oFv2mBEq2DEQzBpDepv1hXLY8ayB2hJYLFZiFSd7hjtGAtc5jp4m2wi
vtMatYrHvXHVs0LReyv/AfKRIXYGwOiT7OYs6RVymn33wk/nFhdu5FqffWHtnDlbDMWhyXoZtxJ3
9X4Yvg3+B/3iRcRMPFPMaNbvN5lqQh9D4en1M/nE4pBw/i6HUhxA/Ay3JKD8hMr+7PwWMjDqhXvy
IwsQZJcDbZc6SLNQiDHrYXzcAcK3FDuv2V6Ubw3WizFqPrVJRMTgSfnu176Blx9+F6xOG/+rZ4dA
IJ9QjCtlDQl+vSS2wAzvCaeqthpHVBCETECzs3JS2AYy94y8310l/sBi/XySZ+/qiLVDxvLNsSzO
CStNkl5LFs2iMlXiE4UG2tfIcOGVoVR8OrNLsRZUKxn7TyL9BaT6EUiTxn5rNKcxqPthViXrHEOh
4bctmr1/XDNIDHvvPm6RJ8CqszGHPzSMGPe2s0flswSdGcoflGID+HKlMN8hahdjqj/S49nxYwpX
7P0hWkYaXfZHg8HjnqPbmXLtDZ2zAoRdjco6HmXR30pq93G+VFaAUoLCOcIVxw6iwF+dCZroXGy0
SSi1HBpftyjSR5Sb3sa3BwAjdoQQNtevPyvavjW1Q4tYzqSCdKEHd50ejmtdaaYA5kvOV/4Xr52Q
FUI+4rZjwFj9tLSZ3EE7MGwyWVKfJCrAoxwQm+UlzwJ947ihZEkSja0Tp8D5TclxcPxw5CFuHrxc
oyj8tWGAs96AAeUXpHax7oJmHUEyRHbmY7DyGkQlAX0CNDExuUfsSACfBqM2ZPEF5ggSaoV7ZFON
zIiU3OGYmZILjKanq//eiil/tP0/U9asGQXfeI0cghWMP4sv194XxuSqZnMRndoNHFVHnOqeViQl
4KXmQRQFraXk5vhuMXjvwDEzqtJyxBMPhPBfWqnK/aMUreOANUHZUOB2vKZn/16CUM/IHDTvXsmg
pdt0OgsKUbR1giSa26imS+ewATlXXlwLvmQVxZl1Nt/mJ5iayrLfh9cwAZEp8cAHGvlByknzZLCd
ubI6k0j8zN2r+HNXmk8zgotfJhrMi9Gu9y6i7KbpVNzTSiRh/n2aTxTIgbkTws4VwD0xvVg2xiFy
aKqsHqcGcw+lmRS0aXDSxaqf5Nl/8uZZAdvlUM/oGDE1bCkj20OOu3Blu8kXe4ago3eSksVphrLa
+GdeXjBl8K42vg24JvoGr5IB/8evGPGjeiL1slx8WDjCy9jIfOaZ294SWN0iIEQSB5sXnPJ9d/eK
wwqB3zNRETqXkHi7Yr/a+7juuEd1xNLS10gVz4MGuQcA4F5JNTFtT6UsTxDkNVIzerOZHac5udvy
2zMqFpO5E+giW4vSSZlNCswTSBSArWOFjmkpI29+ZfPaoC+9fshFbRK+kvm0WmUuq7AWYSeuJQbx
oUnXvjTR+4MKJEKH0deHMDCQX8Z0WygLgu/Hwb+6D/wNyWghWXJJfACxn64OeOr2NFSOm2e1WtQt
UHKL2pyy/t1ujLdLSzBj1kNky3Wq62TgHOR3mJI2G8InnnXs2nUqV7cjiJw1RASg9qcwXnz8/x5A
sAog86guKATiNJxI7edTVs0F9sVX4fx3/PXk7ODpn7rJS5gZN1YekeD5sQ1srxXSMVf6HhTunVa+
cXVJDYbbQjnUwOLZSTm8Mm7xQHR15X0SowXPhqSJ2yANxut3gatY6gMzN7nbx5AtRg4h1KvGisJg
yFFmhzpmp9C7vtYsmHOtEF1oe+VA6V5bujOkCbr8HCVb6Wil7zq5s1bae6RMFRHMf7WxXeHcH4R4
DsxWBRJ4T8eOXqKkUZEtUhr2oZDr2SnQz/ms0ylqFCuaN8uwnnHZp4Gq2FbsRb4vvrsMyiVEcq+w
eG18z/jy+QN2ydw8UQyWalYtX5fPxAuSk5BfmBopfkryWJPNzYJ+y9JZaJbc87Um7RSIj8m8GtpT
UqzazJ3FUZ9LG9o32T9Mjf6Wya9QTWMN+awUskfFZkZLgkIjJi9G0bu7ZvRgLZci805dkoR9b29p
m1/qiFoZe4VfQ3BWnQwQPedm6X9ldnUfu4+RCnCtOYbnmYPeOEHjG470hlLyHN+Rgi6GdbEhIgiC
EBrmvDzBiKDIpYqtj1jbA9jPKJzfl77CJ+IObKJxALjHeG5OUT/cOSO9TL1ty/JVV4hOcoDv8hhJ
ZBFEVzGth5UmQu5zOdwvAwyCQs061EphOqoa25U1so8WIAzDHMRZcuYfkvsTWmNMGae4zEv8FvnV
LeqPemnvWBYoD+r+W9/g08OrYPm8XHPlzxNOQCLxLxwLtgkWTruU2xEWmxFxl7x2UhuPSjaZ+PXE
7DdPGGM5IyMzr1BElK0D2NwwdZMbrbSnojgfTGC6jcjbZ8o8n4seB3s7TUAGQya1Q1Ca4AQmwdoP
P1u8pr2/8eIx6xJiScNhMIZjAxmDPhvfe3bQRgiaPxkYu93sqsM0iHwP22TOcDWNtk6BSpa0kgcd
zB36ImvZmG6ua4Ny3bg7WPgp2NWmyFbnHUx5NPIVXf54dXNJzABwkpgeZCxuE5kNkoomSVMcZ5ST
gX9gbgH8FxWsedE61Kf3elli8hXdn7/Zjeyhfff/CeRKE1YiUPwqkR+Zd+ZEubcDBa1x80OOMzET
HByooFyHvsdrcS6z9YRQrth2cyCdsTEcMpvlOabt6zbXNtnpq16dYXGM+alxPBZudX9yljPWX++G
oe7JuYSuoj2F1GN7hFYECFRfYSgSFv0xESTxR3kN4MBKcpJ7m6eLXHeuazLUtnxpNqjQteVToHFT
pRIxUp99UAGXztNd/FVrYY/jw46G8WzscpO8E1mzY7zjOB0o8LeC31GbXEysOMViA7B1ITrvnda/
ic/CGbMdh9GsOttC+MXt6XWHulGd2HZdv3StH5KEeZkVFEoMvMYKa6GiJNQea1K7yDPD/u/kX3kx
nrciISFPbTb2ffuYAg2G4+nHconXhg4siUFsIfg7bksw4jFKE+w7r/R5pMe9br5xHB9xAsb/BD2l
eUlC82xcFkOaQjFrljCsXAtTjoJx28K9Ymg+kPOCsPsm8FYyjV+4TfTpn17geEL9g6KviUtN6ziO
NppqGASM+96G3nsP3yhwIZBgMIWVtRlaNxAzPnaZ9kT9OaNP8gG0RhUTvZzov6VFAkUHW+UgXk38
3VIJI3TC4Ewy6VAJpy9AgC/6wKdDJ/CrlX9WH7vXVYlj8BtmLHDqRU6jviKB7t5S4yfwGT0BZLJg
VJtjFEPoYR9MJz5fOdQcBuMdWD26ItE049nppiixKRSSe2z9AqrPzZcbWLhUeXqBFMKikQsejeH5
MtwUAsQT/SzuZDP/PkkuXDhjOUHPEYXzsjwdhNqmuZzDWRKYYjD2p8thVxxLWvc1IYjzx7p9Qyj6
qtW/IdozAaEZO0TjASWE1dXpPzA86n8LvqQor7xdOd2JUOn7Esdyl6rd1zgAxp9PMhWbZv+bgtf+
PwadGl88JsBbp7il6BnVTtdX9JklrAU2ce0JaKnphUtVR979F6GGr1hnsuRl9iAC+E78OfHuP1kA
9qD4y/V4O7mWy9ctji/2HB+loUp+IyeJyCtSjGdMkSTVlEMFWoBA2l5TQvTyNQqQXgaKM3quz6kf
XBpyk+ymwKU/Bopf6giwlBjmg8O9iGWK2Sx831oq/u+YPaXTs8HTHoy0Bzcfw7dtGklP8W3IAdd+
JuL82phwSObsmnL4uQsc7k2ta2NQJo0TqLAmgFWX25oWrJpLQejjbNdhGyI+vLTGK6VQ/vYYHBgb
h1htpzjH/a4Z2UYpU85o6CJnHyC0iGS/WUUr720TUa5kv7MbyaD/n2DLEqBYvm5A/18h6MMnM6vX
YUQB4xZvZB0q0wn8P4seswNREvG/sl5yLUiHbnZYOG/Ci7UsxgJXx698gwoqx2I0DU79epsnikCw
7RlhajzsZ2YQfvB6dENHOi7DqXOAoc5STdqGnaURqT7IQUKuFxL4lwIBtNYuwNv3XTtQsKiabdTG
CurS/mecp1arSM4ZfkkZwyju/DYAL8+yr4NIcmYFj90a6n/Gam3z8l4oCNKclDTJ8gATBgjhYGvs
P6wDdkE2+WWzEU+kHXHYv0H+LC26PR7BnDuLWmaQRTDZNdKRxYsgFjsr2bvhBh8THRn+fmpbNXxU
CMOKG9ANwVArPoXKsh+4kbnlM1RHmZ2XpKe4910QBZRPnlpCkZtNGAOCY9J0LdU1d//BjMzzc6Rc
QjPHAfPPb1CEyWe1clfneitiNfZqMlwnVfBgtdOh1EE5jrqlolQaD/ST20vh9zG88+4UjCSp8y4P
XrPlpOguoVIu4anntQ0ZSgtTthBsCiCpmRNvia2tnIo0PPf0pubJake+YZGOr9Z50X0TLQmW2KZN
3UHM3yjuT833K6w7GybUk1ly/w9tONRI11pam4FPicUvm37UWBd9/qCQwe/RkrFMsYruJxIyKiDm
0gXpagpyBrEYQOHkDTyxouIJbWW54Of+Kbd9onssWrlKjbSL4AY87B7ssBPA561rIWJJ13QtKv9T
gT6RAEwaUva5T5NSd0zoj1RxPPEWpuEtOGzkKwqdL56UQklc00BUCLSKbA8LCDsEZ7z6GIMqQ0mD
AjwUcbVKaO5RUnR8du8EOVHQCbKCxtSUHhf69CV/rPKSaHTg1ETbcxn3eu96bX3y8cnxjrG+Va/N
Ahvsj8NElG8RiyrSeOBM+UfqvXGafLhY/5P6lxP/pqAbfEWSnQN3IVELwwzbUGHU7+0J4hT4v0wO
8rYipxOyunvqxwWC0FM7s7kcYqJJ9iUlZ2roaGPYJm5hSSD0kKi5DNB8xHX2vrULFrFlIVv06zE+
cCVjLzq7cXSnIKLRPJ5euyfp4AkDwLatl3eGTc4c9khduJ9yXUayzQmvtJAjeY1tQozoYbXMGQfx
+l4AJd37Sm1ELNTeEEAEKSa3TYQDo8ROdqQ9wmgz/A8PMMkwGaZx4GGg5CrO9cPYgNjZmNmxn3Cg
m1bTBrbg5Rq8TouEL8mgdQ7E+qMfcv9QfQSDcS110g6mPWXZSCSkEWQ5SQmcZBffY9d8cgeaveu0
3TZuNSF2gxlZ5JDAeWVIPXnCScbUkopFDx9XsSROkNTAKLzyxyOO73pc/5WSnhAGG/7fcFw9jRmn
w69j/yh1LghrRMU2gIOrz9AVWRXqhw8Ha1proc2dwSmVOsXkkMl1bOjTW0dlef1f5jN0Zex4fHLK
ojp8IKJtZhsCpIjb6hE2rVGJ3sfwGvFi5CDAjpsKL7KWRaUsbOrn9CEzP91VGCuQwOAQdeEXAWGW
0mk6WGME0JEh5ixkVDn86LVeOwnISpRuEjjuWJd1LuptGFwtGUT07RLj0pgc9CwIOfrH7wC6ftBT
BqiCnjIzPCTrFxNCSlrif6JN4URMsluQbv6XAB6nuHmaGH5b9DOtP2snnVUiWO8cgWHK15XWcMXk
8ltXV4+hUJPo04n6qzaVFZHiAH+mhkkB+FEUUk5zdcRiS2SaL6r4lzcAEIwlZ0ZbsNBZmRmJX/j6
lliCD7lSIlK5DCbmmmFdn6uj0PTSbph45BbRY6isAjsUBer7YiTm1ii/dkBN0oNjon6gA/rVpOop
NyA9n+NE/OEoyPA1bpxf5cz/A14X0z6u6C+bSvFt9JkRy2mtxxF7txWDMchC+R2v9somHp28D8LW
cN+nVQnpV57MYqxZR8yMTBkCTCpFQd5iLm7v+EuKb0srFJmp/BK4zkV+GTi4HjwkDPVKbl+fbpVM
iVvmEfB7RNxCw8gpsPF2AEvB5MedUOO5LAqKcNNkI5HRItkJDEdmGyfMCKBZ/X3nJqKejh8VDPMg
UN/fSZprNPZ6olErhkFenMiazTKlzsAImqtnrU91FJ0XMVf0TV23XyI2yScHfdCXM1H/Kq+JAeLA
AVpdhQQwrJoCKeWcWUx1y10P/tFov94dS35ALcwiCO8MO5ac9IocSjXOkVzfUO2Nl5QCQj5Da5c6
UakD1EETzxGgLVgQl/V04xX32rMphtoTT75OViHbLkXtJfzHMXq1mrsmNL2MqchirkXGCN+wK0sH
UjvRbjRFLrveGV/4cV8tZdgkkG5X1GMekXUAdPPqTdalQKmapCz/RvJ3L90RpxTij08+1H5SH2Fz
cF3pcp9SHW9sW7/CpIJP9zOaF9EQdP/HRSlNHAIG9nv34D1JVDL2AMlPKb736L0Fnq6Q8o72Y4dh
xfOzpcP/T483CdMfuqsaB7rwRQYHaYdBp3TH8MjaQ1IFJ3sHFcDJE0WEqNVkOZ58LCl8HuVLh8QO
WQ5snOyL0kFaQFTNCLd50LKMmerJYPtb6qLrYQFkCBbXtYcQqrC7R3tXl2sVwgApER822ZNNMAZE
tV/gp3MJonc+Y7eMgPcYvY0DqY+67qhG3fpfxCVFu6TxemTNqRxTS8m/zxDF2sQwUf9tu3LOXQ2t
upLYpuGX1Rx3IgKN3wAt8jqb7Jh+X59nkIth2j/2FWT29cgiB6hEVEGx0JCm0E/Nf3OtSR+Rtsho
rXp/VFGh5o1iG2vsq92rzebXivIATmSKg+lfI+wCP3EL2GGAc0002C+MwCM8gl6/3QSr+hqNXvEl
xELKNEfGFlF+77WEj08al8kUChPSALJs2NKYe2T6+88/wAghHeomANa1lfStU3FEujoui4znITxg
cyYn6Af8WNuD3uESppMRUtWOClzFPpffXOy03cvTgDNbRIhChKSoYk8/iGPgXmYAiPjeQdGd+mA8
1FzQK7IePAHpDmquCEmz1fNtY0+K9GdakJrammA2POz2pAGWNZIObSIC8opjiPdQlV5jDYsOtpDq
jcKl68DpCF9CHiNzSjwqrlDJ9bK0O54pCIqmRHwK5yABccQDtvHnqpzncpfgqHFybLD5xoTLXAKt
cjJEDQ4WSgIHA3e8mOLFZWiVWI9/Y3YYkBIBwf35IJynNGD28fIOIfp1DLoOLuzegpZeRXxUGNNW
UwuW1veU3oor0S7JYSJ5NmooyPJTf41jh1/KlBOA//inHfGl8/GXHiewtPzeHgzLe3ZC2u57wa6o
ZD2+bIQSiAqHo8xCrChZqtAI+zTpz9Mo4BSNc9eZ+s6ZqW6cmo6iUfcw/NqlM9H/yXc6aUmNFf60
eADDaryfA+VhMSrYEhTU9KH50GmE31cUWqpuWaI3eYANcGHA9T+aIxIYdNPHGwq7ueU/6NPJDBDj
ki4j1ki8WC+x0Q67B8YvltJ61eD11NcB1G70UIgPttuleaDTC4MFZx49INJN1iknJ3BDxwo6VcwU
Gzzjp+quam2uoVNh1CyM1lcHk2ZYT1x5PGy4kMC9sHKz3hXFYwxlcVI901IuMK5VG3I7Wsq44Nj8
f8rzmpRwEtHl1tsw5iePWR7kqr3oD2R9+eu9R1/J5E2utD/oiKANYgoTSfN7cqXskfUok3fPilEF
Uhvt3bXaAQTnCQgoluFac4+mvi7DBJ57Rw4upUPl/Nv/VCiFa56sW5YRj5UcdHOGCqCGZE6w5IMq
4iUaDQWQdc5392LJ6+FSBZ0bqKBUwzqaOzBTUQDEho/Bbx157oJz3v+HW/GQORXS3Whl2DwSaSem
8rNBpJDVFdwrd1mZMmxcJPYMVAs3qG+d+J6ifQP9HBEw3dgxZbzgNcRo1MTScc2THn0thbi6mECT
aJDM3pxqDdsO3OxBrA3y6KA/VoJK+FHkqwUeUnu1pf2rj7VnMGmPPESU0CLw8CO21q7DiRinQ/VC
rzF03hfWZzEHt6s5wNTssaNubwd9MGNC0QdQpbU7EQo7K4iEQnSGcEVkaDvxehicSv5BJcrGFfJM
1htb7WwWDAiFak+ysSzQdFPOsp4IT4ZGTvbbjE0eViJBxt85nRhvhytLfS7egTIRjrz5KjGjyv/Z
OkZ5pLFoeehsBbLqwG0dI9pcmKBcyp4JhoXkRucfpsoG4IFtx82UrTrfn+QKK/O3BFK4gsqqNhR9
AB3LZ9b5V2rNVWojp7Qq7PYvQEwrx6icxLdThv4XbgR9Bswq/e7FaFioclwmtMkNPQi+D/rQb/ZR
qsv3wS3zXMzZTLJCvL7Km2OYzKjUaZRlgzK3/MuaJb7wR5oTYl16nXl9cqYkfW338HCNVXCGCsCs
Ut3u7BtCT9uxIm4lR8W80KKWvo3hXSz19Fyemm97Q/ovTmltrNmpsvVMNUwvQLxK776tt3KY/X+Y
Myg1jwzDTo48QddwP8AF7VO0848atqVaH9rKU+0/A1vEzC+OIwcdCS9v/kPie8MWoiw3kwxD5iYq
bbckloA1Ejut3dLqm7oV3jODovU7YH1IzLFQvzXBozONdG7TKjVKiAg911gaBSE2hJis2oP/jOWi
cZWnWQlvELA2HC+FxwPn7Ws0vYMgCkx36NGOKBFeEkS2HdcnMbgze8ZFMs0NU94Ou6uopHG7xDVV
Xeh3mVzaxN8FKi/nKSJ+q/XB5/D7oJBbikY4KDjpb8I/u4XYmPC9m/KBp4OCpoiT6uoX9CpxD56Q
ZK/9qVtuoiTy5Xv2pjTytKofgh8v4XDHgzxkZdn2+kNgKTUtGpbyFyfXwRNLAi8xox2w0jjcSdGY
2yNHbtvCiKZ4gzo7J3LTbeaXcyYGsUi++Ly7SrwgoWu95lqXZYmcL2BT0MVMSEohqg4AsyrBO4fd
fiiwQnb6CaxOOrtU64/yXQjr5FLdfkF5ChEQdn+H5VrULdqrFlATetATduVoxGJ34pU+kEMFnA0c
f/WE3ACr6nEtKCUmuDN60CtgaDBWxPVmUubKpmkGuBSfu8esvwojJ4KlMPloRHKhUvhjtOxXzWfy
e8OaBoiDEf5HnqM7isiTRbdcIsupQesy/8gsKZqsha8hua3WgpUFP35spNxpBiipDamakTozdYPY
9eFGsRnycuN/Flr4eZiQAmpzpHrYCBky6jhk2L/vUSOrb4sAj5KokovztJjUuBygQG1ADToRcQ7T
FFWZX3gJt+JgWj3+aU7Z+Lwz5sBYzz2UX7/PPti64tWu3uRbY0eRu7B7jiwCASad9PwmA+VwuLm9
+HlV6vAT0v2D7cQXESNQZejrZe5yOZL3G64zZZyMz9rzhjXnC3rH3KBg6AtTyxvd0IELa26iWjkE
SiTEZ39vPTSUC6BGEKpWZeXfjMVKPBZBZT133SUmgVqzAbxrPMec6w5qsubNX/fqiPObjWc1uSyz
Yf2sELpfIgc/FnuyhsNWCXWAxkfrs9xySoHdRREQrgt390FkpG5so9Sf7HqbALnKNbeSy7Uhkn+P
TYWu3Y9B2/3ZfVWGP64i8TGdKLybVzgKHMHbShmB/SnWCjvS57+5gdx/1oRBlr/aJRWEb01uU7Ln
lelRldbqZsc6H1MfEReJEo3lB2OmqJqLiZ/1JMsuq1rvFYfd6W1gtnedxFs5CD+UeqjMOKkBuTvG
gsqNJfSddWoPxEsiW01l7Wj9gjTeZ+BVro6auui4QxIxihgFQhr2waH1j4MDNBOxECMI9dz/4SVH
osphhYn1jD+q7WqY9oSmqTivsNxoZb+/IcclLPE7GhH5baLnyXKLs5+cN7IyKwxKTxc39ebLeXfv
Wx0KSkvVXWpueKlsUY3tq+WDpIQtGBj2QFBkL+Xontni1xrBfDPk+9PrhAq3FzMx7tlsctEFMjBe
mNCEg6z4dMsAbG3fDe9wrfqlHRUcNOdxZrY0ijtzphGdVKN9jzo/12hnnVICINEs5nf+JUUaZwGZ
IwWIQbaFyM/7GAsLuPBGSFMXTm7M2XAfZtAbraomyQULUjW2soxW/FL9EYR6KaybVG8cCFtb0pN/
inhl/8dXydrIm/DXMrJDlYZbXN5UOT91v6CJacEe80Vj57Avfe8O2Ud+OB+D3NHHKeXVag6e63NU
dQLTC9/ZROXflNYMRruaUMCJgRPJDO6uCte38iuIEd7Vyib00ok5RvK/1PWulvgMIQ5kTPMY/Zsn
xM+n9Xke2U/GHx58Z0Ft86uAmvyaq4okwDcQCuNlLY0hYx+mKjwGlg7mA49cXQ9YJ1L+sE68ABIK
DPnkKV9hdUg8dUywgnkfV7Mm3I6m+isE+TheG/g6Fblj2SdzObZ/ohD6+TqeOry+g+S8U8h75p4Y
7aVnlbJ4xM0E4AxkW4Qb0wtVGWYGKQzwgJqKN7pKqtmrdJNB6m8+CJ8Om0vRSjo6lizdQ6jTzZrU
FXmyHQFGRl0wqqId3xLzqKsgQ9C3kI2yv0DKOs53/B1kwuypcWWOVBO+2urUvBCyyWW0MwPyn9Fo
Bx2iM8W7jzs8Hu3KKPUaehpaFNlx2RYXulEFYIV0S0igg+96jRazIPGhtt7rvtNkLAhg0wrkQr2J
AO+EtisYZx7V3dS+aS6jV4uac3XrxeDTn4DFqIL/dkOIQHuFT4P4ljFb4Qcobg8nnUXqwhaQMLuw
gxp8dSjnlfL1S5rMvU1st+1jVmB9kyfPO4s1KUXGDdEKS0GF1LWBCKK+LN3LNZ6tdMZwj9yRvDWc
M/w3nEjLcUMC3eR16w8lUPgaP164RBemh4d2uH0azBOmJbOttr0y5En0N7xzJ7OEkza8Lo/XG8Z0
Y3S7t2eww3MvD7RbpAR5HDsQjWm4ofYm4ZWqCnP8fd+uKNce45YKhsastdBO5eJkeoshvvcSjdXw
Lw7ZMBYq7b6qq+yd8NC8Y5eXh9e/CflI7npLxrs3YI+UzwxogpJDKS1whmgzb4KIb9dlnVg6tDyK
hIR7df0CplRqb6c3Pq0KED4jonSR9TZeHaFnc7nqvPe5WoX3sA0USo8J+cDLiWac+TC/a/d0u0HV
wb5BMBL1Z10pPY4K5F8yd2UqUz1PSNSKXk6qKsgXfz0hr95ekSjFFC1b8A7GYpCYoA7fd70ADQR/
qSgkvYve9zl8+CwkJiAl5m7LspkF086xxF6VgDcxc8Zj1L9htbVARbL/laDEd3sUwkv+tvUxycBa
OyeY4DVuy/mDXZ0Rhch5I8kNsc5gu1SLa0YzVxcOHZr+Goqm6mu/HR20RyL22j/mdpr4YiOOxBJG
d0yHhsSwheDdWNtC8GoO+Ds/2mGOFvdwIoigrMuKakcrzG1STAKtfc3hUmHzfEgKy9lnxc7zktVV
wQ6HHYma96J/lZMqzFs5sAdP1UREk75SSiY/xIbBuVYHlUm0qjERLkKdTMa7lkq1pAf7XvcjBgMb
KdzbkQLi4liRQoc+FconZqPboTlBShya9Se+NEmznbSQ84hACqSah9WurijJJTkrcWe/OXH0Uw6O
G0DoemJrL2lK4f7i5Ac0KwTaVx7gtMr/f5zd+tvqZYM+DcmoKrNldgae6y1G+r/RRb9JhmNfsvkJ
ZQVdcQDHIAAyxh9pt0LgpVfwp/yubVw846OUQbUYtJ+dtGCLSSRxlogrwkE7/4swlziCOpx0Inu2
eug1ndRWXrQrVQPzWzUHGEK2v/7XHwTd1UMChkaTYrPBom/cSEsN5GJQb5i4whBJ/1aWaxpErCER
EYL/Gw6HOTk6eH4Uzsuo3YTWErGXqR4KEMBFdJhOHeyBXs92zlxyUJ4PAkKv49+yPONv/kBkuz3o
FdCk/uqbQOkqGHPzR36Z6DIRPxCyIPo6yXLl0OxBuiByFtV9zUbcS8CsSYjH9343yHlXZT0+0tRC
xraoiOZ5idBDG9YnV0KPylYjllpJdrXnMhDFb8qmAgTstpyxboCLVRQ1eVnoM9RviqOnD9DpzMsv
fiJ60mON3j0QDNiMLMIlSOviOdTd4vrxsPSQMIGrrHah5t8ccRtHxBDUgczrukZygK+ChpPHxiyM
e1vGNb85El/j1leI3ziAj7e5X07YsFtXuCKbG92vfdLVtzdb1GAbT8BAGgVoJGHd8DWFZmjRARy6
M3/b8R6UmXe6fp049Tj8+aqOo9qM6FMNSd4Ns1HRj1mn/du42dn8k8+g7ukgExxndOMKy+whrcR1
jsup7yJj695kziTcfnmoc+N8rH3gJb8/bziC1KLiHr2AS7PvdYsWeSga3L7RhKFtFzAKZLbDzvL9
bmJZA1oSHQZ+ydt15bck9tAHv3DelpggM8rZvUTBSJSnTnctCoEhw2Y9jIAy5ADD5WjJKRnnxnXf
WQcUzEXUHdDOu/NPLCiS1QHlZoJ4G7Ff+Wdhw4eeKUMenehPJ/7YQgS2Tz+c4ukS/YjfE6piov5n
M3Yt84bNu0Hk2h+B4BmUov9eqHGDxBPN7NT4cHfvn+aKQ1S32FK/Z/LwpVrmcckwzs/UaPeAGY5A
SDYl1kf+p14ALDDj8aYn3zXL1bb2YqhUPSY48xJoNf9OLMezUmVIVMiCos5TKv4y2W1wkGxyD2Zs
Ede0YBTmB95BVRfFd/OZ05trknszu4IBqzUhzr6nFyzW4zLvyOwRGRodJNyfI5x+235drpm1iz2/
0w93QxQ/QJ5AfSUR4ctlblQbPc0W0RJ05mCCFQuzBMtEFdbXh86+qxFTS/vBBE5ef3V489MSaVHv
0xJq/qVPI4yIWLuLyZmxFlnFuPGrVMwOP5PcdHA0KdMi0s7aRqJswdytg/vZNZBcCD/aHp/X2ucR
7un8nvBBnbBvbVFSAXC8YTxldmFbVcx/pNQg5h56liUJAstPYrrel35/IosEr4oakkhRH19H8Bkx
RM18g//Ad5iNoVvVftCcGQCpHsx5vcuXwQMEwCo0ZReBHxP27izpQcdrQt9XONABkid+BNYHQrge
Py88e+9QpqbKG550w4SFZVstONaW4UCgO+2jRHDTjebpYaZ1dqkAoVyI5M38ixVC9mAcv2h2BKl+
/JX5cr0j6POmsi9uNLTrPq6SpBeB2ZYMBGEHB3GfHWc00n6e4sgUI4gbhawmOWnrskjnxZUqc7N5
l51q4xbT0h9lFRYh15rW/tLl5zkw7sJn3bPrgqB8vb/95A+q6CcKn4KddF7yRbZUd9L7v1XwYFBI
1EJ4PdRS9TKWEEt1Pmr8cxOV5MFLArJ7ryksRZfHpEchszXawmlcg61ANzQ0F/Axfhhxxg1d0haM
hf49EBGgeXK64p7iCV8jblBKu8bm+LFouPRLEK+CNXY7AMJ1CdRH8kVbKasbHV8hKlN5nW9tOqLA
Sr9emxmngeEB0XvFeA2hpvPqEpaPzCe3f3ygMjTHnFqnBAfD4fWaCqjVsX7E3rkLwFpoeRPuZnL5
lh9v7xHyEqTFQfIbeUG3jnOAAOLIsDTdtR+W5c0ypy+8Rm5kBlaLSsQfoSye2KfT1TG/be3OrYVC
ka3xd5MLI6zT/8TEXgrSHwLJAZWJGkKJFqbplMvy2NeJeK9emEwpy/uSv5Bd/M/GW6jEhP2MufhO
4R8gwoMTX35jWy64tD3I3oui2aiYrS52ffdpCVO+irZi7fNpBLIvy+HfGWBQOHHHrYWPbP0aOQvl
zH8R0X7MYnqBJGuOY214r8y3VQhXxPaOHFv3Hdcc/kbhG2YLbS0LQaYLO+Ip6A3b7wgiNcsTr40b
bWFxYt9ZoZ+uhb/QAX/vYPvRDOC93Vv2SdR8TwwZMzEtNaqDZH+NY6BoikNou/IHNJxM0GqgtYCk
EnF5SEopsB+6GnZjqmY2uKd16UaNjPiBiyckwS9NW0bfZzGaadRpSzEFCrhDJyGOTwsg7x2ZcjZO
NO96ZvwqzdWuAI5WWXtch80oPbUUQQBAKuNbERJyupBDDgJkvza8OdCYZF8FbC51lAI+BMrm9k+V
4YGJctn9qBukq8HoWY5VxloSx99OK2G5gHubyj9gZtsNHCbEw+SDhew3fNua0la6a5SxTaLMxFD+
5JZYn7POXEpDNT/iXxHzIvQFhKQ+IOa2JmNSyi4qJT/rVAaB8+NIy0J/Zc3sWZhYFYrXEQdZX81G
WkfXiRqkHGQTaHImSvMCdcFaI4CLDKOxbJWqoTaLxmI81gbmzl23Xi0IZB15HHdd1EBIgFnZhRlo
k8QUfSX2NTel9SgulYtZ7O4C4R/N2S99ipVMgMZfL/zFb82ufdm8g7aQXPLab3cprMFvkTjlwHxd
YzLBGEVy3G2ATcriqH9ReAXQ3FwnHmaYARq70ZKIL8H6TQWSdPnOEfXeDQp1GHHKsXobwIBD+5L4
bcLJbkIDEC6F2R3BiU4wiLJT01DN7RCuUwd1Noz6j3v13JOndr1mQKPD/h1DNhh018OV2Ly5iVF/
NFl3mCubJ4XRj238bOudBovehz5FMvipPQJGCMOPW8zvGd29fotE259hA4KAsrqpjRFvVWWZqa3v
KVMukqpe/BS0/HtEnoDnOM8w68X9aaLDoR9c0QRZrX0brAyPnChaU9csvd11JH1Tz5td7Z2LnB4L
Vb6lFp2bH66TIGHXX1OlQEupLflDGPSXN+4RClXS8th+oBeRUdi4pBV0ESJzwlBBxCjGH9CI/Ahz
9AZ4cHDUuyFNDfwd8AXFOoGVQYYa6Urh5ERsOhrsMIQLYYfUQgmRyvyzGoia2KG+n/89LwKB1pc4
kPK4gGF1DEsdtyzVfo1McLDN55TkLl/iOr0VNPQWy/HciB3R1q0odYguDZ19j9U9o09cD1bjYg6S
mG3d3jjwC14TYnMvZp0ug6viAqyqtbLGz56cxOF4x7nsXMUmrtZ0a62G3sKncbsx/HgmChf4PzBf
hmxuNgFu0CAgUJ9+SJQ1l4HUq7GGXE0FhmcaMOVMkdDz4Ki1X4XqWeBVLL2a2fUWHFXIhb04xRmv
sboDGLwyeX3OJd1NBdoCLRE6URsPw17MElb/T1alA7sleYRRlmOPYaMJnel/JeVMMPH4bPzHWxq3
5J7DiTRtLTyi7Dewx/dIWFrikXxAdEgU3Idxk917scqv2BPv9VTs9IaPQudQcYIFOjDLdq7PLRjh
X5kj8a4weOwf2V/u9dHmEFcldjzeEGb3UK8k7e383cKNxzp0KjtIoLCKout3305CYUd0/YV9edWz
Wi1cB1kXiVmbfKKMPrr0LQOhvy25jjC+d5Xp8s30qbUr1z1aHWYuc80tWTtY5AF77MIEyXzPgThE
UHQjETtx/GQWF2DTJ+LvG5myKoQeJDDJNkDnUDmfuw5d22Ak6Mydcu36WZeFFD+mPZyY0VcX5S7E
2tcugAl/7TAPDkM5WtYsaDvDWk4x7MW9/UaSmefswsRrlrCvxbc/weO1P+md1P5Dlg0o2fe5LUPe
VnUUS6AvexxettP5yHvwGh30UQdYZT7526jm0VhrbCF/iLAmYBlHmucuPqaVWSiwBkD5IvU7FsLI
p85nBjkTjhDgkgS/agz+7iWIZn2UxtMXgmgUNOFbJIkdiGpuWIIZzzUvbu+g2IqNMBEkHmt99bpI
qHJk8wT2hm0NrSG8VFmMFXMqKGTR6MofUsjjFt72gO1slu9e858QpnjmMsvwxSdpGcAnQ3h3SSr3
ND3Wq06HjzWZvL58qGqx0n9okyvAK9bvDwCHKznvz53MzJHQh+X4z9EcZJewmRSv69z2Myy/2hfz
anSDdZ4L1KXgFSP7Lsd1OOrfROEzmrnQ2MuxPW8dbzo2XpRgVUydO+4575ZgmYMMlb8RrZpjJKRh
DgdwzU9YrOw5TAVfaOMm+blFLLbZcwUvZJYWXCo1Aea0XGE65xdMRoe6yF+iO2LW8ogMSQ6UhZVq
2BjgZogWxPSzf+YJVRiDn1E/QsihAORgcu7pKN7MgAOOYXA8Ceyphr+jnbZ0A4KEmMe59X0gFR8t
YR79IR6Aue6c2S0kWTEJ5kkV0TuQUJRbib69guLMb8TArGK/HBWDhwgCYJxL32pS11rNmeSJ80ax
jFsrqRJwR4dOvVsUjcaMx5sR398taLanofHowWhmWk/rkeZyUl8dxj81rricNztf17tRtirabvdJ
Rd9eO52wNBUHgHw8lMfkgF6kTrD1KUtSBxuz0lOPYu4QVBHDlIAAiDY0M/rvneuWBecB4MAhRCwj
gR1YwwabVDujq9nfzl1i+qbP2Xl59tNrrFVhwoBbnMCV7fyP9Z4TyuCqvTIDpnCiJjBjTbJg+716
ZfxVZjWAquvnEMvtRuB/Y9W+JK+GpEFsc2ki6Xjg/irsE1ybKy5thHaK/Q/I9/25S9xYQWv8nL6h
RkkwpHMDqNZP6FfMHqxspgOgcZh7ky4JbyBgxXfansdXI5gFsn/VcqfiIOugTUKITtY11zZ85hjf
/ng0B14ZXMfkIcejz/ZqzsmV4nfjgqdGyjdjhOX6+NMC21iI1k/WNqa5cts3+KsV60ogaOO2hNeU
j04B5qmGp4QJ1ddD8k2z1HAx0grm3AFQAadIvKT5AwFQiMZLqU1uJ0fi3/r0kcTn+UZvnzM5Jd+k
dVKEfqNgRFGcIaEqam1HnWbJ4sQkvKu2WUU0CdtkAzLd1pT/eFpGiiGR+jS60zao3nIhSDq6siYO
4P+KiYhn59X3JjCIeQmO5nDQz6XU++tafksuQvb2rl5BzG/kfhiEOdbypQTsrWesiKfC5a9zqRZk
m2AYgvUCOJix8ceYL2JjLHggB8SaWkmINCr0hGWR17muzs9h1DA4J08WXcCMq7y1vjNGqRaPkt/S
XNx42b1L4Rfpae3/Vj7w+fI0awugfa2HDR/1xlMYU4EpOYYvY2BRM1gXshXGRW6SCuNAn14t089F
j1cAU4eLrYmqiBFTGkdUY0dhQCO38vfqJMel6I4Gc8Id9k19bS8q1hMWP151Gzi/GvXDuEt4BCZZ
4Jy7Hms34AXK/tRt2kmU8ebXWafkWWWsIKSzRqwLeDDE6myqjI4zHoNknxZkcKxnb7Xbxt3VqyT7
qt6N9hklOZfdcxlxXKfMVJchdiCgmUnB6baxc8hDCRclN0SJ2jZtwWi3CMQQ8kD2FcC80VPrVZ2Z
QBKQCizqeKmUJYT9LLDIUqHWeqZ47Tu3t25ODe1/UtLgqRpHilyCtFcKHgZlZW3ZfbdFzny3Ohm0
X8KgylDs7bvr3hMOUZ82QqbJ/UUvW76cFZfPYmH2wQj2aDjKDyY4VVJl9VLjDOy4NmRjwLE62QDc
Chx/rW9V5csHv06xZm+bTJaJT1PvwTpg7nPJrQQRhjBUfgMDSkpM+5PpEKyXXHigXDHqmAdWerHB
EF7nkNE/jDAFT0/6zfrxqK4oC0gxLIXU0472kFrooLYLl6NvdUeFcrO3Mq1O5RsaL9/6wioFOr0b
Fy1xe+zrCsV7wRE2B5RT0sYEwKvLoMOUZzL4DA26VINviFJkitWktywsoyQ0UWUlepgHgDaiIQtk
p3Fzny2oZ58b4agiUWe0uzdhcJo3aUvjRXEPJgF6fBf0tm2OT9f8qVdkG8AsrQhd+wHN2L6gn+xv
vnPti++3D6qOn9cpDwjchigePZJzHQzNypVgNZePigjgbTT4vKIcdGDRedCRDYbl20S7VtHiKWYx
tFa8Wb2lN8oLTvadqIKAlU1U3ItgSIu2rcwyeTEEo1NpBBcfqbFd19GIb9g9QltrB3rYb018l2bd
uwfgtAIhLMG5ef9QPmlBeInTNTg2g3Bnm7LWn4wsXVQ5WoX28TkJ58UPk5oLKosI6tD2BSQXUM2a
aWU6YnDCyXkC7rFqOhQz+ESg3Vq3Iw8Gaj4sb1djbAnZtxy+120WdDNiibRacgJhxGOZilbhS2VE
85KSCmHLqnnNrAGHBwE2kivISsz3kSt5ydZIvWC1ZUj5a6Ay8Aetpwlahsue0dvS6MPv5GKlkrEe
9PcnmkLCOml2P5ETz4+ZA2b14mSmPg1Rj/uXU8+BrNcb+hkphFk+t9O3pN1loLymus9jCpd90+BQ
aJQKwIZcFSHHVX8zD1lMXQPx/AdxlMOyH92xUqryL0rHx3r+Mk9HAtftnVIjTYUr9+gU2lnjF4GR
ApGTU7aYZGaUVxJWACSwB2vXeslSnyQCp08ViG4oWrHBBKmLXn1m2CJ3BONEUCibetqEvnsAJjPw
yScjJtVqjhmKOqnD2y/I7z3kh0YEexkrdNQi2d0kYXiBH4/epKzSDWNgg9qmi7QNDkb/5rJXRT1w
zY03JiwAKauZzl8x4CPPT9kF2aMv+cNMCwAbNh0/5CJlWZswQFW3Dk/kpPdENvkADwfcmTy67gLG
Fr4mav1YimKOy6qTiP1DR91KqfAMN5GEQeFtq/aOGudW0uSHLK8evz2KVp5dM7jyS8MYXRkFGcn0
bLQd1J6OoGDp9OwXkdQxznFOe8uD7KyHt5ucqCC+hbSEa5vaUljxU0IqDRGQ9z+U6JIN9T8k3Etz
cahn87Qf+ddCq/6VUqySMc4xD2+zxP+2zGuoOTi+ihH9alH7+tk3+GFF14eKVtHhoUHqeCmvLV2+
6Unwdy/maYBf920fNm+bJyJfGZrz0r5ROO8Zke0liUZB4txMYHOaIRewxU7FLGe8hZAGXzavFGLF
7W9wF4tSjQ/R67LJtg5uCMgCZ6hdy7Q0Sc4FC5MK/yOGpupG7Rm92UZgf+bCsXx/Pj3LtVeDURBB
+SvMbq2nvjcxmbfrFKGCKIKYZeinf9DTJi5Y/Otmt3eeRUH3JLCDM8hnu6az+e89+P5TIKk46odp
0e3WK1bZfE4e4WQEHZ9E9bhk9ngkr4H4HatNtW+mipLmUFAZPa84Zuas4R1UzIfIBBcMqf9U3kP+
boIEANG2qEzTe24Ib5E6yn76+yBhDy5q9EOWV1K5VIVXg4ylApo/G9ZgKVmLf21gFabYXqpN4vTA
wTW5ZgQXeaoN/Oc71IiIyNI9LPtOZI6HgVt7Y4tCqWhwj7/WkH1ys7pfzENXF0Lm0OcNn7hijK3z
RJ3jBvrTga61QwUAy9udlOOjr0W9RgDA/PfDe5CItXq1ZPQqSUbtrQkgldC5kktRWgzwa4McYLaW
BzNK99jUUJsbFAKnaeMlDY41NGLSh/DRvtYL392LXXGfJwUHfzcU1aA8fmBw1zHmZYRlq0OD3ASn
4DbXwruap1KP2iydXaUPX9Grz9s6My+/VFaTCvqCGB4gjkyAYhF0IU11tWfna+K9LWZWpc4LEhQ9
lkA1WuwV/nN7+pVXKYZDvE42ouS7J/kV9EMhSDVSAvJPUi0pQbUbaYE5A8cyD+FSyGuy5CyKvprT
54hcXP782zM7qFZlNDK0ArtRjB1Ph6vvOKYZrLFkQ6/Wrw8RxBV39U00WUMkqgFqZrYx1u2QIt6u
Z05qkqK5ztigrPpwR1Y86Q+0NA05lf+FKkbtOBNdZYik4BmMkrEn0b85ofeeshEG4Yjz1Bu4e0at
S+tsQc1FuMP7+ixe5t5ifKtJ2S0CwJE6oXnEY4lG6PQ8hwvX4b0AF2nswqQTwSSYoJGjJQQS5CbI
FmfUAUGg/lRLfCyUGwVFou7tA7jjJXOi5Vo4K0BobI5MGpIHEe3DgcGR7QEoVwMK5KzB3c2VswWk
RTekLRaQ58XNWt15Ub532fhRN1X7oqaEgimo0b+o23OdQnMd/ke03ISyMrfnE5Nvnfsx6XQVxzlL
sm18BIG814XmLHZV7PGWe51myi6QpouOCs+nwNMJK9tfWUJVCaZbmxwfXiS46F2bqRLtF/l7rrx2
ZCR7uW4DEHjT+bHhnLS4ehy+sf2Mf/x7YyxJi24LaOQgwIx2+jDE4tOZsna00YZyFqgZa7kCcdUA
5XjusrOL7c/epU+gQnJI6+qnMwUSsCPsATiRE7Rkuk7KLSLI0U0mb8eFRiUxEHF7UB70GOKMJKux
uSAH0Z9kS1DF4sC3JROT7+79Vyzo711dPNmZcyj0Q5d+TrzkRDoaHloaQCH3UZYEKohYXgAQceBm
BYNu+GZO/5Afs0XPYm6Opg+A0W8YEgi6LwdHDRW3ANgLy/JUiwN2qLy6+L6O+nknpTnkQsAfGXUd
25MnEIq492W6TDT0xpx1VFBm8+pvuLHGJc2Ys76XdD85N5g+q8bW9RenhKEtW1FFwKwIpD5lPSOb
TRPiBfBGjHriljNpbG1TC5msD1wOdsyGgP69rDqoiNEuCYgOGmupW96nrcxdMxqlMydUcoSoAHPv
KI4SV17sNAq9Q06SNUILjvwV9Gh5bdB5Xhxxg15e3Sx1bkrShWGIg/sliu5Xm4Zx9yisZ92XTqI7
oKAuUzSknPEINY9TUlsCXhEKivm9CCQaNPl5CnvPhAXyTDVYcBBuXVkFITLEBKmxI1cc34wgmVY5
heuieCjNX8GBX8oqZuEETgMwnIhHCPv4dJIpL1Gm8QjPpJlfBoBIlwIihtU4BV1Ty6PLbzGwH2io
nU6QMsaClx1Tr8tZzJIWnz1Heqs61/E3DpG2DnaHA02M2AazJg+DbrOAvuNH0Uot5X2oPbwuAPBK
mcis1O8y9gsVg1GAMSOGSQ7W4RDU1DKwdfaPxFBZ0NVMzWtU/O4UXRYJr5MTuo+rSOLPN9DtKwYb
ksb8/kMpC+C56mylB4IQ0hkVibJaEZMMx5dfzn6Ae9hYlr0AtpD1lNTUZHZcLTnZU9O4hf0D/zDc
XvArZtBuqgkPsYyGBDgyOQ5hrktuIoxLnOltHmQJbSNa6P3iV/ALrZOSqZ0+n+ar4d/e15GQuhLU
xR4P5te0nT22a9Erj0LLpU8IOWeY3XuVdRZQdH97/Wt2gSKvK/D44XHNBlaBUKtA/AnOUv2T+Vib
CnHraX6Nr4pZBfQdCF/n/HuO+bCbNqM3BPv43wXNDOTiCqUDaVP4uKbMHiNbCNKNdgc1NKPnWb9H
BdW3nje/sfzycpYOUqlI0AOnR4RStpiNeLP0nimO2vxuHXj0JuzLVvS5AV5xr1EtEYMZkbpgsm5L
JtkLAzQ5R6TI96BlkrJ/Nmv1n5JFqi1Pgy3ISw2hfm3iM1/5e1htbTYHY/VhwXPDDegSDhVYLJ52
wiOtCz2Ic7iMHTnrag/JhWREH3jltrZKnrT8V+Wlw5ODR45susJ5DpvMsByiGTDhzK9rNxGZHb2A
+dF6iziBjO2uGQabJkgkbtbWsW7y9ZjDK9SilZvlBuwWQOdVFmMpEfD2C5EMB4Fcuzo+lXAkAKZQ
ThJsUELG38jMgSfayFhGryedwY6LEj8Op/geCqjUhZnePRAHrKXepUk0XbJdGJf7PD2MPq3/veuB
vN3nrzKGHy7UUjfHZXzw5fcmOq/DyrIzbf80ZYf/EaMuslFgHW+V2pg4eS8wpnIiIJimg6vs38eK
jwBQ6cFjkcb5cftE20SUbi6V/HTXaVo+aBIQ0du7TaxBqGqjUdoMBz3Z89buVaoR4il/MhnNkqG+
EDdCLbtaTG5ZUiH1H5Iun5DPknSq7vPKLO2gi365BBXMZR7gfTrLQOHikddz81XPXSqaVt0Bu8cT
mTgNvvIJVbDsOhyVNElXQxi9IsnW+43mTG5DXSlZ8WtJfvHs1L1ToDtrGeSuhH/dxCUwDnjDYiSg
BbVqQh2J6QQLIkK0x9U7saVPb+8sXrUK5xDSAHBBnG+c4Hn/za3bHTGcfL1rK2CCwWt/Ow/hmf0i
rUT76pYK91HMPyQ7Gc4epLLMRS2u8XjCsyIeNWFAelGVqMqeqWMoPZhSOGWmx4PIwCqHK1Ym6YbN
PmNoMy+Ci8k+SwmJ30eW34i0UmSaFfuh14Qz4idpHowoHycbc/88/0fX2mCiRU3WufnkpRes/FO3
AsPMq2wzJSyDWDLctB3nYOKXYVNJVet+bTXNcfoAnAODDyj0Vhdunz+Y4Nwp6u4abzMTZa0l1LXC
V2/D32yHgBH6Ml7dSFTEzvpgGxwjRvJerEqfGHrkO8e47galNWTcdmQ7MwvEfKqxButnlgLGvUTf
0BOa1yNZIZKrLP3yrMaM5Dsqomx1TfZrOFx9kiYPR7yiTZlfndncf3EN54e3uexmmY0xxi+7nJft
U3X8+BZ8h3CT9kdFGxI/qAE2PRAMFhC3bCkXiygKH4eT4rKPlLSCdlnrECbc18WjHV382i2MYAT6
Gs7BwnRgerWbtsFOcWcFEt76uhYFcKcHPhUc73i93Vl7ourZ6MxludX2IttcCqoBiwPyH59mQuPR
ytpH7HfR0uSNQufCtppp4XBjOKRZ15kAUKgj3XZScEWhY2+nON5h9e0VeZf8gsG2//Ld8y9CFY13
PNBfa/fs2T8g/6x9Z3FIwtxgSwns9da2/fQaI9mdBA3MeBo1dlXmt/7m6dk3kxa9Gl5q5tt+fvkM
FI0QRxcjlQg6O+QhwbmW7VArBR0MymGAhPN9Ku0SnlenRNBTPtrGINGKNQrPTo1pUzOhVePot6Eu
s23oLtD/EU5hvppMPP95nXfULkILyR4o5oOlf+lHJkzL3j3L3GBez0XMQ2Qt1qwVOe5Z6LKCxTYP
BZ4Qinp9Ufd6NSaYgsQtOVPyl8x5Bebgx5pMLzfVu5at+zf+e3YXH0TbH3uyRPmwWsG4rTkLP93a
8pJ85mooP3V2Fm/dhcT8Txxik/nvvsNZrKbmxugWOd1UhOqlTc2DEjtp9JXvVYcLjR8yR4s0S7jU
k2k/mpshh4FNQsk72RuzYAzPKZnlIijcThrWygLojsq3WbZmh+GQmHgZCz0hEGWmtnyZbVnfv4ed
bchg5ULQUFpoNyghcnCcsYn6aGnWaf4shB/A/kv6l0ue17gG+lGz/Q6KdHiVRa4sHvkmwVrQAnuN
55uLV3Rx1JUzPMUtPA+2zNe66Gpia2x6EB7HtLJi4BTtAQQdYpNht/C8EpVsXun6Ilw+muQ2Ihyx
/kdstPKp4XUxlRV9BF7nWcBcEMQzWizbdTZjPIbvodDn9ysRUfszWbZj3tfYdVLAZ3siqTDyQibq
A/MKSaQqyWWPvzkDWpUViwiWNkG5qsgpshtfh5eq7haeMrl3RJ/Cf5+/R3LKGcA4K78VkdzXGfXY
12P05Ce45oBNvwHT0t1mXMVZXcX8Dw2EKdwJ9wd2wiRHYBwF+4l/Gule1t2v0+M/hsKVcuGf4mQv
Il7eewKWWzWR5f2Cr/ym4OUnX8ju/S5dJ3/QgxaK7yxCQ45g+3uykeZD93m7p6MKOohc2fmvgkCm
b7b/GzfaR1YPDh0OtviiwLKVYbPHfQUE4EJsqEtLru8s2V9t99S+mjOJGXZUFahcsGro8pwfJMRk
yGk+CgEfzaB9MlVjhl2vxBJFCaoNVwxVP5LSwIQfVwwXep/qzQFYTmyHMXKbZb7hFKCGJjEQHGQl
5SoUdqphQWrTbu/cofX4gcpYa0AsFdczlohRFmiofXnQakw0MOwaJJf1l8A3+U61J93Qs0yADo9y
7LlPs1xIB87iVF4h5XzF/tD3N5oSHXvdINRDCEHAATI5l1w1NES9mN42oCIUVZcAkLH58QY2kW30
C00rWGt4zjVdBaVcEqRHVhaYEooAYdasX8/d0VLX/iTz4lPQWHBP3WaPLWBie4pUzvnSfND6zy8T
ikYIzWfr1wVi1lf0aylCrzmt9wbTB4IORwW9p6VNrafF55icw+2BbAtj1CJOOHPzE3YB40qA6mkD
EILGpzYyyKasramejVp9CimNysZhwd6Xmrag3lM+bJ38CwPF1moyehEdka/6RMRAm0zyMVIbjv7u
jOzez6OEbhzB03PffenZknRAKeVj2S0TD3CEkdIKiA6iBCvt0wAnvrpe9a2YYfLBFsaj/um4Y5Nq
UsIoBBzIxO1ydYOWZrzTAd+ZOOGXQLZL3tzNmY5bK5AsxsGkuY6Gs/3rR/pMuGfPLzIzo5ZYgOZ4
Cavq984lSeqo7So5mKny6VQ5imEQm0wL+TtoscYNamwMdot8+yERoyCVXAc7gOt/RcXY9cm4DcH7
zPYyYKNWpsz4+uGnQYmduwpe6+0ZgMnuIJPazlZjnO3lN4VkbyfrOYJ2FbiBZnLPreGWQLvMm2HE
xJyUfx6z2m4AGFHMnkGs5T29KgijA46+b0HHugOBmpYB4Gxt/FfnOt0r7VYf2+boHzvMcDeWB9ig
GIK08jY43IPWJ9t6laQr5RMbGikrb52kJsfnYNLMmP/+vtRVrtajQN174WpL4g2WSaTsqQ+0Q6Ur
qW8JByQVerfVPWh5z/Ndsu1ISyNlLtTEoz3c22N+PcapuiVaZfyE9qgoN/ywjEnQAj+ZRg0BwoDh
DW74fSoU5OAyVzkrGxJcR0H24m/fNAGVda4JEqD/CX6dSmkDZLC+h7di+x9Y7YQvDJ8XjTQ8w6DM
NsUNijcbVuGndIsVKzgsBOAhvPQzVCJs9tyCbgorXvVE++Z8IHBGkRTYkIJQGHMdgvAm9pabTB5L
n92KBJhoSeirKq1YYg4HkHWxctzWIvuM0aXUDM0SEuSIv3NCAgkcLBKZRV/g89k84VQMyOcGon9b
zIY7XyJj9wrATTKdt1v9VeFh5aYZIEa/6Y5lkxmzJfId1c6QzynLiFJMjhTFWXom/ymOZoPHCKk2
EbEfWNlI17M4+qW+RfxhW0HbQe7GL1ZoWek5u8UEL+wxcaWhayQ6unKTaP4SSCnNezSM95FBORd3
OZPBILreS/aMQP4MY9eGZGIcRuNJWTiSRHyGUoSwom8NIViYAH0d4ZwXgBT5gvPqhR+w++ZwIcBr
4QVp/jFSRTDJjLoXHSiEZwLJoYVvlokFl4XLLHwrCW/L9yKQRUxskKAbvT0aLMIlMKt6qUPS0zqm
dlnFvgTpEEW4w70ZvMR3uB0voLNy6wUdB80EsyXapvsufdi8vaPTf3kNAaR7uf0s94rS61lvCeAK
HnBEPzuU3blLPdVvgLDNE7FdcqX4QYIjoQRi4y0Etvv+PkM+d5Y49aTLhevMPde8CUOCpLJtKewL
cVzoNJBqowhcdNZFcQAdQabgv8agm/VmaVwCHtCLJuadrGqIfsKISkHqbMa1pCfFHic8S16eGCQc
c8kWhjDoE3S93/44nhtMM2Vl0hW5562w9xNIWLm5EEe1zX705yFtj9XuBIydjoXoL502Mq08Pd/I
JzmHRDOpyO+MkpaHTRIR7iXm3gUIX2tfcI93SycN1ML6/HZnIHPQQkdKBIdKl/aT0k82f/TpNirM
6ZCPvU5etc9aAgqsYvVgWbIEamT+IpttJyRkGDEEZdhjG+JKgrsmaK0eQXZF8FHfxyZgyKXrzhIi
J4s9YIuYTVM8OoNjx13wm83py4cCw4xtjac07BbhzryH8dkJbcGh0+W3+N0nhCThrBGVDoJB8rD1
K+5iSStBS/sQtrZIKMOnUh4wWJMz7C/foi6g4IqruupWFWihKs8FbrHqmbihg3lWz4QHhXOb4bbF
NPDQzdto58Qn405RqUJqNCvXEFHnKPUc5XepoaGihGfkvzGmh5UQTo1Z1umlIs22+fy8UhFNQ/qx
Vu/LLL5cd94Rx1afDVZRce/8YZkBpIfg3JlRw4CwLah+46G54dSLSrYpY3oBsBMpp3g+ho8Bqq/J
TM1wjItvs+rqbfkcJMigh7wh+fYYMand9GLqviyb0NeWONR5HNyt5C0kaEI5siboc+lKMDTqZ0pv
GxPNoO/bXZtqTNalRUoTmTTNpJHfr+dMWGeGwmRXPkD9byIpvzHsK4oIS7E3t3rMeAAf1pfB85ix
wrcCtkEKKsAtx4gjtXMwMTZDdfXIxjVnNXxTacGKblRUkf0Eap1uwgQnu/VpJ6vE5PbQxd09TBve
f3I8aQhfL6Dy+cRebD4AAjVBueCJ6siBhe5Mic4BkcelcehKQiZ8uys456N+e3snEOaa6n1nj1mE
WhUFIGkh6ZeBcFr3j4XsFyLx+BMmfDirtgvLLZk3pn6pob/BgzDd/90Zg+IVAQ+auI9fkGPyEh0d
vFTNYcknYX683BcdwCU7Fjs8n3ERkC0E13HWsU/b/xUx+ofU6K5mN8RzIloxavi4OJUf/ji9q80f
zc8DpN94Vp8yvlLDe4JMSmV1idC6O6l/fqS25XUfiqZUS5yzbZWPb+ng061IsGCM9kdv0A4zJK34
8pwX3zztT2dp10s7AyuGc2Bd8twpomyX7q5qUHDV3fbXUjoK2QPJcxu8HixVG7YposwFgnsDHYpc
48nN2M14q8o6RSdbDqeQmlzDk1iROKcbQfrGngh/MoK74HRxix3BEM6tPTp99r1WtNWTpo0e62fz
m/OWPYiCYZIJEbdo2CjU1lLLgxEn1PDzkeiNh/U5bqQrGYQYSmNiZlbl1dAdwnD0XN6JoGn17lFW
ooC89GKjBISELYwP5StWjDerRWAIBVyEPkOPCPRENS64RJ1FBHYp5emrej6K0yhS/UuCQebpObBF
1ZwrQ4+YotyXQ0aHu4u9hbSftyS+wpIFguY+SFEp23tZWlJDY8htveeElFRGRIHqT4V9+JTxqBSO
b9RnZmzn8qU+ZXP2m8hxmU/5NAGn5RX2rnZWUUBIfGbZrizrbR+XjP+ZANeyuOHJjyhKU4P+47em
akMB1X+sv0x54WOWeEKDhNQLG2Le9G68JvVEIvCQQ5PKWIuefn2d2tgGrIv2ia9aWB/fegZxC8QE
TYx/Dc/SbxzD3FF2gNC5TJq6FWbenaXQ7edlpk1IfFkxPyrdj4dw1/FYmTid5d5DlpwrhyJxqARC
vUt89pFrgYKB7e9L0ln8I1jLuKS9XbSNr1AZnyScEp2m5f7Y94IrQTTIUzTYME62oW/C7hwQGKTJ
AVXC/hDwODVrnF+VYajofS/826aCms1o6zoms0APZcsb44gtrLQttEjNQ1Cq7cTjmsh9phoOnKb1
eTEA5oWsQRL7Rb1b/1qEYzVt5ZJOlzeF3Wltc9niqmPSeCwh7PvpZ3ZZisNmBYdz7ScW7oHtVXit
ixYctuaI0p9JVU4zEadG6hp7bCfjS/oXaqPj9n7dNQrVRY9qWhqWsx7hpKx7wUPq8MEKDixIqJxr
yZMSsSriFB5K5MmVNF+ONuXg0m/sl0mrUWvMFu6yjje6LHH7jo6iE+RZdRUwmLnh/Mfpp5BRV4xI
UHH/WYjln9A6FV7IHGq7sM9gftVjHexyuEChivg4H3K9halWXtjm9P/aPLTi4f6RivhfAcZHhx1Q
Hc0fbfOkP0HbRuDtGuejiGwssYNZbIHYFuBGWw9N1TeqW2Uds4FrEXD/zAdGoPdDtWi9fGyXIimO
jAN10g+r8Md6wKauagSCYEXK+Z3s0jSYeUfhDQ9+43V7bhqtB5MrbsG/h2zZjr9cMMi8etZhxUrB
1b0sIl4Wjjf8cuPybh0ZIwShxzfNUoss+VlccSTwqqKYJMoa7uLOCyxPOuthv3g/BIJ6ufoYerRc
clXKeAqNgJa57EirI4SUd549qQExQ/E2Fa3noRw2e+nEU/g8W24IYdTtXp3sr3gj5kpLIn7DuRL4
pqL8xDR+WJemNppWgXiBIJ5hGzCExCagujic0fMgZvY759zSstv3DBbvEVYZiSZ45a6KkP/TQX7m
j5cfreduXyYskrm7zK7SRJog3gvv5gALF+bBm18qjWzUSmua01pVHR/3ob4eXQ8Gb+/xpcoy7rpb
I4tb2CNlVUSj8wzwsHQBPMEqwUUjNE8s8RDib1F41W+nfpXun8zsyIDfskJOiBjN6eRvZyGyHR7j
snj63GBYIPT4CrOSlvbwV/Qpnyj5IPhRmDPrtWkbRa+iWXCCK6V6pns/ic9KQc/KmwCbp7+aW34p
jaaLNgi8ubYxFXAqG/bYFzjMFsK/NL5oWuTvpxylmOQF/n7EVmPmjHytUmSfkBOJxPg38x0gtdfp
Y9sjWPNvV6CwZGaltSuscLEnvAs9lasVceUiLM+QDuVT1CouWKIihSX0syqMpnqkNa/3KKYx5SQc
CxAw99TKn+hXGviKGl19gCKC/dMSRSYs6CIdUJSjQRj2lBvKWJ84wbSEBFUmwjHT/MoLZ41zSkMO
ojtHe0dtsvFBQI1a4WvJQTojukCAVVE7QOP2hNJJbHmIG7SFXUV/mUDHbQQw33MuyesJ7uLryvjx
+FsAkmgk5n3VQic35Q6sCaw1ymiklYN5reKHe10KbCM2Af2KfQEWeiZjK7/Qcf7XFKGbc3GTQgC7
acU+K3OfS4AERvCyXrwkM7xk9tBJ0cJjElkdmKW3j1UjMK87Cq6Csl5PwSgmIo1ht6Bx9sF2fzVG
cnG6Vn06sfpprcbEx973grmw6+w5CoW+IA0luNd9B3Vk48Uxmasf35eMmanRiZDKBVzknmIuCDpx
1+bMuzJuYGpuSzf5aHLsW+jqQLcLXSQP6jOkP9RvoH/r9Wqqw5yzUHGwywhRfzrlTErjmz1mIun9
ZKeipcKCKbDhPlBOTZVRIR1dsXHndpR0ef3mjupn6pSJMJ1aXIN5+K9GHEW4CfXWB4DxpsfeLorX
mvEl1xBHGp1XW/VCaQlaHBFhFASLv3AEskg3QdsI6SC+k0HPzJKqsVH0LBodXeN+GJd6cSwrN5Pv
Ag3ZnO7fqmNpnqdPTdNSIHeuCG1ZhGpNHv2qA0OOvKK2cVguwVvjMyCm2BE5hDZEl3kEmjZ4m6He
1NV7OZp11SqoJTQJ3e27YtMpKMtbJlimVcP0BM9f2zkkNmlHjxf7pXF/naQVjmHdCbaSuMFcv5Ev
dderatvBcsxv9TntaGpiaj1jH40mXcBgZeiQrDjQowIU6trCFriGqcqDm2wVqSrz/HdUI7o9cq7n
T2mC6ueAUbgKEytRjvz8xOFwM2CVIh3chZotkiNmYDKEgDY7oxtCVsglM/D068c3g7hsJrtDJlve
yWG3rrt6mCnJ2baQNPAm/Yyj4uPTSX1h/Gc9xUVTEcOlZaWR28uZUWvyFhUV760+1AQVDVHKAHTh
l0Kz48gcB/l+HmwkfJC2k+ToVOeKUjkKzRsjvdjGfVZt+Qvo66iDV5ju3t80cS5w/xYP4HlBfUJo
SA7X0AsCj+z2eWOxtnUHZjuMzOavuhlOzSwxYhVHpwgz04zbq1ltvCle18Xk5n6zczRlYqQf314u
9i/W5o99C7IdPonQ/7h1VXrCRHJ4dknNNsbR2Qf4m9iNexDJULmFddApsuEYZTQF1Q6FwGSprowY
Cd50Z7TztAshVYnb6tkvaWB7tcdoMoBAgZiqralNUNa2iv5JTD9VoaJ0NhozRqVae/hyM/rl/oRf
ADchkh/a9EfLudIFPMhptJ9MqXdg49Af/j6yhNWNbFXfp3rj4wmPcJbxZIYO1JGBp9g1hhJ8QRxC
IQTeY3K8yhJAKKarHWhrp+F9ZDhSS0rn4V4l+HK8auzRogGWOraywh8viVJx4B1baFo3I3qEidwb
SPbAg4FLnnF7j9NT3pJNxKpQUkyhnq+8oN3lms9CkVzZo8nJjryeZw3TscX8qu0wzGsJZ4jXXHQM
UkFuvgWJzwUcvq8yU8c5T2ePlDTSzvEPH0fp7ia6BUdwA2jQE4mnUE7+i/Xgq7vnz1XVodvNZKJ9
/aGmQyeaep9QL6cnmjsRg2w9wLAYdwgoEotoxjZyiV3JyuZv0JXd3744kNxH0KGmIJoV9R6kZpRm
1vQTAjvMAz1B7dlzxzmhBeIu+pDrzHijr/Ub0somJZs2BDeowDT7mY/qtV93MN3GCklpy3SiaLmE
nnJPIncCMVDEQeGzqPC7zOertfoDKZ6iare4On85KWH7ESJpX8fZTxYmFwI5aWaKujmaKMCXySl+
LXOAJwNxL5PT9ghNnL3LM4e6CsVKN80M44KgmOMFBjMtT/8NXu4ng1dbNopqAmiF8SitGaKmKF9a
6YEWiaj9D6i68Vba9sPciOe1fx+rZuZAwnH7yMekCD2RlbmVwmBTwaMMvP90VnHqbg32WrOj4eyO
OEleds47jbfEh5OSdj8cY6CbrNPu4eo3I6lchx1ti/hZj0CFMS6uLlkf/avjRNdeA1tF1FOcLzdT
/bSKuthfntSEYLdZNRLjUmgJZVvVRblcJS/n6E+6P6eMV5nIHDSFTBh0zOXJRR+SBa1LXH5dkIJq
GFkpQsA3RQonanBB7gRc8UQgAYxYd6dyvt4mFTyLLgCprWKDCLu9fa+hM6nWJoeUUnQsG4U/Jzar
rUOnLWVjqMIvU25vM0hkTtSgdjyin2ggNfYx3WujHAQLwjLrsOc/Pi5emcY5687lDzJg6f2nYD9S
Hj99viZmefIZQ5SfgRXnMF65k53geZPYw7ED4025DWiMgGjl3qtYSoJPBYYzb5YvDUs45YZOzD1L
IDijCqWJ6S4c0JBHl3Dy0cWDu8rqXSWgffnGFAnjMC/L9NG2QxRMU08qJvFBVlu+txRekUcGOAsP
7bASC9ccLSTZbBrIsdPW9eySOfyPh1s49UIuLRo9VXf783Q10qSZxW3ARdJk8umUh4tfgf1VtCbk
44Tn+SN1MNhLo/8VMoTs6mjdBgRTcO11pGoS1KGntRvv1Vrh7xKxFvmSjHvWvvrOD5eqYsDZdzam
TxKcsz6iqRqidzRUR6lBQdovr0gUNeWEoyzWawskJxcZSq7BkptJZt2lFSFJ7M6PjXJCWt0Fo+Xf
Igeqx6DIq/9KHi4Ii73Mheg4gxADmrSWzOswOdWoq52Goy0akaOA7Y18EqUlXIuc9VdHYbbxvv0U
yKkyehxVkTtK1wiTKLQP/LC4549mNlq/hh+iReuTvk5cpeaYukKPcusOyr+DxBDvC3VUNZVREjAc
EqzYewDv4heDi09h6U5WF4uyImoxbjsJFYcLybXI/fqBei4oi2JtX4IipJ24kWOAZpxWYuxktiUl
hoyunMqyc4+1sJG8gC0mysUFTelnYk4QXftjEsvKC5nujHUijpydsgclSIeNSIqvt2pIU6DZfTJk
jU7Rq9vTKi+/54k/lUFAgFeBSgTcaOmUEwmqTfoOGSQKzpI6UTNKSrfKnmlRlSErGNyzpA6JuOPM
OlDvwj+MJcCgGBCuGo6RFWK6gllUpoybQ/q65FAV7GzVjz5pXXlxnWsqbq7w4jsZZEC/+bb23ymB
wD5ESLwmtzNgQnJz/hA35iq4rMZ9CzIDxrpczqkgcz6mSVIsZ7VKfCbf8d/rOAcLEVDnOe5a8HcA
tqZWI0o96X119QYEMCEqt1VspyZRarUdlVcLa9gArZ3kDSssfI9tjvwV/RiJ3Kq7FpTX9odJHdCd
iD+lt1DjsFzdnk4eUuZYoz+3I90CvXI8dQtz4noE74dkU/zjWAlh8XeRs4pv4SvTOsPKtuhJEDqI
aQhjsVxOazYfiv7FFHmK+ppuxcXangNpN7aGilshUYdrsOi9b+s4PRNlvnxt96fRSBztT8VjL18o
VjrCqY8g9RLoE06+1y/3nu8bvdhJkJi1S97gb2s7RL8WygrGNqoDrZsxltzbIQ/zEU4XGfeperqI
AAgiegsx17mHTHa91abhQd4hS8OnATFkICaAWXPNDOl6owiG5mqHQN6o9xrbWhzTQyb+HuGWvVmz
UiRX8AesSrbC2zmg66jihMnZDD+6jYEM0Ecw31QAtmUo8esnv+XEbY6bvm9nShK+1hzjUODeJ4fK
4yK6MYO8TpKIWa003djkeEov3lxbkN54H4Rizj9ybnAs4JdRdNpUKH35F/vEfye9E/nyKaj5Y9CH
hDQj65SaDoOROxNvi2FUdTYfCRR5P12Yc4MRMWCe4lsD/uR2GhElT+jg7R3vS1kiQ803Ev+Z2n0V
ihjKUtuCEuR00ul6RI8CsGD2AQjaQOyUV03VXCfNBj/91xDuWPqdVV5WC/7rAmtzslLnAfEemoyH
M4V4+5p2p+qZK0TyDkZtUWFhL02+FyYzeoU5eKUqRa49c5jIc20r5JtjKCinsR8222fu45QcxwKP
LoIEv9Rm+yIk9ur6jBHQMa+OtafSt+EDCLNntjTTOL6EmSVOByoaZBZpjYkXd2G2kRoiPwvet6ID
qlQUBJajO3HxwvioyzdxN2+7ocKQXOUEg1ou4pBCyfcifkGMAa1gfwNlorIxPIO94383NCPp+9Oo
iTEC3IK7BtHMBXBB5iM+aDTWuKSRIwPJJGuYBct07XpGrqLCuEQvHRFswZFRJE+isZGxT7ObwSgC
LcgrJZqu61PEMsrh704Ck9nvHp29vuwPJ6pPZBRxOGezw0Tq0HZYoE8bj4TttU/udPHKzvzecyTR
h431IKkJWfzRppfvhDNBHiEOwCyohf1wXyyH+U03isemojTDo2na81ip8cxlL/WNOEsyhcULfpiv
DlXy8Hmi+XZ4m2h/wcVhrbEVm4cojlBq1DKBKle9BTdda0w3fG8kj+jWWCfe/ktahTg9XSk5SFpN
BZiW8hV3qPbn1ZN6n9d6iHZgNgM5n04+eDRCKpyVEXGlFk3U0psR1Cr4ifjP96HnbRalebouywFV
DF59l1FkV/dKyMPOObvlaZjpY2SABHBUpjPV6xIt3yhoEF9+ixyb4QOXYZ/p0JbtZIxLPp3a5VEs
grOKrlYmjczx44n92hivPQapYQIaYGllDAB9zVvSOPf28PNIfFV1YPPxrCbuze7kazE7JUIZgF7u
hiGXCrOVL6ezzR4wl2bNXB1dMCb1KLF0pVHrlSoClr+r7A8IrXse4Cpk1F6kMmWS2+DRESUqKJNX
/kILX1iUu3w/AbYSdW9kMSHA9MUKccPKhqbDPh8ONqLfGJ1O8tW4bJlxJa1ogTmS8Dg/IENna6ma
t4LRAuumSRPzUrdbPu7ca8GUaHdZVJdmQJMfR7GseTixFMuSQhL/wlpb0kISUQTClPZzQnw3T6/S
/JkXZUMJnN1M84aPpdSav3RTvIfPIZfjq2jKLLrFGMcaHxuo9cORqaF1zQnP1Bbtx4+2BLUuhIeO
yVCzgY0j+iohAhwZRU27yer03sdk5RT42A5tACtiX/lxcJUqT69GLsbldCtTQz+5R273O/eKi6dj
49Oj3bI+90uKXC88Gd+0um8RRnXdDdNpipOhH8k7kkn4Ac+fa14LLf9Ma9cJeoxOEq3jpDwnhHo0
gok1nD0SIxHM9L95YF/Tvk8/OcdGqGxyzVnkxsl9tdvG3fcvG9pEGVh8gYQliBAMLSs2BxTgw9p2
OQEPWSFSiLK+z4kQ6c7vcjB/LO8uK8XuhZfJPCWfoqZKm/4GTux2pULIP6gdtaFzQbu2+fzK0n/t
xbkt5Pw8yhljBxIXXVLJOSy0KwZXlp7fzJtBo+BBLyN1C7P5LkBN9jQ/p9AAT3UJ21Si4TSAVk6/
c3C3MkXk7r7JHVE7iCKvaOslQBHJiZdLZg3lYP7NRbmR9JwhVMWT3BcVyZWsrgL+/krhPNH5+OqP
TlyFHDsFWTp4K6YxdGlZsmQuT4ggAz4CBz0v3IdL8kMcaOkRSymkbrlbdm8CfKivu4IfHeNCvEEF
Kxz9u30Q7T5qAecqQD6qtyvLXhweZeTl9velQ5AauO4x9XNl4bLOvEiqONbjnAYBvJTT24R9y6Q+
5DRqbvc1Zde44tIJlKgyAjhSdIHZ/Wa1f8pZYiZUn4V+r7nY1BsI1sBfCysxL34cRVuLOChpq2Qv
H2iTuiLCs53IGQpEnmAxRJweVZAlP07swPdZCKJ7Auj1nLHN5/Gj/S7ZxCTez/+DyHwOmi2avF+L
wQy98k3GSt7GhXitkGQu2Unun+mZWQhlEGaB0+dCCCHjWjKLJEdepETGUXMviCjnDXGEpw4Bgd8n
f15U5WEWIW7zuOYlO+OvSoEcnMCAhA0q4ndIL0GvwwZZClufT/EL5paCrtkMsp3atklKuMUUyMDE
OCPqVoqRDkiwOHmbkceywws/JOhI7sC3mlCD0wB+bebPEsfrmlBrQ4PN3aubtVVcCs24OqnKJmwx
mi+YEjM3FnBj5etdXGGw0/y0gasb0AKoauQ7NjaDNJB6OS0s1kNx+q+to9Xy+YmPtHiJD1G0m1vP
EhVJeEw7I2KLIEHd4jdR1PVedJsivwj/bZFnXayIHkDpjRDWX22jJ+JCKdBukodiuJyH+G7esnAO
n11zFq4OEvA04+DhlAOBQXm4VtG2YhvunK7rAgUU+uFLpOHJkNXNxpqxefyft3n2jIs1w+Tl1taz
LYyBcQW0DTJradSzdW02PCYV/tjgD7QRgWVfPzGy/eOMSqaiuiY34mMk2hxXLTSp27uaYJpapXBs
iFAv2FTjOQUpK3wC7ND4KlREaaJRl0OscCYASHo19YNgA4NUxvHWaAoxQwqvRWK/B24DeYQ1nuiM
oqWIUgXcUyLFod6mU7I6S3NX77Lt+wN8gQrKy9fuClLsfJGk02MR4aHe7pHcMU8RntK70YLgP4VX
62E/GD3XIqtSGssriSk7JiuqyWuiwleWqB9VXFmZtzxWrjXkVZXUkkyYmIqpmuqL5gk41XIRK55P
4xbFWYA8CA3yjQLjuqWK1fBPxyBP0ls4Hg2amTzkqSU4Ws9FDXRTeerN3wetuM32J/7J1SvXTAgv
niVJollZb3r9Kj9VnVGHFLGIC33jEPFDuZDdsH1Dvizu+AaEBQR2toVKGdKe6cZOqGB44phKNP1q
InDxYTys2nVwe5SPPeklTYCaMm43Z4R6QR5ok2yHWfHAIEsPk3y/3SFFwf07fOGXMVpKlDUe9OPv
2oTiGvq9JLntUdOPc5KcAFu70nOGM4gsClsdvwDL3SDpNtnHNmql6BXHy7pKUazLNJzPsr0QtP7k
dUID2k4rKjGChGQ+9HaI4sZK3GN3YRMcRBGsAojVbUgoIPGXKNl3kxE0ZASGp7zquV0rmp+xIB4A
UH6WnRkbxBdqbUQc8KCbh+gWi6eXHS9ILSWZ1pkGMAeMZHnuG+0724u5uwJGh633bXnMTjYI13MI
+qmhPOwwQONBudPn8urQsGV3zCUgywvNN3uTx0PmLr53kYjrPOQE4vlVKnG+KK00cUIGKNJpmDny
q4WR1qheeKAbYWLlMCcNgUUSfDDdfeJtahro8u57nCMfc+sHAnkNHEBtrWoDYYax+vfl8DgP85mJ
1P2dC6yCOWPcmQR05P67rAMysMb1OpDlIdWsmMD3hTFxBV8tvKb743UAh+17ca1FigaXtN/H4BFc
894k6oeWiZ1putGdLfqv7CK9KvlIz+wc7QHMkoAkytyAmwHGp/5KwKUxb07J+V1ojydL6DFktXub
PFbv/U1YVAPuOZZfVFQp7QdqK9G57mDl37ANqeaJaDDDc2ctm1PmAeGPXjBxLaJy+ZEvoERtO2/y
x+T8ezpZaRamPL/+9x9shB+8L62y2bVfMDBMyc9yV8zOyWkUDqdvVYJnOS2XwRCNXaBctuse34sk
DTmVzc/xtdsVyS62K2qBIpTXMa60aZeJrc6WbHNlCDYwidY4E3OICoQzBTR6L3k+S59oBEiGXY1J
M4CF7SqVV2DgBCB4K2uTrHHuW0G6CRY+qjvA4BoVEh5z693w9cO3TnSRz3IG7+mVebZWSZavqCbQ
WgwNDBtEC/nVNSoKVEruPffcYpClt6zvSvZeQ2S09XCaJTtihxRZ3d+lUYJqQ5eL+pefvF6ppwlB
nhBgR5tNn0zHdy/BM+pzHvBV3Ep2glSjRuJCQxz+a2L2BmfsoX/e0EhSgcuy6XFpBiXaIEgSVk9k
U4bMoA+L6Hc8R2vY09Iew0efIrZPV8DTYdFShiavuH5ybVml7JZ5kGMNuXX1evXufxEZd8gVy/ky
hBH13LoUhI7CjW7PFhxu1X61wvG5ym6SXDhPpbEvgBqqeveHhM4Tc8kOFgbP0Vm+nw9efTlTaV7X
z60KQwTyU3BbXzTZu7Nc85DbZ7W9dBiwSXP0p4o6OD2LkEv1cSJvKYTmXJw2qRUSxvTfIK9SlW2i
ak+Y+BHgNUHCVVRdYDyj0mj8S92ww0F219vAAn/kZ5MHTBqVo1qewodl31h5VMqKlTJ5gRfCD9Wv
sgywFdsNQ0SFrLVdMN7TrCgSENT9NZYO8+XSUStj02F9h2Al/8Gv2Wvj3Ie0KLdhVM82f65Bkfop
iALri/psK82LqyJk9Mos/QBIHuEG0nZmDDjCpC5vjcsTqixHXLn4D3iTP0KI8ZNOdmlSHiqVrpMp
g5oUM72hRAbRT+IuWiqlNY7UeS25wgjouSxEO96YDNX0t/ZDZUUqBAYs16dGwErjUwslOn64kgv2
tiFUdnRDv5ssxMCQddQmpfJlDBzdrSb+m6+BdvuufkWRzKf642Emv0VAOjyypKLX5VMiB5xUtRs3
ZVPg2v3eBs911s0bRikhqkWNbqxwbc8D6PPFgDleXkECrWvxWWkJcmfUdxObdoDTVZbmW78V3/wa
8En6ifm5zAQgQYqs4k3rF2aS/PhtdrE6GlN61sVfetEoPBd/Zd9GvpNXrR+2kjWDnFeya/4sfnRw
eHetYRt5C5RODRK+PV7uA7NwfbFLpsYy6vWKgfq5WmI3potg+PlcqbGppWww7Pcu/Z3nL76l+qwh
9ZpoE7RSH1PxDRYdtg3f+AOZljC3xmj7mSy41fmzlPr4F+dfM6znJjtl5saOj3D0mt5dKBUGsATz
fN+SAZ+VbvdncdbV7UV1s+UIGEf0iP3yNZjn/xI7aAtczc/53EEJM7ofnDCfg4NeBDkbD38IF0Of
RxdEY56RxBe/04qBwljdiPhVbmVBeidiZjtiPO/9Iu5vmfR1L8ATnuq1uMC370C+S+uPeDRmfWtA
Ec6rI/etc2bd7yrZ9ejn9in1BBVpkaI8d91J8N3ybVEMoZP8qIu5wBNDsb2bcQV0Cq9s9O7G7sRO
KnePH+8AFgn0C9XnioelPBLuUen1FNI7itbf9q7NtJEtJa5gDm85aNq44KsKQ0CadU/oHjDbm9uy
b7ig08WYBs+6vGVYNIAE6WESeDDoxPwpM6JPkifilYNxt9paulPxMdoH8rq3JO5XF/J0iUw6rPu/
ZSLIR2Wa9FeqF5JSBWNFiaFR3awaOj8zYx0aLZL54IQYAJ38Da/p8eYICEq76Cj50V/At5fQjP9D
Ae9J5xbYcnCI3BtQQHvOWFfZPN2X+m48rQpdrJjCTNE270Pf3eEBqBuqsUUnXy2Qw2BuMiN9dEjo
khZ9cIj51daRfaNob0MmcVGke7hMY8VgvEaHTDkd11siHFDh4GsgA07UZR4o5yy7//BIZekHxJcQ
gvo8LDv6VlZpJvxzVjf7IUZtNU8QWl+BC/J0IDYCqsVk2XcR++eClkDMIrfeh96xnrld3riJiLja
1Wtu9SzCUoO/dI6use4TGwYkM/xym3pwf0cZBHyfmphzfZ4emysL4XjvbSwGShKSaGU2Dzejk6dm
RcrlCMDQPnFAqrJ4SA+eT8rjHfl0accllsTEJrz4DomkDnh5ps1T7mWrp/FcG+ByR6j5yRmWJsQi
wTjWpTKBDPg88xtwly0ofQWrmqhvF1/fcfdqGNcfM66Xdc5gAW51gdY7IWgvyugPobzeHfSti/vb
vesY4fasLDfhKNpfZ/gLnAJuNe2dYGjxz5TFZl8O79schxZeDGLxnWBvLgpVv4hGOTD3j8IRUVrY
4JWqYoQcT1DqlT74zDvy8OKnNRkTOQ+Ij+yknVZXtDimT612989AVfTbxSH8lQm1hLn/1Lh8690G
tReE6bLttA8Nw6Ori9vLG1Dvx/00y0FQsfoN8F4BsQsKiUxJlcqGLsfKtdU1m25umKelxFTEZbQX
uzeM5//vK2TljRPhBtSX0Eylo3+CoRFCrChOK7I+lMgyZPwyRxGv4rdjEnXdVQSnxPGGL0AslOqv
GlhMsyRdwxmAe/I7KTyZm4Q/49ABPfsGixgtKfRHz5Now3Tz161x/uoJFSotrYlmXKXFJcK+LT52
zaLnpbVfBs9U1koU1p2hgzHDwmupkZGkWW0vCVgRAtrAtGn4kYVKjdCMM9PDDmuNXJy/6Tk/WXDF
dXQZJ0B+VNBwBJMiaG/+EgJ0u39LTg8eOz/wFo9BqdC7IMMO1mUobE9/GgmPiIdo/eikRANdTBNM
7h+lFPIh073zTcY4UHHwAMMVb+C0zs1v8Lwj9v+xaX4Hmzgpw6SQGmahcEDojmf2wQOZOzvI7Eod
7Nf9vF4bahWkCrEwA8i0dY+M73WSzEJWypO7ZXA4sPSq0mbur1U6pEEEq+Hv2u6N5gDeFNGOcH09
WfMLR1PuvPrL7pODhieupeerhPZi2IFtNvEhcx594BERnr4hXSMBUH0BwtYq1AQuPuEW6hIaLx9P
BtGnsOWnZu31ZWtT6zFGTgtzaOroHko6iWC2LKxUDgzRx0JmR3l7aWXz6ZJxM1rckE6qXV0Ap0+c
ElxKkKyt3aQt6oD//og6u0MNmAp2U+C6ad/l8CzO+b7ND6H51SFUInGglkkOAPs47yBUkDSRiJ2o
/UYojbr5i5222bEN1sXVouREOJxRtROwDVsCxPuzbbHnozkFpC3uUXsK/spA69+MREwc1lSBnrMM
hBsmCorDCxSSw/qDMClQmqGimbxE7vNJZb0xekscajajEKeL336IfDoDhgIaeulcDxPFvzbLfmMd
LYKsF8DtHND4MY15w2rsAkBje06f/27yZzw24Vg4EA10qpHGoSUUsiLT+B/hLEhGCrUBaMH0xots
oDMgie3coa6k5OEyMuavE2T1eYJXKHJ/X8YqtHOK8qVPzZ7rBZSyN9j4eJen0bA8tfGcuuTIS4Ro
snL22hbICis4wS6ShSfzxGhPBS72MzERAUxHZcJnzpEmM7geYOE8da4ZDTrJx78Ob5a33G/sTvEd
8PurUeNzFkXgjUo/5jHUnUJjD8KKr5vHoLU2cuLdWRzznIpDuTiLT2cTKmJq5guP0zydNTi/YjtV
hXdvZbyGSK1Zf6F+JN/fdq6/afP55VB9MJfjeZMeDOmIZiEoJwt5VfR5tWag7OwtHFXPPs8itWdj
JMcO+HnxdKZHsTfc+ZPOKrdPTwTQtdIhEE5cSCWhayUOs0XYxr6xKEph/RNHpegv2qRS+cjXyQwf
zAt+r3RMDO83eDyAefOZIOSrnviczaMOfa3WzRf2kuwwQ8xys4K0GXavmvQ2Pd4kq7RYUpwI3p4u
LpRugjowiYJeMlKvwmtC4NGEJBNZx2DatsIYEhe3PtDKK29CxlSMgmPXHzSvHYO5gklwzdzppD2L
eSY5VOT/eoqHGQPfm6ypKJYMS0HqjKzNtJ56XAi4h55r/v2PbFAQ6E3A3Ph5Vdu7VIBAYwl10DgF
UvnCFVsvDMrg/ESnmd6kiKfw0tPW8xfaeJ1snD6fI0W46Rs1W6qeb9pOz+RxWxVGjmhFzMfhWVtK
VRpxj9zoZOIOpldXjh3BdqM63jQcKtcAGZiRUJOFVIo3+PBEVnjHblbgl7crICUCkqJ7qIgxsTFC
Jkr2rz1ZsqOCig2Kuf3lAr6EgExvWKxTx2VFhbxdO/9oIQwVeZazFakwU21ABlSyFoFc7589NPVt
tbv3V4+m9UZsh+7pLFdJJnH5WUWJOxnLzpCdUzngil3T0t/alSFvD1IySs0z2m3rstR488P1rxGt
2OccWgGWcqzwd7M2Mx7BdpTQbQ74jsxWm8MJ/cnV/KO+ybJVYW3RduRKY6Lcs4U0qEG4eNu0l1yc
8GYvmzTks6Y2FqY5/tNIPKhJG/1wGDZ5zilPwApQYa8bvXxSmLCRwwuaatUwJ/nttJuMy9wENIgr
E3uma/DrOFZys8+iYUfJfl7IWrzVHoU90D/17imr++d0YCJOD/uZGXrh8bFhZSN6VIsd5l4YOZ+k
5+RIk853eqgZVfRszMnfz/7mISGa5C20QWjUA3t4toblMoGo7kpvNKf3g2f7qawqll+56280+gQa
NkNNd8LF0FDC56NRle/tDVFRpupxFS9hMvWGG+KHClvwamt+RrS3kSLzGJE9fe9HtRQnvxtOu5h1
Ph8TZEW6IDYA87kFkijsTMNMKJr01WYdsOHwLNbEtZLdOIidE5iCpdiITAzD4QwJoupZ3Y0G/jVZ
Zz3cfwp92uhktAEtR9c7aFUA/jIDPtbhOgUKRMFev/mXtfYGZTh5xPVmOXAbXsmZu2ygXKcMlB0x
r8I4KJw7NLUvbQTOW3e0X9DS/M+ixiYuFy6tUuUy1ch7Tcwfw/NBH7t7jBtPqLHogRtjWJmCFPMj
X79x6H0Xt0P+vn0xT2fUU27g3YboifLtt5kjZAuXJGSmhqIn1RFmzzm8tsKLOrXcbfsquDE/j3Zr
wEo6GCEqNAJ6S6PnAAXmM32pZ4inXHaId+IouOsh1DT9rBbAJgCidFotTUgXvB4SwIrp0AUMoWAi
C5kWEi9rvzAwZwsGvcJ+v2vsvouZ4WhQX7P7cU5je/KHqbEsIGzfDJckpq9KzVNKa0UaH3W9tnc+
7bYOTTwqMaFh/7SO7Ronz4aAk2E7fFNUEk0aPhGd8p/L88fu+EBITOJVqTad2JhoLdhn4cAxz0mn
Hz+cNkinRoG3VTUKON0se5s7kctxhfuujGWNyhoqbToIvZKIE+5VRzi/kTB4+IH6XlZCJUy8C0xc
7/SWBfVBiKtaIdJKbvhkIzxO9ig8sLReKWNy/R0ERYmdUqey0kwWuPmP68kuvhgmXfOc6EtZttXx
tUCsKEv2GUdbMnK3aHgrhoujNKTcCCGys34yK1TVQPOKkxDng9yJ4rDKxrFqgp9Fntd+Vxk0lTDN
4JUauUhjplGjX+E4t2baKQIJhggbEJZwKWtGJQYyIsM5QsIqHxz8S0shD3bX/XRapPAiUq0VQs3j
DlDooBgvkHMsJDGNFb4RRFr8wsUzdyGkuOgmt+uNm0LeVjym8dab8nLPbxrDox4hO8T4IS4g8nk8
Pfd+9eOwETacGCAUHU57UT6dLcCG/v0TkP2sskRTitrHpjbLPvcuWExKuQ9dTvtlFkEhtF3gfkes
FLRzrtOAeGvfpYfEVplmOITFYP8Q28DitQjimEPg0FIUtX5u3y3auznuYLe5EaMOus4DKjI0kkVK
q+TryAzv4R/+c1j848XneX/hiw4AvTWvfsTv4XQlx8IF2jTWVIKV9qJ1oFz7AGRsgX260Q27DhLG
4aUxBjB5eCGzv/0rE/2GUt0CUIJhgsqfhde8AtxQzuLrFstYvEykNtDUxKtD3DRg4MgHr3BBcBu9
4Aa+FtjKQPzbfmLPmQdHTMRaiVZUyEiQyNwX9oblSDXgexDS2dbmwNiWefyWuVl6fWuNlzweviD1
DY6FgRLZj/aq2qYg9oXKVGXTdDsg9kzkEPPpb2OevLNHD5mZ0Ckrrt0rXi9OIzWs1gdkbaJCm2WK
bM+7Bum6oW31M4/e9+mIQIkpsuD8+V8TuSfoSqi7Ba2R+wx99xnbDXWsGO9P3OCrYVwa93JGIKDr
Ajk21R/Yuhg2d98ifKR2av8w9Ivvpz5jVblcsZk1XdbuGL3jz9ObeRKPiu0Lx/p+heSewIJo3zjK
pUV9LRKG2sT48g4bB4XEb7HcEVNzQUCCWeS65RKzXNDdrddvTp4US9v2tj7D3xwZhXK/BejrRwa/
c5EBGhcYziA1uDZwo/OWb/9hgh9JnxBRxvYMj8c65xotAJLMu1dmL6VPrkjBoO8/hAiVG/XaRNDR
IV0ed6c4RVRos605TmKks9xHKS77d52LohQ183xVG0jKUONDe2U0QMY4W08CE1Yvy5S9eeeXj5Ax
8sFLODqqGfjM1KnHRrX1KR4Py11C2/cg9sPWliHB42HAeS1I2EMwxUFe3qlIX0xw84K8dkvl6Rtw
7xfIQX/oneyfVvfQmqzDUeUYg+VrlEyxmjkd77842pmEdGvWVuhWtLVon3H36bPuMSR9K1+k8+Sg
DaOhbNEG9WB7QyL9BydWrwUc3Me7fsgKjG2uGWYHTPoDzLGV/Z8hJot9p5obDCs26E6u3xnTV6d+
MH1EFOF5L1sCcoH/wkayBEJH1MJMas/rRAz7n628Rc9DPR8tcj5rccqxOWCLidghF+azcmyr4lIB
aduEsahuoMNJx+1Zef2ISJJtJWIrBgjak/glRGDxEaY2w/OwzPxiitrlE3kgnbFOXnQaAxeCwlpL
nJPKSbFSNyg+8/FZhpsAL3oqs61H7KME77VbubfceDLcDTsZRHRy50gSJQSAZW3MXxcgdC4O43l5
6awM7QFBJBgyPnQr8mglTRIkvka8u5fnEnk4CBs0MCJQ9KwLviX1AqXIyxeLg6gsBvaH9KurusXl
8eKowB6pL3y878JXziup4+3n9yw0afN44H/3d/HQN+b1x8xooUCcKn/MFvVmE+bplgmNQupVmQrL
Qib6SU2Utfo9Lj+Tvo8tOY+n2IBndIAsDWmRCJcO6YvC51G8QjZHFsJ8tvcLAfjIbZriTdkwFAyr
6TxIrA6xdICtp9yq+BNwNOFr4CgKD97J+hyXdrvceGS4eALTvPfeDQ24Tn1H1ru+P/Qg6q3AA17H
6edeEpv56GPwD69HNusvZeOV44lo6+6n+eOi4F4on8duy9UdfIMnx3lnMup2jbRQP3byAFIEZnO3
OvHOzPpt5IOmVj+BkCplpv4kCYgO9+jsZ7nefdBosl9XjL4+CRd9ozdjujZIP/+beRTRZelMxp92
90BdD3ktPlBl2xyCedaPVoM4piBKbcSnKGza0DMioncIBxnnIUtPZb5E/NgoK+ZlV352beMyNlqc
qyDOOs+fPQpW0r5TztrnMwiC5LPlBfx7p7dgpriaRJKSbCON8fX0IvPN+kk740NVPCTYGZa20acE
rasOuwtcQCpsYlD6X3r0fARKzex96L6GUdG82AN8FERmC4r6hisAYPoqTSa88uET6LRNot9Jij6I
6wgzWSVCBMQTliiTdOctN2CPvtKAqpY/M6DWlP/m4lkKr1JUW4MSDQEOflMff9sYW9+zl/XHTfi7
noDfXmAqH3RYvmtKMaRZQ3DhN+CPIgBijCcXjjbre1nD6MtbAB9Qt1PMDSAaftTxBANOGUnyCCv1
OSTQWWf012PKmmMmj3RZd+QCnELRAtV57hUgJ8Shnq6q7nCSc6haSi76LGliqzOcngdAAqkpQHZx
DcL58HQGvDeGX0GhcVPNgoHcHzKf7JRrgEgxumFdTUuShmlxoZNcOHhrlVdTWoT+xoLKqssbSy20
A9JY+eg3hdvUTvqWqb15BeuXMQ1Txbf+L139xgAM98RonziDKOfbPv0+BhhnfTeWprH6C1rpiIoo
+l33Q69Onlq5o4YML64ToE3Ra2VjA7iVf1fKWPEBGnpe3VupssSrfaxP6bvZg7SUP/2/fdaf7Jpt
clMNM79tYT7AYhBwl8R3kJNZ2D6Y5Ds7vivavpZ2dvn+lPpoO239NDYqznvnvWc+xvaUAB78x/yC
CqqdsHby4JfCDoUjJ1me+PSuU2aDHBMtRoRaOHQlaWBO1N/K+JfPi07pqsiD3OMBO35vSAU8FBHp
Nw5N0NsOThXPtUdOQwFG663G9GJBEO2SAwSl0pzUDddxNgN0XVRiHQ7dfMNO4KOytfbY7w+HRmr5
fyF1Lx93g7F4x29OMEvo7I9SgjDZ9aRKiq87bT3BG1AsfQ+SG/NrL0uwzgMvc72Td5R3HQ3Ey6ms
ejE/v5GGB/7kJ1WseSbiFI9oi5v+OkUofk8RLAYnH/th9hyCnf1zl/guPFT9CaXaniuWxXARZjn5
JhxW/nJdS5YsxL4joeShMj5Tgws8VVkBg53aRoIpeRAW2QyFP8yA2JQsM49RleA6p5lnkcS358C/
BUpjCXLv5j2jbqSZMtiEgUnZqyMuaETsiTxAMd2ljtAl6DVe0EKYg1JfaJ1lpr7ZyUKDrLK8Sd4E
qkUHN4phZDvrt39lH7xpGGHQojpoLOLg+sE38qLsZpVU/6dUNSwPBqevrQ3JXy+T5Z5SMqICVlIm
zrOTLpy9M1vmahD3TxZdzeDgHa6hX50Sb4yHP1lnYuiQUhBJj1jnEmGZlH7Wd56h1GpQOLNoIwsO
YdC5n+VVN1IQ5yWrcMLqH/GijppbUnQlLwA3PPu9V0aC2bS3ujprOqtdAMoagu2uAksl9VqpDxhm
7XBMLHRNaUFWAfZw/BHOXsSPp2/RstPFBwzRBWwRVRo9/AOd3fgAtwjK46m7LspzZKUBZY4DAHqZ
NoMKRRrWKznvlJwW24Gi9scW4VF1HQbm2UOUwwN0S+WmhjOXV6mPqTtKpXu10itjgi7TQxtYAq5p
a/oLV5rSFiAK1lEqDrCLYVCTocRqn+YM6yFG4dtE1vhq55jj2YiM3cfDYvq1K6ytsFHuJdRKQWLN
F2Svi1HX6JjhTInQCn1s8+J27BHbrI0Y8OaQvQdZumIpn7g6yv+TdF/m8ictcSJGlNWLrdSbZG+Z
MWmRuQ1+24guPnelGy7Ym+8Dp1wO2+VXi7JaYE2UXpZpmPVXgfhz+cYk6zA/3Utmgwc0763FqJ4h
VbgwPVHys3dN8jbRtXNeXKhl3RKWoTni9/5Cm6XGLmW66oUR4x03RtQFMVTht2cwA2lLOYHp7y0L
/5AUhOqhmxNTXbI85964lx68lVgsdi/r94HRHtqnPj7v4pbONqomCyo2CPIx3QbWNiAr5hyrfhKg
SIZtdFoBxsHT8Zp3OR7vnc3vm//Sc4R/64kR6u1/KUZw1g4Pn8UCC4U6OK3hPXKMaR5klDcoA+Ps
nOj85/bEtLHX6zfhUZnW0ebkZ4hbQgRTPXQFQ1jbbwOFcIDFvWSWJXuOo+XcZoSCTUnVM4wUXcGr
JQDeb7BgK1GzKAgee+E3KpBE95Ukwx9iJcM33cxXtlkPrunnbeHOqb4gsKExADfLRVljOt0InJsW
RAP99Wkkn91bs9nhGnkEfcfQYpPv3MKp0WrhM0kR85n2tupik3k0xSoVJtC5Nks2G1UsFMivj+tF
KUz+zLf807gDcH7mMwF5Xold6ng6eoZ5XmN3qpYnbRycup3v0A8YqNYcECIHlKD9XbxGKKzGrR60
0M1jYrYlLsdMe56xzSZg3BkNhkL3XeZU/pNHeLg5rmwtmefYm7RSDfiBcxcTGTWayRmMdFVRnKrj
XefrtJEJPKPkhHBx+SFa+F4r6Ouw3Bxpaj5MOILhOSh4O/S9+9A5ZwWS4QOvgapNBQiWwQtIBrav
nLLGpya7vqm/WVvuZlBR4r8wTHNDdZaPDki4ty7oAPfVg0HGgTTGUvcNcbUxo7NhqilBJ2lRUwIL
LTZAvymoJGTGp3icARZRVT6SYqznFfh0ZRbcpTpCv30F0tl/RT0t5i5MtzJqiWx8bXZqC0g3KJB/
JeeYYvWhyWqNIQoqy8W8fOPjIoEgInaxtSjeBwB4UYxPqgdYGygcUH4L2WMoob39nBJmQ2G0kr+O
zwc7avMu99jKdoJ5bBAzSHWrfgql0SleOkYbqrAs7XxwwGVm33L7WAoeoeNlBF4a2UBLFgQT1M6u
4zjHVxGykeNtAwgQUfL6Lou3+43azdc3r0FfrNOrIX74FGla61IFTA1m86v7VyNZK30Y3csFu6tY
KkZcjnjcNzzhocdsTqOEo1djWNmAF5KWsCqcxt5zJaugrJbcrQ2RETNnhcxTMMnycsX0YRo0LY4g
sO1yT1avADSxhIbjl88xbAmvw4iN8zNYjuc3c+/O1+Mo73qnt1394lBgKkU/nGdz+ncQrwgNnARl
4KwPyG2DHH8kxnKjOUsL2OAK2hj7nuRYEkRMI3Gkj8jBBY8zrXDFeJaz20MWojmooSq4ok8NThbg
mpmmNzy5dP97Wfyucg295a15iPbeMN4TkXQ32dX8/PJGkqpaktnxHz4Iao0SbCF5WAVSrDMLixpQ
7ajxn++TZx4G31AshI5X9/YRMg4HNaBu+jPOwCQRycFCXskYbOILrTE7BeKRH7vtsCVSAh7noUrj
YTEXN3BOF2Zkgf6wbQ6hvtoEegwP3FKlANG3r8r3TJkjYU1cOh/di3vTV6NTdD6VGpYq24kCiasp
1wgM8VEYXVAnzD5HeJq+pdOAceWWS1ryP+wZb5o8oplODB8zcQiWnNpyAm1CjszmTDmU0YJ0SHkj
Fn/+a7cttSbXMYLZYM1mKYgJCCzAz3qXPpBTorpybd0ge1rtVUEdrIykeqOeZrO7eLL6Zag60S9U
82vIejYLdDInHGbCkdzs74GSakSRl0k86Rn8g7lEAIoeGZuerx13kuOh2xbiKk8BGiu4lXRsELs/
nDaJMiSQe/Gs8H6kvXG4v48fVcUzeNV/VgeS549EwGoL9IyLv0IPHks/ON9FI5j3T0MweZoj6bZM
tA4Cu5sb19TYP08kPGBan5iZ+g8wh2ho2SIJa0LBoezhg0DgV3SQXiD7fs0/LkY19y4fU9b7Eq7I
9+1l+GxHxqa08Jp/V0Ju9uL97agvnu9BFfP2NzAtAIaLBCpUAw0nE27Iwi7h5A13FCQOqGpKj2pC
/sEANsNNACTq4qFNoIOpYBRIbDlWPvpnMXxoewT3BQZEUp/Kyf+g6TCBF7egMm7qMPhEoJSgbhA4
EAAwLsH/6QJ910HPqbpxIVjG91yk9p79VBw9CuQR1fkC5z6n5fVJbOQ3ql9pqM+nghRNbkY64RuE
B5A9tJT1c+4DcqZ4bI/cJxglhRA9H6HtMC/UGxRWhzbJSgGzfwFD0FWaUNH+qWdF38aCpz7GSMXe
JsKmkxy/SOAEeucGOMe4HwJNjjNcd1x6GP/L4aM0jAUZ30PaS8NCO1puU8IIcZek6nnWRk779n/F
5FT9k+LZbJFOymCh+tSk66sioGROg8J/ilPuhBgNjn/lwLrMqj1B0E3VuLmm3hrawQGefNPfQWem
qgOVOw4nn8+FJ/o1DmUawK1vXSUG9cZzn66QQUd8bEy0GKSxmtb3gdQluHIngJT00iIM4SjzUySe
c6eGo9JlxSKfogLpQKQzkTvzrkFeaR82lVFqvqkjSTrkWSKXyqTeXObFybnjiWBTkcuABAAlQWOA
A8inKyKySNyjMIfXGgA/ZgXe/y0NjnFzIRjMuQEoRrxLfMYujYq73TTrpUEqWyHF9j69kTEn4yMr
IWhPI4bOfhiOeHgvQE5YPzcfzPEir79Q32qdF3IAJqYcz9aWM6X6bFgYUZD4vNgciZsuLZy44Xa+
3TOWdl0E4LI8//zU/KkW1rK4Y7DkzS5BMSalLpGIkxHauV5KVsvZi219nNZT6B7VSZz5MDzHI3gd
8btxlwVNnmoyICgKrcyoyyGO97SLeZkN7Ln8uHAcL9kRXL/M8hM8BikrQbJkXUurmYJjUyKwtoKb
dicqDPeluyuLJJkH1QSNejyUH5rrTZ6fRMM8IMljsKnj2FCf/XOj7kaRAmvwo7KYMAIhJ83/urnz
NpSQaJpOFo58zpnewhAgztqrcSuz10eJyAttUxuP9X69ZcuzPADhb0Ai1WKfTdvIwXvGTbc/tp+e
JRverQNu994Bga2bEs100ZKhYsGTY357qZnApeYdqE0Ak+7fXXK4f8fEFtyo0uC9BZkwXUVxEm8Y
3EdzHXW/IW9etR1iInYvnFZSZGtIlqrW0mpC+kGfdaW9mCIEO9uVSWQv3PkjaCRiJKp/uo3Nr/zX
fk7Q2IRhIG3NPW4Ggik/NGdh7ENjgDPKLT5kLD4Z68YVSsEmF0SIJjzJmvnzAJPnvhgO2b8fVhKm
LTsqqAf0DN6QnFHTmuELSsv+HuSncKmxaCBUpIVNRjh1LbIg2JxeQhZDCCEE7h6zDZRfocKSDuN8
r/iPJv0/VjDz97K7yhrX4L+BLQ4lJjTd71W6ZzbGQOZYWk/40DmVuy98zlfJK3OoES6h3b262hlA
8G6QA5QYIwmy/selcVgOZTZGua/7V47DJdhO6sNqp93//g1e9ItKmiXE67uI8qgTL/nF+uuSbErG
S8SkkwMTWNHQ4KhlsP/F7rNl85bDTilLHXCOfELKRuojulYBPuS9IqNeqt4t4LlKuiOQc+Vd95le
NXoFv0heRd0qMtsWYy+Iih4YrBrdh3wl9iV1l1hVd8mVx/LVe3Sejfwwg2AGKuWnBrzEjwpa9or0
5MgNTA0SCECgJXd089Mh7f9nereRvdpYZb4hS0jFrVYcJLoq8M5Ge1+CUpD+/F1pD7gz5Tvkp7vG
PcXdth2sl6GqZWTbDECPF01DQ6LFqsts6QicslYfqkyQO044+oWNRgU4MnRD2gUqBl3S0j6yzdgx
D+e+LgM+UFu31ZKr9qbNaWGtGqnvFbbDLCvTnIsApKQbUm0Ud/x7AnFuH+dhfPbrDbqPmgwK6ibA
x8NLe8yaoZYWbLtIpbV3jzzFauNSWsKpBuxnG8xWZsZf1tdK49oSCFh9g0zGc7v1BH7fVvTUsHHT
Pb9HPIAKEWiUvmaRqUIJr7dcijeKDqTTfbu5qqYdXMEo3WshxfQr/GP4Pvtpmk0YfrOnn+Vlo5/Z
of5x4L6xksQjxO6gH4mLdYO+RtHk1H4t9jdbFleo55QCi0sKw6swrekS4i8xTtloA3/ajZw3aOBu
fpriFWqTDoLPSEf4dQvANyhdqFqweF+BzlL7wYrnYeL6jY0WHcgCsRWJATyY9NsrEarpIKldCWrD
DvFPbIWZh75/FvCPGIewx5ua8il/K8GPvU8Mm9L0oCXzmvOiU1Kctu1M5TrnPi2fU36uQaZ6Qm4O
zURmD/Mfp9b2lQ7glHUB+Exej7HO05tqOYV+p3J0rz2eovDgrHYjnBm3Gf9XAgWShUNhr2SjVNaO
nCppDrw/xH0q4X7yDzPahVjrFFx6mIEaIAq3hVQVzXhOsxwSsa/+eb9fz8SqKRMfHYm3yDmCEKgS
lSK642M+3Jqd7VkBtxW7glNZ1dvkTYd6lFS6UiGowV7FSpHW81OEVo6MVOYzsVr/Gr1cP3aD0juc
lyYoa74RwCb4vqM39czUcwuwygvjq0Z/Ovz8nhZPs2kEq7qus6vWjGRpge4r3nf2oalH9kRpTNYT
V/6MF4h4MyBO3pEX9AcEYDgqFVUmitP89pfe9XDcam3UlG0YSCj2bkmqckzfJLcd78YcY4r2fH/3
2Eo05d8xud2oiMQqktWz6rSELObruK5uZdHlMj5vtdXGOfPxlIyyuDzLKlMdPoZUqnsPmPu1uKhx
q11RiIu36ZbMKpaRktFlyuI84VAfbJ+ErFVK0vQxNuiZSgqOf3w0GpeWwkquUWn5np27ZDs9ys3U
pUJctXJioohCQYYMZfpwHg3I0zvwLw8GfrwhrZuXxgTMzZkD0IPkoNYpvSOmqDPPPHxZ1/5wd7cJ
osVeUdjOLKlALTkj5OJ7TC2b/xC8f6Nw1cbZymmdQffnYqiXqFVFQJlgnCd+T3ZvW5WCELZjnx6o
7kKxViWUfA5A5fg3GLAlIaOLNse4CHG/8H+CN9LJ00D3twzre31F1HAfHxJuCvjIzS1LXmXBE/ns
B5DwGIwCUEeNMtwPOIXONsmdJT3XPfJbDB6AzmrYbaQTM/W/scZAKXhgIB4XvvH/y3fjSxzVn/LI
q+b5FwAE6Z9cKWuks0bzIkCCtUZZSkUdd7lexOYEjI1mrZImTx/fke0RaqhiyAd0mVNDRbWIqE62
R7k/99urKgFAq6O7MnR7pnIFck0ynS53x0p3BqHWV+rXcWFuV81hF8j+3O5Dx0lxYxD7irojC/MY
6TOYPS2tneJC7M0QxMlzvZhcpvlYL7bbowIQPrwta6zS8YU9+cfPszODjO7zZpgZOOZ2G2tq6pbv
KWxyfLNWleA52uqkuMdEtKSyXa3PJVoRfTkz4Ohn1CpKz0qlS/MxX/hcZej6pMSy9GrOOskmLpOm
3cPmVJ7Qq0SEbuF4DUdL8xh3dsSnuJwSKVEIP+gzswj2knQnV/kCD+rYRxOoOb1j1rxwNb0gXU7U
zV5gjb7ghqz+Th0Iha0d345SNoAThPQ+BzjXS/I9NVim/gLZg/Mkf1wjT0x+2Xiq5m7y7OlgcLv7
a08r4/i9BYVGp00RkepCjn8bjRGyvL+V1xXwIIYcaEWULssDPuCjcG/Z1ZhXzORMIlp6Vfq3AZYt
+pSL4fhvhvcuQsaJQzpju7GunV2kVil+eB9InFJBmcsHECh9sphwDGVJ/zOj71i2xO39xgjBKFA1
lLn4gAiSeqvXKFBolMXlITQKF3aFBVA0pQ5h/E4z39MxPD9BD4hPuCcl8PtOcJt64GHqvUd+0H/s
X2R5kYc2x1b72qgFXbpU3PDYKyl0AkDOF11mqbE2s+d9gpcdFX8nrDMLnJPw7oTnfW7bmucmQmeu
JTqgCz9oTf+WeLYjuAmpg5hD32MiYrSdHlgCs89uEUrWck+zMGMnKCI8Svs13iNxM3WU+TCULeNo
VUrLfkWweRErtm0FCg9dmmwehL0ffgjcCfopL9RwHKBHD2WfEHGUkk/xNedL5Un5V0WLATRkLV4m
sTXNopjv0zvB/H2Q78KXPXz52w1UG7+oaS5gk2htTDgDIGOIgqenafSLJncHMheB8KHEobDHn9CR
1gEdzSLckDXMhAkaB/9je2c+ckeFImBdXtZu9xnRlhyyI/bsFMkkCtie81zx56plcZy5VkyqPeFL
vvY80GaMT9I6UUjG7xqFjbmYq35J55p0jHgd0pobKSMLe+XUk9hAyzEoRPbuKN1MR+soewR3S1th
KpKRkF11Rezr7Ax6EmbEGzRXlVpi/dP7QYwmMuWb3zG8NnB253V92CdJ36S31FbkhbzvDE552+8y
95HJh5oDE31Gu23vOHn+v2HmfLnXKckvQg/t2cv8pIKKq5S8wGn9D1qIlwBqmJBxaceda9nq8WmB
BValx7RbSxrMpV8+vTy7OqkNs1EEVtcAueUe9PqNZ5htYDJR1izg0leCmLJ1rgXIZpk10Fckw79Q
bC9lv0G/yIuVA0LzGeIKKV+GY/KmvK+egfpKQTmcubHW9FOGFuSPKVn+IqDHm5yf8L3TC6tJ1H1Y
0JCpDxFmGR/Lfixf+FAY6Eg8YHiT/14RnDUMTf/A5S3SyS7ddF6iBBxAgcqAS/gP63vPKZZiqIjz
Nw/IvDrH6Jsm49oZflcC/LKFhdJo3oimNOPkjt7TYv11APVMNKjaRl1g6xHusl7V7dO4eqxNfVDn
7juKVmN5o3oO6hRWp2BEdVXg932Au/l4OcrQdVmCbZS2ZvaEHBEL/1JE64mP58fF36k37jsyrzga
a4rL6JgDSDhiUL6bmIf0J7qvsJ2xTooftI6ApHcS3Rx5g9viXCZQRSCYwKu6DjVNOuhA4UiOP+Dd
dsSUwT6yqk64vYjQc/LRa0mPyaPwuesy2fpvOix7ly0ACmCcggY4n5pmz7JyqpHw49DeYTD1Ijwu
b5bps8UMF7ftnYLSXCOCYa6H0KT2FIut5evg/FVOh6wHuO6I6Vthea32pP18AsMDOpu4X2PsQlC2
nVSZUZySCPliionTYlDQz5ez25u04PIELAXHWNyCcA8kN41r7ujfERUx36XoClX5Vx0kqsreO+Iw
JEWCHRlF5Ph+dz2azqEAhJc0Kg4rOrO/AUcgvays9EpGy0uATfZKEvLw0SCyJpeRs7VusBkRjfcP
4tT3MuIVPP7FDtKauevpg74VRVIRk6OQqRiHlyASuFXlvSsVr1DiYl0XgGrZ+4UYaE5j1l3FF62E
wAtPwsvI6SzN/7SWibIvgTozqwKqmYhMsCZK5xC6beBMCbilBW6vFC2vLarhn1bL2ydAlcCShCJQ
IqdBrzoAvB7YLMA6/WrgYzg/AG26pHu3nI0w3UaE3pYa5WemEiqHWhtp48OiMjL9k0lMobDqfdse
rV1oZWbG52+7BmnHF9yW91R74UczSVSfQ8qfMSjIKaFzrv5KnwiUxP6iqyMyzI4EJ5n0KuGTMJM/
U3r4MlrYqdxmMdJVuMuooNo4a7GZ6v0JvkD+n0CvYlw0lApEsO1tY0Wr6kugNBkT+4hv3JLe/zS6
y+OVLZpVsVn08q+veZKa0jYbwVfkvZ5WwHUMgcJ2S2wOWjdtFa+YujJYgud/pOKbf+MCphzM6+CV
bBiiRJUxm1dFhYkRuWpdcvmkwDyM7oy7D4/LRR50o8N8MByTIc28+WhewytjMDBPIIPL+kCM6rvD
CbMMY4HPjXqedmqKVLbhM/e5YzBXhqvQNexsEtpnOV0Ycnzi6HAkFmx/9zCIxKU0mKMCIfPkOkrM
1+TlA59TtB2/NA7CSm64KZ/b8u4UB/+Yif2W2qS3DDVmZ2QhZGlf1SgZZRQDJEx6dCExakpM7L7S
jtdmyHJUQf7kpzuXXv+QP1Ad/VZMUr7yuQQfmg2vY3S8V4aQyLUH06qX77AMgJGYCIYqJcGAKYEQ
NeEFFkYE9MxgXTXiyJ4+5wogyGUPn7jKxLcYhbeSkNlSIDQWB+mc3dZoA3bFaKnKQx/qziArcqr0
tVol1fW8vwzx7bw5c/wx0jBS4OrkG0MkOTOqGhJOp8TmDLWivLJVF9uTV0P6drhE+ryHmG5Wi1NZ
iiRvTQ85rVnUwp5lyxixEdt4GfcdqUgF3FfwCoV5JC9XNfvQGXeCpFYCdIpTCss3BlmcsID+vc1G
xwLgLVxa28IPCEPk3giBWL7NT5LhcbyHjgVBrd5xJs7wLypJe3U+8ZhkdcFcVRiV8PtMMwF5ahoa
cwKlHhqpWAq8tX7ad96VeoqnzD9joYFMFQ9Y8aaPNr5MJ1DpdiWEq5Lx1jMT7NwARuM4G1gEknln
+Jdgq2eb9QJKAUIkQezJNxqb466B5wbJmnWzIZvdGn2Fq+Kow7DbXPjDmnfETly0e+o0NzDXHyNL
wA4qvOK+yBUhSJgHarBazKLfl2+o19lIm0p4WYG5Ta+AwsPQHepXzpKH0Vvo//5q3s5xNp1RnHel
ef8wlIAg5FPhDHMLLvFNWiMyXZ4ocd1hwPg/GCoSU5VmBUgSP/SpY2MYcVpFnPJW9Mw0r46EPK4S
1HJo0kQyzGnCIjkFUwdLceZsS5EB85KRQKMd1mL+vu4uylNpRR0LRTIl7BMZRGUtxys7MD5aGhKg
I2yIiVxMWXX2CiAZNeCZyMH09eL5G6X1IgYIU+vl1BBG/Wls8tBqaqx6xgtCzH3bncYrEajvs6xI
cGfCrUKtvLfLViOcWu3UBdHci5/AvviBmXcgII7Fr1qOnr5P3xJdLrzkxYD6XrQYCgnm5vtFI9lb
CqZKhbjptkvo0ljhIrGMRRS0JZ2Mo53GI8TYqmN4sa46+6JRM7z5a8LGfyL8asUktXbeaLRtQpwE
CQXcPrXTFfkRL850xPDzrBKvf+35JojTetpAXuO0TkyHpB7C2ablxFBR7CeT3e7iV9WOistkwquE
3qAgI3eBovyjWfqbBpAOR//e3++Imxrj5mlEi5916elzPixmIQUdRgxMqjBLr63SOLrC9bbovOkF
Ohb6oYCK0Bc4jGCoOirUbADwqeKDGcWy/9//PtvCLX5/FxFpLFCBv4jGeyDDLQ0IAkm64cO7EOSc
ePsggaSgB7HTh0XD0weHsn/Ao15FBSaz+SU8dmLqV92BQxIRan5AXiprMf16OVDUqq+mHNM+oVzq
3IcjqqzsNKkVCp1/V1psEhKs0VtgAbhgPyCYh7CsOmd9X9Ft19S9XizZZe+O2XDLEYVqhCRU1ps9
uE52NYDZE/Fd4Ln/P1q31hbP8vKTePUjHIl/W0ZZkxaBSX+kJTcmTGX5VaWV1HGb4B8rLQ0R+n+G
ydpZRN/xdkws1boQI/mtJiPlKVma13Jt2Rc5GzqAxA761w/5RZQtIcj2PeQhZhSDM1QKOMrn0jbg
8TAhTvDmbeOA/wNIO6+qS631Q23lZlLKdlvo9aM21yzucUbsbVhhmhnrMTVqknF2gAZXd3XIp29g
Sh1olXMPO5PasX2NtpW9Dh9V9+51fJkq1HI5Er1iCwIpZ+rJQowwfvb/gfVwTLBe9FXc0RsKlmzh
65EMQyIPAsuBom1tARwT5++on7bzZKC+pXJ/nXP93ORcyxLSf0kI9DAh41R4RBVUA7o9OihH1izh
IuOm6yQhHaihnN9ONmC3jXHm1815+SZk8oI/snAHZjPjLfpRGKj/y5RIeSzte/+ty3BiuYrWU9Wv
gFdQrjQIRghj3oPSs8XTGMCnejtJAPBZyRXwWOQRVK/N/JtxTzeG+3bb+SQxEVZcjlojZJxAFfQz
xDsdmjOGAHCYd9NPe+DmN8eTLvcN/LO3g0hSGSCXKeqqQRckHRJ3mA7gXHOKrdfpTMx0X/gNxM6w
kMKa5A1LjZWQMyfC9QjdxMaGBCLx+D0mywDb4giGdV1oe/eHj5ATj4w34Fdcp9X7nCWTJW1/ET+q
mYf2SuTT3iMGIpAeUjN2T7B07Sx5tqGm2fw1qqQ2gn9ENjfpwmp0Fex282NaDaF/QMhgxwRIe4rC
TYh6vMBwmL4h6p7jzMpEsgYl4IudrhMuDNiBTp1NA0Yt6tw5Zq73RLssrUehUQpHwQ/L64il3HoG
81Voev+/c+uS4SUMoCa68rH4aAHDJE7BEysFJSBbfOFgYnmuYph4Qdp7bpexYish4+ZwcMbvZbWv
v9nas9RHeTTzTUCpzh/I4z+N4TK9Uhgsl+3utBEedlCc4EQdRtmrWynxU+sLHH92UL0w+rvJAaWV
k2t/74VTItRjLKIP2c2L3QwwVphG06R2PTYC/jTjCuYyR/zYTs9N7IGcwsbiyu/0X2mgKLooXHMf
qQvJ+h7WpeDSsjQEgg3Xg/7KzRWE/Z58fvKxwoHCynIRiDX+qaRhk9PugVmA587wd1xmDuEZuxB7
Ab6FjXd2pZCJV1leuya7yYrU0B+o0069Grfmu5uB1lqV+G1F16wqP43M1gCvdSbrCLkLS+NET52d
s2Zxmm90V2pCsLFCFa1uMbGclJx/Ucd7nf0CZ0VQpTFtE4lkTrysbQ6/lmQnhjwm80kKXMRT0jqj
X4sKKP5AhLoVm2Km2m2bZaKp8Yk/lgAAzynQAoloZDWlbG9NuP/BxeWm4ET1s9geOMFM0SkhNWKR
4ftRz0SbGfqfiwbqGgOLUgk5LG7T6uOv6gAa5i8Ol/9nwO60zt1sbyj1eJp9ybBe6+NaixE/2iOl
Qkg7rJDNgctYmUXu0O3KlVeX0JZ2/bjiqjHCVe6kW69IMoT7FgcIIj28c5IeWVbJKZ6DljcY/MsX
Q8cc03Nxkgd4v115tIMmdB18Ry/ji1D3ev4NMzfN2jnQ2jUm0BYpyUVJyylv5TykLiLA8Fk++L2v
sMUagiziShtS2vV9Ehte8t9zBuGCxtmEX7Dx5LfGn7UVGnsVBbZ0Ufc7a8FNQ/EMyE8Mn8jzAEIC
EXRYAUR4eQI/Ph8+lwLjmEWKmrzO9M2PDh5QrXdcPpBbJMDwEtqfxgzLNXkuu6iFiidIOHr4Ry7S
7rFI7dOlTTGZnHzAKq13JIPbu983ySHqvn7zZK6hZyYqvTcj8/F+w2CtyGBNyNFUSmGegRH64DST
ostiko8+fNGzB5Cpp7o0HQwytTfFWsnf1AjU/rY4ErP1xKPd2/0W2HmIM/MWblw8mnoqXbQRZ4Pb
Okp8l4DUhW2h4C68CF5OqPd7ensEFXCQuhJSMFLqYDsrN8hfJDIzrSCM/6z2FXc88OUz98TEZgxO
3AMJ2nI1eaMJhJ1ECbA3/3e605Fdyowd45PGFSqvGwWgyQPWb+dRKfUR2EihSV7ZJzLNNYqWvG34
gfFAVa51g7ZBoReHWQUBcuGYujZzyb92NBWzjEb2IwEVTmFXjsbY3jSekx6DqP1qp6ccNtSkjMJf
xJ3C9WQ4hpolXVw81qIQRkxxLmKfOQxSE8abkeTLRrVlJ1DYuBw+THkwx6IEZC+myukOiIRGATme
v9+qU2g4LNF1xipCb7kcVSYV9f23odUZRMfx2pQjDp0lmgBMt/vN5wY6l8tpfyUiBWjn+ffc735+
qwKpL3kCobjHgxu6GT2Qmhb0sF9Ge2IMqC1hHuQNoywadl9UfM4MgBYc83NfJCLFd5cRP1yheRWr
CxYEsdvtxZ/jwy5OduXoalM/eQqUa6NGtSHue+7nJFbA/VcOiNAPGiQf18144RlU86RThBgKet13
MwVH94hjdMYgEBxK3G3MeTxuJjzxWSKy17LAE++FIx58jtG/1XkTTHnRAi2eWsiXGFswIaynFwa/
cQJX91TgbKMKFhvwkbrZ+mDc824XOIrOIdfKl3TMOFPKumkadFeC/owvroBSYWAg6MWZ8ra+jBip
OSyrrz8shJzGK6D4dbQRTrgxSZVuTNzVmWXJtWung4kT7WMc8WqZ7B472xP797mWI10DI+DGH06X
9BgXeDglQdTaXBYDaY1GNo0z157YeZ5sfjidjee31zj1EB9ahQnn43vVhvKiHfc2fHDl9MyuuODT
QprOSpII/DPNYMGiOEL4p9uCiV9okSFad/BATCj6Egd5HcFqdmgRsTkjb3fL4lWUspd7KRwCoxGK
hLbyBvBMP0duhqM37owUhYdNzkxG9Nu4rFgRavbmt7QVzLsFZD5pq07UHlxoFRdcr1/MWnNUDjqb
pxOZXSZ7YxeBOp7WXs0wjEfhh37Sn+PPrG0XMyAY+C8nRCM3+2d5i+K9tEbMbnhOQjqDQ97vEJDP
vYbX7aFJLWFAKuIZA+WcwxboGqg+20y8Cgf46WVbktHWLRDiLsNafyTNTTktIf/dbgSJKBOVaOqf
Yi/sW8i6ejG2TThsexiIlCSLAPKXS9EFpPA1QvR5ibFTQEZ4D2NjDZt6q2KaL+L+RtfRdl0n+fSv
ccSYgW+PCgMlojmmTo+iY+EUMufAD2ORGtu1YH5f48qPrhWMAWdG5EzULQ4TsHYwDb2gp9WkMdA4
G3zV4L+pEJg9gvDnDjFIsNG2ALgVMZr0rxDp9HAqGE2EbWP1juuh6Lwob0V+2Jd/znFTy3RUHNeF
OPe24FV7KWhySSl4wkTCy6Os7a6XpsXixxCaA5SqDpBr/H96gUC+efEJONxwSkXG7cj1RJwsEiPG
0qMqm11vMx3g0EmkBN/H3b946QvqteII2RpHUZpOTs28wt9EbnZ5c3GczYv+ladtN0J9a3dtg+eU
TEvG/+CjK3SgdlUbUNKjdFlEdA2tW/d2UgcaGg+TaedcP6hyWpVR9CclrnTBSFYHpzD0F4F61HcF
UwsgCim9h1Kuo1vmK4IMeBVB7ha1mvJgS3xkZ7qht7WX3m6FEzQq9vvihuF6lbOWF/SpL2pyJVPa
Yjaf90h5zZIrrlSx9HGdUladX+Nj9huxUTgNMS2aPmEb11uzcdtCG3YZ943iCPBGSZwW3m3q1jRg
ytRxNuy0OSTgmLz5AhnrilmRZ8DHZLWGBqcE2mqA71cUDTVk6QZ8djfk86xeDKs2bWH4L7DrE9hx
18dUVEdrDv/+YobJVxf1vlZWun6TmJZxjdudzV6are8OkydW1wDxXJcjiimrVZvpfjJeygpn2HUw
qk/jFeichpoJoQaL+4AQ0cPa+zd24GdZ5OBQf/eJ7KAvwS5eY9zDvC5un5Pw1UdzexYsWBRhNU/Q
crs3cPBVM8fKR4FazDIDHR1jRg21rrU2J2pE2kw5f7Rvf74buoc9qj3+Zl5jaj/EESG0aNmp0XyP
o5omc2mgfTR1mAqJ77YRG1P2wtBtxakFcz10zioC5cRZPGm+cx7qEEOpE2ppdlPqObki5Qasa/Wz
uMzNd0aQLVZssGU+r5coHV6EBFolTEpBzGdiDPfkUrJAQO+OXCumDfL2c8VeH6gTNA8luSkSDxwQ
E2f2ktQB8wykWoKD+UBYZct5POQW7qlmFCjw/vga4B1oRtXSQKF9y6E7LRqmH2y00N3z7WINn5XC
UUnzvd3hJHuntEjPi1VjIzYVbj5L5m51Kfb06yIIL0Td9B81gnroQEErW2mHuCYaYKJwObw1ukY4
OKNswIoEReOS/Sc1z4Oy66oHYJdCMIowL3GdkLXHc7WZG1iP1RkkTLMgGvrKYhfhTMBWE6QXCxT1
uAVmzOE8aXJ18udvy7YiIWulzWwAPTiufyYXJgJaoLSrtsZK/6zKzjn+60FLhLRJqRbQnN2JX0Xa
vN2eEZ3p56AJkxLfMRSYG/CV85CDt+f1u0u/ITi0OintlOrcKRqFSBb2Sgs7kwaRHr2asKP08BCU
o5lTqVQb/cJPcQrmclMw/meF55ocnF7NLIGhJjLpMSl7/BzG1Xlp5JgTRITtrtgPAn9Q53l+Cajq
6BOOm/quRk4b9yRkwFnhSfVsTglXJqJ6Si/QUlgWfG/osTDRiCKZppmpVkrM6BJw4I/DM+uzDVSw
1gdgyEL+skcVSAk8OVjkARUZwrMxodXUY/QyuhiZFM3Bgad9wr4JqJq8fkPW+MPkBgqRdz+IpF4z
GtOGZve9Js/RgNgj01LvO0MXUL7iQzVgq8xNvqHd9u7g+U2C50f+/6aHFT4mLVBkIOaHY0TLTdaQ
kO61yHhbIqBDLDFWD8TGgEePbrtu47BoGaNjJOh1KqHA8PTCGKdP1zvWMnn7FFV8T9oIxgvrmBBi
Pp7LK1AXMaSzsW+RlYXI8H3W04o2BEYj1i9hft5Y/V3tg1xqBLMghHFBynRZ7AWg+tbNLIdGJckf
dp5mawpzM0TW8AM1uRTCygFHROS4vbAejApqlIyKESotz2XpSAh4tyD99zZCWF9MWSF4h50g8Vdp
jWZKAK3Z6OFdRYBBwP7DMGjxO+6I8H/ckeHCzrnODGEpfq0x+LwiEoe2wXbdCBqSWvGYP4Gn0RI0
DhK7xHmW9J5rMmf8ZuG77IcvUFJq7jKI7H9Q1DxSR0zWpMJpqGj2mPQ3d93UrV7TV0uATa61a57W
xyqkXPaxQ1beRfgX6iRSr6BdrRgG/SNPIgLTrVA51s3lmlNpXnueJHI5AUV7qykG8F+ATt+ptnI0
CXo9xcLTA/TYqpjXplR/NtKHYEbGP1xnFtu1u0oNEMJCCmJkkhWUHmsWBMPUVJrEdy7wypGxW6XM
imxvR8vaGpPF/TpV4j9ZK3jF2U44IPTbGkl8koMFSEJdMm07onyyU1hcEbJyR9R27XySkyXcy3oq
iBPAymAZsMOX4lujh9sKDiryORImEeHDA39WF8528e+oFHjn89TPNviOOkx0TH0qPbrpF5ZCYxhv
RPyg/pNc6Ioc8W9XtnDBLFhitx/aWY5yt/2jYohUrxbbSKHvYjPQcLwejPIGndpVCv5JyC6YxuS/
/R+actI6PdzxNkIerFGx+LCP940k0RspKSUv+lMlETew4jOT9OnM/owHA7cz9s9TQE2vR1cb34uj
j4wj+td/SDHb8i5GOicoZrjKa9XKrCkGf6IKFIzAxHLWtnbtNGk+Sff57w+DTazGl5SvemkNwUrb
MVrZnBdhiPZNKDUDfSt+VkXBamPC7ONqy1LMEjkFTlLU1KSo3+/WP1TLY8yE+dLEqQlRALs8gT3S
BzZqSi+JSgrw/C88WoeiKjz7HwfNXb5Oe8E26SJAjQj1gkN1LRjblbpK5luNKGOhWXcCinddhN4F
0r8wsrVdXZR2GQOyL9k2CeI1YK3Ll5PgLGXCPqOtomYsuHDXloCGJdELAYUf8URO7Oun5SraWfLH
bQr5SvG9LKme7/tTu92JRMDC2j4na/RAVVxwgHhGxQGuwFlGGAT6hkXwd7Fh4jYZP8CURRmuzwH1
NOezetmdTKEEyP1vnCo00OCQg88HlYMKabMCtpkIz7AiMb5gOgca/k/mN2O3FknN+IVaD5AUpAMS
GA7M9rKJjb0zDPmWIqN3Lv2DrxXmwqpThYHVnY9YsZevHOFg+WYe03CjjFcn4+6bXbisg0urTIYV
cLSHhY4Ej7tIbSizR0k9fxt62l5fj0IhvTapzvHOML/WAkaIbN9hCA8DJd0TQqkdzzRUttPlxY8k
XiM1lNasTsJL4xHFwRKhqn2uZICZATToyxnDeU54VKXlugWiMlZ1N9abKgRoplLfLptu+K1VIfl0
L+0IKC/GlRBI0UuICFfGxXcmg5lbFz5JxikM9XpxQ0VxxRpMEP2SvmmzrxDeZjvDTXhagi3r9jgT
i1Ycc7TBSXgcxd+N0GFSSCjwDyYOik7DNr8LfQBS0r6HFyCh/i/GJxu/adcEyggGIVMbXS1QUEz+
QDDznZVN2Po4T98fzAqEKAIFSBQW0tedd7Ulx9HBbwTOeiXc+rf0yolPy71UAOralY9CmJatJyb2
u+XgxTI2wfXuUcUTVkL/qFDPi93C0WSgWiOvViZEf2t1CX+2OUN8fUmQLF67L7XeHyo5tJxQgrnJ
dStIarLE9Sm9k7/uIsIpuhtbtnbAhRPcvhLxjGWsUir3vyF4/8Jhq/rVAqAdksLG1XXzjdqMX5Dk
S5LLMhkYfh+wVVxI/mNrcOQLRFepv6HQNfL/psS6WjQT9SN4G+gfssZIMEMCmaDm/b72KIJbghAV
kwKPXg8f/ZdWk8ld++c32u3kjqNTfMA959dwTuX9J5c9Bfl1JH75hsO3MGm1kNvwsqjVXQGEjdnc
c81HXhgEg0ulgEiit4XgMrUBkwSGYpkESktVLtIoIUzSoPip4p7aMMxaTKHqyNzF+EdiQzLob55O
wP2lydG8NouYnQPiyAaqsXIfAapMBdR3/BKlbkpYJEQiF+MM3Vu5g0a+mi1BkLgLvwWpsMy5XlAD
elAvGFseICxP2xoZEjsZcKMPix7H3UQ2Y8LfQmFCT59dBraGiCGKLMUJE9nZsyJk0XPQziXvz/uO
xv7m9d/1jjzgyUazXRi/CTr5bP0HZR77cJHRrF4ESVW0C5zu5lpWWpkTPTaK+BhE2YELDFC4vjBZ
/8hz6gzrlwO9lOh58gKUOvCPesLn6pddKVZbsht2F/6mPcHERA9Rwm+mlcKpgf0T+rhifJY8KVHQ
zHpxJLRTq/rq3H+G+DHzZLNeGdLNahiYKrVDD6ZnENyE3LO3Ske8m27/gygYIhBtLO24B5RP7NEO
UTNVVoQzLcEBzfHU4VKaVwxhnSj03ap6Oj6BaGQiBUNhvJg8WpdheZzdqXTqYnOVNG7zim7sGkIG
gMKmvfutu1Y1ftpRnYfmdwpueJQ0tkjF9qZmVsVLDkHMLtL8o/eZRQgUfS49UOU0HFLAxW1EqXup
a7AkmGEB6hLjoCkdQDFfxdyVayiJwPcXGWlHHAv6F5Vbfqw737f1Aw+tltzZBeAkw/y2A9m0ZEUC
rlw096eX7LPoGr+AA1ivs2QHdfFukHehszBVxQbCxWRBkyf7PtDV6SN05NS3ogoPByWYnaA9/SeM
ux1zEksl6Urh0FA/btvEcD43hMyzuAuhK3vS2D8zVWSQOiVP0h/7c0z4XwHej5NQDtwWFv2HHzQr
MIfHJjdO5EEPxyYCiRSopaEklYY4k/KJrYxy9Jpu+TlS4FMfk7LhVMiwx4X6Hc1IEfGhTXl4vQVU
nHgmVBf353W+0FPj3hXMSrj5KL7M01qHt3fTmhYqHg376Qsn76F/kKsFfDxKaGym4SY7bWRqhamy
jEQSY1GoUH9J+jWijeQFG3+wTQKVea7F1O7gjvZaGWAmg8NG5Ikr3IaHkq0BvDIgw6FcdtiWV5ll
NjuH5UXeqyjWlZ4VYNdV0yL33ZC8fTZ3dVzutl6ZyU7C5OLDpsl9tutD28kqtaSTKpzayKn2kcYb
njvfINnAjdUCnGaebaFrwf0mroTEmJAXJJwJ0rf4nHYa3o0NtveHvJICYt7JQ92arlL82Ij9JEzN
uAWFcU4zNZunkusti1CukdPnn+I0AJXNhIwmwpJ3q26joADUgbFxy0H8Q7GHgsmWuZacUUTrqtxs
EJaoFFeeUGmaMysujEGZZyTzEIjsfw5OAOBVL18Ol8TzssNKIO0XM35T/dL3W59ThpWivl7ySq1Y
GQ6H9I2L7SRpqlPHjSP0IOKvuVlQzpZ6mSOdaz4AygTgErpiesBDGvgapyFTosfBx0AeF0ljIm4w
UQ2zz+IXyXDkOEXtw6HmeYYzTwrmWvVvykWGR3RgZMm0wYhZ4D43vUp6+BFFwnYO1+S28YJ4IUZr
+dncTgvcbBIeDDDIuBWX/hGDM0hELRnJgU9CPHWDoDMQ+Y13Jp2L4gT0j9O5QOzENzdjwRflJvb8
fVs4fUv//0uvlsg/apPRcIGBT6c10ckcxsLhC1Yq6s6Frf1mzMeMTAG+H3wYIXZawfPo10pPVA22
JNr81zXMcW2ZtZRueev3MfkOPkLSX6R2k4tDF8MuhuF3901TRwBgT8PRd3CdoTlrlOf4q/KgdAog
2JUvmw+vA7AqBsNdNa3WERwpusasBQX8E9twWy/IyC4Ivd4qC7EfzofihNSKxjJrKyFo9TXal4iZ
sO28thVglmaXAoEeZ2VWHDdAwGv8iPZNyd0Q9jRpFYo73YpeSr3aJAUSxCYNyuISUbK/7mCOKpXJ
gN+JADKejBoEw6WXxLQxvuhfmfwOYQSQ7BPI7bDyLj+InS7gL5rjJtNDP6p8ZJQSFGEXzcYEcPVn
YTkfWR5sSR/IYZhMM3Udg/7+qgZIfd0EHYJhMkZNCxlEpbVEdUUsCxjmf9UUR1FnctBOc+OzWCjE
JLnAG8A1uQ1h70Vwynd+kaY/f3vnnKMkGKageFgMCKPMi/i93CkX49svczt5awxBSnLZ2JuSrPQU
Ll5uSsX15raSK1AHIZAlORkktv92jWCk6q3Be5H/qSiQvQzfEqipAJuVf4QEYoL5E92KOotuH3Gx
ZOePZ3PGD/HqttPM778/x9twTn5GzCK/1ISt0JfJxfxYwO6C7uPWQqNlXIZgQm0xpJXyfGu14LXo
rrYnrdow+AHPnRibfVE4cDTL40cHzBn+3uXaKtbViDMwSZrNu6dVQeS63qSXAjYK8p0/t3Bm8qF1
yxJBRytJkDSxd9LbpqVSm4MrUWpwJOo99LlkhqVAPX3+af6CbJQhMjTGeTHY3xdrnqmckgOPV1Ch
yOrztOlyeTCZLk27usgfPFwhSjOTjLlwHw/2iexdPfnWunNvVknGJy+P8kxLE47V5yP/a7mNg810
EC2lNrfjIr6KPaC7IqolO9fB8hFHZo9nRLiOhQBoc8o7MG8bjMiWG5rSpQw7YHDAwJSmozPeEmol
m8VDoXjl6Snkqj1AhnQbzKVB/IkXDo0/o9XKvSA309KKL4cSw7F1i4VzSstjA/NWf6fIGsp1oo1Y
85QM7rO6unBzIKJQAvEMeePLw+3vLGb2RAQ+JGzVcyb6ZH2m8HvlHBod8eU//BnsOnyNBWwYtjAc
9Wn66Eo+tqql3/K2tMozNVya1qu+AEwJgvQGjkB1ldskYpwjgT0x9ZBkaqKJwDFYdOq7eAWmt8sI
Z3FI1BhG6Qv25vMvGlnU+LQHxhhOLX0u9p4CUjer/yS6IbGlEnrOX1HwVTcVdvftbSxwZUVjMhDw
Fta58qvS3xOFqBCjgfIjpiB2ZlCvXnPZWHyc5HPr2z4ftCwjEiZJtJKQI6AsuuIk6GzJVJDKsCXN
4FJvrtKV9Tq6GhhpwYC+8QMcBw71j+TFAI4IoiSodOETMYgC5GkXOJWfPEEi/lW5EczT6AT6RfEv
ZbyLbjVediFhwkhSivqfWQmxZORIb4Opoa7SGZizQm4JNlEsedbdAv6SaEMS/JMeh1kd7/RuqlFn
1z8Bado7I3tHsFi7EvXdxN0+EpG+Wo3DG29zT6HWv1WMFTn0rMSK9+tXFfqJORznwHr2Mzq8vO3W
iFTroMaNvb4o0ykaq454Laxb3ceW3+/TeZ5CsZSlL5NUhDYjZJhDdN4qrKhlc0D7OPvVK1s4fhTY
fOjjcintFgRYqdJCNAsMC7qT3+kHCFwv1/Am0gqqGavmbdNc9XlX+VirsiAs7+wwxOSVcvCSJtjo
dk5N23R2J89wMIHdGHH8p+/rt9pqhSs4Do/Xc78l3nVfozfasQ3jWGqP8YRYrf70wO8ZEQQOpP9j
qnMvkJdra3XFjx0B66QptxG/06uZxDIApEFYWTxZ8HmsPCp7pufmWl5kjbXsGrJ5Uef46CPoyMQX
Dzmwt74KgaHNfQwaNFwgkM8+Rt4SIMDYvyza3Re1CCbtOMHWeFIBh7FM6ogeC2p/lubqtiQbbtU6
lkI4w8PQ37i/fm6J3poDZHhw1MRHWp2RQlA/f3RLYo3tDrUURNwD4b5x6+xjp206aCEGButR7P4e
8AtPHxFtAJaKQgXlrlr72ZdYxjMgVAbY9oPf4d5Dhb3wXHURfTLVHjtO74rn+4arRWhvkr+Rdb+f
qx48Zi7EJb05+PLmaQskEZnkXvjjNYubpJ22nAjNPSUeIZTxo0jjXTAEZJc6u+jQSOwiFUOr6j86
0pR1Zh7wR8s97XoB5DhbERIAq7x2sbkJ0Z24XhvqCtSCJMVwHBuij3qvrsH3BaTk0/n96LO8Nn0D
0wSB9zwqj40TyCOAtwMLUX+3cr17YRbJBgbY7BNkZwpBO/6r1Hwn0/hgT7vNXfY4lpTiUkqlOJuQ
/AeYDE0q4tuOyhWgFjr/imtmUNbev9mAXDgoUEOsOmjzncGKbttE0/jg2M4qTi7XpUSYuCQTUHMi
544S0SqKgcRtwdf/pRkFSwYC8Ugf0Za5Qqh5rkKibo45zLfmaL58s8cfUxpUtItrmpsdBcwTHNHW
MLCgSLXnb0jtBlEmGTS/KFP+rgQ2TSpUfz6GEqHev4TZoo3az/g55Sji6aH8LTAbBuLl4UfQLCGc
3PkuJd4326w8zJIG8dSLo8gZ5+x1EVfv+NIucdZ0DQXNVY9zFD8TVE6Z+xVBnVfMdXHLDmHn2bq2
o18H8Irl5jN1P3MNR/yA+HtHsJuVIaLFGxCsukSlrRbuuHbFsGaSm5tNBS/MQgSpuD5ck7iatNjq
VdJUNdlVDSTC87WHLXUmV9Q2K/WdG2BwbERZTZa7x92CLyjYh3spRST2jOLYFfjM9KhCWasJgU8l
t8OgBOhSzArhDUiJE/btX3Vo7kN/kk5NaQPKOcwGGpk3K8bJXyCEEbDapq9BMbmfO43DwWI+//Rq
m1KHhjNNvWaMpOXtsZdcNtUeKjjGBPqq9A7o1+UBpnrchLPikIi5eDAtiaR/3u1CmEmY8pGypUqo
pikmJUYsC38VIVfQWnzEFuYyKxoFTjjZoG+TFjaQSERiZ3pqLZXWR22gXS04eDnN5/Ebkal6/LGN
kkmvzo2jbX9w4VpfmcJDdOm6nBkzZMb3qDIcFrXXts8i8K7hJBykWIYarweXx6UgqadNwapZhB1I
wx4sL2McUjnnvcvbu9FjEt9WI2Q2W0FTbYKS1/izY3MleibMuJ1cbR3GhxnmflY4bH6K35wojtPK
JzjjaD2N1+/2vQHRI5C6CCvXLUOot7zNqSraYe+fRxNfjSCIuTU4+b5efiphqxLz7Sr73J6LXGZ+
EyuOpY93bCyVCgH0YvY6DrAu/kZwxJZ7Ru/efoHRGrdcbhUdhx5FwtF2j+jXrIKl21fTdWGHRdod
7cxmj3CpK5YUMbLt+SbNQYBCBs5Zk0pz4sS5knK2aelOrIzIuZBHOqNseO50GM7HWrIT6ZbwiXR7
aWoiD0AlXEKsnPKWxV93bSZJerHVQkGRWQ5KCq8dTKVzOr4Vwvip+UfgVPBKUVuHcHtxYbHp1+a4
SyQGmlrJM1zDLr7TMZDTsrt1ZhqIviWX7MSXi4eBfZRA247sfkCyyZKRjLgS9YYB6vpnLjajQWUI
1neicUfODxGZJPNLq3WoAbjr3kZgyQB6/kWsi5ppiIEAgcJh3DLqrLbRwbAd5jd2ZK5uCsig6TAE
tctPAUCzo3725u6klfhbk16dFYBwBFkBmJJuq8JzInjO/YEFEbBXzAVr4GHkisaba/I9YCpTrsNc
LoXnYN/3328PeHUn9gdgSXS0u1BT9gLy9PRBzdn/+TTpQtYaVis2z2aVQtUiq/XnftwYyyQ0CVFg
53fP3jjhZxQO+oleL6dMpq0wIfAta1XhF7ou1WG0sFlUnlmgUw4Yb4yZOrnDEJCxU6uUPqgzgtDl
JAL1QnP6dP1Ql8WPUfSUndNy4kuwwhV4xhrz/AKfSdR7YeN+WhKRhWiRaneYN29Lw6dQMlJWFlre
1hEJQLjHhmiAqPL07DAeW4QUAM/gLdHv+7PDWMNuBRLQTjO7f8tdz3rbkhchB2ptihprderi8P3I
A+kf9lO1uavcGR/bYtqzESkRZpjGCocy7jK4PPyd3rHlxZ81hICg9DJ79uuLZwDtI49JYu09h4Tj
0+4uMVpaMsKUsSbkTMcUD3rh1y9k00mIGUkDa3dzmNVOGcYKO2oDBuG4kASGiDE67Od8MrdcxBLH
Kc85zqbwrkTN/RtXsPgn4c6YA7FPIACMSIrkIsNYgJ1cPb/rki86BZi4X0GuD0Ce8fy7RdmPwDBI
ax/9qjxNQLastmWjFORWhMirsYIdR2U3Oa1n8IwNPiaxjG3jYX13AWN5LWfGtu/jsAqfZOeh8Wo4
Zn0NaJ2A4PlPHke2QG+7sg5NIjm/by9FSBYrGHDCzeNQ0DqjcC5eqhUFFfL4lZGq5J7cr4kqZGGE
gBgydFwvbUpJrUH0are66PyPt7JTXNYUOS3EoI1KrAShQ9mN6dVuC3lmUoNXO5dROq/Hmrjlweae
Q66UlxoLBhrOaMlHP47lnIvx2odItW5ZPrdIFCw9rVXIqJae6XAIo/SQyTLcxbJAXALxhkMbMs+p
SlWMhqNRVcOXxxydbK2Dsoj+jrzHRlf9zkfdvLClL9orzfQrUm+QNg+9BmEeQw0pn3Rd/S+KirgV
xb09QHKSwIsUdHvs2WrQIAjlL05Wpt1+hfVRrdU7IiBrxX6PsWDbEZa7zvasoGMhBZNLSuD+sQQq
BWuWAITplSdYk3MP1GlrUd8GWK+MeZDwN953jfioYPc6GbVxLR631yb5SLVEOMyzA1C1lLIX0xzV
H7+Kk1XpPdBaIpPfoo5UnAIhyBXjd1HMIEWRL1jfNCxUNhDHscSe+YfLOoSKssxrIAtu+vDzUV3j
497rEQPjtEjFB0RFe/MNYEZulm25QpQo0y7kgFOMZNmkOxNAxH0c4kyYkJM/uylef+mXzVhgb1Jn
b0PJFDXynRqjr2GixLqrgvAXf42g0buFHC8x1FZNe+tNfyCz3gHPVYlO8jDCaFkTw++03+ybu444
zctzUDaD/xsZFdocbS6DD+npeWE9M5Y0zuXt0g8aJaYFNIU+vbTVbG5c56cUEs4KH9WmQwgRavss
PyvNzyh/oRAuzoa99qp0xUmiHc9tiy3V3trCXWTCODr69D+nbgzz+aP7tVVDa4m/PnRyANkRZCI6
x9e1TvRe0zB31IOdV9KLTiWpUb29OfOw/60Lzfz+3ehivc/s++HXunqbU1tNd3itpvInrstaeNiJ
lUITc4vvMXASuQ/jGG0/WzLOPBwo1nYK1Ha1WFTDcD11uHY+UyoYDIXZVzyYUOziRZ1k74qkiXqq
6EewRyb5/xaWKinuVxD62cBt/Y/iPBA3wTwUdmFltUD4nJhB5kzw6eQGwQr34FozBwZJkRFnq5tE
7uq7l0XTtYMaRDAtRuax9UdRIGc7yfe1Gwgn22b7RNJTM6CQEtNnG0HyYzv1mqhh+mFqWErRlNNz
X3z4vtR5B7WMFytHmBjqw/CErHRZO8NHgJzhtzCA2HQq1JmaSz4BUKoq5doVJrYBG0N2U0nINt/T
Ejm4JmV+D1onjKl98NQgipa30APNkR2ech5d/b2rMffmkI8pdxhQ7MY3yC7oVM3Bgo1g71PpWZmi
P3PuG1Twn+DCg6aBhjlbIzmtArRQdePTCxSZK7+FigveLrqc7isAaZxVn2Oauprv8axHPG01K7YV
Xe6Vi14aAU9ydmBqccc2//Dab2kyElYNWpaH4lmMb0miug1MFl0UFdABQBEfvicWzNfh6SqJh4RC
/uFL2kySJAyWrDtxXioaqs7g2ytfcEaVbJY4T1VqA+KHRSfBQ2iJdMSwKtzE8KMSPcpmjYLg1JRd
oDYp/sqq1LznwHTQUj4p0gUrwkimBfnK+YLBBE/SzkXs//alsLuv9adcQNYZ7vKv/6SutZmqbV/m
cXOhIarFFOXPVzq+jIqJCdLjnv5HQ6zioN9hwHjx2XyyQcyBv34VPy2SFib+qqUhfZ7J0lHvVLn7
yPLuZWvFa7T4HfUnCbzpYyQN9/4Nr+0pF9haOuC3/qrsNrAjfh8p3d670nZn0XCPNZdWzMXbL0e3
bHQbkZ2stkcH4fSLxHI3muyVPaCEWhLnggwogE1cdi2XI/yGZhfi9SUaBVo1forp5yaAGLN1kg/X
XVMKybblFS45Bmurt7mU7Sa9obmRWrdYFFeMjQCxuunOaQXh6BokkvhpssaIQ1ZnAmKlG/Or2AqQ
+z36b0buZWobC/DS3FeIXMTmRe45HSOdKAKRungz1ko1h818Of6K9GLOQPJppwouLvkLvedBQ4me
KgJkUMNAE2ZQIUIpsYvKgZ4rPm5k2Pp4Qj3DB+hfLonE1v/RJrC7Jhcfol7nkFi0a2dDfE+ZKHg+
gS5miLLRivPGNCGl2OLf+CKi+/Rqebasma9dm0k69Qz7jAUrtFCdafHr3LAdERYxpYuxdsJN1IXn
ooCYq9IwjOfs1bRLSNw0/nSViO1N8HcockU2323Jtu5QpPAxuyvnyKS7PcUdxK+8TF9v5h5vHc1K
bLCC3mlMmnU+BGIZveDegY4lkB/0c5+rvRQ/8RC74OGNipxS37KZ/IyZuT2a7iezP/rQdKkXLaBZ
4xil1ZB6UDi+mz4FSPAN7ThgyUw59yzlfgcR3OFv2Do7VS4i9uM3RXsQOiY61f54wFT9MR6g1IHZ
BZhLeJ1YksxXyYLMlFMlxIslPsw37cVzPybVQvTFoG3tXmJjd8BYTCBCnEsJ0tIYa39Y1VFkeY46
3Qg4H/fjOXIUu6IuSON5aC2CnbaY4oucKo+3paVyWNEeaxCACsNZX4fTO412vFjjKMV3i8sX9ykD
YyOPmbfGdzKkKtW8QBsZZj4sAC21QKz/+rfrR6D+acaDeeykb9HcMc/drKNbbIrMdtTlGZYhlvPs
fN40ftoDL2T3IchKN3hAxQ6k5703CDOYErhvq5M0PpHsVxfVBPOPJhlTgr0+tD1XzksF8xQY/GI2
4zlFmsmS6cTRLs3lzzLlHUF555fm6ukZ/omk0TyFnfjjjdMWUCUTcw+dG9Bi/mWQTabjYekMUNNU
+cDikM74p+1AKXCBLqXVtmNSjGPYo+8ZYjL/qbA4paxlbGHcNKiQ49anzHK+0vfZEQtPlknc1Tv8
otVC3j7cfcRkwsSjD1OflAqn/1kPaBns35wae+O7xZGL
`protect end_protected
