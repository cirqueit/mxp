��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���y?HUc֪�Eq��&ܾ�]�r�����#VM©�"&�!C^�����6����z��9PS�OD�6M��Yi~Ħ�1�
 
���R�|:;� �࣠X�9�tTiY3�w�.2�)�*��T��6��h�'�Tj�Y���/N�͕�v�o7�p��EU_��8}@O���b��!�~�i��݉c�7�0mB��
Q�A_����DOuݦ���(�W~��C�}䔆(�Y���_3��\)��
����f�.�BЄ��K4�f'zrB���߶P�:�Ѳp���d���2uJ)�Z�ч��S����:{P��N?+0n�=ڶ��d[,��6�O}�?I��Xk��;e.\�diHD�~�2l0��Vz!�b�M&t|9��{lYE�e:������Ie}"f��������<�P��S-�p��
��2$q�94O�́��#�ҋ�ЬY�T�RM79J�OهI!e���Щ�Y	�L�,٧�J�Oq+��w̬�&_�J�S��y�E�6�a���x���0U��Z�����Qdb�Z�:0^B������m�'F`�Js�8�2`�;i�4�݃��e&Ho��Q���?�B܃~^�B�#?������q��`��W3:'ϖ�n�a�y%���ٜ�G�8�+��L$��m�ԩc�_��b̖����}�)I�T�s��Y�\\]�U~[C��YZ��4�i��E�OQ�+U�b�8�a�O$FEx�w[�_�s���t3*�yQ�}�"C�$^4��xpW��J���k��`ψy�� "���R�E���8�ë���A���w>NEY�y]�c@f�󚹄!Ii�͎$^��)�dfL�L���, �S�>d`�l�u^Ut6��@��\�6 f��*W�����I$WD9=qs�^�Ȁs��m��gEP��1��A�?���I�Zn��3j&`�5��K�($�g��;>Yԥ~���w�y������8P�&��&�'F(C噞j�����-���/f�E��"c�\.�:���4�F�D"�W��|p�H�T�s-f|�	e{�<.cd����_������CT̵���c����fѸH�M���?6L���j�GD�'&ĺB��V����u���=������������x����K9��v�V��}��ʱs]$?\!sߙxM��p��Z<��z!�w~�wc
��B��*\W����p硆j�"�"X4���9��� Lt��O)�}_���2
�=w�� -6[�7�<�Y��.D�n�
�B�^<2p}���&����ES~����%�&W�[$l�'�o�1-��4��0|���Xc�Z魔����M�l�����#a".�`#t]v�9��o�8�U�ݰ21��\(�=.Q�N0�P�|��'����QU>LĞS�^�>�ϖ�_���q�\���$�s�v�p��*h��5t<$e]J;q�����ըϒ�O�&�T���GA_]����j��,f�H�X��*9�����1���Q;yGy���o��4:�}Ñߜcji���o����[�F��#�ݝ9!�񉬠��DYj��
�S��6��q���r{L�G����!��1l��-��(��!��*��=>X��>1�㋶�^�mn.�z;e�4N5BS]��[�T�����}��[cl&�og+���g��z�>��]���w`M��3׵�%K��z����%�9~|>-���4�(Z����>,�c^P8
�o���m�E�����Okr�?X�n8b+��Ϩ�
�l�5%�V�Zk�5ޠ�W&����Ĭ A`������vJ�QӮ�!햸\���-W/ֽ��Pɨ���r3���5!ۣ}�G	u0[Bif���v}�gSg���������hd���M��+�δ�m�-� ����t��3��^C# }¾X�������{�?_�A�tz`�g���6];btW	�x�����}�$���bӌ�|B����y�w\��^L���DҎ���n��WO���1S�Rr|�G.�1T�8>��2���3c�M�L?]>���鵢;-(�}�����3�Zr�v5�
l�rL����,�0pV��9�i��]�1�+b�f;�{�S�٩��2�~x�������/ i�#n�m�V�/�I�M"��)��?�G�g��# F*.���fb� �~�#�@1B�rD_t��j�h�<���5rYd<y���<��9��\�`�żh��jN!��q���V$�iQ��$���ݕ��	���]�ǐ�u��s}?����nNY�*أB�b��]�|�|^�U����^y�vѬ��-�wIJ>�7.Me�_  ��[	�#��1�vZLj�^Ԡxc��b��`�s��_��F&r��nȲS}lȖs`2"���~�% ]�;�*��4'��>t�t�>���A&_����Y�2N�������B��& k �8���H�d+�|��9��I�~L�U9�ǠC�0RU�'���{$����G�J"�#R�F��#�#���b�]�#�l:#�iOGH��D���{;cXӭ��tI�W(S+����|�� �.m`L��|W"���n�"
��]�8��[vN���eZ�u�5�.�*Y%�f	��S�䣮�bߗ#���h��Q�t�5��ր��������;M����k?Eru��9�]s�p�x�ĝ�>����d��P����.3�� #�(�C%�\}]tN.<���r���Lp��|�c�!����@�Eݶ
�p=ie��ޡ�����Q�K}�;Ve6cS�ZV)��؎�l8iz6	�}���R�t�/1{��ѼE�e��b��������g�Ǚ�9)�2�ԇ"i�8�A��˝��RX�m�
�!��c;�(+�E��79�&�2�n��"�����47�fL^o��:u�'l��P�bc����� ���s�4�ź��7��a�z�	$��J��a/A���Sk7p|i�lث���f7����1�
��+1r�h��Ҍ�<�[�� ��P��%O��vT̻�0�I�E
���b�d��Lrc�H�����>��O׿��W�sh�8�7�"�Aa� �璂p�g0X@S�Z����~� d	�T�r�}x��b%m�k�����l%�`
�/Ma���C����!Sf�!(����eO�+E{��@R���exxh7���#����+�! �@U��Z��9��5�W��v�z�& ��̐Y	Bl�.g5���������U�7�Љ��%f�^���}v@8��3Jؙfh����P�т3:���B��ȅ��t���юH���@
g���@�w����ɇ#m>.�x_?a�DñY�ǿʹ�g�>���������?>�.�����:C�)��m��e.sn�齗��}}��p��A��'�ە��&�}�2�r����Zt�K"O�N5x�g� ���Q�@�v@O;��N��qC(r��s���m�+�>�G���X�n��c���ua���K�m%�ŝN��1�~G�n`�����Hs�;[�X�@�:}[G&,ƙ�i<� [1q����.E6���\m�)�S
a �.�����K�t�	PL� yNgP �GS�.N(�e��3I�h�?=V]�	"�Z�i�m���@y_.�{���1�oꙞ4tI���;�Ʈ�p5h([��H[�G}��7��E����'�uG<��Օ˪1V�X���\@rB%����Zy�<���Ea<�����俱��SK7e��~[��i�&RB�֟�����������wL:|>� `�tS���e��Fnญ>/r���Js�!�<�lO��ZYi�rxv���B��(�M�1{h:��i�����L�f��PkɶqKxo��>���!��?4����% �!�>�@����^�D���+kjݔ������.7��n��T����8���p*�T��=l���iI��>e���UZ�\{��iZ$<zԵ�@�$0�B����V3V����ِ��s��7�ť��!��EV�VRn�i̝����̊]�9� ��C�,��7���ك
j����e:��dm��':�XdK�4�Y��B%�1���|=9�!_��&ҵ���tx���j�;ّqX�L}�=�jB�ak[;�8r�̤�U�2�W���u��y�%���2�����f�6��;.���+�Ӄ����b۪8�`�E//m�FY����(]~�w%	Jz�����_���Zm��l:A1+?Չ+)ic���Mn�<q�<��6o"P3��Seܜ�x�V����j���eI��;��s�֎���$y'`�]�B������]YMzc7_Y0�A5N/~5����i	��(ʴ�A�j<�G%�`W�Q��#����7�&G���������
aϊ?�7�2@$��,�<	�>c�i�r�7�����|�����2�u{B��Oy5
:J�F՞8I�).a���3-S����z*�>72���$u�tm"F�U���ϯ�;�,v0�d�-��'"�p���⥱���қ2W5�m;��5����؇��[]l���ĐH/i�lq2gl�D��ɷ���v ql�g�0�{�з���:�TytF�ё'���B�Z��6��Y����t����Z����X.қ��U���I��Y�N�b���W�@ɶI��J�V�0;T�`K}�f)b�������@W�����)�G���Wk'J�Q� K�|�_��~��0�R	��� B!�(�]��B-i�:�_X�Ni�9"�3�*�q��:�iE�!m���y2</�}�E���j�� G�Z��O���/c#Ÿ��]�9� %J 0=��Ql�J>���±[�]�tU��$���/�a��B�����1K�p#���DqĪ���8�^��3*)���D�e��uR��sv'���e�_nf�YC���2����1�T��u�WY6�n9��3�
�_Z.F��C�N�4��P��ﮈy�G|�D���/�g�Zϸ�� I��Ba2MY�:�Գ9b�������S��\��ұ�w������ܚ��q`�D���5��/X���MfΝw�Ak�Q-��,~Kg����#��c�]vǌ_"�Gɉi�ʁ��D��p�'�ue��}�hE��w��Lwa�M��\�`�-�*���&��w��c؇3~��"o��i
�wފD���v^�9L�������V��x��:f)�,϶^p˴Q{����,�q�I�����u��~k�O��DrY���h�O4C���0k;���f�[!Ki}i�Y*��H�@(�J�UFpwB�rU/���G�;��wΚ|Th<��l{<�Fcq��Y�|��=������=�/I�5�Ӗ�ݣZ�3�����2��μ'������l����b��L�{�F�4c���Q�g2�7��d�% =b����t�0I' 	/`U�J�Xt��>��z�z�y$a �5S2�]�4���,�����8,�%�-��>����/��z+�T�?;bY����ʃ�&`y��L,��bv"=[�X��sB����21�#F�������)�8G�ʭp�.������C;�l�7N;M�P�y�/��q�+U��j|�u��F�˰�!��y�e©q[���o������OBl$u���Y����o|�����Obԑ����.DJ���$OY��*�";�CQ�a�x%�'����;��m���j���#��7�)ҶR.��~�en��cS=5��k;��L�|�K�e�Z�����)��ꕂ��Դ�]9x������NB�E~�z_����L��G�E��E�u������TlT�{/�o	ьJ��~FR��J##��J�N�..3�A��g���#�0D���6{��@PT�>�:N�p�B��M�NS$����cO��ª�;�{��X2�t����r�{À�&>?ƋS�j�����)�Vb�cx����6� 6��=Q��"H�	�ү5�����6�5�d���+���5��5eA�őb�'�|�D˵3l�O�;t^�*_�%�ۂ���#�8�V&X�r�o-v�����zBL�Ѕ(^өpū*r���=>��1_�4�2Z�&D�H���ń$��)�b�𹤏��>��u��m\�OE�����%���̄\�E��^��3K%5Ӫ��n������V�[H/c��Mq	�j�خ�]k�4�E�"�}��n�dn�l���δ?n�kh�8!@b�ԩ�)�so�,��<!8a؃T�O\�g<���S�@��W��6|�X���Ԡ���2:vJR�#���YP|c�V�<���s9��T�PԞ'SQ�(
�oj`� lh�-�Ղ/p�m}sHlYxm��cvI���ф*!#Ŵu	�܃�ZZ���r��PD|�������K5�$���l���=�H��l�Kά�kNφSǈ��\��w-�E��:շcVBz���p�}��S��{Z$���&=�g��l��{*/�w�Ƒ�p�K7����J���A�F����KT�x`��>-�rz����b,����G��}9o	X��$������`�\�3����� FY
������fvm����X*-� �j�, ��%��Ȳ2�#���4���FZp�(�����8:�lY�Ht��QX�4D��\�.�84T¤-��3v����h�f�-�Yc�/���ۊ�D��; �r+4Ηf�i t�;�V.B�5&����Q#��[W�#�2�?��Z"��g^��:�4���;����3P��?��=^;�f�W�F���<y^)B�!�[�`1�&A|�j���� ����Tu��A*� ��?�O��ߔ�>3'������)�$��`�vs�SzU�����2��;!��3��� k��G���(E�En�%(�@�5�ønW���f�wI.C/�#t�Y�7J2%�sa�[Jx�}��_�"�n�vE��^�w�j�<�S��r�͓8�f|�g�_>�g�焃��y&��l���p"�п6��>ls�5 �DD��@[�����H��Í�M����_�{�Z?�P��r ��Nd J�j>�=�|�҅To��
fʃ����GZV"3.�n��I6R�@Eֺ<J1����X�
���Rj�߉Z!⿉�'3����T�\`g#��8u��~n�OYP5��T� ��9N\��ᖣ�����O`U����j4���/��e8BН55�ف�0��Jjd�e���^)��ߘ���	V˨7�3�4������x˭	�u��@�D��6kH�D\* ��A|LS�Wg�yR?`2h����-wN�����$K\�TOOrr����s�/'HA�5o�1w���FT����z@J�4��i[o,}"��O&с�������������vO���z�BN�YΗ\�+*na�(��r�92k]���$|klre=���"�8�&[���:�BQҘWH@-,�B@�+�^#��lSi{�\�/1��݃��"�:P.�*�f�����Ĥ�c�U?��oP�p��ti��qq-�b�Cȸ���f��׀Bgq�(��c4����� P��԰;�Q!��xXӓ��s}���h�ŘO��N@��9��A�*�q���i���/��~�6C�������<o���8���ߢ�i<>�z��ĺ;�<~�E�%
�U��E6���ե�=�t����3��v�h�+��.����N�����>�����5^8��f�2wѕ�JC�Y��/�/5+�i�K),�y}�Mc��A�.���b�ҚZ�KUn��g�
��n��f3�&|1�C��]r�)�C�	uYmd	�,�����5�/��*�c+;�R����-�P6=�och-���Ɖ�
V3���
���AS%�5���H��Vt�c&��o�w���+��E��E����F��o�V@{�^/~:�w]���yB�D+�s�m�
m�o@G��*��jo��E�`Dlr��vhA����i�J����Ғ�� ���������\�B�8�����J#j��hK�Cĉ�����N���<�4e.��
$z�퉸W�e(�)8�C5��L�W�����C*�,p�=.�b#`O��7�+I�����;u��*��� 9`�k�@��?FY���v�v���x�+���Գ��Su	�'��H�>X����Cn��E��~	ki�Ov�ˡ�j�4��|Dk��9r4�Avq���.���d���}5����%�����lf����O~Yj[�o��g���"z?���*E������ݒ����5��z ����<|�@J�˕�Yvб�K"�n�����I�b��J7D|�{��L`$���M]�������z�F���Is�5�N7���UX�����d�=�֩�(s�hG�k5��.�R��_��x�a<ؒ+���k��8����9�ʧXg�.ӼO���irZ`|A��1�������������С�怣�S.	i��u�Ĉn�N=J��f������I;)l�C0�����M�4Ǔ ��{��-�!� m���< p��W�!��2+�I�����!u��`���zVmq���v��b�!���608^A��>�|��`#巃���a���]��J��:�	$ՋD�x�4+�W��{�N5S�O�����;�H�aQw�܎]���I���YT�=�^"ĻS�z����3w�K7�b��]!C���|b)������m`��_�`���D6�RTE���%u0�U^��@ׁ�C_���5��ΘhS��3�z��fd����`z�T0�S����խ�JM؀�;h�~@�83����49/\H�j�f��n���h�Kp,����:,��0�A,��.���=G��55����
�U���?���J��)��6��c�Q���TƷw��%�FP����}Gh��l�?Y�\�̨�w�Bނ��q�� }2����ކ�;�o�,k3��y/�+��P�	͵�V0� 2���{���@�rD�/L��'����U�֣2d�Ӥ��Br� p����m{�2�����>kJ�69W�D���(q�z�0C�#������<M��S��(r�17]MC����.�Ć7��{-1l}D-3E�\����<�[q�[�k1�jR7�2��KOf~�A�ף��Ć��+�-�-��̂�������#vt�Ff���ɭl��������?�M'O*��?�e�{�U<m5�V �/�����s��(?��):s���ۈ�f�A0�����}P'渢�w��;sرy����A�@�`����~�g����<���&��=�@h�J�/y2�3��3���Զ��i�h�C�Xm������l���r��w�ő6a��E�ف� ��4�!$����v3��bXbEX�y���T6�b��P ������S�D���Z�1�p6�] q�[�-�=���_x�ʺԨ�'IX8wv��!El`�P��ċ��5e�;F�����Ft���R�y�ev�OI*�뽏����w}���#�d�q?�H\�¥I�Ӆ�����Rv�����Ĉ�K<��Bidz8fR��0]1����n�ʲ�Pj�d�r��r�#* ���Q�ꦭ,�m��q�J@��*&~i1���e5֖A�>�W���J�eO�N�n�M��;�^��|�`R~<Sz���s�o�=��G/b=1R�o����4ƨ���
h���a��/ʃ�� ��0;����P�[&�b�|ݝ�V��������e0��Q>U�s=�_�j#���΂Z=��˰���G�2���/c6��w2Q�qL�C�6,���5m�.�*g�	�;Q��&����e�.^�Ʒ�O�;��Ή��B.��H�[HȄ�!�59�ɾ-�FuHn���FF?�W���|G�έv2�w���3��,���S�Z ?;똳	_2�Λ� ��5��{6'}Lc^B� Z�=ѽ{����z��͗l�3��
�>u5�9��h}v"\:&'7+�z�����7�	�U�e�+�^f��4=���7��Bf��������|O����*�Buz��|tA����04t׺Ʌ�����Y⭷p�����S��d��Σ}���G�l\I&�S�M/�v��.�F�u�Wq�֫�sn��$����n��t�/����r@	�1���;�&�H���x�9�u����c�W�l����l��E�?�U�L!g}����!�ϙ]K�~D�3O@�vF�.��q Y�J��Ʒ)Yb ����	"_6%�˓QZ��8��`�:��k0X�LH�����O�/`L���NQ�7��\C����t�fpl�
���U���R-$Ւ�YI0�� �����gWѠ��v&W:���[&\[֗@tP�k�%+��@4Q8[8�\X?�nƃ��H����=W
�(RCJ�ĩ�z�G6K/��M�T?C?����^lQ9�!zƧd��*B����
��(���?<�KMӪ��Ć3�qvlǹm��+�t���������|���i��y��>�O�$
'CV|#�_���i��9k(��U5R�JC���ؗ�|قS�q�O����!�W�|�Z��S��V}���#����X��p��3K�_�O���=#usn�%���[|��R�9��%_q8x�dt_\A�i<H�!ܷ�K5�bd	�Bm@9���=���Ԥ-���)ߞ�ߧM��{���%��;�H$gٍU��#1�����h��3p��y׹����' @|*��b=��)��Q���Oϣ��ñ�^(,u���
o���pjx��'����ET�K�������\Բ%�c�?b]i��v'p���õ�Q-fb�Ǹ�V�3�p[��L�x����p�*�
J �S�Gg�l��� |LOy�C�*5kq�>��`��|�dt���ӅnzV��=�[��W���x;�9ޠ�$���Y�&�o���R� ��o)�� 鍣�:P��xT�~��n�:Rj�Ѣ��{0�\<�т.�:���Z���L�L���B�ҡ�FÉ���p�Şٿ�����@�-v��-���$��:c��DM�_ł|)\HQ�$��%I*�V��'�t04����Q+�$R��X.y+��ȣ����>�x������c#��;�lz��t(�[�Od�
�3�m�֯
|���L�G��wv$����񄯱'��m�=l�ꂘ�E�,|ͱN4X �U
�O��돟�,^2�:G��&�<LBr>�P�u����m���Kq�>E�V���'��{�2�xE"`"AzU�œ���⣎�F���PW?T�՗���It����`��e���[fMWM��Z
�����y[�=�b��^�5��nD��� �0�y����z�m�����ǘ�O��i�?�p���q�ee���_�J���h|����bo���x�pb�R��q �Џת�Ͱ�B�5&wM��!���){3}�Ëu6���s!�L��+m`ƍ��V�Tg�u¼�8���׵�(��$�21��8���tx]"={q��cZ�i����JW
nݲ8b=���_U5�ø�N�z*p�������T���1"#�(��>��ܸ��b��5����}�;S���z=:���?�w�� 7���x�dO׹�Y�]��4qd?>G?�+�m���̮$� ]� R�Փ�>@nä�@vF ��6*��JÂg�`БucM�02g-f�DƝ����D��>���>3�\pO��H�&�Z � =��˂\r�'']ٵ�;{�53�}\.�����r/\�]\���#�,��]�8���߅�f+9o=�ٿ�'JS�/�+��yښ2�B��s픱�-���`���dsJTB��@7%�@#�Y�����o���,�(�@(�L���~��#!�{̑`���bV{��H�0�$ޓ����7�:�n��Z�"���oO��[%���v���xrn��C���,���P2�5NȏFR�uZw�* O:?F�"9V?5`e�mY<`�r�֠��t�y���s���ئ�W�'�?��V���:Fe�I�+��_���a��*�;���O{�4"yK3�y~h�ѿя�rى�Pw�̺��ͽL�O]W������@E��֘�O��� '4�����Fl/�ƙ��<�&iu	���y��,�$���bO�����,�t���@H����=����u�QGqb[y�e~�r.�Ŧ���i"�":����EN�|9�?��{��R�t?�-�J}Z��!\9�o�kR��eOK���m)�]	f��5���#f������hw�ߵ��.������
S��-��C����4�	d�� U�q�lsG�ӷi�H��&����{��R)�9�}yO-��)��]0�l���O3�,�� nX6�Z�uV5%�@��}�S��gTԣ�?>��]�����<"w��&i�#�Y'P�[��Ȟ�<TA�V�����3wOH��a�˽{�o#��j(���_ð`ɒ�C��^-l���#k��z��ȰZ{L
/��dQ^��ö^m�N�Pa�K"�C�KHL�C��s�S2=L�O(�U=&o�VeM��;��@A���%ƒ�?prLiy�>�1�"��f��֣'geSߣ)J�"�����5�#�7}�$/7�̙�G��\�VV������<�O����UUj��/~��+2f�Gk�+��Y;����	�9B�|,�CI^�2.O?���/�ۭ%�^�}�Q_Q߉#�T��/@%�l�	.p͏�#R�ҩ�"�s�l>�����i�=�c*�_��ly]Zv��s�dkZl�Ө�Āص�BJ92Sk��ԃ;D���-rk����c�܎՞�I��i�l5���G�2�Ȍ���u)d���ex���ν�U�Yn��U��0Ɨ���F�Pm��%�Y"(wP�I[�����ը�8������q�u������f��=��!ݝ�G�}��qB�zD�������m6̠�T���d���j����Y �AE~��/��k�[㋸Aeyy=��$^���ը��/��n�IʓE�_����`��	BY*:����Y�[��Avb�9�)?ok[���q�K�BeH��:��z�����.8��֜h�R�
YRyb&y��F�<2�O�C�� Ae�^����IP�]T�1��(R����$�Ӻ���3};�E�TS��kur��OP���HL2j�dd]��U,M�$܇�=�4��*��b���;���:���
-3i8�qp��!@ݢPs��Im�(&М����Pu@�t*,D�)�9��\3$��-2@��ZHz�~%�]���	�q�ӳ����7�L ����;����¨�G(�+�RՉ��O�ă�wq�R��?y��������k^�o�Cߓ�~Br#�������������ifr�}�T	X�8CxO��z.����Q�i������^"m�%�>+�D�
�����x��|8v�0��Gb #D�;?>���Cy�Q�����X.�!��Fx����y<Լ==�%���h��hm;�$(�����G�~)l{�4؇�J��z꒘���L�S��l���>ZCu2٪��¼i����)��p��䍱$ng�@֥����,₃(��Z ���2s�I�G�p䴡8�K� ���RG�� �A��`��A�t�5T䮻k��@�xL]1�x��U�Z2>6``˔/��e�>?IPƨa�U;c�{�.�[[����B�~;�οc�"k͹���������5\�9��;ȍ�FDJ��%���ҵ���Kv)�L�j`�J�ab�y�BW>��+�uT���,�����Z@�;s�3�=��ws���ζ���!kU�3�V�z����S�{����p��)�O�h�	 �
P+��q����X�|�U�倇 �U6�X��5�_��X�-�*�=�B�
���y�/�zV�l��*��*�)!D5d��f��r�3r���~rnB����]��>V?��<7voC�2�� Px�JC�����}>�o��wD^�v*�nZr���;�UxX�q��K��劜�e��ǁֳ��n�	џ�� ��$�)~�*�-C�=�"�2V@���{�� �ɴ͘I��l�~��΋N�I�7gֆ��%�LZ�� ��+�%�&L�aC���Z5`�K�$i�f� 7[r��A�u�q4��>���2��@�h݇��(K�q�`�?��U�����ۄ�,��1�1���� Bg㡌mY���0Dq�_�|��s��B�ʳG�	1�jR��P�OTM� 3e �W@���N�ǆ.�]�1	f�*��ɪd�)�qɍ�, �v�AR��[!R�M�a���28N(������5#f�/TP1��j�o,0]�fP��?8���0���È+��<{��"L3�\�
k�*���-(̿���y_A	on��)�~A�$�{f
���.��J���c���>Q��^��S���"�`���|�yߢQ;�Y����YH�U;E��o;������ �%;GD?R��@[$�_�N��q����J��ۣ8��_/�����B8K�q��ΙF�
 #��'�R�v�G7��Xb�Tt׆�g��U��������������bJ/��I\��i$gh�G⦆&�I����w�5�-X���N��E�i���+��:h���(���-+h�
����%&�~���������J�q�Z�1ӛ��V�o�	,���6b��Iw���N�-t0?�F�.���`�ͽ�/���nܡ�`�������$����c�x�]oA4�Q13�T����|8��$��%��*�Y�����9�&���b�Gd1:���i�%��k�I!��0xF��4���S�6p�r���2�J�4�������H�	ߪ�~
}����"Jw��Ri�Z���``��3 /C���\�^ô�P��;q ���O������q��ـ���p�C[���Z7� �Qx��3��Vt��I�5���J��z]��y��T�M�t du�4���3ށR1)0%�}���c�s�<Ft'0��Z�&Y�Գ���c���U��HX��j|s�"]�cq͗+"ד�w�v���p�.�Wdwc�ŕ��6�+3�q[ߤ.�9,�,ÿ����"6f�˿���D%pM�}2���QG�T��4�Ô05m�m���÷j���P3��6�}��#8��=�(a�4z�I/2N�V�����P�/T�ۖa����?+:H(Z�S�.h��fK�3+d T]���Gf��-,7��E�U���Ae���IB���C�pH�s-N�T��H�l�ə�5�k���O��<_��Z�g�j����ޚ�F��N�-P�fy9*�t}�*u���o�
���\�� #������&*�>×SLN�e�A�>%���5OK�ɕcr��:�c��!��g�i��'���ؙY�5q7i�>�L�HU���pK����{�wo���(�\,}�V�ճ�2�Z'��j"���ǰE�.C�A?��a���a����mK��/�	�
t��#}y(y�:��?���=f�t��&	1h2a����5�J1)�׏md�D'�g,�Y�)���5˚k��%����saK�u��b���J|1	l��s
338/�AsU|���Bݚ<�'���<û�R[���2���r��U�X`tAO�p�UD�C.·��oܑ�q�����1��Gޟ�;�%�����XS���%-gu�_^�/B3URG�m��Ԃ�����i����2hTܠ����E�u�.5����&��_:�G85����E�Bӵeo��1�p�%XҐ�{��+)>�T ��f���.`�m9�g������¿�B�������$���Rh�ݯiIt!;��	z���&�	6]�T�E5�F���Od����yeb�%#2�2��{)UVodK:Fµ�6Zi���,��b�������k�)�&�-G�6,u�t�6aȐc�F=v����c��T{�@��G��n�>��$_c�ȡ�&���iku*&t`��s^���f�l\��m44����Y�Zrf� ��hS(�[�\�h�XK�qKuu:���BB�I���ǭ��ԟ�)��h��*8'1�Uk�����m��A�s�}������r�蹔l�@Du檒պ���"����`��@�^^~�z�ܤ͓���A9$�17c6�Z'V����)��e���@VH�R����k�KꁶN�]_��@ǐ���]D��	~���5
`�3��*��FLUJ8���r�5�����n�\_	������@q'6WU�ci-����Z��p[2�,"�h����]��ՍAM�JѴ�Zzד^���p;��@ �꟣|7���!�Y�)c6�Y���f��? ��>�@����t���F4�(*�����+�PQ�˼�~l2�l� i��J �����n����̓*��t�� ��"�� <Jv*�C�m5�����d;f������/>X��P�ݸ�r�A1l��=G�i����7f�*�j�e�c��Bl�f8C�x�R�`B�������bԾ{W�Ϭ#�L8p�G��m���i$�eIU��#X��i�G �Q����">"�^w���e3�q_	 ���b�L������iRshc�*w��p�}P��N"���f����Qe%y���^B���ez�̥0���gpq���aӔݙ�hy�Oh�t�g�����˳`$����ź�c)2@��*(�(����b�L8f�@l���;�$�1Q���kp�.w��C��Q�����:Tn߭u=۰-��`]��dUf9lЖ52^�3���n���i��S�qw;�VM�^�H�C��D��@�4�r�����䬷$��r���XM�zM���o��p�ʴ�6��V^H���?�Y�����8��(!�S1�3��<��a!d�o��6[�� N�ݡ��f��7�5�n"ÝU!�y�.�Γ��5��5�B�3Z�~�.�[?+���<Wr�I��-Pw{���	HA{L���8;� � _6�t�+��Ἀ�"_���&�K]G�n �A];]\Er�čw�؂(���5��ϽYdy}�=rI�3$'��;v�,��f�W~N�s�OOB�t�]���cY��Ѽ�S���Jڋh�dm�L���a�:��H�|^���A{3��Ε�G�] LU��U�U��d�qP:����ot�J�X��Q�C�W,(d�;�����%�`�.
�򠫖w!ѐ���w���5�E�o.s��f(�o��1m	Z�wv�+�w.����^I���|�v�|C������t*�V{��!���r��f�o֢�:���d��/�`8{�Ht@����]s�h�;%�̮���1��9�1ُFs"C�f�����R��U�B�,�<1��i��
4^����.s[$#��
���8'n ����o�aeI�U��A[�b�L ��]q#�x w��n ��u��҃��#-�C$~��U�(̹A��.7��K�Rs�op�^��[���Nj�9#lw͝��]��$ �����-N�P�=�|й�l�͐�.�G�
4]�](�Tʈ�)5���B��nBK��<��@�ja�(��,��c#�M��̠�.[ʤ��@��sn��D�B�U]&P{:2ޜI,�4L"�w.uB�����1A:�'�dS'ǐ�fK��h�I1Ǧ[J�ٛ	�Xb�)Y������c�G����ݔw|���xs).��r�ڂ��;����(�̱�i�0M�l~?(d{��\ɠ�4���H!�0�ӄ�B� �^�=/�;g]�w�,2=��C�K�u^F,$53���!�YF�3klr��#K��$Z��d�1qt�47#8���:c;��H:��>{2k��������X�#.�Z���´��U<�X�a�+�0+�:�����p�R���'4�V��4]���x����G]���>����0tj�y�Ő�k2O䏏���n�%����?2f���20y�?kj%C1���F�YU���2�
uK��Łs���M��+78*AC��-���'��]I2�0;�l#ʨ�^CzU��@��2K��؂�/� �-�|W(n�|!���B)S��O��j�0bU@��\�g�)�T�X~�5�L��R����Q���/|W�u�](7�T���?q8Z��|�r�1�>�b)�Ǘ��!�/[��P��}2�G|�KE㰑��ޔx�%��O���$��9�)���V3U{F�Ov�?'n��׆C�h#���:(\�Dt�\����篢Jٰ\��F�-$�1�t*+���Xf�	/q,$*��Tx�>ʟ��@{o�/~�[�����V�&%�1(Kb0���C����	0˳	����Lx����/���{}ØY���h���R�L��"	@��y ½Z����v=�m���m�^�K�؈�_�i�����e�c(\�\�@�=����B	�S���ϴr���C���j�g�oK�7&]�����D����aI�����ZzJsk�p���H�p'�9�L���<,�\ZU|� ��8&(t�,�z�ԫ����(����a�����r���vd�F$����/�1�3�����hB�"klb~�������-ٛ�waYl�r��.��`e^Y��#��vOŻ�n��XS��.��'���%�=�-�7[��ְt�]�0n6l~�w��::�U@_d�s�E�6�pʅHg�OMxc�@�:�=�W.�4�x&)#s#%��UQ�!���ˇ|���t��15�q�6^�TX�=Z������<��g�R�5n�t4�,�Vs��^�����AZ�K-"��g�K]�~b�ӌ�H~�"$m��}@�G")����<�lp)���4t;8��g�Ez
y�F<fՅ�w�\.˷�7G�����lZ�V�am%:�ߧuH�k����hc��N,ɇ[���7�(�}��>;����"�Bb��P_l�cɛ���Id��[�;������b���Mf�va���߹I���Wn,��$�?N4l�7�/f�>�|�F�. ���f���4�ci��/���0^�Bƌ(@�||i�Wv⍫�[��+��z�j�q�eL	d�q�Ź�TW�=��Z׶c�T|� q��n[�"�g^	X|�j�`��{+�}2��Ȧ�_"0�����Ca��{*H
-ɼ����_�_9�3�ݫ�h嘒�j۹ַd(���������VLVp�=��N˜�m�b��mf����ۤ3�
�nXZ����������I�u�_ӕ�Y;Q�F����A�Ѝ�F��i�پ/�2��#��hI��q,x���(T� ő�d���	����(�&uҭ	§�����\6��CC���>�4:!�O��@+\��~���!4����^k�D�q3I�^�٧J��Ɲ����F=+nc��r��#!2c�?lI�Z*O��Q��(9�̲�ê^���b�i�s(B�>W���5o'~Sw�d��dkP��ॻ��Fr.�4��!�ɞ��q~:A�6��^��pH��5.�������!��'	*�X��V� /s����D��he~����I��"�]w��0�]�ãO������4�,^ ��.:�#��`������W.+�yMk����8݁Zl�˒�a�>������y�Õ��Qe��3��	g��צ"��N{���K� ��\���P�+a�H=�U��4�+����	�h���(>.vA#�>8�Z��DS$m�q��A�I�w�mb���܅T�+�Т�<bS�7�u6W�(©�\H���l�UjJ�c��vD������-��"�}��d���CT��Xk������|�$�����*۠7G�*(X�8ơū��Q����:'$3��'��u�"���ú�7�g++�&�mʊ����z8*�������S2��_�}a_#%(5	��O�Ƃ��FFC!��k����sZ+�1�g������-���&�V��y������)	\x�ͬ�:\�u(PzJ]bB,T�&⃺�VFޥ�8�{���:G�?:��P��ϻ�JM��3�g���1�x���C�z�m�La(3լ�����C��\��=�//X����Xv��[懯�C�zɑM���\����*^��㊠�eD�?_��F��H�������z�T~4SK��O!�-{ۿ7�����1���SO�~���n�Z'����X���n{V�Z��Q�[�����ģ�d�g�P��S����%p$�H�G#�Ne���%&M;y�|�{��WJ��<�v��]s���GJ^w�^nU�6�<���ɓ�8�s���	Z�Un��[{���QO!2��h[e�VR����i�:�r$Yv���B_ <��ю�����U��=�y��L���Dϑҽ�.+�^ȼޞ�J����{��	�\����j ��V~<��rㅑn��A*��?ko����V@��/��j��������A鯈<�
�W�p�)�:8��p7�6uul�3s���������+.�ª���iU��x�{��	�C0�H���#���9�2��_3Lf�Ӏ�J�l���k^�{�YH(��`J(t��TW"4˶D��U�����tjM��x����@�Sex8L9I]g����w6�	��R��!O���cE�=��f�����C�}��[�.Jau��0�����D9k��\("-��u[�ϯ�Щ\���5�ѽ��� ��X��8�|ǡFF4.K0u�/��N�P�� X��3�}�A�G麯�]{ ���tD�΢��Au�M(��R�A�P�W�y-����S��/�m��f^gGbn�7�����:Ҳ��}� W1%"��EG4��Ύ����G��Q�1{PU�0�r�ܜ"���o1�5�_�h�ɔM�d%��Κ�;�Հ��w�VUatd��&8��ѮXK[�r���1����OR��=��AqԴ\@L0�.�L�J-�BT����ɌV�1�E�x�Ž��ぶ+����Gp�$���~�v	M�5O��(1
��+(�,�0��u	SsLѻ���Yeg9�o��٥�y��ל�_�@w��<p$�e�F.p�?�f�G�g_��c~�hj�O������k�:��:�6�O:H*��M�n�f��+Е�Z��) ;�4N��o��W��t5>�N�M��U��Q��U�J��� s� �nR�f~�eIxY�t��=�+J�ʲ0�������O���M<x�iEɈ���^���ۓ�T�
�'�[p,�n��ۜvx&ꪧx:���g�������2j��S4��[
�+^b0&��.�q�GB题�jb�����Rej��#(���Q��V�x��G$�� �H+�-�I^̵g4aF�z1%B��Y�7MDo4|��R�i~�Xz��lb[��J� t�U�'x(a?�]	[�n�Lɔ[c�:L�]�lʊ��Yz�Έ��:@��&�����;>�P�+�o�74g}�g~H�X��h����@��o���ѭ<�	7FL�%�3���IRP�;��&�����{�S#r����I��g_~�3�G.eRƞoL�C`�ٱ%0G�E4Tz����fm�D#�/��	���Ģ�w�Zd�,ȥ�-�z	f���Y���ЍU4�Z��ޅ����3.Iiz��)���E-*s�����S2��X$� �4la�f�Wj{���s_�ڑ�8���P3緞Qy�E �bw���6j��<�`x̢�&�}�X�vG}�@�3�ͣ��+��
t,�:�Fw���"*އ�'������;�DM]�9�Yh�=���\9-�3]j��Ӄk?ݤ3bDRH ��O�釤����P=
j����WS2bІ���{DL
kz?����P��G�(���	-W�Sv�����Ĵڗ8g�lT�me�f��J.0� �+`u_�?z�α��q5J,��
�P�ڏp3ɯ�$��Ɗ�N>�e��a�,>���3z:=~���P�c9^�9�|�����3�y�QJ��e}%H���'P� J�e�7�r�(OF��sִ9&�ޫ1�{"�CZ}yG;���M�����5A�KN,ݐ]�Kl2�ʥ,��lxg��rhg�^��M���D�2i<���eS���Z:s�.:�}9�FrGf�<��w�-6�Ut��#)���%v�����ވ\1Ԝ���_�����y�{:{E����M�­�VE@�>"��n͕Ľ�6���f�mv�ܺ�+Z{n_��Z�0v�� �S(�yU��GER����.'߲����(�	���^�Ԁ��� �C�M��R���BD*]�����R��*O����]y����4)�vt�
�ѷ)1�0��Q7����Oj�3s_[�δ0��\@\D��V��{�n�?�A��%�����ٱ�XF����)%_+�q$���$��U]2:a/�=R��ʃ.�8)�aS����k�Qޙ�r6q�4�C4�+xr� �D�Q�%��V�+��vo�Zꅦf���D��>�QZ��O|��"�/�`0@�/�v5(SӺ�|ݱ,aF�9����H�7�IGO����6��.�-!]���y��񊘶T�´c�F�4� �-��-�٭�uM�8�ĳ���8�I+&������c<l�{���4���!6��3��\n�=H�Pt�%P=p�W��2#|G��[��%�w1b��M ��X�����{��� ��2�/¿�R�z���C}��������>E4_���]ϭ�$�^9_oZ����aBPk&dv5����ϩ:�)}9�hW�G�@��V5�sQ@T��09�R��u�?�=+�k8�Wn#��B���c��������A^X�,�-��Z⃆tg��X��?#U &�G*�=��)��C%��)�5�����(���;IN܇�Cei�ZT�[���ֽc(������r>0)�K-�0����VIըD��U[<�I.�Z�s:���� ���D^<^;u�$Tif�:�[��ıY��${XJ|T�ZN��)���f���2�����8u�U���l��{����o���,� ��1���d���f�ߵ�������5ӭ��e%�<�l�i;j�9J��Ӎx�� ��%� �'�j�`�+7{��I�	T�޼���#N�&ކ�J�^% Kw�+�ΦQ���|���?�_��j�T�|��S_DHq~А*úl{��C�����
d�;a�ƶ�o# �I�8��*$I���P�p��B3�j�<���s�@�P�jn�l�3(o�gu���d�蚾G���C�Th�t�w�75�ջ��u�_���|I�(��������bǦ
P�B�]�ߦ��S�y�8�*�j��P��7�(�)i����q�ǜ�9�x 5DUj���M��>� X�~��+o�2��[�)�7~e�u����֨�V�3wB�խ!�8�T�}rN�)|��Rt��=���+�|t7t��$��Q�ņ��O�(��S'�Vvt�V�CrBޭ���Y����)���L��3�kބ\B��ke~G+�aXw
ۡ�o�Px�)4@ ��� R�糈4��`�V=;ۖ�sp.�m"�tl���vϹ���g
�4D�͊�N[���͢���=٩B���2��}�[U(�!�P]z��m�ϸ?����=f@A�bC��S0���l,�V����/� ��~�p��=�[�A�'�*�S=$�g^ɞ�p �g����m!�C	S���!���q?ð(��%�5�H+g/ێt�0�r;6
��9ʏ��H6�vnu��S2k�4�"�t�J�©�[J�d����J�&-�0��=K�J99�v�b�6��lf���LԂ?��p!Cl<I���;��|�<�%�In��PGEFr�=��	�Q�	AW�k�NH����9f�����H�Hw���P�?�!��=���P��֎	�s����U^.}��5�zU�"T����d`<������nsۜq%���b��~�y��ͧA�ȅN�Ƴ�قX���,VC��a��I}��#n���<hj�����Q��Nm���K��Y̥�^Zc�h!���&�H���n�o�\�)-ӃiI�xƿC(���G���m�\��?�-��u_{8���Us�����	"V���)Uq�csn���8^��4]�:o�h��e�?$�g���:��<^��-�r�i����~�r;��Ze�']�7T�� �bnPɁ��5�����U��V�g�eZ��8(�|�;��H�${��%��1 �^�n�]���{Og�L��k٤�;��a��n�u�c#f�'dc��Qœh�:�S�Z�A�;Y��2S�n�n�]M�)���Wx����z.������4OU�M� Ϩ�$* ##:��iډJ�M��ڑ�7��àngH{��J�s����������k���H�YC��I�]p�]Gz&e�5[>�AX�<�{z���gf�4iE ����ThxUE)J�iW�W�Y�<�����1���;����th�Q����YU�hǓh.�����8[e�������Eb�������Cf(Ȑ~�7ې\!����8�������Ij��Ov#$1�k�c�P�dq{�hD�W��!`n����v�4�|<�T�ͬ2ƶ�KP{w��x3�d0L�q2?}��|ml�tO��@���)�G�+� [��>ƿVC�hyp��,���6�X4$vN����S�%��_,lM�V�0��e��x.j�\�5ؖQ����˒v�{��}�p�ǈ��'f��$������)ŷ��`w�ԣg�t��PN�פ�5Z��8������칚��7�lͩL1�#m��*���e՛x���A�����Y���zo��K�đ�|
}0..�ER)��3(�[>2f!S�e n��c<��3�BoR9���^���h��<�w��jh���^�ħ ��d���8�x�teV
û����i,ӻ�e���F��̅�G�|�?6�4�'븙7�+WʿE�^�h��ޤ���OtG�S����Q�:*�j^L��(�w�i�"@�p���ZW���dgb����d�ƧmhrZ�[n|n���E����5�ƙR���=�<u�L���ArB��&*� +���g-�Z���4$�D��O��.�_u,!�:#�,)�,��m�6[�1�txv�Q�p�j�C��@BN��Ð0E�Yj��=��
d���}Xod���RQ����L����nߍ�����C���]Ǹ.eK�=���j� �~V��-�;���![595}"�΀1�Ї���G��ѯ�-t$||�q�<�)����x���F8"&��깉�W(�J���O��eW3[0H�����27C��ʛ��{�0�qL1�*�e�!�W��b�	��sT	�Q%b#�J��ݰFKj����r��{�kV|��<[���U0V��������,�SL��܀i���!��(:ʴ���|#�p]m�f:yu�\�8:�3X�)��PG��F,G��*ߍ/B㘵�\H��P�8��}@�Չ�.���n��"���t�!MF�_��������A=8�F������%�O�=0/�P��^&��/��6�Q6j��~�ڀ"f�~}�$��M�
:��a����K�ہ��QI����,M쮫���mx��f�IXl Re��P��+�"�]&u�U]���)6G��-,,S�M>�����p
��&�jd&�S�p:ǬT9�@\Ct^Y��&1F�����he�|q[Y����U��J�Lܡ(:��@���5ႄ�#2dB������%�+y�&�u5²���Yo��<�#�q��:-��t�!�����8����7��Hc*�T�)}B�W�h�mgsG!'^��V�J7P�����8~�F<��٪y��$b;�~#`�*8�+���e�C��iDrH��l��Ů�*�'�쐰 ����OL濚<@W�����8\w�^� � �5��̑��C�z��A����^���3���g�SKz�yJ�ޙ��^�����к��I�)�iW�6�h�評���.�\f�Δ d���_���+�.UC��;�g��cg�J�=�zZ#���_�u/Yu�S��h��X8"h-#"Pق�-!����E[�`�[�#D07�l}D:�� -��(�_����ʍHP�h���N=),J�L�3�ݦ�r�[g���_Դ�v�f��Ћ�rm%i��ݛy����Q=���x�����3��~@������_�Bl�S�&�D�gŻ85$�°2�~e4P�/�E�T���ʢ���#�MX��x;Gu@u�$"BI`���ǒW���j��@�f�� �S��#x^��i�4�f砱�b�^��@��z��}m5#�-��YRƤ��s{�^�aH�a
C�`*�#/�	��:�r�|�E�n�.���d���Zip.��x����Z�
r�I�l<҅A��O�"�� �Mc���³�z)Ma����F�V~[�t��^�+`Tz�?��hN(�_�O~�#���R�S<?�����r���'�A�G�(0�����*���?�X��WE&{�߰���#���q��i�����D�g�	6;"����X�o	�=�Q��}�. ����I�\<�+@�]�C�e�9��{����K�� �6g��ꉲ�~<+Kic-�y� Nn�S��� ��`�@�ԍ��zS�˻h�wg����aF6I�ww>��
��+�Tq7�=N;�¡!c$'XO����o�d�j��o�\>z�l���=�
(��#� ^�J�X2ɘ�r���^?__%��.�u�Ī���Kg����{V}$nP劫��`�2@�c�d�3��t�?�(�
�����<�{>YS1�]��\����'W0Ǿ�$)4�u�?�&by� ��<�ɫ�V��1��$lV�RB����c ����@p�EG�U,��t����:]��ޗ+W7Y�=f7(.�&ѶE��{���hvS6k����u��TP���E��r��)����X ��%�