XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��cf�QD�Y�go�)$�g6;�i*��c���Ԝ���)��Ap���+�֎h�U��c��'��h�7�uy�W��JKZЊ��%�^h��+O��lw(�03��bױ�>��Q��13���TTޯ�T�i��[�K�*����no�dZ���F�������Bu���`bp·d�{�a��p�����m^W�Ez��`��J�j�`�Ӹ : ��ƾʞ4АB%o ��B�P�r�fl�G¿7̥�`ވ��Hq�,!�(�7�L�����4�D
goSm1Wz(��W��ڿ���q��!����'/��L�M{��՟�8Z�m�
#<
���_d�bI�u�@7M?T��{ՠ���#0�����¹S?�9��m�Eƭ��Jum��]Ef�Ǟ�4�S��o���oi{Y"]u���6��냦'[�<�.�v_g)��R���|;Y{�!E�倒�V��8�$pX��Lg����=�g+W���`���x���q1M:6 �'�HSGD4�������\�.��03s7'��
Wq\����rS�Ԫ�`*�Z��Σ�Q��o:&u��:TKIG+����w�81��2�zT� 
uL�.�;g������ Vf��9ջ�"�5�oA6Ι�m�U2(g�W��Ьl�F��B�"�y�5b%gp9*�Q���]���W��_� �K�0�J�V[�0����Q�}n����z����ː�}2�y��p��)�G�Y/b S��VQ*�����c����x��"XlxVHYEB     400     180i�|Dl!Ӽ�v'�y�p�&��e:��|R�F��<��$�%-�)�k����,9.�cak��BaD��5�.o$~%I�Ҝ�� Ч�k���*�Zk?e3�	wb�ǉ�d�]�F�@V���	|��O������P�;Z\(^�I!���K�l���(�sn��+�fY��l����� |F	�T�"���@�ְL�Sd�?-�И1�Ϧ̬7�2�N5���n�g�
���6�~ti��j��~�~��*�A3�w�ڞ��u'�L��Q;B�d�	��8471�h�.| ��2'Z������Zq�X ��p�;O]�@J�����j=c�&�l�����Jw�I�GUU�o᱘SL�	 KZij9��uz�RcN���J��XlxVHYEB     400     160��ז���(���\���]m:	�o��n�k�W<�^�avᾝ!��C�[�������={1#)�O"ƀ� ���('mxV%*0]}���5�����R&
���T��fAa�7�)_��۲<c= t����R*��u�U�M%�F�RƳ>��Q_p�7XV�ě�"�5��$}i�=��iL�ҿ���0���ӭsv|�����o��ZoS��;����xr3z��"�̳L&��7��ԉ���<��)+;��*=��`tv�%����B�ұݖ����##����T�qC׍�yx��SL����n�=�\$s�iЌ�gBt�7���G���â�$p��XlxVHYEB     400      a01���A`{k�-�j�x���N>\�����P*�r\+�ɒ��#%bM�
K#�ƚ��?�[VEԚ�X޶�dUpd�ڢpv�~�`[��;T�br�� ���굥 h�|�ռ�T� 3q�?�:��.����<,�c�XY9����wY��g����
g��۾��0XlxVHYEB     400     120�IS��)N��}:`��|O��?_�uqD�mM�2�dq�˚F�i�%���+g@vu��pS�e
WB�[p����D`��s�*Z!^{���j���z�����1�����O>\Iˈ� 6��R>�#�%�$r���y'$�����2)5+}�{7:�]P��1�C[���
���7Uer�
Ɏ�����Q�h�m���z�du��L�kBO	Ro���\��[�ЯX����vy>��yt�ѓq��9����v	���Z
��ȝ��9����I�o��4
�9!�e���XlxVHYEB     400     110�!]GM�r�9)y�,�[�����n�>�<Բ�4��C\U*��~�{����������0�V�W�Z��A�Oq{g��ԫ�%�!x��U�*{\�d+��gV͙��}Q�Ke���Q� u�zڦաy���s,jT���0����e���;�-������I�� �]�B������荤}���;2���?�є������8��6�7�JN�h0���� 	�SO��)lMM�*�q}j�'!*�O��b��VM
�G=j�qh�j�@lXlxVHYEB     400     130�F��~W���ʚ��Ͱ���a�oM1[�h�Žc��}�����晪�nNT���
b
����ds�l��i�N��%�"vɉu��?U�����hx1aׁ\�Met�����E��JK�P��3 \k')��pg~{2'`#���R2�u���5'g�v��t��K�gB�Q�G~��s.R�Ҥײ,�����.�5��$5��U$\�\�٢5�@���N�2^���cz�oc5�8�)���y���kY#�ѵzXBjfg���K�.Ixӿ�z��H9�WJ��k�=JЏy��6�[�XlxVHYEB     400     130����]he� i�X�����^����:cU9�q0F��^>��Q5�s�Ī�����XQ^� ��ͪ
5��6�<���<_����-�y�no�\|�䌍 �Itr�q2��w�4'%��$nRjgy��!�̋��"���Gd�a�r*��=hq�A�5��cm���95<I�p*�!�-Q���I|�s|fN �Q�c�6_I�#-܁���P����hd�b̌\ud�Jcn��,so�1;�ܺ?�qw����J}i� r�]EѺ�d�	��#�J�7�x'N�9��6�Gj��BCKXlxVHYEB     400     120�,��� [і��J݈	�Ӏ�`F9ڹ@����PS�_��·��3dMI#?�I��O-���%$�G�!����(�f��L�+��F#�ꍪ�7-�E�m�㑗�IJ�+?0c��N�*�$Sy��J�0]�HѴ��7��Ŧ7�j�:fW�Y�����4�/N�Բ�/.N�B�����$`8M���9�{/�H�)'�����=B �Ө����6=M.�JL3�IT�L2-\�ܰr�rQ�c��[�e1��<-������kѶ�Q�k�~g�++���H+&)XlxVHYEB     3a6     180�܀��K�z��Ap뗴�E�����T����M	��Iz�����n�{�c�Z�xA.m�'V�1�R��#7uҒ70dD?&W���-��iR�a�Ț@��ڡ�7�l=���i��w*���]�/�'&|!��$X���5�Y+�zk���Ό��3���|���r��j9
C\�]��o���b�C��!�4�\1�:�-=X�&�*D7�3���d�!H+����ȿk�����w�Ufq�/n���I,�3��
����%�>�"��I3Y�������h�^���N�J�_�2��Z%��	cjo{��ےgq�a�-���nhſ/���!]���G�Tu����QPSk�2ýګk'�\#��N��