XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(tA�3'�YZ��dT��+Hv�f�B�OE��済��.s�l��6#hTzՂT[�v9�q*��Z����:?��Q�	�w<����\� �\EE���� ]R��J(\#Y�4*ީM�G^DT�^��Q`U���&����BO l�w�zy5{�U��\�6�Ђ��йb���ܳ)�S/x�R����k�iq������Z�"%����++�C
�[�U�t�T�c��������8bɠً�8ڽ���;dC���(HՏ��
K7��+�]))PK_�#��HNn�ڝJV%q^��k��U�Q8V�QZԿم���<������:�H�$)ޮ^�&"�6u�2��Ԇ(h0ñ��ΐ<��*A����l.���E=�M�me{{9�(��F�!g��,m�����D�F-�ve
�ƒ�Ỏ�����m*��;�S�J떢Y=�՜�����ހ���M,p�D����P��m;"䇄�:�~�U$=�|aE���4 ����o1�4��̄=r0���:��O*�Q�8#%�>
?ol'}�z6}���ج��ȿAg�I���c�OH� �ڐ�U���AJ�>�򒓫әd݇��*P��L{`@��	��)܀�͸O�������^쓈�?�@��!��/�>�{/�C�;�j�w$_`�����G4�֩���c�(�B3�G#	���Vl�����Q=��r$3{D#Nt�}��{�Lz��V�VB�D<�y��,BJ�_��$�}��I�&XlxVHYEB     400     1e0���%Y
��K�Ƚ�mP�`�y���'������neQuF/���q��<�h���N���]��t�G�10���)�29���������H�|x��|�����d��jӬ�`����ťC�<�f�`-Y)s
t�������%1�d=�8�nm ���֡am?�c$���W�(1E�M�kH3xZ��>}`��	~30���Yh��^|�'TJ��z�� 9�F,�o!�!8����Ǡ��hΒM}q
��U�_�_�#�9�a�˺�ly/�H���2�GRQ����ŇX�kD��q
@a<[�1��P��e�ݞ��������	
7_vWJ�hʹ��*����<HIR��AA��&žͰЧ��o�n�"8��l-�U
ST�N1��sF��.��Nĥ�>���t8@�h5�C�Hdj��S��́BfU
��s
�
J%��#��������ks����?�a��E��'���c'Jp��~-�wsw�XlxVHYEB     213      b0�.��z籌R�q!|F�0A�y(����[��;X��� 3f,��i��[�O`^�MZ�lgR�^�őJ���͘�99��0i�@�eϚH9�7?��j��@. ��"y��!�8.3��R=wW�OH<����l|��zN(u?f�$�2p�-����O����Yʾ�зT���
!)