`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74304)
`protect data_block
JTfejIL7HCccFok9m18LrhtM0jZsDjgZHnLsCQJJTY10FXGHEbnlnpCAd7GqPfwIPPjRiTtuYmx3
cxovO3e9JoqxhnnMSXI1TdkDQJLdPhKfrzEgWDpBD4EOcLqUGMUztDe6+hb/GrZTW/kfqdS5zz+5
LhCPVi9e7XztzhUzmxiuOIsptzGJ0BJkL7ASSk6LFeCf4eg2pZy7qman3jQ/3FTjsLQ5QdEqcP0R
XVdYtopXaAO+iT17oUOa/8AYQxUW7hNuw5b2B5g9RmT3XGTp6ZL5bGa/DCXPgPhL5/QkBRY5GNq3
8lPRB9EcuZ3hxREZ5GbeyyIjZHBrgF2gR9pYBbgrJqRzB+CcGZdE84lwRlWlDADvWaNtl7+fjVa8
3y6bR0Sg3ygJi6ISYmxPgjWb6Ci/TyxGZvj7CpyDCnwFgOnaSNOUPqk/Q+R8B6Zdh/Iyb3DQzMFy
sofDFD0DLMVJajODVsY2c+jLnDm9XW8jEVB2G+Cj/sax2M+3+A63nIYt1GV/kU0O0DLfWBvYHbE7
7kPzGZ8umpnoF7pv+oGox1CSttU2Syc3rM+rBRb6VjguNd90BZKNLuSH1PlzG1QvW9PBqyDad57I
VUd38wkhSV5f09sIvQH0IWM4yksldIjdsFepxWMciZvjUu3TCj0ynyB/E/AFxTaBQ9sFp5L+RdUx
bbnhfg7FQm5SEs0lcTA8RLGbh3dSECJvVawGp+/+XoKeBCbantcubuKFUhjG6Tvx5sMy/3g2z4lz
+M7qMum49lMmekUsy8sgMdM/SSZ4mVOcEcWmZarUMNAnOm6o2USKiOneFwmgnlmnJV4T73gD+Bje
y0pUAvnYlvwK+K11mMZ9pMGr0dneiU5+ThBrpDwvb8HC0R4CTYnzAgsf+2lMlnoHPONqNqVJ8WaV
eOSq2NZd+8mi6udN3slbcpEeIdZc7HMv8s9gGif0vjYd6GmLcXUrM7lo9NodUiUMICtNII0pasP7
vqOFuAyoeFcHXt5oI2bVMHEujy3+jWAvQUzAUbAj6bz22BTMQlaq+ftnJETT8VbsPbdrRiQIaOVd
2NRi/lzAfUfcsuNNjuQJnOhTS/6xzCh+by5w1EqYup3fbVWpOOuFRc2zccwC0m/iAOS5gh5XEud4
TjnlfcdN7BCxvZ6xBANQRTEEv4Svmjv2pUg6nZy0WKWey44E+obnhX/ncLmTG0Cr4wqRwKkhmtsQ
CyLKVi1cznZEBYfCUqwB9/jmjB2L2vrJcQ2lIUyKC3Msr11tBPvFXOPd2ytUoHorMtLXSppGlIz1
LemmnGKpJVUBi2qFBTK+Q0lY7eTgqshPEvxUMndfPNeXMY+hWCEoHS7mADUcjw79GWhG2Yy/+2U0
QrBpR/7tRqZpD/AV8y6E/HkLlrAFGmwdoJSxyTz5O9ab2RYRy0lYr2DXJMvg03bdI0ILxg4lNPMv
MHUx18TWrWkWT4bcjVR9QR0oOniHOFjHJvYVtKadYiP5VtzsybEY+SpmeBNvesX7MnfAepWw6zJm
p1Hdme0WkCtlSgkgP7GrcuN3aU/WNwmUfTA/zBMur9VdcrPi5XgZAmZrNQWLg8l6e0PvI8kaCAD8
g5wRfsxKzwxff8jA7zqgKGtfnW+qafGDDzJ02R66boQkbtLvRFs9iZnfnUXzl42SdIb2M7EoDtks
Sdsr/FiYKxrUwlfxQzXaxXSpfPf03zg3Na7i+qOaQemZ4FlvtJIWMU2vsp/wStwCskCUoyMGbO94
N3mKqaakfm/iNgW1VNYMjb+8BMPYweJ3u4v9puYbz/tQxtHZcpujdwDfe19Sa4Z13cOQ5e5gDRvf
/ZGpTH9TGc9arme+hlocPC21gHYVtNeEUnsIB8QaBRPos6plHW6wVS0YqgUdF1vCsDTwP6nCtb65
Ug2elrNIdaHH7OcjNYoCrCuSKF83Vbjkm4dqhmOVYgK0YtqVP0ZLSy/gFsLnecfVK61uGBs/voFZ
/h1eBHUQ8QQ12MLCJDOMc5EAUT9VMIQbKVu4iGZDdv5crWkgZ27fU+vR3ej1g6zblNoqXe9ZB7p9
qi7Iq2ppmT0IMFDfsQDfC3WysQgOJ36u7gcXtzgJdITXDqmb4jrc6DL46sDIDHkjq6PvjdYej8qp
+hOiyQOvIJxPByYAjIl1wyD6S9N1ULNYAngspndyzwN0DzPx7sH0Yfl+0MStyozjbmc23uwgwmc3
Hj5Hk215A2V+hq9RcaNQVO4agAvARJXgl7cUTbCqVfD/IRhhLHqLYNFyDYLtZZXBMqXmd1Tyb22h
TDn3N1KOEU9BTVKaNHaZbZOdytbcy4hg/cvYkz8+G6RksJkMacJ6JKmGU0hIoxKEpMkYc9Q5nuLD
7FUhaTHbXJfzAEkt9B52CU/r/ORVa5MNpx6FVSvVOrgt8GKN/4PFxN8jU/tDrreGZbN10qqqxLd2
pCkcTInJQDPMbJlfKXHEdxx7pJeQ1J/7lQgDZVJk7PbSBn0pj5JoIq/N1yI5gtslaG5MAcxVqh05
i6Xl8slHew54JQ6/1OcfWaJhup4Ck8sVuHPMgtKrSP6cqhJEn1QSaE30FWtPKWl9JY5MkJu5SuXt
PuwRYk7Xrqzk+hs7kGfDMKE9s+0nByMkdA2cYaV+poXYZS3sfr0zic53whSDhRti4SlAUx1CmEBH
5/nOLe+Pg+Pt/H1F6WRYT520e9FasAcbDu8MfSu1T/w2bLBdULFGkB02eCto5GO1ZCQqMWSt0HUz
FZxtR7et8C55E2vEBYaAiP3N3aEcULCcCjgr/Fjlp9pORjhf3FeABXvJMpu4Z9eTYsMmaxM9PDJy
y67qapniR8f05XC5N1CvyD3nXODMJN9w1KWKhObL3aZ9X3vx/aEoQpZEjbeQHsZxJrnMZpeuFHvF
56CEmK+3bSjd2m0kncC3KpWxAMHlkoGdAgNm69MZrQDqkgg/AbY8SKUs992R7pJR8FywYfYRLbK9
xsBKayOVTYU71rjD6YyOVpPJJIHrj0o15QcJfKU1IQAkvI+13l+5RtNbIF7FK0ukNypHLuJD+ijg
YFMizKZA5FANgNxtMDQ87ekIkAZL4bDw7GHKoAJyMja88a/FRmm2GiYs4Xtd1Lp44VtiDsByklFA
li/nkl2HApxt2ecychONFifV5sPSl0YeXIVaTIo5vggiEOk3UMnq27woTfyQzeXCiLqwYSms9pEA
7+7hua1GStkyzvufuCY6RXQimmS5ygLpKSnOA9Yx1DEWIVlJUf1ABET/AvSCqxKQA+M+9hMrXFZ1
Dk5e716P5hKWk/P5t7LDiCyY52iSGMUmEHZLc5bMfafjqqmUiTQwIGCqRqQGwPQ/0QgpqOsqmLQq
izRbIVAYqxi60y7xlPM8rwjBKq7afPfnokqG+ENJrArdiYTJtQ4Y1OfPzC0pcy3TOToMLRQq8h+/
+TMaDiZjXs/fGCQYGt5wbgMtwYHKZyVHDiA0rnGQOxuEIfcgKIoUNLOZRZ0ePpPTyW5IcKqlTX0K
wxsoxwrTQ7Qpo4z31jm0XOIIHUNVAxc/51X66rJe4FUIKYs0A/s/ttiteMkRXG5WqhgkQBXXadSi
SmgzmvlI/PKD3jEAAJM2rpketwz0Payaq8np7eQwuQjHEMGgyMAoqSQh+w8KhO0OqWIvWWDHYZcJ
BGuCGM/P+EPp9bfsrsTuvLklASMG2AXC6voU8mb/RxVuT6E/yX5DmuR4VvLk0lV9mqoLNgcbXB3T
sr0TkVmKpWbtLCSqQ5iCoa2Sth52onuAuRl37Ws8oei5iRJ8M0SLZC7j0KKa1os0qood9WXmIy2f
4JauXpTaipcUjR6D4NeCLriBG7zzoQ4UIRm2kPmhyOY/o+g3UJGizToXT0XvX6BjgAo01rLEFBix
EvIouJBCB9dIW/1DB2T2ppB1KyrRGpawhkrWREIBnkY9YoDjKZ0fhySCv/oVneQa5bS+McNtxSYR
E31WY2tFOhQY0Ytul8nRwpagj7Y0pl2tMitKhuVzNeS3hqkaBluIwDMq+vLoDSayM/uQzW/Ftbhl
I1H9NqZV/pGP/4UInORS9JL5NGTD0CQDKXxtTwgMSrmLNH6ZUdaaWXqmgZTRbE3dinbyfq1cV7co
g0RGQKUWhBlsOPj8+7kqsITtdot/GbCMf174Ewws7kk3UOrivaY/j8cejcnwT3DJ/EoGYMlfv8rt
1kFLcf0P8Zlcu617DirTn+qDZb7nZa3LeS8QvV8UZcw6aH0J8j7DV5w8Sg0OMG37p27TzH3v4roX
5sM1VU5E1pGpCu6kK/dsN/U4jByMPcJQ9UN632EndAWVyLvd+R2BLnu9v/47Dx8BPW0RWx0Ii/zr
T0E1a679MvtyPQuT6MrHnbM3xc/pSTMTfhlAS+fDzH8tvp47RnNoF0IvcRo/7iDXTC4NahKuXNat
QST+tlU9Exscuv6XSjCLMvdEYLd5uD2bMrt7UVuMlk/B5T/oebE4VtihfnrpNf4lfwQdOkI+vM+w
eJaIC96A/cesz2NxsH7EwwMSCPmhJtC0SyDe1W7ky8f56XvIf1bR69EhG4DLVFcToJag0lpfTRXe
yC6l/I/1fX9+PqHmGhynLUKBJortpTYbMP+6mCm8PUP2USH/BLfztbNzf5+yinzH62R8aueGYaVD
iayI7p54u8mafT79RXksLEsWRE9yX4ZxKjVFD2wnlCTI4cwaAGd1JwEW4JjmL+i9EJN88s7Ef9aJ
HU5px2rmSNS1cpqTJQ86K1wPLW0vxKFBb3SGyRT3DoD1VmhLhpWnmaHgUV5Jmr77DEfyUVIzxM0P
wTz2ukfKAT20XK8JutYQd6WfKANt9W4FymmcVjM53FWnGxTtJOkm43CQpvEtkI15b+juAcCul2Vp
jEC5jUdpdTTZCH1mOpDFQ77fxHU2mvp1Ar9naVBPikuS2/384HEJ2FluDHKc7F/rdViHNSkeYWiX
w98ZMHchp6d+I7KQ8KVJ6+k1oSaBwGt2GYkw/n7LKkvDs9jdp6xZNd/uZE6vgOVYudZSQIi9NL/F
KCMNQRcngJV7F+iSMAeK1vJqZF2FFw2M66HRJ++RlK8G21kIlq19pABTo3cDrYNuDbc3ZgxMk5Di
q5DlCBeqZldG+SAqSbnAc5SfhBBCJijCs7viMSzT2imZ09kLe1Np78rdt4r32FVoKlA3RSdN8tYm
km7dkxTQopWhts80/b9WvqAy1ARIu6UWfk0vwMjFk+CQxnPxWxxxAzDljctoh4uqWTHvgCd1XmCf
5PQbVwhoEiKVqGtK7K5qJBCFAvPe33x7qpi7/6kqMJn9a7/d4tavT5Nsn9fbL4g6Br+/B2VRqPb4
ciTmf5oPfD+bzLtJukZAX07uvYdLIMgPpCmkIBMbxwmgZj5uuoJs8BvecSjkvstHGqsehK8VH2yA
tglWZaGBOU82nywgT3RZpsWnjvX1mD3UPL0K7A8jmC+xe3AL1NbfCMcHNeANhwviu0pQOvSuG3ZV
2ZFKmImITDR11bEFeJ/MF7RFFheuYZIvEzmlOJJzDV9mF2mBQMITM/xLv5UpZvigvVAqlfe99J7u
ZVYHfmFTJQFoz4OsjLZwyIAqlmE37/aeAuXjYVX1Bd5/dKrJnO0qbEvTvcsAIfMBwVvDN0NEjpJA
WkGD5GiMqf/x5sDFTK2Jy1W3ZlrYjljjeID7KGVdII9eQNfdyfkhJAn3RZg+jpkv5wYdrpe28NHd
dpQ9qAMJz9LXM5HXCSTp46X29DEqP4Is3sOHqqG0ZWpqkl9Xn9zqf73yOY89l7+Vw646ozDBCK7r
rppqN6/IHkOQUfWDD9mI48bW4ZQWVlR4voTejNJZopdKUKS96EjNuwWxhk1ObVuKCGQP5w2iyjJT
4UiZ1nn+TDjXStOs+CEJn+/eMj2JU7hgMWbvoknag9UEf4moitVxndAsXeDEpNsmtNHUB1nU4Y0Q
kFNpQ7LxRFDHn1ZQzIy5FB7jz3mD1r77XQAi4HxXqzlmxQTWyF6kx1H2reSDO6w5shQNGg9SyaXA
ZPN2AMVeh7QrMuau/5Ad9vsRhP2eZpGIdR7qX0a2B+fZWbF0Pby94E+HJUK9ysoPyJDvGh6jALlr
B6Rb0yqZqNv+DLuNFu7Q6lHQKTLpGlf09UkXs6LeKGZL8iQcMHjguXP3MdcGOut9Fg/m8nDC/Wm0
EnNGqq/M7m/dO828r4Vbtq8y5HdM4eaf9JGIC2fEiouzx11HYVhJNYYJhw9sYKDA3l1FJJvUFcHd
2VxoO7t0Mb/2P2wmqyYcelKPGfBV2RIgIeT/pJNB0qVLYPunZj5DQIcsoPYPZ3cx6+x2BuoAhxoC
J7HDA210oat4wIjVl4cmyxeoQ6EMsme+tKpSG3KXfGgYFpTHhJbdyIpLj38madfGweC+cRZiVeAL
ELTLqa+A8i6b/K2ZMfyFQM29PoqxldG1yyl7J2q9SOSlGS6zVWJ9cvFfNAkAGMuRa3VxCRFfk0Oj
dDoE+/Wmiog+Kmn7b53b0aUkleBrWuDwi4/IoKQ39uTkxhzZ42DDMvQD+XjTQkR5OLqVk23b2AyV
8cRWKJwdEGlnhq2LISEJyn4Hfzd50SnspwN3S8z90VZZEtEYY1k+a0fXh0t4zn1vCN+eReTOC9K1
lDqUR1UzQ4YcnhamX3MzgEYfRIQJWQXc1JyNJ22kEoilz6g/NpXDbvj2nMzc0tpuhWQ2hKzL1jOv
RKr8Hd0xzJ5JF9RM6ZqIQx/wS4NtjJsmCVLEPg4DNc/gj1mU1eMk7PyazqklfUQCEvZs5nhP1qeP
BxvSlFeWq4FUmCSTqRuHUCXBFCmjJXWILPmSMq12++Hd7+Z+c2fYYHs03ghGH+QwyBjvo8lwI84P
K2StLx36y623weukQdujLCbsSXb6HvXMAFiZtQcyKxI+NksHiMvM2Bz+/DF6ABKPsDBagC3CprH0
X2XpS46g34bOhFWxeoLtwYy6Q67HS4Ih1r4Vt65hw2E/fXlfiD7T5U3a6GfGroLHacHUUpS6LDId
OxLpmyROfr4DaY9osyMW1ykAmpGNRtogOHJo5OHuvuF9oSxzybhlsdWWDpbyJgw8z9RGmDPGVwi2
ABGgh5H/DQUdj9quqRw+AX/A/kQzc1Qt+66gr2IwmTmzWdsODDwSLZS9OObzHMslppQd3JyMR8l6
h9sOTdUr3JpTEUTLJ5UEdkAt2GxwXf5ncuUrVoA/IxBZSCj9TfH3RKYC9566A39Pe/a9Dy3p4AOv
qQ/oiiur0kUQTp3ufsE6pZHlvfadoxLhYLmLqLebhfKkAMZDRFOVQWB0kpwlrLAacNIUqvOskTcV
Lhlw2jE6v4QAaXNRWQDaAkE3gJD6BnbmxIBm3DY1jXdfhLy59Sf54ESqx6BIxu8h3w+SpfSYa2KZ
O0Y+Ye1wYu5drZeBW87BDZH/mE3X40a/MkCTqL2W7Z009BG/4InS6Z8ZKITkvCLVMGvI9RjP7E6w
Q2ZZnvgHNYz54FNfOwL4ua8PQTj9u+1W+v9CPh5CKnp7EGWflE+gbZfVFty3rtGZG8UTZmlYEXPH
e8ANBYnysUcdf+yIOWmegkiXzaff/hF9zVpxUCYBqZttwNeklH5d2VblmUWwCEss/yAdGgP9igNt
93sX9uAdu+85jJAl+ENT8M5pad6/EvjvCWeB0ZggKfD7GE06Po/C1rhq5MQhKuDaHxVhNHoow2v8
ujH9vUkwhyM4V7gqnpXDyT0pyhXLG1f87Ne3NJsTfW3A0hzRawvtaA7JjqBdSOQEQJ0fYvWJg0MI
4fStUdMeckLGHHm3oF5dFKTctruFpBZGJoaBaE7gTs4bwCUlhx6Put1wgWcjfdtMEsADnQ1TRdWv
zSGjNzrgfMySHu5FMOfD/O7bLSmgrMdzwd9/bt5Uk/CeaUy+OtN2HMh4ELrR55AnSL8xM2SIVGTb
Fb+pFT3WBQGLp66wRre53a089Z8Q+8iTzH4SN8jckFZOG7Mqc1iiOFkMjHZehePnA8xT5n+Zk52g
y0PD4OexZgMEwWbL/s5tOVipPajlcVrmfV0DHB2Ar6hWJv7n41BWMbUetDe8sZbvSe9vC9FEjEmb
1LwdUt0VoX8YkOxeawNG8PBA86kyIx/M4TkQ2mCXYQQN+VumYHrb+u0xwe0u66magfCXIt5u8sFQ
iQNQ2zJztNRuBz7Fk0Nm0gVU9eUdkNhxfFHMThxWPMbf1I3CdE0E4PH9AFypXBg8hJvIpH2n6Msm
Z2fndpF9k/HIyeAk8/aKSfFnhvwNTVCw3wlWU4zB4TA8cEjMARGhCUZYEKqdzuow6LnofWpKCMeL
iJNJL9pnffmgAHO3liZJr9BtVwm+96jGY0hycqzKKlN7bHajAVA3S66CmlsAcpnvYL/T5BDXwUj9
XGBd6Ja+gB0IN5JBdaMClLO+IKv9wPGiA677VlHrQphWOUZ4VkQI3uW3v1ioSAmyxdw5y697Z0j8
pAVH/4CbhulLcHFO/pYBxW+2GK51fr0ZF2+EpAdZW/O9K0WillkEpsAe4PZMk09l6llLyKHa9KPQ
iTcU7Z+Vx/D7TQS0VSD6vbjSoi6wkaK9d+l71+EwqZ1fDuSON9lcEjHIYYmuedMD2UgQlpWI5OYh
bBxVTGLWhKFfQZQjHfYlOOBD0DDx1v2LRLVg6G9CF5U7AgVlKBZMNHib4BsN/9d6lKeZPDVdfe/U
0BE0duqs5G0kOMV5ae3TcW4Me2uMZmgj+wb6T4c0FOXNLhdyWgXFGyUlIHbHBZyzrnpQIHI3e7+Z
c4GF4NQfWLI07v8Q8EuLS6efPWmuYsWhCXhEeyPGULv2yX/HdX/wG90VMSAdSuhhj25qHNn5C93D
X9ZJq218B6GfX0tg+B7iyfExwzMbnBdP9t2d56YBPGy3N2My4ie9YkR5Qw4+R6mJuCgJQTY5dvSy
q3TbZvtJ3WbQbuZ3a7zJ/RSImGQ/9f3+wg6DlS0ZZGv6DGue6b3huJZoi22XIgoOUV3KOfyn7+Ee
GZt4V8aoTQJtkeQDoMDUgkQp/mRpxPT4xv7bvgcwSSXY5Q5XKQvW1WT5I37/hZXQ8bojY6IqH7DV
lvs0v693W63Ic5Gr0zQd0/wfnSUVcgClQCsW8WRJJMvVEAEUMuOEczleX3hj3hLzFokY8nLIdt0e
sdz8JP8Ax1UKp/9/PJUbCbNqd1PmwF2zsU+4/my0mq8Agftw924RqL3814zoU24L10PHZfS6h8HB
IYXMnFKjkdv1vRhTZMw3rihuuNQY/2xassckiUbK2Hjohq73XOi27IHmLZwmEdRR7ISyRwVriz2E
PD6HpNa7XFQNwKCO5MDev8M7eY+s5eaOyCvOLeE/tiKsatChWIPagVjHhCIVCBImxD2NmtwcZpk7
KU4fmFFyu6CDEbk2lNWDim5uWmA+9McgMYQPuDhXYGl/oxhnFabH/Ej5rHopx2dgVii+E+YbvnI5
QogiVYsab5JArqH2mKeuIguUIk4l/dMCi+11rtCYgqqYWB3WlXyRmfPAqipMi7q9MXIGYimafybI
KRw53vhV1bb3IqkYc0htnoYNfaIx5vYAz0/hJoQEL5gmKhe4Kbt0fWpPaB3D7rL7vQmEyTlRVtlf
YkY9CkjLjCUv5skyiPjP/zfaVe9GYcDYXQ15e21jqvY2oz79iYUTvZ+WVZmCgyQjMMa0L3JaUtcl
Jj5mYAP9kZL0y5rJYbFWJQzJJzmlR3ITYnl8PCi4Kylfn/Rh3sbZoKhXtIhPspXR1Ku25T2QiMpG
cPIzKhRcuDhQKkdomNl+nFY6RHerfNRLUESneGGAOnK4TMGujvjqA82eWrNo//MVNlHHjC3u7nfG
7lP0c3f0qrlHmDHaaeoYCUMkhygvDWR5Fd7I2xknWIYmhs76ZUaG3PVF8rtPr2lFxvxpnn0lAucg
jp/UM+93V6016hIQN//S1xmgqO5anvZq7NfsUj6bb6K93GSk4oP4RDCYnP7sxfp7sr1w0p6xLmNO
HmSOhmErmGp3X2qRw8QZ4wSseJjnBFZunGNX3J8E1Ya3iNxdmzTrYeZ0+Le1EJGj4SIJPVBpgm0U
vNNPvny9eZwxtMWuGxPJqLr4Rps0IwCBDICR6iOiVMTW5X8kD30fWzMUWhImWdJj1/3VyIXRP4oQ
AsQVc6HSK916j0D8Gq9R11UShZ+q6by20giOyOechVrGfHmuFGZpUuMD3HGGigkBxqC8eB5nbI8o
uj0pUZ+lFcf4h59TUWk34I9ZtcxgFWS1ysU9PSvRb0Pi36423T6ml/kM79OqOmF3xjOUPTmKF6+W
uM8bF0MWq9O+zANdIOg+SASFzpcK1Fm89+KSKWRQaXfUjIaJOMisCVlqPX3qgWsHPuzOzWsJMk26
WrUYLPzk/EQYTO36MPA6dD91At/hNkNceRT/R4wf6pVGANXm7BVlvdsaZwTmaqfFb8jBjLhPSgCH
RPUVyuu+vJEqg5xEx5o7sFSZ366QWc4hDWL/fBLKsinORcnRVZIOWYg6cccwlmHbWxkax2UG9gfO
M1GoI2Uz7SfoLFboiQqIyxWQLmj6jDQ/nG4V79prc3VtNsJI6WnYpeXbcteeA2qpwjY+KsAOiHtv
zaE9mfvCA+KkgUITqneLDEKP0TeWflAp+bYXXX/X0fIKKwP0wFcOyXpBqbH3a+qkh11cE+gNAAfF
ma2QvRUsm9MJHRID8maIGM535+jIV/8vDZ/y2E6N+03V/GGdATWxq68bQaDs3Jd58y4s4zp+7Id+
rDo07La9lIRXRBLmKDGTHhG7bRz6C0Lkk7MicuU9zcUPiouxvk+bpimeyrS+vNB3gD4ThbOChwDk
3HRO712e5ueXQ5iNGHbUQVQ2moz9mZ7407/z/Nocp+XRYIL1ALlRvZubVNyuqg2j05ZyUOKxwQ+H
PZX9uqhfdax0jLvH0ep5UEjK3qKsgvwJ/xlUTBdf/dCwlIyDvNAs5hCYroRYMBA3dLClSiU2KGkO
5Id8roGLZZeteBWV78pIfV+ahIFj+9w+KyGxrgat5QRE3kbHI0fxBE+cQgPkRjdIm0sXGhfOt8kn
0SNen5Va5joWtxeLba99TfOsvQYNxyjWqxhb3G2Irr9CWqKijhLF+oscdytHIL6bP9q3vrv2vJUL
4+VEzFWEslOP4HNk5/0SiAKZ8GDGQTrd0cWO+9lsGVJUyrsXVHZmumSU8XacF/6A+CQwSqJZcIVa
ZzgzkdehIfW7rjxOs7VrWa5piNukR/TIe1yS/HWzORKIUAmVDiybrg2Re3Y8184pyAufEBEFVK3v
GTHZXpYHYvvq06ogcdQhYu5rr0dU9F7fg/9/q/Q5OdvI3UHVeBXSv3DEkGEj+Y443/+NGwZd1rAw
spetpkeHkFyiejjH9oq1TnmcvgE11KOIqtkXInvQRToYEwXkcBHgBQ1HyZTRguD8eeL8/9h0efgG
2veKxVc+2YJ5nmWPG8ezB9nX9Pa0VSHYE2nm2kvBJtEwbSDV7iexd/ozad75BBs3RaYRM9Bt9V72
xajQuwSFjPlfwOaqFrUmAMxjYfdnvwmptI6tpUE3PzzJtUVkKFJTpQPZwRoU6HdL7U6OEw45mTSF
y0Nta23JyXeCrXfRTjP1wzB7s3Ktp9HXRna+7cxd3SldYd8kjxiS1CiuKh1Rr9UqMaL335DZ2ujL
XKTjhFpxW2ulNasWybmy402H4STirfK9w7TtitWt2Tr5WlNn/FyQ6PM8Z9o7fKnyD2DLT379K+jf
Rxs+9HA0yVtoxV8/e3PXyMLKyHBxugOFg6nCLp+Bmsw2bw+JPmmOLtfsHpjxvTxq68Xe/bKF015u
/viQONzI7FWH56qb/Og5Efp2FIP5nAsfym9bkemJ7XQmZ019nCvousnwMwekMURhifNDC11DYwUZ
rGXYTzbFZLjm6f6TOJEAo1/rK/IWdk59pMnW0KxELJRZYMpVjKVdsMA3Pata/qMgGS7wkqGLu/l3
Y2nf5D2SuGmrDxiQfAAEmO/PpNg1BR/B4PvyCcLK+zgkR7PMNUNLT9+dq4F08GJAhhDXLJUTr+Xp
/pn+W7ITb3BUkI0OqojYUzfagZMQSd2l7QWLzTqWGehLzVqR7l+qJLwYNuXyBMCypyDVXpQASfqM
7mrbP1RbFZf4L8Hdv9uxWBJhVuxzXdTvonZG62Brx+3MLM3evXXsEWN59CW1fRkFggqmz8HQFmSw
OpzlCSWBsz4/qBUsCeV4u0CkYUwoFblROX0aU+qFXtYQ22S1e3wBmWeaCCYatpV7834+IL2wi2oE
SE+Wn4Wq2Rk8ANCJw5OBGSFuj2wIWgswdXzCH0DS/l9NNHEk9LEdeZDdyQZYmI2eD2gvq47sQYH5
cYU4sSaBT32YXWYdk+sSdEV3G0DbN0Er4L1yHCW2W5e7Epe+ZYSicvO3HZgQMvd1ALJmx1t/nDoZ
CpumpToNQ1S12ADucgXGAnLp+EfUr1e4BJaASEAKIwxEuvC9hFyz+gbi4vNHAqftSyELeG/c3Fws
BC1L0iwGshQAskDpGKeOchf5nYtiWYFN9/p+WVtvsDnmgnE7Ry85+fiUtSxB/OBghjhaSz8vFUKz
f3QKgQDC/Ha9VHdabVFIj8aGLgYkHzwRsyw5iZejBlFuy1uMSt4xRX65UKDkc4Iv+vgxUq7U2vjU
2TFCDK4gQsqkt6TK3uPkZJ6NYvWtH9m9tUkcuaNhH/FTf7bDXW/qsV78X8W1cNF+2zEyxyWumjtG
0zRwv2ctUgPKijwHaJuWHMMZ6FwFSAB/Xt6nN8MXW2pDOJHGTFRKeEq7xpzREHjm6ttfHIxF8vJz
KfeW0p8ZutHFC4m49t/PIak+2xgU6Oq7qjgghym4VVw6fsPk3jla1GoWb0ZxOH8z+kJBkubxSxp+
VdeBj9k9VBEWfU9R+0mWKXT1AQedNgIuITuP77muQvrSM/2ajjEv5GznbQ/6YMpWoMzudh2RRBlG
K20y46wV9+pHhwcxm4csQxVichxafovqQTBAZ3HSHUmUPjPPakRWRWpy3s7m05APUG8hkV4Q5vE0
O6CBGon4lM74JqQO7GUgpdACFgrVZWwvgvscT84usZ7H5MYsd4HsNo/MktGvdta1DxJ06YKbik/T
aXSZeydbui+LZUXpu/S2PjHaQdLskIsVtSWolm+xMpegF9+magJVwYe1Fys7rt76OcxcwTSr9/zV
xqZ69/9oExGoLIRobna3MqBH7c/8L8JJZiECkr1bp9Om1eg5TRvrOLd7jkDNKQdmV5e4A1nLhQ5i
jNCA7c+Qsbg3sl+2jzasKEbDxMxsRawV9Nq+6j/y1A0WVjSogvn1HMggWTXplsq3sORCK8BvBzVt
1xGdQyGeF+Y9bUpmKO8gGbzcQW+wNpcG44huDB6SdlGM5nIfC1ZM7ptqZXtg0O92+u8N0RZhm5/A
72j21YNFf0qWNwqhLzz4RatZz2cogS5rCo+sOqYoYytPQGx8w1xxfML6MMSCvzYOmQoqEVjL4J6j
cIYcisHyPRzpfeHJKkLj1PBNrPMxaXmL20Vnjt+k2nhmg41HOFaV1b4N6Pl9biBegp0T6GvgXCjE
ETO+1YMsbgjLgGeh7m03cDUQ7ldItDbTuXcKNvWdULkMnqI6VoOTLbRNSBcXBVyek4d2ep2PtD/L
Cbt2rUSBgmtsLqJwLiM1icCITi1Cb9s0wX74TnEg4XaIFpnZ7AzQgvzNfb/dK+Vz7TUyuK0qh1Ur
WO7EEmQ0Ljdw2QiAwuGgmuk8XF5GOf1JenQqfhyiTMT3mbco00HX+fvWLyvWYhbQQlpzbbvukQGc
882YFMJBygepifKV61Z1THOesqYtNTe9qlP3vLCV1brPGR5VeFEoGqaCqZDOrQHLrwXPMiJVyJvY
0b0NfpvteJ7znYL7AEM1s7WdngoBkFB0osuxp1e5otrRvZsuNW1IQFS1jybsTcxaYwcEvXspzN06
FiVkCDzxRl8Jp9BQBKKT6Rok0rlbqDbchZWtZEffz4tqNU0r8jHb2OtqT2CzKU4YCn4NtqGzTHt5
z2a5S75mNwQXodq/jaOme4S4G8TsLEb0ndC54ZgiP5TURz6MOgppzFi0pelgcQmA2dr/Y1RVLEVD
Xp8DLG0Lx8XwFWR/DUD3WpWbMBg2sdEKxkbCtp2rI5YjHW4M2Uylf8yBB+RUnfT1Y6uI8tNx6izc
B7k5jbJrMpE4q89++ZWy1z6xvkxIvs22cEP46rfWUMXTeFMRogsZuZPp2SQsqDHGX3XivJN2kpFR
4Mn2G1q4xxiZqk3tn2X5/2Xg+OdwY/ZPgGQJjMALiR8T6IhbHCZ0CcElG61gLFF31j0hvFrWBwqN
zkWmyh+i9IrNJI+wCY5Z4m0A/vYdFLA+uN8D+4EwTx+pOnm3tweIaqrEqOkA/NMrYmG+9/08Av88
qvOg4ZQNniQYMkLmfVNTfnNN1i3UeFN7Tzn2eswO4oN1bE9Z53QvvOBgVjlpcEpHX1hztiXEnUOi
zg+NivGItqThOt7Rsq1qLaQyJApM1UBmXPgnFlEKxVhWteTN//URsrtKJSp0Vy22RQqvJCANLfih
YjA9ItXtapJS2lEpzbGWcuqvMpfRUO26EvQ/+co9okKnyNCob97oE1ZH1ZpMf7wzLTA0d1yicA/G
PiWqAnreme23BmMHuV0JaStG7EOJK3i5uLzyhrSqZoSpOw/S87DyzmVxjBMsJG4rNp42cLcXkyKW
NAamD6OdZnfeMXAvnnnmcWd33BKF4mn7o7BgtyqfN3L89GjaJsgVTi4ORe4fGXoeF/8vAkcN4iVF
r5EAJoim6BBg38RzWylGsFjmwqRU0h1balz4ilLyer9GpmgaUE0+p9TupZHKz+ytT2RANiner2RQ
yLVJ/ah0tE3Jf42R/Tnc3s7QbhDKNzSf1XgJngBRpi/Ytud+X5HaJD9bfo0xHfnazsJxPKyROLhP
1FOXTmGsFRfc2KGxWMtMtqI88qiHVJghSzIVAHXeatPAdnmFC5GTTUyn67GSRcgK6HfNB10uAUe5
5kK+dK/rFsjtwOYE8NsU+mOmRJmYgTW69FYXPVCj06y3HUFy3zKLwTiLaxC1cIpkebQm8p5j5A9w
YB7LxGhY/dQ3VMThr3FWiwPj7cITz1XsmHvgZ1GlX2F/1mU/3/Tfcx1TCWfdmtXghv9TvqKBR9Hl
ovKgXaQCPUfyrMAfb/UB7usZe3BRgwHRmW3zxPecxauhXpnztGFQOJsMdKvsfpdxtc3gW9aNFRVo
lxJr+AHPyOykqxS4aoHMw8kzerGYZJ1YlicjpnaTBz2fz4eT/HvGyD9cV1G1jfPe98AA6aUDq+Ft
hp2Y2S05l2N9ukBvLU0ewaIs06IUf8Lm2iRnUkEzbs5SIxd5zCf98bdkd8uv+4JAl1ylRzBSfdl6
3PIYRCmwpMoPC2droXq78HJHg2jg0MPuUFo6Hqp3LPqIe5X7XrGCg/tT6w7WKUky8hIvYlvVpfgg
5PT3AZFPYJASA7Pu4oAgv4GgZGoWuKDoedeERJpWxLZ7QJrUPVydOlOJlIgZ9W1rG8TWiJZBbngY
0sDwk2giUfyZZvwgZu8wxv9xQ1QJ+CUQnmVOQloTyfKOWg4nyKab1KOBGJjPzTgmNNMKa8N78DzJ
Zhr6gs4+Fgof3II1wVVnkKbRBhl2ncnka40bqlbcX72tk7DqOVjfTCuUjt6iar+UOVa/z+uWRBm4
3CiC/1D6yWgYrNpAjUv0+AF0kd2FHRlm9wfzCXVlJs9xlDzaZKp1QjA+FVhJyTcn2GSD4PyygPEN
8yuVuwOqmScmQbfgFMBKStGYxl3c/y4OogHeChNelOe3s3gBEaz8ge5UWHJMEzsE1pDG2EmDrhSx
s2cDSWgl2I5fIQmfgnQEJU2OuuTZ1XxcXZCMe5ar/yXoVsOx/hvtA9pWGg/PAOHkp3Bh8UZP65KW
WxOjpSGZ9/tx6YUYmVFNa/3W/ts/egCDTG4sSxvxduebYVoyJd/9yyM2IdfasgRwCqjJspOMWbir
YnBpco9/JgWBuJJUn6bOCPdOlkI0q14+N60IZKQeJtqnx3jalB8nJLJRgSVDakFajFJ/+s5bhNjz
WJ58qYit6soUkeBJWTijJ88gZSJ2K6XedCzXu7tw4BvPB9PMxYVUkHx6lcCx2t5Lk0OyCmpta8YH
dnhQoUzSfeAuKLqEyccK2+WP8FReRYFFAV6rJuCm8xmz/ZNbmH42K/vk22rPkxWHWkvbIRXZ3BAl
tqKv4e8MQoZvqrTuTkhLD1eoPqEg0ncvfXWWKlZf3OSvXpIkO6GmbGJugdoMPyZ/KqmIT07yIi9p
UDMtJ95p/uYDugT0EMyghXrqdpk2HvlF+/KQmPCp/uik/PaYcLOXRurCFgIQIL3zUxlUgc8WvjSZ
ENKfpsKB/cqR+r63M2IAj+QBhqX5I8iV+yza5Z4gzRG65wc3jv4hgzIlqM+aPfl54RoanjyyFjZ1
vbMZfigAO5eA+1HeOSKAKSUgZOqGqVnps+z1PK242/tXbyZfsOz/g1Hvp+2g0+NVih8R1W1fnzzf
nNgy+F2rcg7ziTr8xT6cOctUOrIk8l6tbEp3Ic8fqes154C7TUVcJhbHaONr83ZEAGg8xKBfKz0y
k8iy3h1N4vpCVKUGvw4I1cVPvJm8dffTeNg4LkjYIGZO2dMCbxdyMNfQtoIMq0F8oZ+osIWjotrJ
gJkXYCIrspJtB+SgWf1leehPOBeg91puFGxmNZJdrtF5jeA/AcKj5pkGoyy0Tj1d3eMdyL4+Ww0A
oAPpPvWmKSYVjug2ZK0lgljgjif5QZ6pdO62z26ZToSQhrnrDOECLgf5OjyFdS750WfrIxAGj7Ok
ef6oYY7NKKMMVOzbBYg3jWLZv8/rgXxegfzMDgzpwpnjeFF2dVCp7SB8/Wlbon/tN8NB3T57GNdZ
DeJhAQer+Y/MuoCZFUUeBNYMUSLE3u/Dc5/JVYUJPlw5nlVgKiHxRb+JlKAzpCmaThgxVp+jJFlW
LJ19JJlxO4TaMTtmRo3oWIdu9nJf+KnZPBcb/lJ/poxl8GD9GEXXXAWyQwUvj9R5KTHA2B4ERu6J
NM5snPO6FJ/xj+cgAFeqews+m/k1HE3m9dDio33lZBNYgcI5lOKJN09gzGmCEDGzzWdyoeGDe0yW
b11W4D1TX0j+hBB6nvGntbLN9dRIKlNnEuE5QDAlnGb7UnbBCE8xSdRjpR2nfxb1Sd9Gcxgp5NbH
Set6s9mefObEeaO2K8Q4yviw8oj0HQ9SbORR0QmIlrz3WLXzj/uEAKDwbpb7askhRY7qcTPXyoFc
euk3BS9foG05vQADEyCM3AzK4kyHku/59DmDIbbz9hMm1BmYiNzzSf5OYJty7bkQ9y2qRl5kfTzk
FDmCJ8Oo8IeqZ4fKqNfwO66Nf/95ib9to8kFIipgsT6BhinzLvGuopLOAQSoCi2W8IntemCspBrA
Qhbc1peG+aaMZmmqLkxAoNSolLZLbMpYtXC62aRALRvEJBlsZp/x8edi9A9TI1MPv61QqbqYvn0k
mW9h1Xh9TyqAEKgLkLF8+rHmW1hklPV9k5pkkyqiVS62dsgCHzxthVmd7eQQ5MoTtIar31ATaWNH
Wtlhrix6FWZOjdQgM2ZGDvrmsMksDkBZuBbBqrHwBIBYjNrh4QpFmNzjslsklQTtb0oFcmLBNzue
pHqwqQaOmHeio1WFQ7zgtJ7VF4+PSxbXAxwrCN2a+v+DVNT2bKqDAfaJdxSV47HB+yzj2ZwZJFuG
K8x7kewyrsMKXn1dSK36bXxlS8IZ9xNxImAtOFUrQ71zqalBdyAqrpbwa+1whiTn0oFZmDB9npSg
6qTEAV510vamxbCTrN8yV0NyQWJ6ZEiFWrgqZ4zeM7awR+FDrutFemlTnm6CTgOgbYPwhVzs6KMG
MTWAnHWbCbHN+W0J8ybhvUYRPfmMl7lPDHfnxaeUg53SEHTT1P/6iWB1coP25tsDv1oMk2c1YGLb
qUidZ3VVGk5fE1qG3+rJ+1nlzPBiqgXfoJf2tb3peQWh12b/5pNyOyoARRaRrS+2dCbwy52o09Ts
0MJNyMGn/5T2KDjmbFy+GY2SVAI6wltB0wDwd2B119WbfCNvu5oisTlv++No0kbpCN9AOtg9utiZ
Ce91Md3JDVgCxlCv3pKcksGGC9C+7RE/KWhv/hYasQ2nocztxjBDhhTAFbKLggQV06NANwRO4WsW
zgGWW2zhIcj/OrZQ0YdlvK+V8RDE3wcbRohrqm7ZPTI9G9kRW2GzfIuJxm7TiE019Ry05IrNab+H
7xFRAlzSYG+m1+kCpOC84kQw+eR2myKyDYs+SqlSViUlE6JwX1mu7q4/K0/F8WRuRLdAb00FCKEl
ZM5RkSEI6tWdydTV3vPtUHIZOhbMcqzAicBZbDv3is0NMuS9HUc5WTIPixmaNKDQy7FZKiwBu5AB
XsGTKdPiugQNVn03XbZ3VTHW8RzvR+6cqYhSQmQHggEIZci0fSme8Rtn1+tjUPYTzbjaYFXgJ8ZU
Mk1dgNEiuewuF1mlc3EIGz2wlMTIKmE+ICZGe7YIcCpYyp2nVx1qJKsyse+dJdgul1biJVxsKCPO
hjNpXcnWIA5SX7PMUp9FiIwg1/ZKPhsWzZghlqOqZWmtAGFu50MZD7Ua4M29no0knn1Q4t8QVmn1
rOei26O5/Iy1k3C3J8+075JENNQL1bH18sKhw4+AN2YPxzZcglvaOoypl9lCTuYGoIEqswsLehZQ
9ALSiCclS8sW8bUMYnuG+OOLlsV7HRIPjfjFoHrfcnJo0Yfd82NdlvWekWv8jw6MpOXzk4WVNMcI
qAKncsTixu+w6EwQVi/oMnZwQQloDN2bcfW/klZVBUkM0R7/dLLgeiz+r/UmvhKs4VsqZG6zXrbE
d1/HQbXqnocrRaBqqCTa5v2k5Vhv1cEH7p4H6xbBBpPAKh+RzNIQMM/5H09iBrg9qv5byhDhlyJp
T8k3SZ6dZ5YB/twxiUh0i2MDUr99lgx5n9R322mYQANv0DAm/l52eeP+yC8iXsEJqVPvlis2/lGT
WBdA6s8ZRM4KdHEK6WtCLVieSuaMg7ONXvIYR+vGi5BEhwwYVimN0U2V++5H/G25VsZ8e1OgqCPq
V7qDEZBTOcYOxr2Iur2AeJ/1Om2i9YFRXZR+4ym+VXZybOsj7KWgEFGOGWCSNUrmK+73MnSq01lr
nQ3nqQHMhGV4SDyyKnSKATeXnXj7usnUJgCpGWFBJaiBvltiHaQF5bd4gO9lScl6+fFcZDlRZh4f
bs7M8JKr6s8BnatpC7NKB2wLH7e7rnTNJfyVHL+OuUlrsOGpd7024RfQLzUMWy8POsLkQ5bhBOHt
JEV63hU8/Trl55n/iobPGobdPi0ncsdr8sSnuIoP1w4xJidLrV7ApsINahxSs1pyYXLfVRF767Ps
qIxSokb1btiRSFndmvEmxDwfO4sIsNdxH4zt4aMubxAY6x9ZxJMYsEfTCu7LOkH6EVhLTvvQy/R0
duLAWLGznAOEzfkMun1F+aAxFvlP9K8nHtXBeEV4FH3MOeZx9k+YBKJNNjCWCuOgeERgb3XF5vhC
VSg5bl879tVXF3dJSP/tLCkwElUs7ipW5qBh0ZqVuJJHCxVlIyqqGMht6ysZQA7VAHWQZ6RW+k7m
MBJgtdRixHVNIUAaL9Rj5ORp5W1zZ7tYC3NP1akDfZav0tSHRxdVD6iDSGzB+LYitJ5sshROgugP
q9BLKwVu1e43uXNONHVuIsEYE9w1iLl5hWB9GXLZYgslSoNEKB1M/ZRXFsV2+F07gW/fKOlUJ96q
cIfzjNci7/gWSPNTEXbzcY1iTTdP9AKJHM5HhTw2j5abXCsdADBVakMq2Q9lrP39zhhI1IzedHpr
WKqEx1lj7iEaph4cQLJLMjgQ7wj5c2XEDudW8ns3dxiA9OK7hdmOjUXHDnjfVkvaOXfS7gkDZS7K
8TO/yqv31qtvA10GtmTson5bOUdVBlSTxYQbY/GnAVgvScD6NSlNwBYj2oN5TTlqnZGHsdZKOS4q
TQny66K3G4MopEl1MjQVW2pecYojKBpI65tHwSEtuWgOtETfyBe4GDTDQnAirSafBh5ouYRvfpW8
/Hbf5Ex644xFZoYkmkYKcKYaNoQrhqKUkTgE0O0k6X4dkmt5VERAuK5oi2O50Q9/zPEdkclVhcxK
9vHyMqVg3B9KothhL+dJh5UN4XrWjB/g7yvs3CYREUDWB0GcyTLDORGKE0CUO6xvDFF4riul0w3b
q3iyBfqWD+N5IMnAkortDFu23Ne2ygp1DjViOj0TT3nR/JMEpf5t04VimCx6j+6RE8+D+svOppH1
sJnzP79nZtS9SVoNBDJTFgijPPpwSDRSPvwCFrh5EXDB7WmJ3vBokzRqP647NMHM5XfWvJwmMVi0
N48zTmifSNFU6/9vtj5cJO4Ul7YW23RakgbK0uGbkzR4oPh4Hloh1qhFhFDnm6/L9g31CEeh0k2h
dvah5gFE/H5AgBslk7i1lpynx3aUId+DEMK7NJbjsDY7hns5JrElFp5xMI7qVDCDRHpjSZt2CQCN
M3AH+XxswAVk8RpsAScYVBMlGIq8dfS+qSvthdbbwGYjYmPDVjZJXZ5N5gCw9050tKiOKHtJxM9S
YZFp4OReds9oKXa/aOwg+5huqRb/V2hin8/tmKARQ5L3gLJTFFmz0K2+dR6QTEus+o/mFi/1esB1
MLlSlmv1kB6QhguT5gJ3ZdD0M6YqNVJY/eH0duUgBehLBlnHgmA7oC2JfVghbmlVQuHnMb3jNscF
zY52WUslIl37HG7QtsPIPzzTLJFJvy/ri65QXp1AvKAMDzQuJcC10cFDe+bLXOHK3kxyXUtVf7cP
gjyKAYi53UPph4gp9uov0wopexL3k46puxVw3XIlAjfpzzsjo0upuwrrMLLuuBNfbY+sY1hbJyXu
6RRCBjQo8soWqJsSAzfxCR7ALlzWMJj71YYjQ58LPtkhwC0QQZQF6QMFBznEvFX61XMfS5V2blsZ
aGc9s42RZWc45qVvs0ZObh2wTZR24PSCwgZmaDt2XpbIcjPgaB272ALFa5Y8kEZdIP0kC0TG6A+k
1Mu2HBl+CY1prgPPq+Wh0kM0kluYccCA96CNys/2hPnX0YsG9DZ4pWrEzr6kGHzgR1NEKdJ5TVQy
ZMfC7EmeLSgdsCQYSoz1MTkCIa8jcHy4upV0CvIgL+oB+Zc2rIZvqbqI8yPg8xqxk81of8ZG2v30
el0Jq80T2BkVyMv8QU1PUafpStr04a6/UmHZAlaiU3zTdmYMbR0bp2glSienalkolMn5er/YdxYo
LqGKqU5IIm73PnfS4vJ3++3hakgm4u1mLX/zUJDmymC+B1A1CdW4FPRi0gqHO9U4uD9ovbGT2TGb
Cki6VB4HinD75FEj8aMyQMvAUer9OEEM2CR+GQnbOG1cFA0iIA4KbuYnjllqYfflz+rnecjPZuWV
jHmtGhKT5vNcP6AdZaAmdtCNpdvlm0hrHZSWbjPcblf3dOe06eIz1hGgZhyZEd7psr+ZCcLNukQb
zBnvgMczpE3GasbBSnUMsbXm3N0ReP1fTA/GsNnX2MEB5i43dtohpiKelftG5TEve6OdtISiUueo
6dhD35xSviloD/sjDjqahBSinPgZYLkWhnF3C3pkEbsaapPrwIQF7iVpB8nLfSwB8jSSZWatDKTk
n6+6D1snY038D9YYNsPOH5HjtVbej8A2cHp0g1oXoBZS+b5pD4hWWMQUdiim3bW0yCYIcK42hGgj
YWz8P9KuZWwk5WWrFylaKcfzuWkqCLCWJ3whltl3sCYSn0GiUCu+xjQjWSE3d3Ns9Ez7MGpBYUma
FKWB5F2IHqULjFXm4gyw7jSEMhYH9rU+6kLDqP5G485Gg4emLYpXh7wZ+JIzVIZVXFPpHY1yBVAK
pcZbcihkCASFXp7tpIq2bAs9DzjgFCj/HE/4mm/QFqAsQiFuEx+SI6ZjpXhvMiTJYHzoWhAyX8+g
9ErQTdlqGaUGTQd8I9kjsjkAXGo47GHr2drxyvudzzSv/0z/lRPS9J8ruqbgRkpeLdy2JeUOZPhF
Dpg5WzqJnmbtF8cb48mxd/w4+J56+3EXfs2Q9MXCH6Nozk5tOunD6gFrvIWTaRZ32BhpQNzsKGK6
PZcatOgzUkBlVmgzdHX7b2MLpMgv25K3miD4Bnyzr3Dtv3TIIm0bNVS0bLi2PphiGEWCVlK8MXWI
VsFVLZz40DoSLe/hu1AqKZnzeP7pFj094PAolraJp/n3W/o1ETmMvDhWCjAtSh1VtuRPmZxGG2Eo
bfnWj99g6oXoSuq6gWHchniyBs+Or1ranWELcNbgapKF6vop9zMiRTySdXpbuLHOjUHcMe7h3eqY
6lB/eB1bq/HQbyZ4ccLc1lclezV8QHg1nVFU+X18pfR+jHQhXtVnb5pZ9MRsBpeWLCASyHd591LI
nx9rU2Kca5utxKH6PMyGwezmHymIxD7FzubfAybbLAG85/V6XTPD4rMK1NxBWVdfEUE77sW8LpZy
Z6moVzrpNrqBXNC0KMTAP/iLbBzPXYDb1eu/TEjAVEiDGuRebNLPlF9kXSRfqu9uVQRgxyAozH74
gc+fWIe/jkg+wEYtmycQs9qYaPqIlNpH7uDHtFJJreBkZGigi3HInYxkHTxC34OQJAea8vOilLEs
1UkDw5alyWWCYfHlmXzf/2HTX/vg+D7Kp0lM1fXXqOeTqtpTpp9WsDMlZ+Y05IJsgZJKGj1dOXB8
kCku9sGWLBY0JPIP1vO/l0N2x9ybMsc2XjrzelL0SIZj39x0baXW7bgzD6tTOIR7PZsaAcnNwtTJ
i+FKnHgRea/coq+klaqkAZV2F20Ztzg8C67BwPWse/rWGBM8M1Jm8HTxQy17OLYm3fzyAC3R9tEE
iTKYXa0ZG1PaUjPGE92xAO1RTS7FspP6E2jODoOH5u5aITidVKhaZmFsYSH7/YSZ+Xtyo941gOSw
Ft9U2U6v5SCJ4PjqQa7YH0gYExRDhfTV39TWbLJ8cyjEGCawKocn5bNbEPRsM0YBlrt419wFjNzk
0IR9Nx4ymMkDR3VNzr+td2UXNcXAYO8TuaCgyMt8qGkOLO9hZTq86IXRh/xd69VA1u2Nzv1rrskD
DwFW8J1A4lbV3XNFSGyhNh39YNWbnZBFL+X3nWEewa0rVDlMSFY9dSE1TW5iDpLBIohm+9ZI3h//
QX8PyG9HH58eUa08HWcD/T2AUFQs+d/d9tw2RpAg11eAAC7NzElkHoqB2Hhj8T8rUoFdmV+J9Sm7
oVuTaywLbNqZ0+bjFUcDkLnNTzOiHLksBqmAKDRBEXHPj+sQFwD26mo+knJ1OSO6P905MZh5yvdl
kTDpdPh6y9r3g/Abn9Cf7CDxBBlFcTVZKs1lMQUDoC4FwQTb+62HXFkLqjh6vTQ3RZkw5JfTA7hg
xYwvggMR/WTdIA6ZzK0uJgm1PxPqwa6m1A1P/yCOUnIO0r025GlVqojYAqJz5zlCnXAYF3GlTg7l
7Z088tAaY8/lgL9CIq0ICT0+OneTqUQwI7hJrITBOc+EQIck379ENG3jzvyujazLktDsBezvkPzf
LCEn+ACc6MoCiBxH787IBttzN10At+j+lDjtR/N8ZZaZgi9MJo9hrgKaALjlUqO4F2u6eFWZB+e9
ERNFTDH1liaT3zNVA8JhItzD1wYOpMQetxI2LEjzRzx+bMxdvmKsfKCXdg51Hu1mp/YTUmrytNbI
0uSv+ehAVXcr8sHAHu9BVcn5hiBEoGyFNIYP5p0T6SNjuT9NZxL2q87wJPyQtCAYf/chajlnIFQX
aW9WYKF/QYPXYfVyPVO/s43UchEKPFZCComBJ8s28QPdb1woavwiSimcFhptSVe4okM1rEqfCXFa
qNK3NYOOD17kD8gMF3zd29qPa0w/aYgJ8yCMer5a0vzu/KRdn461NJ8oqoMpJtyAXfswOQupAbNf
mWyMQJ95udHRHslB1mXXmC5ovWTWPP2K5XXdCmEz6eleOzvy6unTFfEpkoBKIGFTj8Hx01xFHYRu
dys8rV8vj4LCTy3PYcZrNgtoYyyeBk0cgFSTcNquuvGO1mdyhLf+CGwHszmBH7X+w6dkLvyT1PNi
3m4/sOVxCimcut/+pmlJS/skdTsGfJWOGP/vF3NeEdpTuv4ZS/LPJkYvANFuiD8BcbJqHrSl5KYY
eBvjNLS3vGR0c8S7FtbE+Qxgsr4PaVveLU/TzArbQ3hQTEgJuw2DqrqvzIJYrSkCf2jYkLuCKvPx
Ffm8G1DPfSNpf1JntEzbyM5MNOIwMMPLAZmDq7/K2LpJuYYRf7MjlEeZWmfGiSJo6966ilrNz76v
AqxFXSFFg/m0+vvvO1Dv74XC2b2nxyyOw0se6+hQTKDf8fXsD3r5kTxHpy/sXl/tyInSkLeowDpE
svy3V3ORtBF+whEdwE2icCXZVCvcjXltxpJr6/2QNDisq5ockuybilhVjP7KXeU6oQdFriqAIaHw
wWpkxUZL0ZAgyGbhVy5CEBHT4qmZsHGyPxohhj466WmBQEECXeybVGXNPi2a0pQzMCTFTy0nXu++
lJDAeTidJyBBXxQ16HtDMuR/mBvIPSAgVauTRl9o7Xff9diJRXJKK4KPpxH9ulswGQnu/hTDQ8Cd
NGal6nlAq/y/yuyOQqwIrkK7CEpz78zV2qJ+z7G1fY8pCfsLb+S2sb/GPGdzlI/gNPeDY6qbvYbU
d/vtxBO3mjGkGDUNjrasE+TZ9d94Aqzik0N+6zZKsP3M8D0iwWlpHtdLj7qhNtqGLz/lbTpcKusm
J80QgORGBPqkxQWLgo5HFmX1YmeZsIG5Iyw9xFpbfp+Oe9gADX/cxVvSxPIQZBU4lSV3dyffZAmC
wUcRtFr3TAnZbwbFdbj94OQ5oFteBCyOsZNdLaFO5N9J6p37vEboY0VIHUHcsJHE/do9q5BSS9oJ
2tdYYyYss6FChUm6ckT5Zz9OKJEHDEIldxXSX3dI94BrgmLnYOuqXHK1epW9LHHKgESD5xa9E6fS
HsqGMAKHkqjc9JArKznLjW+Nc2MYrBn+hK2vVo7hPrwwluxN2aqAuGEs355ePVB92Qtb0wrF9g4T
gT+ZTjNyAGtxQid5JalE9FF/mGN81Tf+pIeeRpSzcoYYvs8+DGCAg/+TsbCvkdqhrtcFvAbpOTLj
QcmhtqlSgZfg6wodGyVkEeqnK5+1IbmE6PSlgc1zmqvrVrKFEgc1fVnHD0dnNK8sh6Ho0pUj2ya+
5wiaQJRI9aQ8odDLqjRzR1nPlB5SrLVwrMUz9BymABVA+jPiDpFgIQWToWOPz+6NnSK2P7g3tdsQ
tn+octnan9ZlHVt/4/BjhTD4PdFeKVMbUXEvDF38v3Uf1qxcKv3ijdAmIcNWYP8eLpJRIfbddMYH
fDIfSCaOJW3qQwrOrwatHeMfxS+ScZsM2r+2iBkuxltj0yZqUCtwwF1vNWJAVyRVAiBX9Mil0CT9
fgG+wi3dmPBGoFY0EUZjb4Z0uqJHGaTKpXwcLo4/4zpmpRR06S40EBRjNHqOLxbvxeRu+EfE2aO2
R7lxpsPQRyD7wZdlMSwY2T7SIAl2p2huyrF7mpSOzA2776h5XjSg/WOhNZ/bKG1igy30SnEfB+vx
SNp6KLsSIVr5iUkx/tDosrlgKH5eT5Jhuz1xcFM5SD89zZgvS1gCmHLtg/GjKe6eBZNkK/OqVl5R
hbBoR79i2sxgcm/TjC4goYL2MMt7s/933o+wQO+Trik99MJkTjsXyHGUBnaMq2w8OQBVbZev9lF2
JzdZ/VT4BlzVZ6Xhfi6cqYUURGoF5a5HXh4UA4ECdXX+bP6Q5t2jUnKnldjlYXzcOQ162BpgLEzy
Lg3HgNTON5tNjRKwA1ILXbHd5ygMdT+pcy0M0b3KdDcQ/k3DEMg+VI8QorVu6vX+28RY5/ps+9xe
O5svPUqtVK9fMlh1LfRdnQTZR7VA8OqcZj9Tk+xbmptD5Jz8nZaGmECZhplv4MOAWkS6DzwbNElL
DDV8lp8bSp+8WgCVlEQvDjOD9fuDh2gFh4R3R8Fbifmmj5Gbd+CFoFn2FLSVqP0cjTbz0VQt2k8w
7YnqWyziExIAofoEX3Me9k4ir6BhoPNCFYYvY+R4f1O5v3UGoe+AY0fTdR9zeRaLoVj2wB1PAtZu
nAzCqQ+xu7bUqii0YXcG9uwfK+SJSDBOXHYxqp1SI/ae7OCzNIGUtNspZ3EfuNAlxIZZPEg5ANiY
g/8h3L/PvPlEqYSQJ1ekqkJCSodL4LL9lWaqux3HD3ZxShCNdJdxUnJ+yx0q/bJPWCBmtfonZv14
/3z37EiG6QhnlTxyxAi/WS9m/W02JV4zDfnp5oPJ8+bKelQO4KSx6Kr4aF/fTMWql2rnY5ccRWfC
w679/jhpBu9lxCZY7H5H8rCGyLj4HZB9Trf/y5xHJfn7Mgf7L8nr1MveD9NRuWJSnAIfVH2nQGmd
XkoWHtLBLKH1Gwlajp2ALIo7G9a38EFj4Hh0PhmQUwCIsk48ER0MSjBqNjpgiAVeGZGoqhnUHVEq
So2UjstZ/YxipTTfVE43DB+nuXnwEn5pAYnYFyAWtPmHW1rDwhmQ8faeMvOBRuTTaEKUz0/k5Ywo
0Si+OsyGWHM13JbXPoSxR2aBIq02itNgb4IH0IM2tkpamlfnvk3Kqrsbt2DQ+Hef2htFfjtX0Ui+
Broe8PYrRwaTF691yBkOl56bbd7YdpMAmQRWpzbXWu3IpzhOuRhP0cPItF+R4RHU++0yC83wZT7T
sJrr603kqOojbgz4Hs3Nez20DdsowmgeEwoXV1i0BEPy4/os7uDiYcACSNDENo8/Wiy7gUhci89H
mtA/ZKtgdEtQChxmWiPBuSH6Grt0pZuIEypzdbnptflT+AKZRvezGewqMO6GdAHllAXT5kfiseW/
BEVGbz3d3BE7Rz3VCOyEtw/4J78EHOR2Ua/8sSF6P1oa6BcNfT3tjCEXIriwh7Gd574vVJ3fCu9Q
JK9K6xGNdoPyIMalnldiuyCr2JTldDxTwtjRtaPX261c1FmN2pRgCJJWaLp1kM3F3uXxnpUy2qJt
Ep2j89/KIiuI0awgWX9DAbszB83BYN4k1V+aMDZh/foTW6N5XsBHlhK90CvEb7LG3FoIN7CTcU+k
2Aa36CEAZKrEfgITRWeQbDU7DxGH6JZTSlvrPratI9We5aVmoLzGBjZbqdCuk36etw/59Pmr6/Ip
TPVEpXWez9PBjxwUqjDWos9Xq1cctXyvMwmRsEPFDzUDi+TRltDaLFmCcn9p0PdcmE3ajxj47zxJ
YlfCtrRqxWj2xFvciFKMKaK3eRwnCGQDome943+Dsi47J1ohLx4YDYZfQxcDI4T4oL8DxMBeiZvM
+IxM5qzAkk5o8sWVCitspABiA1fhdAyPBuiwcnZtW6njZ65lz1Fn/x9Tf+aKUxe2wRh2JZ4rFl1+
/gVhNDiwaAKrIz687dr/8BmY1uZe9z4rgQOSBYN+3YSydlTSWJvJ1OvTJTLRCP3slZFl+0/48ywJ
CtwDn4kJyvV8TvLzvz1I75VEXS2idBWaT+FtSChb2KjwhQJLzMcdgB2gfkGJ6zX46W62ScE5wVsr
cWDq9OprxvP/kB4xclSN5j4zuT66pxK3Md78TViJvzi+amVdHLxDq8MFKM3kEtsoLIG5b5eEVi4r
inUUj1MBXlbBcoLNp1h0B4iMwSPA24Yv1XUBSpa8WyWEPZUtJADJDF54F8zP4eQJ+iQOy8ZpWyn0
TEJQn2VAajM1WPxVRqehIET5OO2BG8r0waOac/yaWLOJNQ84BXAVKdOuBamlI9iI25NHUHAeMqKi
k9A0bZO3X47ryTquniFadLLQiUeo3m2mmFsXRDq5JcCgvAfSFiAA88CexrdcS4DpHQiQF96ICPrH
/XFd7k4x4Cdsbz1oAiqHbXmYyWIVBOYM+ZYcTcBtwdU2DIqPZbGElz2tKpiygYe7X1r8SB9jPFNk
n5fTNjnO23aFlz+Njossd8x431UrEl5ZHl6njBWuBq4kAkO/aSNvlk8w1IUph2FcKww/48Ujii0n
ELshZ4S3sMvR4/eKjaGrFCIG/DCLAGb6CGCOBRqd8DxvO7Vzc7TMBvjd9XJg6RcMve8Exy9ikF9N
LCHFO0/6nFMjNMXfZhU9W/rWTKieNo/5iGQz5GZ+93qAkPLo2/wO0QR3msvvenRRbce9nGgdcqY8
pbTKcUacx+CdhQ9nVkFwGGkyz7zm9sEQLMorOcXz4CBrCq/f7ui2BM8s4u6o/6NAB3NG2pOLoy5X
AgCCOHp1EVjlisiXovFuTuF26roPl+2gOldzig3SmahM0Ln5m3D3FGJclOI85S9yc7I7X52ZonxE
5qKUAZY4UKTaFuPcCDJR6WwN3F3DErKUfzhj5r1y2ewUXwSlcnOFHb1Ah7gmYUCBy5I4Twe0J4mu
YCXj6fh+BNqurAihWjHpOHCXXYvs97qnE31m3AZOB0nRG7+cVwNRABkmrrkg4wNxQJtuDqidoLno
toh89w3J+San87zpRip9Eoe8TExhNfi5t54UGXVWU46CixNNdY3kAncDWrAbRhDOvxjLC8lcqOyE
tahuYoEZUHsIGcPkJDTr4LB9Hc2PgI8LvrWXMFtwmEN+lFXVm2mqBZzXuyYg4XtCYaRN5hr1sVr5
JbiJDgCXmVgkGIclRLaVB54KifDHYuJ2itp4sgwERxvLJhafFC87TiQMfF8L8trOFfqpEjIovRU8
blva3gsttE8mI7SkUxIqNLVS8v8O0Z481zBN7qaXvNGMSKp7SFdZyEChQoGFYlHPcjjATKG03pWX
Q/Pm7EhCmwaZkpLhpfwuvHETfKKBcGys6VcAdUCISUAQdEqPVcsVjOBMiSNhWrXaEQmf8JNpZLyq
dEf+Cst+uOVfcdMF2xKEbwGz3Ix2yy06pyUR6XlLjbt2WEs199j6IFmDoPGyh5s20h+xMWoMphqd
QeVlx5frkr19PDfLV7TqTvNRvuI/Rf4MiQE0OV0EtczoarDS+FLOWvjRQWYZwZ0xejejwXaTXIim
fWCQJHzfElfX/l0Y4aJudSiMTnuCzJ5HjZpzLy2AGcn3BQcm2yEQpu6+4XV1Vc2KyhJJ3WV5CyF0
1CqtC97cWT79bSi89Wvm0sdjLVLUyqDe+0WPgTxj07HONHErYCceou1UihhjVI0twJ7HNtqwaff4
VXB8b/KPUiAy/f7MyUq4HYjaL2y8iHcV1Kcp9xee0gyP7ujj+g/6DI/AtDcYjTvd3GCtxqASjesx
yYVd9xdxMTYkh89wZ52WqCPjfyOqEtJgNEdXmgn13rXSb5J76CI5I4LqXmVkfzbAOR43HocofuZd
zKjM0P8werrq+xzC4NPhwxBfGe5cfMH3D+Kt3HOtq3znq565I0DWfPY+eIjj9GTxO0KDWiMbjS3G
tTgzge+UpEIxXgZDk21GOIQdCAnU7PyIZfdbG9mg2CBcSiAqokeWX+V3iaFJt+gtWQSBFic5Qr3V
cSEkEZXlAE7AdpT8lMjNPtsWxVq0hpd6+wgdeLBy3QFQvuLrZ5nDu5Qk1pFP5lnHbcK1wjuuua+N
Z2/HmsNtA3hneOTZ1hu+HZ86WtwzlroVotZ46MWTlGy5vmdifkfw3jmgOkYhHsOBwQuTiNTBD8oa
8+P+jJcOPM2zWKSshL6rcuK8i5hQJz7f5tQQnCuK9mQ1zYbZS7H2ZG0wOwWwd8dpfKcPo6wpmjWD
hlukR83U5mGQuiH17KPMZDnggD7mukkbh/aeJLsc3yU2Xaq3pHzuIosHMOKuErN54wlFcT1Xe51L
YcpKrjzIIDS6puUcaniueBW4cml3mYrxeY3CO6XeEVmfFVUdV4x2UGS3eXLisU95/1UjjtpCpIF6
5ik7bVw7uLYsCsCI7kIT9rP8zv7Dp3/x9y28z3zbv2ofWXcnNSvSkUA3VUL8Ick/feRqWCwMatPJ
VdHBy5nlgCuwtxPEAc9Tr6pX/QTjVbZYVuWucX0cci8hynK96w2TtgU8Eg8px7qSYNzp8tf/baAv
KbURMR2r+aj+6FNa5+hp+N3hd2Y3hZ0NoXTvpKRcxXN/8Ui7IDVTYaUhEabydzbPbr/blJXDRGD3
721OXecx41m78wcUTd+8St+N53roc58JXYo7loPsHFrMW53uMiK7ZllBsIf5Fug0awDBDs5Twru3
guIXZmVT5JWFJZZcN6qlL6QTdo8ot0lmvQeQrHaBOlLZYFX5k30WSQzYRyVX8lrxOZC0OrwRARGY
MZPEM8YVPQssvsiRLSSwpINS7eziNKigVZeHxSzSftZgpvGnuenc5bllxUCuxjUXRmRE6EJTCxfR
M3/gzhPbXBXkldjTav2C65lUFblSYje4NZspxnntcLP+y2MBq9CtPxGZAgNPldcfIzQRLs+voT/5
lNhk2Mq5ou2Q5uFsgaWr2pYQdrb9UjppfTACc+wdfeE62lz+P5XB8LVTAqrOiMd9BH63OnUNSuWz
awax0qzb3UN3loZtqK+C68e76YCKYrAmdpVbg2DAig3PssIg8T5jbCZvW9oQN4RCnQNSK9qdwyfQ
WOk052WsF8+9yETyqVayVkOk2VABaygAtcnh0SEjcxRgmmjYWtT4FkFeJqxbMZUXkyrvViM/ce1w
mJzVAC4djthb48uQp20YDavCu7WdVhH8jQFzsB/DgLfED66QZMHpc52h8B2GmeWY1XAuSlJK810W
oQxeExMKLvTgeYqeryp315qLzCsYWIKEanevkTvC3A0bL8t+wQyqj6jA5yhnv7ogw7lZ6YvGNVeS
qXpGTao0gJL6qVAQS10rDeOzetnOQHjpCgPWgtDf2b8WbOUT3PXdaxUKTpO8UhWs/H31H+xc9sZ0
AEix9hFvGMqhhVs+PgIuEmg6EBYE3IX8ygN2HHJcHfUAyLUbO6/PrEzE/TS33hQN3npf35tSl/SK
36pMzPjL7DkWOepg8z41tUiXXdYOQxnKKZryNSnn6RFA5GaxMV/e8DUVa4zJsxG4sPawVEc1cq+3
QSYWcOeh/1VSIyzC1dwVbOp98BeQ3EQInK0Ajb8f0ZYIxr58TDxw33u13igIoIHJCiAqU0xtj6Jc
5rJszxD4YxW36LOYwv+N1z1xJRJg+gsSCNfkh1H5Nel3mPnKPpK3Q8fwPjMky+mvtXV4T+GPLq0R
nu7Lsvib1Fr88tf5oMSi+0l5lil46pFPHmKOhJCBxTrthXNez8zo2f//HDHLVNqnKTzwvUucacdl
wNM0fzYU7dXxz6GNqhIn25YXO391ZjExdQkKwV85Ha45tJwMwEI42ddDwSVo6qfKSsbpbCHZAUfs
8Ss0Y9MLGtqOIHSIo0f49Z3hFSNrcHnkl1PQK1am3mQAWbLgM20oCEYuUOw/BgfxtFEAgVhr6U8p
3AqVVIQ6yOPfe0Z9o5D5BvcC2Q29TRttnPs2PP7CNF1yaC6S6UEMKcsNSnYMhhdI25tPhZGW56eR
9fADPuVK6yeUkwNzeFjve9eN47enXCkCwc6sZA1XuFf0fXXOnxDizBFz5QwdZLoKgLePnL3CZm+a
eoFpklDI16dapP/BBq/U0GLcsCznU5EOVSfFO75fNKBQl0y+l2pzg1tyac7SHRxSXtboZkzFu4Y4
x+nkmV72piS7jXCRx0lmrmo5y3GmmtiH1zw8DWMfE7tw5e0qfFddAexN51ZlCZuixT0z6PRNWfYW
iS//3UWhTB30deygq3GcnULm2rZL8XxBIW3h3z7DaEA5QBseNigxXBUyO7rkdJ68oZHDaGbp61kW
yiC/E350zGZP61qrTxq9rYzY6PRbsrOm6rkANMnkIGqkWzEporzKX9i2W2TSRVARDFtHwAD+86x/
q0dXQWmOftEkLSzuDHH+Yf/4rpXGy+PSojvJ+w7YofysLX5HRUOOfM4Lu4Dmz3FimspcKZ+NmkTP
90mtPMoFNWmV4+lH6vHD4cRIbpGmY+4VMMnzwxZdMTpakM4SYqRBQ/LJqRQdSCxkSYeo1dz8TfhQ
FygKje5EV5kVg5m0aqlVYLnNhATBu6pyuxAx5A7F0b8o3SEkYimj0gUi/VU0R/5IdCGdrt1W9QwZ
LHz7nbVkkJdKeR9a0M9a+TfXVyFWOzq6WJgTMF/wfbU16kYGyPyY+b5xdqFrnige+1R2Ml3xI9kU
Ddk31NyiOMfJYgpsEvR5qbOpTCLvzk9lBgFMkoRY/AagVFirLsdiRIXKi1N2cY0sOFu9drrBs4VA
zyUjeXat9WdwmcPFVjZHIaB6IcNqdMT7hPrzunfmYvuSCpooLVVJ5tQYozjfUwcmI7/J+hyOGlvn
A//tfxUclCykJZhtl6TArxsaCHVzHKobQwV/3Df9WmXDQxQN1d6V6m3u3KX3WtYI74fRPPO6WJ6R
XOBbLWJR1kyWQ82s8Eph5WhSV2FtZZufGRR6jtuB36xysrhmrIqoDkO5xPBKjZThHwiIkmkIgskR
peePtLC4M2UBkoLj6z8jKNhd9/EgtE2Ojv0NAgdWYgCIaIb1VK+LM3CgQWDPUzE+gyIRvIp+tW+O
hFCzFQMNyJWfOILZZq9yB0fq6D5pbJLDRsWI45DvzN2/rFDJ63Tq3fk9zWBrWsNsO06Cbquvybpt
N9dWnHwHOLQ8foIzrAmWOcCUp6pERikfdlXLfRfgg7ChnW4XsHtrCF3uBtBlJriliPJfUmqk42hG
kFJFiWUkR6/w85PqOpl10EJ+cNbQEBRwkslvl7bqaQv1DC5hwQjreTWYhPwE15yoVIqrOxj4kHPC
5pqfYj93+FBkmtSKF5hDb1ORClq7oZHCd3Kn/QYPmnylyN0B6YV7cA2q7OivbSc4JGb0q3dGciIQ
aYNhxrez4P9UHvN4tYiQiL+Qadx14J0n+QVl9X33niO+kIiazwpVUE8iBgragJlbC2hJ3eqkLlO4
tn4jNh2OjPBNzgBB6XVJtiLAr2cWpXm8Wxx099CYWay/9Rf45o+gVb4eFJQPfHkP93tCG1Erdj1K
mgDNBHaUawZ+JUdUQKyJr62S+b7/NGCiiiyUUKesVBI9KLswARyPTK/Dx7EGzriZaKxKmvngpPwm
XALJasCePH6YRyi/8x3vdmte9uexLMMs0DrDZXbkAA7g0tJ6pC9oVqGiF7yqQ2KEo19XlYWKm+Lj
zqH5yPlmMk995L6q/LJduMnPoPO9IL2kbiFDto2S8KBKz/R4N5VDCQNvjPtxHWKIyTwb4kun6UeP
RXN1+VWNwl0pjnOGKG1JrXPsf7X1bCsQ85/K3H6Fvma/WPx8oonyW9pHefa8SH2wp1itHCwvWre8
QwGvDgOZabis8vE30bIk08dX/hK6Qv7I7sjBPbeY/98Ja2rYwZAIopMrRCvT/ttWVpbDMv2S4UvZ
6b7vmIcct/sxjDRTH527JwIQjFeoumbfisiS1fXh72uUqQZ8xsN6Qm1bJ5vfJPSZtYU5H/Q1pVJD
EydcSzyhEcVljn8IZczblE3yLra7vAOvDKx+VzjxLEDahhC294zedQjAATB61rQ5ivNkDaWP+JHh
vSW+LM7r0fDSlbFT1kA/HVfM6eOX2Pb2VCp7axvjLzWjbBj4I0qyLjlhnLcgACkRQsm6IQlip+NE
kb9dHhNN1ueRfXrlwrhok5daVz5OFbgpwXZbzRqQkPrxokK1qfNBeVvlJfW4vfz6QcrQDlw5G94P
naQnCT7k+L/amJ+puHlTIZUSdbsX70NdxfsSxPcTwvnpX3kon2Bf4ZS83Th46mejVrDJpSUTWMBK
t/p9g7dnCwNudvaeDYrhqkJsT6RR4GMFVhisK1sztmZT/6o6mbLftvwSqsY3j3ORZBOH73hMFrro
Gch5IjdUvLMWgNTWf+wCbjFEdahrJJv2N6N3xcUndGhvvx3DIA5qLDsvkvbvqo2YWVh2Xe1uVVsL
s6tYTSlH2fAsrNoT7ZYS5/vCVqMoFy1LV8NgfVKJboJThzzg5XAJx5tgQsCusk9NBCK+0q2sAur8
dA1YfWt7llkrWbFqp1xuLmaOyC6x8e1ZjztbhMJ5X4VUgUqOiVgtYTdzeAr2wVRI+LZs/IqCFgvj
/BmwJe6g3mfItleQnAcvNCkyf40PtU3DHRDRPNi/0AWnmp4+6R9jlltjg2dTXhhkMwWw/clIGNB/
g1C53m3I7p0V0RvVwq3I8AcFnf7yRtwdaS/06rTqF7PGJ7UeNI3GUWYQMRoriYZ1wu1jGzY7wWBs
WqMKMhA6fhv09EOSYTScJffzlHzPX2ZiIn5QKNTHAw4URYawL7BOq/cR0Ve1XuFbcCnsMXDgGI33
mRFYBtKKXapkIy3w/QSgFCDiKhfAM6Zpv/SdUoIp0Fc6HU4dAD/E/QYISMBm2ngFM9n4OE/O3N7/
2yZ2VtJWNDGYm0BcbhXCv6lMXlfjrItY835s2fWxYNc75mhjZmTg2kmuDIzOXUa10FOjB2ZnmDiA
KzfRZBy70Fg3lXMdfoo/yDPKpLLe+716Y5D821baC1j100kl0ep6jAQYur2YGBRj0btREO8+W8oj
lf35IYzD8lrLYUswMXm1KLxi/g7GSNz3g42SU54hR2F1XmaEIKlRuXiZF/PsYE0g/oyy4X1kVT2t
XpEI0IBY9Dkb9vfcCvRGOy6ungaNZfYVRxzqBvZy5Re8HCExT+A3sV1F1R3PNt8RnS2NOvP6ezG/
tH0ZEmaQpmtq17atzHlVOAtrWN5+c6hfzidnq8VzZTFYJUtAmI+PhmvLjDrnS29jopg8jJ6BUeRe
ltun0PIPkuew6y8av7cjRM1U5FqrmrUNxbCAi5225xpY2RAvSlXJcD2MezzVZCzHqOn1f3+mk3Uw
qu3a67AX/vPxus8Dvs7hRqjlfRxClZv4qyLKJ4zLFaOcnLJWea5IHJxWq3qJRMF5k3L/7fHs5T76
ErRkMt9IeHISu18t9TjojPwc7QyBjuVMEWOm/hOC/swG5LZKrx797QmRimaRzkoZp0OXn91Vvryg
xEk5VAaYOdfUNWl04dDIXMaMbEjdQK3LHdCcBojE9D/g7nHDUaGrS8eA1Iqd7BSXU8IvhaGkNq7t
9xlv6R1E0eoRhNP9MiY5bj6EpaDSPGUnYuPbXoE3zyZqncdns7H2ubDT3jljfpgEDcBTqmlt4wev
AuqoUXy8I+C+nl9O1rDWefBnajlNw6MAj5P/7MrHMCDemgNftrTVDO0ASk28asUHpuZANl93LrDk
a0AHkvcBlnWrOsel3g1vmKtyst+32ToPH8/El+Rs5Vo5gPAe1w01vgXBDuxvheXp31PBBG5xDBnb
667EJM8bEYAmGMnlFFPo3AdvAP5DLxSqWmINf9ZxLKS2AUP3UuQZt/4WvoWIKj3isQI02+nbr5aK
L1lPtoz4xpuitn10jwtOw0K1tBM2UIbiEKUYXPHhN3dAIdKG2SbZW0CcPTFv4Ll7nHhZOO5Mzpcl
+E/K4bko7ZpYBdnel5cYSJLSlG4qCX7lSNb+V+X47iXQIS/KpNIGN4P8pOG30WiOm2iEy4o9+aqu
V9/IZTFnNwPDCWnmlj9fMzttmN7TSK/LPFDctDHyfh7+f349B/zlLMlgfTFj21bzYhOA8RRnbu0V
i7KVx0rGrgy+tjuKvNw4VHgby/0QCsqnPRQ59t4oofNodfCT8NpxVARXUQGgAgwqRwykcvRXDV+4
EeoZno3Cp/m67rE11vTM5CM/mdXC0jFq8O6BB86QKeUTy5ovxXduH+CLzwSWfaNhcFlSmt2DfhNv
Lsbu1pQDTnfRC8mKvJH/JTbBO4HhLFcPItOya1iD/rGoMik7AX7mNW9haJBg4ZpHWmrZ4wDPikTu
v+Em5eLTzms1pZakuarq2nKMZXkxllsboHbVtC2IWu0g1Aoof5+Zb0AhNv+f+rBa5x622UBKyMez
RtVL6S85sfDNXDl369hdOqCFTz4B3WfU4UYA4BipqF7Mzrxb+UMQsRMrx94szLFk8CjZMFL0YC+8
5qrJ3E1xPlv4ZThbL9QNFpq9vfG/ec4mEq0onGb0SdbDG9q53vGYi+DvJCvqHPI50ASWd8T4Lrga
V9pCm4f1t+eiyJ8lGFBcghrydXaA8ejiLOET68y4AuEjoMPbFEPTo6BUcoZiJQfDVBenFMzMiP7N
vZNAC76Lb+WyyIAS0JW0BUFAr/fGOpzHb8Ib70fIx0lHNZKVCFE7YA0lC+fXeBwIpaCJSobeM8Cp
/iKyw8AyzMNXQHmaw2mfcdr+vTSUgpC+SFCSehlpe/MXez22bQQ+wzXtAuZssLqj4ZUzcp2MsaOU
lyrZWIOl8vt5N2iE8xbEYhQxVPXU8et4zBh7bboTo5aZ45OQNOYPf98rSBdzahJOua6IzG8uMJdY
WqJkE6NA3eMzuFXQJJOZogP0jMxq96D4i739IC4QyRj43wFhg+DMON0hUKr3E1HvEYpDK1RUvPYF
wfdU1iiUkWnivmhLDHzMoqm+LmuLXAPkaDOI6We0iPHTTGA/xwWfwyI0CHb1UvI+EaeuOc66qhZV
2IItWoSmKkzjVs9SqdKWglrASkxw3haQo9d2WUg9oY7vygQTCjuqTtAuxdWUwhCnxuokuPpYgXAN
nTbcyyjYocLvytetZiLUiN3J1MdO/TKZ0DTAaPIKXinoSjMfgjPRifc9K7Gt7TTxB8RtFvReUM0V
1DahS+cWDSur1w3+ORirvnNxR7irg0ecqaXJzf4GwPIYnaa9uTm15MfFltni0+QKMuoSEh8hTIei
sF4z7ujOdzu1dsqq6W/DcA6tiuSFvmD4O6dILKA2RuRygxs5xpk9nRS78abDA2X/523yv/Z3B+JN
KTM7NWPaAx2bY7f97/IIP7y/6f/30qBTEPWn7sLUKUTmlxFWAIHjWZ17Q913BN7aRwx9rfQk3wvr
RGWdlgdDOU8Of5rR7fddAGVls9RHEGje2DYRR1miBLjKbggrUozsj/4yHzoNk5XwtjVE0aeC0gIC
OOvl3TJ2VBLsgm+7xNrPwWwasyCdXMHggezqimEsQgldDtwIuZVHpE+lj3YoTEEQ/B7tgjggNFvu
RYCUOhOOwHuIpWEP5C+sv7vx7/NFNKC208RliboQJEXxvW0K5ecGuUL970HI1AD4JlMmmlyh2OIi
S5MnsWtD+tTxGBykOyHAuOz2du34r9zFXjW3ohCDGCAgNsdH5Lw6xyT+cck4K8SEdqQbO6UT6E8K
VtOK7fzVOnOl6KO6slO6U8Oerdh2kYp2oJfo+YUblO0rEsl/A98+bl1pMucoKqddZlNoJSrW0Aa7
tihhwBLwOOX0vaMNLJhDOFv2pZNPh0i/GupI5GrkIq/v/u6g2GKUNczyU3QAKmvfzrIC7Dkt3Rza
Q7YHs+hMmK9azORE8GhISh0CnjjeaU8Ha/fO9RpqzciwuNesr3O4oYj0BaB24yOPIoLwyapd5I9q
etQwc5bsCKo2QeenkHqemBEo8C2FcAZOihCHwJFyqtP9jy5gmbsdL9eajCyd1UJttXqAUwOkTxtJ
b7NeB5XLuKkn8s/7B24xWa85AXDJfQOpdYDy4qqm+wpNq1VGV7fSOwz7wITF/xUlF2t/BZ+tUoZr
1z7RSA5TyMsZQqwwYP8a1QODyHbCvGJt55YSIZkm+3UPS0PIgnJ3YbnIkX4yvRAagIjJEsMF6ysG
R8bW+8B36wV8/YWeroJ0VoOEQHH2IIuFe11PpUXIh536n/o/S0QWFOEN+jgoKFeePs9Flu4st+2J
c5csqdWWXTopHdBfHZoj5LGumuOx2dIXCYrE0rLDUYLs4t5tNM3KHWMcxEPl+YuxgmMKu03g39Qp
PaE+O0+kK7aKwvKmCYB0BNHVEQawdkcdtxajpulrVUKXgJYKhO2pd1naL2Heq7ze/tBKXuvMik4Q
OLRo47nApKoOO21eRdD8RmTSeGyCjDydjF33fnggziVyq3Fdfd464shZzYHIrdyMn38+WU2enrA2
w/szPnsLGmoERYo7DRsfvCpFgrmakgdrjwCNyz0TWG3yEAKqkDbt5JG7JpC4+32GXHg0wA5bm+UP
bBJ9SCXRoTP2ul8Qs2s5rJPcyeQ/7m7Dr85vfYh6chUGlQZwVwlMFD0ilgRaqgalaxtwf4E1V6ek
dcosfZnB9jVCf9XSX4XoyBAcgQq0+Z0nPMDyHmAKH+0ZiaJBBoTb8gfqSGdt21NQbiIxxCiyL1c+
wtHby0ulMFSIoQKbEBbwCGTpRz1+LNlk2k7oXp3zpifxO+891dWsu9z4ASjdm5N5RgsqEh2kCRh1
JWFSKhrNdgQtDg61ziAlgEP3t+bOzP/tyzmJdKFgOQeXEhj6Zc9JP1Zr20wP5RnNIrgj/+DJiwyI
hi/rdEcihB/iOxkkLmlqNs+k8QDZGyKrL94DbXNVunJ0csAX88vBaBPIqD/jUXNJ/T/vMxnOa8/a
FbSQwI8PjH3AiJQIj/h6hPZ351+VdDXVWXYgr1ynyx/ukf3oXOA47FMCb5kXECly2AWW2NSqpB70
oMr6HCIX7wZe5KbrnHqHqaRAtVRMVvAZlIXr/VoAbvMPvdQAhH2wfvM0HuyUmexMAwvNFNpK6L11
YE93wba4ROr8YZDFpteIRE7meHIllemL7fPenvOe1u2en2m1n8bB/pvAr08T5vncSp3dEr6uex2B
xHw+S7O7Y/LQgUerdPMXWQtZY3CLcd214AUozr8tNphNlDZd+pfHFRAJIJ00DPNg5xLXG3ukITqp
czHuvRhiv4vGXW+X5DJHyRpy+rOzmAEybIcMDAw+3vdG8Oe83IbP8th2QrN+K/ZSn92dWFEpMJJD
7gl4F4NVUY00OHrFiG0rSLk1n/YDtbqw+FriLJJ7E4GLHe+uEKMNsjhPIAsoyCeIsGGGuOL7PUim
BaEav7DweKZBa99AuLKgDolRwEAdt/f8Zh+PNVm7b3psEyhOhg3UWLd7zwUGczr9g2BZ7X4t9qij
q6KMMhrQaHpA1KZ1i0juo00Mey75vRYm41+XeKSW1TZSehzYbqvoGKA6Al5z5YpJyXsY7PZfEP06
X4ugccI3UOHSPBRDxBP/gNUDLS2KhlCLU4X+sIEWH1d/EO1c1elSL4FXx54ZbgwRs3ElmT4Kw0Lw
TMw+TD/BtZwrHd0Vd/xwEG/yO8nXl+QKUmLJLGjukOmZNtvhppmHt5Zczd/tjqaQ68z9o61H+gTs
FOILGmad9i2ohUEKswsOttLlq+Qa9qgFebFr6eMoMrOeE4ZnI5T9E7elOpqvML3BEdVUJnQ/g10u
zpiielyxOiTJWrLxJKYhk86a8T33HR4+DADVr5dl3XSN1cbCvW3ecLzEuzBW+CglJ7guaos1R24P
YgY6ayEJKrnBHCKJXF9T4MJogPsqF0/RDdx0X3oDObuOcYKLc3Q3hS2/o8TDRSFMJG0BBkG5khBg
XirvxTncN3q/FG9WJ4MzhjGfiA3ueBgkH4YAm1uPLIBxb6O3s4RM/B4K+HuTxr6KPznkHoTIB/KY
hcsHYQAKLhfzEY7Y6JfOyxdCaWryK7LrZsxj107TmtdPB71ra4XuQtlRNdaC3GLrIz8Rd6B8FkDJ
mBzluYi+7HeQ+Ve3kDjJJEJpe0uets8tpDa2tcrM10jU3oHr0lmf425HHtwLnxcOhz9fqmxW3L7s
L1LobL6ISVtT+sDIrE4UluWBo/N7+YNqGD7rCEM5FwbL+avN8OdX2su9QnMOroe0v+SI6cFBaPWd
OjhZ/HCWfHT+L54HezwGcOqqovtOcJjkNUKkdm+3rZDNIbuPKNc9lwXHHVRUNpxv96RARtrq8SLK
Ct4a5sxARHqet5ZBkG+LvXNl7TvOOFaWhHGR5jwUye1RklAFRpCWeSV2dxUCk+MAbh9Q4SL5EyOn
iUgbp3nSTu3MB3LI6Y2vUeyArnjRXlQ7QtSD0TtWBWvJ8OM3bvesHQekxuq9oA1uMcu0yZewvqEw
mRzC16M0pJ5H9CGUd3T4OEkhBTK+58yfEUCVaXdspnEonfpyQiktaPS7I0McnxmKh3aTt+qiotcO
WHNkjfzbWjrjKsp4VR3sw0TEWXGD4Jpq7p7QlRMF0VcpLMuh0ujd2av5loO8uqMlVsm8k4+Zyxfl
a0U5rHjZoQGG0WZZF/0Oku9rO1tW/tq1VM+OqXv3R2Lph0Ql//jXXt8GzCuwTeY8g51npzGXOsIL
i9pQf05bw29bMiVuhN2c9cO7lcU1xgrjL3JAfVRKIpNilDfIvTc/19sIvxX3T/uvQE8f/HZSmmnB
8JloZbx0l/P6ObNCnzj7xEFOkHZTVz4AEPFsIMb513Zof3dyzRbCBds6GqALNykrrYar11einyLL
bVuW/2exBdpXKM5HYbQQrNKXZPqoXsJuzc76KyZuMY0BJcNb4ZtfKGdR+wIUgA4NAvIVtfdjDD6P
Q9YXEe1tqes/RnoXrtJ7VYHINfRhLxgpreAB6ddUWVu0APnQcQprzyUiSOw9CnI6HleAoyUZtgc8
8R7q2eP5aaHIz+ZKbRqUaH6YOGAQbdh9IvC8lBu+jLFtMOXrbWRlITzNdA5KljwjxQU8r2nmHjol
1lzR9aAy96ioeLQHzycdcWcuh8t011KbraEmRydECp6mi7u5bSXZ61shQJW9miSQ9IfHCKugPy9H
c1zlz6J1TC9xCMbOuaQiJrzmNKZ+BOxYisJkGeL+4Ar3nWILqawDSUmhJk8BzHIMoAqLxEO1NPUA
dYq42yJ0fHtW8An0Dz7NX+JBR7exOcDqxOxpASi5H0hpWMx3IxkE7D1fqPoY7nCXeG7tbmjlDOLh
JG8SaHHGTNGtSORbj5wr/GObTIeKhlbeNbDmAKaVqVoBkUBR1QerRW/GT2SrWxi+PvdeNpu9s2Zb
aBRTQSU9e2JeS4jzbC9ezHuyjbsbfmI3t0vN4Pb23A0ZW+AmyPXbgTg4P4vNnOXBQnmMf8t01hBT
qVDgYu0FZjiI4hKskgIfZkB0SRZ/PCg7zEuHugRGTN7d9FlWYJxMgWnK2X14ApkYzJpHrnyyZinR
Usutcc4Lod+ep+6+arqBTJ0i3UWujO/t4IGe7BKGVtbp1OIpYlpQXX3L9OYFS7rucOqdxHbb70zw
nNwdislMIJX0KGDTSBupt36oMGyKUWSTY5h8vOOxo/IZv3V0ldFwte8TX1dbKu9gl0/j2oQvtfHB
Z0qxNd4BEPQ0fkft9uwEPY3etb4AyHmKxQqNBqdOqHZeYY0KtZ8f+nAzKsc1wNf4joh/B6y0l331
kDzO+aLMNmkKHN50qsBbzR4bnsNRqAhjq3TJDRwsp9y4IxBKSj9mp3N172kAckwHi0Ju2srUNvKS
RSUu+rDvjLlNClrhpqGjurdy5Qu0aKtkP4Wqx4eK7GLwHYI7i/K2aIGt2uS54gw3BSMYVAn0sbf5
VnA2+JDtvWSRsWcmdIt9XyEd/y0LuJpZyp6dhtkObDxMIH4tRuKAmk2YyGrs+MZuHG6fChpuyzob
E22yf2gsPDEqUV8fA38r8AV2k518OE/JS4gDqH4vHqICHax73QKB0Js5/bgfPrmzyJ7mxV13bEmL
Z8q4UbV0+QNWxB5AmU2spWLiEOOY87bEzrc8jkrsNdmJwVBmzzle8R0Xjw+sVXEc7cZVQO/Cp5cu
jD6UYvkV77ABWAUC/ChZKm3RHrkU0ka/veLH/PlmfsYQNuu6Thypw4f0leoQ91V5z8bv0oj7j46k
wc8uvbQR75+lu3nVRDBKGZ6UWey59xMD3AvXZKm+j9NMcXtTg9Lyueh5ELoqgv6TNQrQU/xeMm0p
3KWZO1GivrILIgunEZTKiPU6ldqUHI/bZnqidomCrDP4pUnxQ9YzpAWsgPoq3hsVR/Qtzw/pVACF
h454SmBOj98XaB5ZCE/4oqztjGYiJIyOoiTAyoSuErfHISw34hg7UBVrrnmDwdr7m7mrgHqAqTbZ
Udphxb59hn3N04x4FRgBRgxbcO163Lhsn8zvi6vLYHsjoYPpCNa+t5aMSwFpcLY+jteaj65GefUF
fjYgLlv6lD9GyFgUMAth6x4pWZyA+LB1edO2SuhJtpFXNPU+QMGIahByk3FFGJAMw8zIS8621c4u
jjDdZQqUR+Kw43XwXPENT/j4WmejvjacTml2muJJUM3BTAyGHxltO/wV1rB2uKOvWdpDXOsM6r5b
8L7fBLPyt96yAYWMS/YomVpG0B0U7GLciacSEYmfPQsylLg/WKfcdjb5M3slmuOg50Wp+iSrH5U+
FQ+EkOza8MEkRPkAxwWbAyhWMEB6FPHprxbpNgT84+Eakn5FZwDIF+rf7kcqDSRbDjyiRUAkpPmp
2CygmU2exa1Mu9F6PYUQj2oq2B39lJShUrZ3JeYU55PjN0dPqhFtUdMwI3afyCPIFQ0i1Pzeknjz
ILCeiYwOw41DuxVVgMpk3JGDGh3SC3+9k1eobCcKjJS+AUAuwA7vqTMz1VthoDD7pGXta7Osbi8x
eCnS6gH+LQlrjFx0d/SIpU75XvGUn5xyegoi33sBJZkEyD4Ob9IldP2Sw7FZ9G6x0WZpaCXG9acY
TitbBUqsf7r+3+v4dOpkpAwWQ8Vi3xYftKs7sBKUjgG+teTWbCeu/KrfaYEfvwa8m2SK5WE+cT/b
jMnEPwmtpuhTYz8XFMCSRPYiCJxjSwkjzTAGUy0W/cKMrMvhhp/+QnBDST2holE9g+QClG3JeRVP
YvzCkBURI8tOMylQbrNE22qcjqhbN+evWXkpNZjBEm6ZWZ+QrVflBWM0YmrSZ+0aKtY6Nc65HRn0
S9lMI++wenrIQjCqlYd9JBpxpEIK5Kf3LwbG4u3iau9fBh+TB/GQzW097FON1ZRxJHXEJzuuyqGg
dh3haAcR5GcurzODRUti4hh579mO6daHVQ/26pmV/qBkCITcqQd6e558o3SimJ5Z/g4ngt7Fd4fJ
KtY5/iOtK8QKsPgVaYRoAw4S0Yzl+CYI7DXkx5s3xmvJkXtDuOhTUBXVEcvdkO+2topPEZQv1DRp
GF8QhOSV+xMUAQG0oTJlUke0XjRqVsGWNlJDQWHt+k/HwF8Zca8UdrlGJVK9SBuwVu7PfPeqGoiF
HS61q2330qTot2Gld4rX4WC73yOk2s8YpcimLuPPn8ICRiyAcA5DepvpQweWtSWPznlj4wInQ58O
vWY08ycsRZTt+8oP/qsLiiu6X2ufUT4G/ypg8z7JWhYIzvnsIlx+fLpMATYs/5hUMZjyhr8taZTF
g1r6OMo/TU4lA5m01oL/HXCiST2awj1+3GBXks09QcVQYPNTzqWAlnu7cEV9W1YZ9pwnVq/r9w9Y
8CPhk475/K104lI6jG5ky5WkptVJ1SL6RJW4ZLJQDJzjumu316U2+GYJwfwuj5aLnMxdjbn4r02v
Ydq/CMcwY9RPZKPmI/Qmf0+w3EBKQYHypoTTWDAS84w+QujK76s/OLTnawvw0di5sUtcZj9I3XzF
cpo8KVta3zbiBJEK++Gaf/37P+wQydlrtQ+7z4W/BtxP1s09cCQks1yIR1/Z93XriK0lj+sO49y/
/MTygcjrJUccLuXxd5eKJzkb8WfPzKamQGN6z2PdvXPrp94wJOVVNDqOQY+dneak9TVy2dXBhWfE
L2Ukir+wgpk9c/Lb7D3gdELG0GRFLIMKD+la8Plqu6KsqH3ishL2Js2DRSao650mZfuYV4wDut+b
yIyHWoKtPMWu5W0yhT9KPu0sPbGeHxAh465clYznOeDU+vD4P70SEmRi0t7cPbJehw8VQ/iNSub0
fkeB06cbB3Vs3RS7+KhF9zTwH9NrqqkwO7rIJMVvbPpJd0ZXpjmnQFr2o2F8aoPC/1ghGpBd+JEQ
R1mxM6yyr99ZU2jTQmBHN+Ibd1O2XF6bdNCaABl9gqc3LGaEU0fO1WoAX7bqYlA7wrUYg12IqhpU
tUK3lohG0lnD9en36517/g3n7XntAoCvi+6sRWmaNWHtSFWEIfg+Pv4u9oB9LOqx/8RL8bu5wrHR
Tw4sqoloRAjy0mwJRtl53g2oMX50rww6kijyDJK3gO2YTfj254xVlvYdnqFio3AlLZzwVwfkD6zU
64UTkrL81/t+T+j79Dn943PMsuNkOwvVNi/mV02cmE6bHJlxuUZozpb14whxAOKESdMMxBMKZwSr
za+KZoSiLGlZaeDS0u7ODZW1DtH6V7TAntHjyuQP21CAjyD1OlUMuO0EmSuJhw++z8TbxdQbQs/Y
tzXDu3tC+1lwhml/UAd7gMQiBdAhbfvtEbqH3LgmdTUO93kDPaIebdv76K5jwIq49GV9CSHzeFmC
zBGr/PNhZ5f4jKLomb/xnhJmjBe3vVk5XcN3ANyzIJJHvmxiDRsrxaif3K6JFyPYJjxjJBjfz6Lh
ytjxwaPhh15L+9KzjYkWAXt5Dul0p7h0bNtQcRZOpaVpOT/eP7kF8xJ6GasU+2O7pZxYmiN+UsT2
5Sk7bpNy+ondUQ7SGujiTAN//roYEPcfOHk563sJ6P83yPCL1VuV7no2alTZyouV8i/b61LbVtTl
wmV197e9K7EJF4Ha9+CjvXwKaG+RNIhXZLxkIsqA2M2qMIXGP8rGBM5/ElgaA9+PzbQjWUDwXGqi
BxcK19O//QAtvybiqlxbN/327WzNMUhoLRXJHISKdef2ZmIpTkRG+yErS52XGb7XprLyl91PXEoD
CxN9vLdnG059EvxVII/pmGC0UAsgWFuTQseFJc82ZvBut/iqaiPqZ6el6/0Iql3Bn7nVggKgJP9W
q9qz4HzYkBwMYPhtoYgFgrDkIuh8GzP/iBsAOSn4zN89XBCIxBlONHD/cvpjNb5grVGYXr+BaIFp
6AWDa3xsihdR/zaQdbUKSTPPpqHpug+2HH8/XgShS1sD5guMpmjStrjzm7ww+d5eNeeqzUIap48P
2w1HhZDK0RY+jg0dpvEAW66CRcXfWdwRlIi/94qYUeIpxrxWjc4aQ1Io2m8hgrYi0p7qVRuVbaXY
lUTE90Pr2I6ubd/qcI3muc/mAHKfOfGf14qDwfS4QgjOlfc9PjLSSsHeipnCQCo17naDCaU5MeRw
WR8G090vAjcBKzsTlzRSC+m6gcwHQMl7q2gEKoTSVtwGpK7oNd4E6e+Ia3zMNOBNAHAC2wj4FVef
V/ASNYKJ5b4GTcmeDlD9FoaSAzFm09jkrX3bUQeDM9uTvtSBbiTc03VgCFT0YhvuAUQ/pF8WRR1y
odAOjKQjHSqhCcdqcR/rN1H/8I34f0TzNXMPHeniexGs+yksAZbfqf1FCQek8IB0alxoHmmWD3Do
Q9CB87DRL21Zgbbn4RmCZVN46bZhhAXPI9P32xPA5CAjRwoKYunCDA/HK/WMPx6JAR6kZIIZrjj+
G962fNme2Eofml0+Aw8vqEEkIeyfRLSC4nCASnJJDLwS4OnSgzSmN3JAiMr9IOJzXYVbP2nFkyRv
UzIy3h+AJuoOf84oKceE7v8He2juuVWGyn/X85+bSjDG8s6EIzzHM7Xx9h7yoyKz3FumxG4pk2S3
NJDvFjk9nv3ugOwQ8jPN8ttDUdhkvLjxrgiDgB2UHOWbiy8Ly8tqUJHioU6DbRS21pL+JLs9tW8L
XVKfDOovq4npGS7DREpZIaN8ZNOHmKn7SgUIMJtFcDZ94XeUMMeyEciGGo2zYgH/Us7SmBxRs3Hl
/3BqsQEHWXHHjiCN8FzN3n6dfVNY7jKfPJ1JZJ/QoOK4jspqXWGON0JyzfYOzf80UK7k6NG+bfny
NnbM8WCOMKuVXqyYqWS+qtOObAzYfMDg/+y7Rp8FRgZ2xp6L0dhinPgvoXTzgBLea+gEnW2hgmE2
WpCp8Ju2+yIGfxGv28MB2Q5jRhGDViiJjzllRHzvWr2q989AmGW5wKUIafcfHycOXKhPTrXJGwZX
n8ArlGkgUkXjUqwLOAU3MI9jAAWBKADh5Y6H0utc8poq1nviSi1NhjO825MjSCPU9Wx4voZK15tM
ebUuPTMYd/usCs+E202SSpzK4HKTD+X+9aS/23wKY/psRW1mvI4GmjlN+UbFxaiGZhEejz+HR2vf
4AP2oKVET5PybmYAfpc9nngdaJq69/1P8oBb9qgIY7NTtUF8rx5GFx4N3auBoNXdviqtcW5jnzWZ
fVOHbEwaZd+pDi72/HJ35ZZWBM+jHFNJ7BqnnRWmB1ykKRwbGYbJEBNS7P7zopiD6rMboeobtKtG
BCp10p9BBmEM6mlawfvRp8MGe8Ca8Wpj3/JL52wsNK3uaeq0yo/B/11Mzd3zRalv946EkMBQexOh
lXjBfwOs31c06DZG5s9Sr7/Ket8H24OyaDeph+mmXat4ik4dyLp8QEpY1s6GlwdHUvZL+BY2XE7w
8/6tkG5dl6VVoc+qr3/rOmei/QMZBCvCfO8Yjd/DWNNxICEtrCAa/6Lnns/bqPQiM6/6typcxf/R
jUME/ZpITOEKQTeoGFDIiQY1vkGQrU45nSJzgiqMhdYS6bU5Mq1P1ZPxW00JrgfUZ/l4wWuZjPjs
CVMLPEYH6qw+BIlH4WXCfW41c8CYRpgND8yJvRKEfmW9yaQm3MBH/N4CCQ/ITBW1nAcuqGzAvUA+
tEspWQnr8e9D/Jyn8za+OoM4b8stuYJobXAo2D9CCIBRlwMqQtm0LrcL3mz4pGunA7tmlo+2XPzM
Dcbt02IRE6piZLUvSfUE4ODbzMLdJ15nIDiNeGGDPUwSsmKcRwiyfFpmxSG1qET817FzJpsfc5Jz
n6zQCMNXT+kJTQroYs4fQO1GwE2sMitgv541wGYSg2OUCv1ebBSgumVZy2e/3z42dW5iH025pg+O
N08p50Zh8vt19FP93YWfPq0f/VIZHwxLQFaqXAAU5ijSeom17hwTIUntg0FUAeRLsTJMeGEIdr01
qTC4fvluVWuTnPmCcehE608Smmr9HmiPHu8NTxI9GDFgWaIfa3IUxeUslaxIOcs1/2bPPh0zMzqw
YP6nBlk7Cr+xHyexP20GFvi6sbbEwnEahWdzb2hcotHGRvhSlNQzPlR1hMC0pEQXzqU+C4NYS3JU
zXw6bk6QtbYlDqyuG0P3fhDhy10SLcP06XU7w3EbL8o68iGQjtmFccFbVociafF/0W39ZbQxYVjA
hdTb5NrqWCcIOCfqSmbDO7evcz6iYZ3U58cnqYdgECi2ATw6rBVtDOi4B1Nk3Bgc+/7P49XZ2jv2
M6vQ5+wuUPqyT5Dju43Wi3W0yb6kOgGhEj9V1xQwMBC9U6Lkhgbm/LnHdwXDB58aI+xspyi46ERA
ywgSnQONQHomVvQQ/huDYT6X7XuFPi2FXCn6fBiznxNCFE3yN0k7Fm6gAKtrfO4nDXmV3463lStw
BkuHxu0Env/7CSJ0qGSlCMhWPft/tf+xvw98OvsQaBYGwTBCtOYUVMyFDRehq8gXH9ef6a2er/X2
icNavpbpLz+TEJcTHg52gZK1H9NxwVCt+L+eMfrPqixPBt2ZJSjhCqWTG1rSQJXKqNcCJIhWZrQs
8bC5fjjyUR9ZgOZYzXq+k3VAyJSpdBcOEQloxR/nfpO6Ws6qgnnPbqVkeTBRAD9hANit9+wXm5it
1XGXRrpTydWmQGivBh9k6FHijBomq4kuMTGvnE9bRWprq1u7BaLmEWQwFGYLvkszJOJ7Fl/c6JkO
nMAY8ZFydVEG0VeQ3/P4/aRwxjHEoURlm8+7Q3U9DRV62Wcxn84vwfMjQzX0pE9Mfa/e7iYnXC3P
KtVg82YQWeYAYA/85AryO2kK1CBWC9fjtTUzTVNauWuG0rq/rrRSJ+qIn0t0IV2MBhXhFTbtI+sy
a8HnbivgbjdDd2waGGPQwUigF8fNtxE1dJdB6WSYKFJ9slMhI/x7pHXy+O5cqxJGePJ+bUKQn/+l
Oyp3H9O6MMGs8VElpekOae9uIwZ3DSe5DFxFFSwxvZCqhnp6OPgpEZ5+SgpGsDxQYH84ofcHYoKR
HoNNkEv75J+Q0pnE8E0QxNItj9tiJFH3eDAuLRIVAasOJwDkxanMeaqBVVoqqm3bFRzw901/sDAS
qWCQFdjvcKj2RVYFEvD2533wakrDtm4P2GH92VGvI1eRY0j70Q0oke5/+6c0sTeRCYrVbTU9pDE0
jEIPW0h5HSZxaTdPP5k3GusSjeNLe/FJhmVlmA0KKdnz6rs9wp4QuC8U8Iqw+b6dcdDU8h4G/y1L
d0CcN5Wvgbej4/EIruza+Qvea+rokhuZjta7ls6MyJiUwtQaMEgvwhzLoI2dMQKomDE/fEqC1UAD
9mhYIibnTovndOxmJMYUfhSxWFBaGXFMx/KjsvF11HNeKMABR3oxEdVtOs9GRuDRnLveoRAdVgA+
bBXO1it4h7j2m+kZRnAo/9N1FYNfsseySz6DFiqlurJDBwas1NcFkrrCfeoxEoGHdLj+c18nxII0
UPMlj9I5sglamNjAqlkgc28EPkQjsuiKU2JUGtyC7Q0M+/VAeZgPcLvQMpktC8E1Y2uWmQqVQcjP
3qudBzFRpO2QqCbTQbsig1BPwlSxcvWgJcGehgF1jbt4uQsrOVfLoM2+XZc1YKSO9d36n5Aousoo
iWeRXnXmDFCnxTcu1whF3vaNkkxCdksdzCsq1ErdvXf+E8/Ft4CYWRIpqEl07KMC47v79aF2Xjss
s0sLYuDChjiycer4EKnNdSsEau6zvMdYi7cMEowztjmbpdzR8e8xtrQQMzyCHLcvbPx70iddqcay
V6Z9qyaaYo2mY0x1pGA/VChHh10FFWFCC/lnhi2e4M9fez28Yeg5OfJ9CqPFgjAIP/EjxVqvj/53
QrmEXDaHtkaO23RRiLkGd7aLd4qWdNN5zM4ypIGrrR7IOVFdrjyJliiWG35aEC7KE1pUVlsPdXH8
1l8E9YVI2z6Oy6LnGUfX7B3XMGm2ZKKdtunipPXD+yLRJIRJiJ1N4Er94AMplti6VFzkBuurs1ei
gLJBglSe8eCuloouC+3TVjYXdhZZ11fbXSUGCdnIXpLE601TUYrKgrjODzYPZLdBPv6l29Iv0M6B
TKrtDUBtEFLrRjGvdlCqCeDmG5B7uD8r7k85aoa7ENhWYXSEJ8hx+PZPpiY/GQ0ChfSmJ5lc9Swn
0cj/szMc4K2tk8d+kc2SZ711kxioVIAjBTB8ZGrhlBqtU88BkNn1a4CAZpQ7VeE25r8Yb3j6PVgB
xNVt0SL6WSiJdCPKvVYgE/HzgN/3xqC7Ja29CTChBHqa8zWhitgG9+E0CceWBQF3Q5RyopZ+IBKI
W6NKc1gqwaaXqJSz1JVmx9VgsFCKTJrm2NjFpicDSRvW6AD3y6NseiGdNE4ibPTINPkVRBtesjgb
IxEigHxUkJeEToeqRKk247E99ejjJEteLMhx6SqWMn3EzHKFJATnULGNkCIkkkR7iJcMJjQCGzu6
KxRVYW62iLwBkMjIYWOJxRef0gK4pLpfc5WPMpnicncvLjf8d1m+C2pimmOmHCD/duDrKke9bt1w
qjwotlHL13AFziA5OrquRfY1q8zNW40N4jETB8U4gdNRlj81wJOuLtpj7opCXlkkCPU2HUnVJbeU
5DMyC2277V019iH/TgTpsTyCHYhw2gMgIRMW9U7McAxgIQO2/3Clm8xut4WG5/yRZ/oZtFn04+lk
8OVOWU5KF93BXlABPX30A0DpQVkW8aQRk10+vtxcMMY0ycZVKvdRAg7n1DR8ccAo2Q7A6NQT955n
YzONoE4F0j6NA9ai5t6IZh27oldzhgJPyaFe5pSmcjZA4LYieH++QghWN+l+itr5Z+i6akwP7yke
hnxHEKtnN48Vvy7ZNf97sYiribdfezyV54h7TmgMX/+D9GWXaA09DfV+LF68haywKL9EYgmPekTX
zmkSnpmEj4As21U1QP4Dkcd6B9Ccle+6j4vveY/rettMbSjm+Hw03HGSMC6Ee8aHhqeF+uk4MOCI
wSM+ouMH0F49sC7vSI4iViHP8E8Ah1e5WwR6XOhAEGlcnY8ftSfMk/anly08S8fnzwHlLQlRDneT
eiI/ELo8kQHd+sCMavPmuWMNGaOcMJrb3X2QNK8D24XiC4RlOrYyJ387yjS3zTijxaBi3K5sJHK0
d96HkvaFwyCjnanusc50pknWsN2EolifTALG/8WUfkZCw5VcuMr5KNaYtwJvBiYl2gBPMaWTbqyF
0ce9ojb6LMuUYtA6N+qiE0UzMbhlLIXYXVAorR5Bmm3vn8E7wWQUlCuJlYt2SEwP2CjqSquEo8Yw
vj3keD80GoOZcopJxfGNB4WWwrxpnz7wYxD/9ExrXQVX054JkHJJq0LonwxXP7pc7CPfCxhdKdzD
RwNb95ZtBQ663bTMlYLzojUfPxSOec95ON4ihZqZoHrbsaYlZOyc4KLzIDtsObGjn1nyijEl2oSl
3w/DnEvy2JUb+2NBgvcrdn7SY/DlVGjcsB9fbaNHVoRfbk2IDk6H1uynmzpwoBf9gjWtEWBDJMwl
r7RdFZ3kf91VmVtBG9+wPlF6FBFTXa+ItVZ9tG8mAHDeE6P2xgmyau674gjjSBfwX3ImHu5vRpfl
YeEeX6+h1PA1Yp5+zCOarrUAihvOQHclL4gbq+AnYxTzJQwLkmfSwSb3+meQ9ktZJs4yULNDlBrB
/1Y2cr4o3KlR1SP5XMT0pI9tiLiGpf7RfOkhgTuB77GtNry/XyeBC53xZm/XtpeIIAInBREfE4rF
MiJHnLoDjKFJ9JlkwUBUEjpKbdtNr/yJq0TjakmMnwnrgp5KsBA+J6raOUGby1kheBz+G0h2rdpD
S+X6cxubmd257zFBiN4uHhvbd0YfIGUN4CtZduAWzAvttBFGWh0TNMraBIfjH5KZ828FTSzhnTlk
ULND4reyXFc1UcsmVwXmHuX0VAp5gHmS5RrZjs3Svstq1dHAv+cbAoLYh97ivEegKFYwmyMHhibA
GfCUT/VJSR1sNCFaCnuT+PKrmZXBUqlJxe8x4rZKMU9aNdJAY+wbLS8or0JQQ703xMQxRbvgldzw
o9emcn0PI/yqdB2a3QrvQ2tjn4hKGNZ11J9B5VHbQFTuhON430hA0brreitdQ0w0AVLJnozbzzjb
w1v2zdoFMre1xWlUOFJ4eoWZbQJCeG2MaVYW+iYo+G8O+eiMIxFODR5JaTEu5j7C3Y21Bv3csxnc
jk0jVXihotz5cRU0imPtHIFnQEuxzH6KfatFNplBgoww2pkpPLDiXS1k1NYkyrPAGjQ4edjX+RS6
cSsyOLNLvii1bVmNRriJDDpFUYRYtIssXkM5FStIWwMcRs70HSSXT1bMB7CB9kms0r5Z3Ufj5Hww
W0y7VPpNA0I5EMtavYQmMcGMXHCa3mPcO/F9T9IYLfpdld7m7mt98ktSLeqxSMTBVE6nPKPQ82ZU
EmiWVw6Cyy+EjAz/DAIHAC6gza5Qkp7J7elBLKsLOznQyU00tNFciDH11aY+1Qqi/wfcaDy4iHMH
Liy2nfH5yy/FGRAEK6+jAYFWz/mCAQtGIHe0KiUApzETF9xr+gHC/O/9VrXQ56dvuWTAE+TgqjU9
03kB2s84IQizF7GWA5RT+q+12cpNxn0n9a+SX2lCAniSz3mSKl1otol5VpPrdHcG4cn6GnANXlao
yw0EL/hvUL4POgWsfNftjfOPKwhFeg2kgGgDVdUF9Pek0BJJPAON+ahQoOrVGmTpTnQaE0DaVi2R
uZC6LWv0X8hnOjFxDoUrat6GA79NAIE6eB013L/865GbYi9Z6MgE5lSZhfVy8HxYnGw50RXlcKTw
c6wisq9xPZT0EVxOu/232AsvteGzBQnckPVfWA7MxkjJCS1lfQ14XrHH7+0hOcR9+IzWNF2Kkebx
NYfmNoQ1YvgWN+SZTxtbIqvUYoW5mU4tYfq2xpWIoe9vJZ+F7S9My2tMXIUuJ6jiw3+1dDG7bfdp
eP5LeVtlz9XPahOw4MaQQKnqZs5uQziISjBx7xcC36q0LXbx5dGXHC+FpO/mHdNFrT/Ks6hZcdYS
Vm9nfRXxJNc62oDyqll6S5ndZlMQAaUUVtHlzlIqQdtZCL3sy2nC5IdPKUwBL51N9OqFLrBN1mCU
1sThrLKCcpcV823JceI/aUH27lOYgEVBz3Rp3shgijULNtM6kNp87X+qlSrM2hqb36Ke5gwf4EGK
Y3AM8/9/Tb/AiuHeP9uOJb8xv6kV/P2TwEb8EjVWJj0FMc8o7PHdIeZQhyAaZUlLxsPEi5lfgGGj
sAqGdKctNZt3xWan68L6ejnTtPwgHyKIMo+E+Gzif6lMaBZNg8FAzg59274GkcKKhGwI0o9Gf7xV
m2Y0B5FrzhCLQqQOKK2Q22KAkn4znQLBK6eFe9JTsaFF4ahyW8PvqtoJ976t6/t8XJN3yDR4yXsm
7hR6SYNwww5Y8yBtfTvJGZyVLRZSptyLWt2yoy7Y901IxEFzIF6u9Kcm5S5z0uwyVaqysDOiwFr3
E6huLQbEVrjlOebABVYNrqA7RrGpyfVWsMAIPZfadOl9Nzo+i40CbM0vTe5e+Te1UWscAhUXfOMt
eVw5qUHVmb1D6glPgIg8gPGAHbzB8pP+TfxN81gy8hvhApMOsyRkUhmWfmhMxkW1gfUWlZwply7c
kdwPmBoJdQUI4iPou8fembojN6qkPzDZTnHI9AszDv2LQn7ImND82jRkDwDZCxBe/D+kMrsjERKE
aiCv/x7W1qhatckd/fbOqbJvZkJiSCPMnAdoMCzTkNsC6wque5dF+etaCoMEdR0zozVLTBWCmdqC
lAZ+/mDr3uvXC1e0ni2f/SsMGZy/9U2/2AUQ2TZ/1RLV/WAI1cBMQ0MTMjtQqmf5eRdWnJw1L25z
OZbN0SbWAg1f9QTAmuZ3Uu/o2PUiiz42X5riz351tOo3BZ8p1vk7ePMwHq7XK2wSZNoahnAWa3Nh
8AILXxWoS86kK5Hj4HZFLf+JLUwKGXw3JP1dd/t97N5ld3Mo4zIJmcZeJn8W/proMO0g/xCLsWrL
V80RYQOsfddQnSHpeVVZny70G2HV2jy+bUOLDvffu4v/OnodPPv5QwRAQUu0F0aUwTXtjKHHtK1f
85tD4HdSlFDGHb0YVI5nu+OYCyEz8bN5bd0VqoCfunsn5XJrKidu3p4yt7kKRlvx65cXbR0oU/8w
L9/go1kxUo019Uy+ZFDPk56+jNIS94QVlurUELDGwhbECSmyIZuUGIdQ59jo/qhXvrmaM/C/i1wq
zymeuYGyxnwqI3bwObllQhwd0C8x5L9qiMT5Uz4JJJUPYFPdBEycsJKJ/9erWuVr5ZNLO/JmVsd/
G+HqW9e+tBYJiIqHKMDa83EiZv4x8035VwG+nyXptKtANm2ejTr05IrzHHnR4mAovS9uDR27cb6U
h2QNvG/3B/8+nrwXITyKgFrz3PJphXiHaJQL4BmtxmXi5NVgICXwFAQVHjSiAgIQvyHE4NdbMerL
ICOfDVtwgtn7iPjBCKAMb7UkI4YWLYsHrSh/05lMmKFZi91Xo12iCx45Kqu6Wyj97ESsIsa9keza
ZXqvzzRarDxljOktyFBDHVu3tZFn0AUdeaJdgiAbfNuibqrJy0PISVp0l7boa+b9mrpEPY125zS/
v9ImqISQeE2nfAKiziclsLMFhzloQgfp6QTJ81+kn3/XojgY/QVM5UkRBwauAGun+h4kr5G/n7Eb
KqolpO18/YkVIjibH0iHPKLrZi367aU+QEicPw0cF1nOkhRq8B1FvPgWY/jMwDpkfx2hHlHFclpm
8hCd1AIutCP46wCMap9zbPF6tK7wGSmINix80FgD0vBjE3O3NoOAW0nirXsEn/oWwjwETjCLKaqk
bTz/dV6od8dnsve3ZukXM18NUirm5wGLKkLnMgA15/D12hOdJg+m/3hTxF3H2Ti+P8G9KROk031q
3MpjKw3CWJ6twlzzvzsybp0+5TSGaarx/fwX2t4LdeIGxoVPziY1bEESlNXP/y7m1d+CXIn1lGIw
JGTJoH40YwcTCldiFXLt2oviCbvmqD9q0q4sXYukFaaNdiIcUXmmgimSBD8OYJWVC7Q42ljbFSeA
jRQbDkhGojRFnsS66kuXKS+a+VGaKlRt+u6W8LPVpOKlXEIyty9icyw2q6CIn90HpF3xsM3ehDqW
36w0Swf4vesN1H2BeT3/5j9/vNi2gR6MbpvMTarEhbNjdzZip5jKGVItVjAFU+iXdt4YkQNGKaxN
IvirlRLlC2K1L0ePEDgJvd5KuyfmDwg4uDbr9TLpU978rE6ZFiUjOTlISkbl0wI67JF8v4AP+kWo
6XJ6IXAZwruVkf3e555UL/l7NpumflSyc8UpoFtcBw0vnY3AgGeOO51pdhtqAQTNH4FLvWDYP+8q
zMgIPpvew8/jAqrPvGFgYRZegxH3YoiF/87sattF0XqRh6MaoNHdcy9F4YzzU6mp8TMzTeDuDGj0
71RyStIJXx8/yppcsnUH5xYnX48PqnSYZAZlT+TMWS2kNhFEkaTfWNjTW9iU7Zh9HQenNhQWU4Au
OEyWnhN+3ZpXJPQvB+llkfonS8l/RaNaQXzpF7nVikpRGJDXUIumuj3dM9LbFUEe4R6Ymj3QOviG
w2pQn8eN9M4/ve5pplqYq8rL8pQZJxpR+TAwSBnGfoOzjTccugBMta43frHiUbunUlHOqT10b65M
7wiYtYGsj99jtNV8KhO0+RNqShU5mSitvz0MGm/4SEziNae+AxrJ2S4T3fkU0Dj5vj+iDKDht7Oy
/TFUdZokYjX8UGH1l1vqpkl7Wyc6/fMXyTsW2Vegz7wGz5qWjFN2nb3GLRbvtaB9ZPLdwqU++Zlf
TacuoL2sIO7NhzBzI4ELLefaT1KUCEqqmnqZMBYDlHpbrUOqSqrln70YhYBbyPCn1oU/RFmx5/Nh
zdNm/9hlsCSCLPqRXx7GtxbFg2WJio4THE4dzn1huEEAZ0BxmzG8oTsE05GWhLqbK6oEpcvU32ZE
5MNxx/TnPuK/WxEJKfr6tABxoeKG4TaKu4WJ0UB8XbuTZX3Kx/GMP6Vl9JQeYeMktt9XYy9RJ+uV
RCMl89QqdUqod/E7LiwodaGW8VVDIK3WBkBE2gu/M34N84TmJ6Cr1aHP3yKttvuYVz4MwKdxadgS
iWPPuwQIvunPqMPAlYQBheOjePEY8FWHc5o0A5rDveTml3tq662el7/hYkz9JoiVllRVoCuqR6aO
D3FRXUop0Un/X81a9CUAXL8vOrOHS+QJc33jy1vabPkdPotD9zHXUiY7oQUjSX2n9QjOi33vFVlR
H0SWdfq0Y1wdjdD+BPJSG1L4oM/JaOhWcobjMj6Aa0akqqTo94Nbzp4UE0b5arSKTJ5KszKhw6Z5
U5Xot5JYp6GdbZp86mHmlgzR9QEGXJlmRLg0NGGcV1w0+3dAaNXnKn7mpvK5KPWfaVJBRT9HYKEF
qnYf5EG+9kcfNeAvxAjMO15qiAP50X0QIJ8TvCPIdGZGXjtaqBQUEZONOGfUMyFc/u9VLcNQxaBD
CyfzoxDsrn/szd7AKbs4VtaSfGrdjR+6fom1A7bqWRDCGgmPXwJX5Lq3Kpnm0DywqBZw2RGBT17F
jtcZz0Vq8cUI66SrPQNMlbkI8/uoT9EOtcu8LXhb6Td0Txv4vMyJ9YNs9nIlD1OA/wxDZJawwfk0
Xv0DF75g6NYYw26QNPDXJKzRFTbygY4URQgn243fZfgnlgTXEg1w2CCwqwH4mC4Ylrf8UpZlkd96
qePn35qa9QfGD7c1EOTC8rldBNVquyLo8o+DtLp2b3dUAoMJ6Ae8mIbNft0GpVFYwVgXqaZIFiJv
3ta2C61aahYN32kfFOuibVtMLy9wpgXZQNj86VqsesngDLg8we1gQd/eTL0Ey6buHf3I9IdMqc2k
tXUt/Mnmg5caKvkvib2oUQBX/Srjk3JUelkEkOqvEAv5cluHnwQ0qPCkeMll4f8G1tSujSnfrlTd
gws9sdh9YSlp2dAypPsEvSvdm/op0EDW/azJ8t0Aj3uB/MttzMMZbnLiXGXQHSl1uKURJsvPf9bm
xVttlSOuXj0MiH8Hwvn6tjSn1DL2QCkLi6enlW/ROxx8fl/cdjOVhlUQFALJv57/HEFBPaz2ax1E
JZsZQ28bomgeP9qGpKRUPw+QbZlqk/ZPoV38e2n8rFEo1iyEI42V19PwfERyUUhxZUQ02UgbDRKA
edwmoYIutS6Mu7KYDF1RYi9F5PN9yQ+PumTMoHjRyNUCa0uM+YMKTfg7WespDDimFFZ1xyerXWbD
0bAt4sP/AKBUvCJhPGtyvzeOD8x3HQAEzdUB1lFvsMqAfsnxs0hO+AS5asxM6UE3rFSspaDcGnsF
yRXyFrjrIV1UQOKQ7A+jyWwDLpyQEsxAdJd+Peo7EGSoHL9xOGSndfEfyCoQyfK4YaiiVhF8H1tc
bZraZlF69F7wlqcnme14tSSx0hOzGAF20YeF6fWuCL581d1Wg3FU6reLQUHknOltX2ER2oADjYvt
bRtKW11WaKS9w1tngwe+3ocVCfIkDlBe6m0P7PgvvI2VvonJyy9/WoPY9pcgmD1hUHpSM63Hn90p
o24L6xHtD168J2srCBDPElWAvP06Z4zOVG5GGiUcC+/pYhSnXPev6jDaX1/HyoDIiV7P4ey3Nld2
ZfpSrFXtEAW9uXAOQ0xXlnCABihsc/Kccz0xWiFKWEUMZBin6ZJDzi4ngCtlK7dBYTUl6Zxkea1O
GQJuxG/QzvV5YySBbR6fSkXpK1XZflPL4DaGTb/A/ceY3l53lUPna/J6+nIjpBuoFau+WyfZZJhH
2cMZBhj0ok5tIhWRxE48xZQMdIJWwI033x+wS/XQbTjp/fpapR8eirodqRraW8nbbITw6dz1pwax
oHZbrtZpCOOy+n+N8ShnxcUqrBnmzEyas+CoflGiiBY5Xo36f7Ys0/bn5EzrvLRYj0ktXxlAjj7n
2NdEG/tFwUxR6w+WvuwB95jJ1M/2IJzJjBv2Dk8V6aHqMaade6StPsGsAMNOMiwoHBKujd+hS4oY
P3EAOgTQ+TjFWHxw3l5XJDBrA25xMShDxg+19Bk8og8HpBmZYrxbQT/QwzOva6NHKmhfbYSunCin
MM5vVfZtm4wZsMRS8b4GsUeBr5u1JGjs0gYpq1e2FQcWTV7pM0ywTtDBkJRWCPNFaBUkJyFcFnA5
VEJQ1EiLBTfs2HhMMS0MGOEGauWAg0wIbNbeaBEyD/D2p+uVBjHVk2a+n3bvxcQwkg7liVMb4GYp
sQ9Ung777GzwBBJL8l9pEasbgr0fDcGA3F50aVVI1jCDgIgD0YYaf0QolD+N4MJr1Z/uI4hVXJT2
o2E7/MDWxrzDFKIiamltPooowuKI/wEIgIK9Kjj5UTra/SqEFVK4F8pO6hUNkPrGB5dCGS7yGJVo
0a64gaPUlAC81qnJ394VwlRwEIhvSmCHmMLbz5LEzU77DaqqJmQk0VbFOaB1ft+1ilVBszM+SjAM
i2T8DVaypAy8au3G8d8AwzcRYoIfrTLWsoZXuC8DKaRZdwP5L6n3bdZne+qG96Uy8tft0vWxIqnf
o4+AQ2U+TJLTZY/l4XhRJMwa01t862ga7mLbL1CjNtYnuYfgpH+oRhxemu7tH1IZ/iblsNCqR/We
9I5cyR8tL2V+gYHjXMyAIJAa7oGvu0C7rUJLpuB0VqdH4NTpdMGAK3PoSOqP2qt+W/NaF74LOQgt
FOQsWzs4pn1kCul9dx0WtnjIsXo/mKfmzGyY+GzYfFJzMxjnzqkatDYkpDAyZ+1tM4jOKgqDfjeN
ZxIHN25GnqOOabY63Xttac7bFrAjfZEcOZJAFP//wgQYz/2w4KH8I7Yv0xDtTT0wD434t2yNFJFz
AWFA+47bp1oN9l2oEpYXdguNtr4oYBkk97ZcpvvM/fxDV3HV9fKOPRbjXKF7TG+bzsK68yP2fmRG
yXNHSKNeX05E3UmL+vWQZR14RsuVkwZfiWQplc7m7EUe0Vg2KJBl6LZNTDTuFzjnqN9AknA4zIDj
zZTgojXYQG1TF9cMxLbsUFO3hUoOFzbssCalnUajNxgH0XJVVBMWOmWe4UzMhEMFEdRnoHpI2zTk
CnOcmT0vHQn83SaRlIo7/0eTzGp31TveoMtYL3XGzXqJfuwA7JiKmKV9McvRhsv88A7l7MNtOJQ7
VZnAYV733DMabr3RhI7Cd/em2pvneLG/7lr5XLGeL5Yfw7Bas3iykinCKTZxpVcL3ztz42C183Gr
kNzA20WZWQ21YL11cZgIi3t0IlSLoyKRPOCNDeijDEdziT8gv4VZRrVfNv3KDjoBRGNEK1OlrqWs
f0mgT1XnZZa3RdZ53yhsp8r5Lft2z6RxepibnDHKRQJV7mgpkLVrKKX7QKdFEyP4EhUjTPOnjnJ1
rJJQQEavptq+e68b0hg0kTlPuzdxozXZIgFocgMaevcr7YTplPGMkI2uR/fq0FSa4Xq0TMuXTpoE
H4aOdGngfKNZZIivzN7ex+0pXUGcG6L5vWXr55v1jRBdsNbq6EhfeDB4s76XfBRG8FdhwYwJOAoc
XRuNr6fMn02QjdPAUlmcNNsSCIAQ+o8Bclyu9FG6JHss5FV1B/5/U523ueHqIJjyguJN6ilFTyhr
Ng2WrNwMovreW9a6V2OtpFHgAnG9ik2DvIKglOf6s/vxKI59V/MJX5/HgSbcgPj1uMGRRORmI9Xo
1RAZYJLJC5gwTD8pVTDjGYdZ6NM2xCqXsPp1Q3Y/HDK46t0qhMAM1e3sEXHIYk3WLGEAqLG3dl1k
fl5IHk9Ye67rLHu5+Zk89sIiwuFgxyuhAVVepQFywCojbobD888TPGnhoiS9OKuyqAIy56axiOjH
Ad6ZKMN58+4YS3wqB49sxmm7SV1ykuEa5yd/AOjcOzed8nfil7O/mRNss2zZK1K9wKZAP8J0ifBn
bX8//ncvrxs3OZ0CmJiDVrqoSoDf7HetGNbT4KGNBxSHr2cexTjL5m5AfFh7o/H/D5d1DgK6pSOp
ixUzf3x8QpgctKzkolexo+8zVgD3ITUWH0nyZkSy6okVtKnlENt5p2MpId2ZgADRbaeF8u77cRMl
wHB92Q2s+rO0pMY3z52zI1xxHoSpfGmCM/u3ebAjwNAQJJJnJpL1qux/NufRI7S7HAn0fa+QLZTw
fYO2dQHVqG5sxoqrQebA13NPYmCfequrHIwy7KJfWYPMBue+78k3cecdf2qG3rxSwwLVC3XS0oRk
T8aZZGSeZgzuw4iglKdvMqMaY5kAPBuyIEMqmwsxLb3Dj6SRePaT3RkaEedVMvV+FNAO/LCYoWfe
sG73CVnv54fF1TrmoqSPJCsILpg2j0qiFE6Ox962Jp/chgulHGJtgxAvoaQCk1sQ56eadXnxoNj0
uwpCwjeF4LtJuvegAbexqv4gEwbs4BNQZMTWmsZm01tuF1iIcFeU6yUuZaOV6Dhgq4z8CPDk4Uw1
XUURWulFfkKrrZ9PaZbj26fOYKvBBbg2YAmDx9qxMuMrlquW+FZnfl+p7Y/k2aCETxJo6wVhledG
zjl7TADlbqdeU5O/D6lDInNnM+sgeXahJKoQu7842FTVQO5gJC3hfY0e7nmJ8XIP1B0FcQQ2gn8u
dkT4B+jDZLqragotTIP8j6+SqkqAzeO78627YVDVrIZMMcMaSUXYgs40Qa7f8IDmlcDQgTzBqIvV
LCJdbF3pO8AGCOTyI0A88XgHRjkIapYCkg4hWzDrk9tj+WOzv6PN/q1VZvaJzU2+wXfeqHoiIQ4n
XFi4+5IGcROD5SGXZPth9NH5o0WPsx4JfSPjH87R5qM98y8KotPqN9xuFV4VUJGrqnjoAjI51c96
Gz4G3ApxSCHaBT0uuwKCwLwF5q1i9MhPVys12lKR4S8MOyHdbhzfhgQ+NV9VeqgwkDgwoof7yvUJ
wGwZmIXGfy0Yq8xmcSupHVr8Z08ZxO+9ciP4z6fIjnL+wcwmnubmzY4zHIOi8Tytvo5dNRPM0BtR
gnWCV2NMxzQoqzB28GiuVXHryJ7QqDpWUT+YjTMMKZOd/bIdKG2/c9UVtKBxCndsK8bMEyZ/HjDO
lNzQPWq7I0LVonFeeREUNhnUPu5Ry3I8p87pRpvPZJH3vxqiJmQc8yyDhxp6wdIxK6JxCx4u27dZ
m+10rglw+s+/sRExg+D6ZZ1KsCOnGIeATGkUJgTTa1lw0IDbLKOxYLHEqLnL7O7ANEnmhqOzA6+M
UHRC6flA1c9gBrNtjOLe9NCrnfJrnwhqhRXXQotObM9Qs5PIhOIcW/Hm0lRjuyHy6qPohoW/8ume
VWaEkPOl2pMTn6HO0u6HkxLSvrHFSiH+tB7ZI8QDKB+e2G0EhxvQ7H43tgJCe++7XuCq9KPhJyWb
9kd4VaiV1WDs0okgn2Wd8JUFfyxo1+ayo2aMrQ9zY86NTahk5G4rimAo6tQroBi05+epCfDj0VSW
OXHzi9z1npdEYi6lNY3odzGYFwtMEDLMO1GtGtgRpYJaYxzgAgk1JLd9f2rod9+Qb4CjqOQ2Blzp
H5mwDU7q4D8pJpzL7pWsg5syjU7aUCvssgtjP0NzQtHsk/VQOYLFdB0lNS0gSPrxdnbNUMhD19r/
0z5MVbztbyNnqu2Hqm3g2dER0lv1kk8KOkKkgFHvmBcB7vHMBSjX/TTa2VLtUwA+kD3IEDqkkMMq
4g/x8A+o2kyLUSVfWvGUwd/Kjdtu+DcKbAhUJS6hwxMvlz+qOlaPWwUfU/+PKPJoxSFqwFY7zo7s
cKnVwgKKg0ZKcOEI0+ySrIt7zg8mHMOiASIVO6IH+quEMTbOV11BHnKM4f8sdckmnpT0lZnNDa02
gdRiO+EgoM8ZP11wkPPfqd8OtTEgp98ucXCiDYYSDoYTN1f8e/pXHTGE3AGGx+f+k3NpaRABtKIV
1C8Rd5+YmM4zuVb8ev6Ll7nIOKphvxv+25U4upgjhXPtbChgEj3iFlSGsA+3jUqIVg9mNj1m1FeM
QWurb8VMfFmRg6QnFTaBgPbWCwtBK5JOKVJSw7oOJ+yDmgAtDGZYKt07yK7fOd+9onQtC+ee6P/e
4yWwccKGQNveDjqOpNRvoIugUCHdGcS/XgQGXVCEbwz11K+QUEnKfP2kLvffiTQakhn2hyGgAp73
L6XxAZEpHE7Pa/y1aFJzzE9DNCZvA5VDdcCHdPMd4tw/G35rs/szZ9pPk7mhwkjto8gJGzb8ZK+J
TIByo6WSWwlkmRdYNV1W1iU9jf2e2qs7hujM75AjVAql4EDysvIktL96bz5tCOjQFW2dp4rI+hAE
gd7DsULpWoDiFl35PzcROH6k86LtuVa1hMaWn0zezkU6jvvVuV9iYHJyyBzwDha7gcFZog8tQ5bc
ag0dOdZWQtb4g9qi0SYljpBqaoYlj9uKNP8D4MMOMxkk7F1fEjZSgXIvAbjM+hgavMIIW8X3k58b
5rD3AlG0hVCPLFZLBuYg5U9geGVAKhgXDYjdKjQL1/RfUYE8JX0D/2FEGbet2NbACulIDHvmv4JH
7O9HKlov6HRtmnsuKi01WO27xKSUuKBcU1nUDhTVFSRpjxU9qbe3GhZbM63MFJRtAw22iomq2G8x
spmTll6+iLQpeVp3BvQ7ZUr7zzQxDZORUsQUVZMB5SnaQ14ucNwOm3kK6eihai52o0QYsyn4WEjg
yD6GBqanIXDVG4AhEcm7Ac3cQuCgEhPVjegDJApooJkCdAiM+8l7dOSdsLbtZXgn8CjyEUCCc5WD
PVvFMmJWdncwGGxHnsBUpR3SIDEb9teWFO8XE4Fw87iiprKUvndC/+OFYfsYqUoLAG10Nseex0NX
DJEn2RHyauhwlkZp6UxdPtVGUCvKhaQmScptN5FOrDLhRLk743Mq/aSnizLnMbwBq3TktZo1pTxe
tasvg8eS3NYamlNMVQ0k87X+9bhYJtkNKf5hyEKKfI3BTgpjGoSwEAZn9NjtAd1CMV1pCDogy70X
l6clqmk2Ps+wvVPBKmQrJGQbwmhDJ/vOYNsUW76C1Uf7doiVpUNgGKhfMLJsxDztpMRgP5DORF7E
Ht3laXzZojEosdPNFhBlP664qnL2xXHhK4W3xtBrwAhzLkGmZo4Twd4PRTLgpv4v/ucRJg5SQaOM
OZDVIqPMdPvHhqioFvVWh3qLVQmxUx3ZOtdaXzYGdyizUyD4GLjjVm0+mRH0F8txyTZojCzRDKos
CupxNQ6N+Tvx+LHUhvdutq4RtcV4GWhaqpCXPNPWnmm04NxmwERUKhPZR2I8V3EinBiI4QeysAqd
G+nBNJdG9tbO+6oJbO+9RHHmIdyfjfid2DEHRwk86EXD8OiZV7pzKSqrwY2J26H8PuJKeoC9h1aZ
Bz8SfQhUjdnj53ogVr21VaznmtvhUBbn7rsk0+GL4vNrqv6yJ2gvdQwZV7krGe6gMX15fjzDoGw1
97ZgoNpX+BETFt90RYPS5xrZEVRvD0MvtcFkPs0Hgb8EsqiAxgDpvV1K+IbAdXu79+6l8VvUq74l
YUXy6Mwxe5WhGEMMbBzjy7wHCA6doGLgXWDt7fSvB0xjYX7L4s28haU9V8f6UOfgmD5+POrMzf+W
edF4LICqAWx0PGQb3gp+uvLgNwCeiFjhwh1ROpmCBC6OqYoRBSJY2rY0apYHguI1rWJMSoAieUl1
0sAAR+zlgmnVO7/JGZMs6VEawVP3OiP9w8OqDig11MnNGxIxyrl8EUGWX1g093ds2tBX6p/J/crQ
oNz7R48Tentft6euGb9terus9adhUGxYKTJWkO16nDaGQUYel6gIMn5yUOHaRIccvZtfIKdcue1Y
1S0XdUU3MICW0RDB2h+ccbIxHh2nH1M2QNB0klZQPmi6xzonudc8xuMThIGXpeCJDgJzRmukUF7Q
XR07Zb0ohmnCf5p63cCzUKR/7K5B5+j0CvVkL6c/EWTth6ypC7EKRWKsMVV+K5c5vtB1ZRbmN4rB
d38Xw5aIpsP0btv7o2Uh1PE7cVn3pvDIUFUXAQcbL+UroOnBY6rwm06IccsHr1XRuo+WMhC4dOpP
Z4e0JF9IKrdPlXLgXC1b0sK+AiLhkVSUrL8hIUwfuLPizQvl1ZL8auOvunIOhTY1GIIXWUkzaMWD
bP3lJ1+cAXSSgHJmJEgbG8/R8LAKkXigiQzlvofs3wtJgB/krmT7gZPbqoDLf+kAmBs4yAgKa8ZO
zFdxM4fR9Os9bQpdj0IswwpNOiKIZ5MKvifvY/37vx7AvpwJ25WrkmiAm5cKmWTgAlGzbtEy04Bu
83+my6M4GfAxfACG3Z0+lY6vegaA/AOKZ57XMbyJNDP+otDcchOfYXJ+LAXc1ySlR9a5tWGayHuW
A++vqXuO4sMUJqhIYvZE4nJB+dpU32EPOK6xP2n4GuM7C9XKJ+xV43xYoCrZGR20K3CADxVJ0umT
qwmcGgf96BDEJRPES0SolmnPDKXypRBxq/kIlog2Dz8hvtU+QZYn4aY2cA0G5VbllV1pwdyEo8S9
Atjy6b7vxPFbCIvfE3FRleDAJYfm5q/no6pCsQ/iFoQ99rv7GmIQzET/9MSny9UXgkCcVWppkJ7I
UwmpetVPIzGk3jO0cLiAyQmYxhQBR07WO+PH31ZbuoKfkf3vGKXuTIMEoSH1xGwEUM4KNi/2+OcC
AmiGLwCRlzU+LDA6RfyNLyqlLlNW0B9fAxgDAh/j+y5/T7s3ZorYXritMNDK9uKJBniwg7YDD0Rf
KbIj9/NmzRZhfnH5bFrC3ZjhMl4qXh5n0kpj4cWGpSEGMPztPm4OOTtKqc0yDgozlLLj7jMLaQaJ
j6h09LApF+RbNLF5lhqy6vajZBnrmkQ0K4sNeu/rbpsg09sUy6QpEJPuBYgN7yx9lLihXhWq57GA
IhXfNNB51RuEDrt3Kag6NbKAQzXlwbzsqcepbmIXDARl/Bn8oXCTP07a5zNvZSwl4lGd5Pd849hN
rPCNhVFUpWteOke0shnL5WM4xzwyOdDTgDF6m3Kfmx+CWusXNSrBS89YqMda3z3wEqIfgkjKCDr3
t3qik6i/7TQ8apr3J6JBFWMrPHbwS2aMt09W6ocmY0KUFxuJttWwDyRM8mDdrN8X6OQKYjLl2VzQ
WSnQPMZuk0G1uvxgf3EFKDfzqvUtVTqEtuD9ILEdFBONy76uxxX8r00gMiHiOKlfdzm3cY85rHR6
vb0pOubXTfQYEG+xZv8nkieoH4i+ikQAf4z9dj8VuC8aF7/5L6GAIO3yor+/Tw1q7x3aaJ+ZvR5E
9FLSJ92myDbX8JiQk4WsOjWfxKmU5bABsr67WoAPKkejZZxvRXw/0TNP62+OdzzylON4rVBiUoOl
tVnXmtSiL8NxVSn+H4PCbWj6CiylZTC7TdWtMcGK7Cy+1MEyKTChA8uyj4fdoHubKhzOEJ0Ij5jJ
vJlpmpQn4pIG21oduMAo9v4p9SlCUckH5oJaYpLqaigPZFTr/LD83dgA1W5DEaAQ9jPo+omVkthd
qPkUF5jSgBtWfgHmNT9X3Y1bnaYuN2+wbsGOSZw45NLtq+0NEfu5jtD9G32NxFccsE2h/1XkAdxy
EcaVLJBD9RpLjnsGGmc54aJCrfnatbi0KGcSWSiucHKydo4/rYyUpd5kJ50Q87tB15ZcbPFrdGph
vOU9S++sXLRIGVOpSvY5gAP4SWTl2a85Vu5NLziEZr5eF1DJYMD1KNc7VkLVTtWtTykxb+gSVZDc
KC0uaHbzMsB+EhzHTsAqEIKao9ggABXGFUSQNK/KhR0IxN/AySKzY6xxn7N1DsYYTjDGTpGQXofA
d7bS+LmOckG7UrcnR1wX3o99BHE+mOVhevlBlOehkgH7a675ytMGs12j69oPL2FQNWMIbQRbaQLw
yxFpwqVcS12sRpht6O9MxvP0hxsihLkzImmKYccfC1O5nSKFPabEQwhMZH9Noa6CSOKdcTjBcrMc
rgohovFc0fbZuLv9Tsa2ebpap5oK8gLzcVtwVSSu8rONPrMn2+RY8uEOP5iU96A0DZAMXED7BoyB
7tOxk0hVtmlkdwHUE3MHQsPedtY0dg9IkkRl5tjUwjByzRrAbUrvuL02QOIHKBFxAIc2n+QkyeZL
1qyynVOUlQhKC/adE+L/dakba8ITt9OtIbOtWgvmBRKFF8CC50jX3jZeuEb4EBLfHfib+nzlPmGB
hj0U2U321q1uF5pdqxhauYLf+Jn5PNpE9eL6ejkZglmPJ3UCSVfkDOe/soh9xfD0y8299QYmivn9
9ZYy/5gfcjof/JNUNjOW2gF0430nSORGXvNVHVMyGrLgRmQI7Uy8iopQLB0aICJ5hCaGq5Zi9Y2L
nh3PjnQn8OwG+qIYwJZ7Aw5bhHoUGkzY7JBzBUN52GgKNQYOEq7K7b/0/jr01mUj+zY/2UbAhQiZ
WcYniEC+/GM71K60uSzDrMVRa+Tpj4VN/uIQD/YptGAF7r1yO6tjdbtFwYUeFiGdvOlSQ3Bn0ads
5z8R0JKbfmAlTq04/FFS5wJApc3g/9+bR2QMbmBW+606BoXCl9IQN3jOWLfgw4j/yksComskWw5P
JE9O/WDs3gGlPBSsE2zvHGFsoeAAV/VeZw8F+Wks4KNaB9KxANDk+T3RVcuGYKrSCifppt38tZ3J
yeCcthHNbIm+te8PpLpiDmBBs/A3GAWDD2yVr1EcKCxEEe0tvybTFicF3LwxPkrXaENnfGV9XQY4
gEFGJ+e0pxTCB1IlnjRg+T6IGt3NNES/gRpLjDmUJDo/rK09MOyIsUmK2TkEMBfVxeEDpAns8WYU
m2uHOn2IHNB149mGDZ5S5k602W6u5YFk7Y6nk66C2x7iUvW44skFU4CXM/IRQzkoZViDhWv0NrhI
9iDQdFg5T5MF4tIIN5dwUgzoNG2m6lMqGG0arga8R2+zIQkNmHNdE240xyIfEM9dH0l6IbgbhgGk
UEzmjKNMhRXZxLszXybZa9Q7tuh6WvWl8H4SvPnz5VduQfZzA3F7cpF77zosMLwoGJFjqg9wNIxs
glYzy9rKpBH4qvVQw5v2RqZhJlccblqkPkPmlNicUjI3RGoQkp1wzNPu1uB3GP1vLVjzeJ0okj6n
FdcsG/I7V6eALvrT5edpKe0IFEjaCm24yYKgaERCqnghuH94Fbk8dlzjOt2ux531/RH/j3QHzR7K
ACxcW0rIAqFZF76Lad7xQOh8BqIgDgdOQjV8K9YzOIAR6v3p6LIcncmo47YJmlyt2r0gKVK8GiVn
B4xmS9kPyKw9PwdqdZ+OG4f/DVCPeo4F5OTiJ42orV4uzzHvB04NSEbEkUwZGEFJrQNX+P+f96Vy
8gHkcA+V6HKiV1mi/uWrjA1Uu5x5bxGBxSaE2yCxiZVt5lZHYoV13ZEUQF7ls1+Dyb3urZIsJs4Z
5c0Ukxf0uM0tC4Qy5eTqBN4VIGxsMdq9pTmwpdOXupi5HZgMWrNYUzAOy65I30laF0/tAYKQvKZt
BlRfkDV8LsRpeJwIoTntITdjm+aDeEuIdYV3g7CKWQCddZr5BaYA/VxPqsPHGXtLl8t2DagllYvs
ztFimC3w/+CsO3K0iVRT00ftCwH/Cpa3nlmoPoqR8aTVs2cMEr5kbZAjD0mzGgnv6U8lvZ8ieGcV
qjMNraB4OYZoJf9uOCe4ibacomtcwtXuQA+PfXZLLdRmqiL9ahTCckx53IcJVCytQaPOy7yff2OS
ufc7Q+SKBc7rs4XZ52aRnpB+aJ+w4C4ngv9fwRfiRLo70AJWjsHQIsCafc81bi1iA4pbrtLCtdb+
NDjVPWltFBhomRQLTX8NawAsfy7qIIpbkGYYTjw8lkjYU2uzaElBpDMj+BDkbFLcuk6VoiLz3QOw
6PUmk18Ar4PZDNt3f/BfiTw26N1RhKG8AwS573C9D86bBLUtL0CgdCppQVWS1uz2fJ0MULKzkWRI
QNOeummrnecy26MKsEVfgMF0jFV38i9fmCQFISqiwBYh2Te6oMh2NwLVRGTF50NKXd6U9bOMMzHs
yqfJ77OSZKCzUddYpjmfNaxsHxZrDkn5swF3U5fbuImG1phPwidF8OZpxpIbf4C4iS3qn4uMctj9
SohsS1Lj+nL2UteYFj8rNOKxlZwhKoiDUja+/xuUOTYQrZuvwPuAMGB6go6Q+hdk7tZ7DLTzL26A
5NerN7RILag4rF714qU3qftgVT3hP0qpVrMNnwFaUUS2efZZmrPj2tERXOrL2eQADV9NKa2bswRT
v0Bqw0gG0+R4W1KBPzaOkPHS8LqLKfkHpO1zkLG1cO113NajDVaI8DcRvoGVg9Ehty0NjWS375Hu
vbjBndx7OAqhA3lB2nd/NtAsWeYA5jPHMeR7sbEf36xC8u4r4sQFQ3NvjDvu0t2y8si+v1xF0sr4
L/2H3ECClAKt2UhMXS/plKyXV47haIN4iOX7E1ps5xEud0cBrnTRtgDI8LneKSzDX8N+Hu5VYbIf
OnYJntUhJHQsxhuIDJhsQ8ival4yYn8yj4kSre7iJAzulGNYLq3IiuHB0zBVA4LK8m5SilzlkQl5
NN1bqI9Uspya2U1jhYOBVVHfM5047Sht0pZXSVM51gzoueUHR5DXfU7QWMa9YTDK9q7iagajX99e
xP6FJXDdwR1Qu11WFhdttklw+Xj/IVqmgv8SKTxTeBtxh0YiT5brolSjY0yTLQCfqzhDoWJp8itL
9h6lnegFNJTX0a4tZZPLAaXI0pubIxLRfY/a6/ayFvY2MeQXZnmgJn6d1SomHII/Uc1s5fWsdi8S
0dxsh0lxjxzSWgiCoAhxzzJN2C8QRJeCe0/MNHFo7mEANs9TQ+KWjp5dAEcG4L747x2uFsTOO+oU
ifZMiuNvP1o9bxXyb9uyiI5dleBCeVMqTjYIh4yHkzJDSj0jFc6nYquO2gdaEGLJSJCQlhXJSQIj
P5YiWsMggzXXhyEcb9/tDhB4SP4H9jiUKFzURdwu0O64xdhIUyMxEDAYaJEwXGVn4u1l70DApzzm
LWv9/9ZhEKuWoZbMaA4XVu5Uzo+R8QKd0QU++JyhAtwSS9/cKdOPc4c4acqK3sk5fu0FX9pNR64/
hHgoW2ujnMlS+a0qOPH+C+l8WjG6KOK8sHNsMY4IDrkygtEo5MPQZ1CSA8nBhyvG0Qrs4EHzD1ci
oKUWh0NEk/J9k36qbzfJS5T8zymYj94cE72G0DvMQpZHuGIPGahKaveYOwsn4bZrGwpSejbaRxZf
qR3F1pX+dkJzRqfiNZ7SJFPz9gp0jwqcC1njA7UhhsNolWGXEb5ClmaGFG7Mz7fjMSVC/v31NZyA
k+8w70FfuD63syYhj3IjWzHEEDaNBpONOYqPcXRYXrZlQsz9mAzhE3HtvwaLYEkDy6N61IuwdLQi
e5AlyEaG7DZj63j1UF4mWH5ZLnJBG6GjhP77hCRZxSfKN0rxdsRhN6pXdRw59HeBNaAXko7sP5Yq
LVYr6ydocd/OQq3BjXIIn0WOeghJVR248b1p8lk575SI9Yn9kqxkyv5yPwUIioMyhHZBYUZI4lLl
CnGvhXZof1cBjiUWpLIFQuFV4vakZLnAkpzP2DCKi8emG4vbAzKiAllOAF8G1bSqL/4M2waOMzEz
blPrcHqR0FQO094MW4AbCXdydRCviLEvcHoMm3TZbcW479XGEVAWIxfofgKOqY4jq/3/mmtjQqZa
tqImSs4bwJdLIen9jRbeLBFxuEfRUNfPiJGIGPg5Lo9wfC85g++Twm51gzTT8DS2XufKq/hwBFdW
1cUJwE5ulb4fh2xcz8po/MIeI01SsLGylQeDC3XBwgRiwbYfBDNlOwyXr8OTKYCosik8UjGDXCEE
naRPWAJrouAqcBryrxhh2IATp/c27end6VATQN27hCotSniUzOy0iKQDH49rnISLELZd8fu8PI0V
AstjmXjpGnngp8i2lt1HEfy6LMZ9EbXZMt89k1SMt3Vk83O1Q4LmN72zr5E8j2cAAbYhH1bovIql
NmkXDOI71PT2tZd/XtVj1Q4zRBBw/k4ZuT8akEBT6bCG3rdZr6W/Od3aFYAFKAg4XMve7J+bQuIM
yRARrL6XgHbn3vM0x9/3q7fkGTp5RlhFAs+K5k8DL/nr8WhjQ1Pmasw4jYbANVCo/tawuKeF1mg9
STIYHFjQ6CHW0CMDmtFmqWalJAip0rdlMu6kTnu0ojGw8EjI6W2YIAHJFmiIJLBVJBlwwdVK7bpC
u2L2Pr2w2tzUnMb5xF1m+RTOJ5AM6sF7koxbWvrnRrRoDXMGzj3ixSxMmYykbVsh25C22ryt4iD7
7Qzwk+QkBVnSYv4Fz7YwUVxzJ5syVJBo5w9b9mcP3gP47Ue2BFLVt+LPBVPkIYrJGIRFpT5kvHhh
/1trTfRBXwlgR3HlafiP/PlhlSahuSft6ifs1hjC9CyrMhc2sj1oTKYk3GlJCs8L4kjMZ5IP232j
h2dZ7FR2WvJknuwgCVOenbkgXepKAeRu/7HLjO0Rrr1IYjpj8ArJKds0IYt34KscnaYiqPsuqdlR
eN19LZU6Iyp6btGinIM3qjHxMWao3sMZ2grUUDoZr/+6KGNuuB4krbjx5GMJVcDSEDH5tqZAWwqC
oUQ7P4hIT5jmhy3vEFWlRgRc487iN393DHmM7DkjkAMWCXC6+yAvLYSbPAlhG3mZX1hOgfk2ag51
hJMN3vZ5i23Uix85fUyb5QGpOuP1KLzxovKkpmbEMDB1ZijzYlLtph9JcvGAzNC8GkBP3GFsSWuK
Q+LEgafMy9K9H++o+xB89HehWEHCdNB4nkyOeQdVQtPfcvv8lv+yFsylH7qw2DNgUcfKY35G4iCH
5JUVeP+lPCJ7CxPQxCc1bGdno3oA2LzI1ihgObZJB+rEy3+quLMIMSQVfjXFNKTqnc9ujeKJ1fhx
lCFGROuY6h14D9WqumtFn9vk4eQdhU5eiFvX0xKfhjq/np7qjLQR0KtqFleA6K6Q+4wBN0ArkAcu
feEYCi+UZhA1z+fGNplFMSV1wdkMS5kNQjtMXv9qcw32VDxrBWnlfiX8j/E1dVAf8vafns3w280j
LasqXAMipZK5W81u+X+oqOyyjxzen5N0U5YwVkHNovh9uPCWii0lXHfGXY/feN2weon87G16Zhiv
h5iPXnzH5/jexfTIWGM3SP1Zvr5hm/nD+qROOZnBX/CVSGwT8nUD4LtwnVqjqI6Z0QalHLr9CNLN
qlc3wqg1ajthAxpmeOtHh68caTQjfjTsPnZRchsNTCtIdKPrZuF6th+S/PY8hurWJ9QFP8rT0ANz
n6DGijKvA/vv/Tak5ndp/bJZ1PeKk7mPuU6CClah9trcgh7DEhAEEcIP8QgLjYRzkI7Qtv8mOQOK
EhHM+SqFrvqew3a5lIXV+hM6LCMKz7l4l0rm5DPt/byT9gMOb+r/bqa8Nr4EiMna86kqWFP0AsSu
dPNeC7UUJJYjxNHGoHLF0SxrEOtzUMjWbolrWdnocOWtq3zBh7iApO+WqROeFN9YmoIQp0yYaAj5
FtewsYeXVv6PklZxgZuowflRHNEKhkIlAD+qu6Csffr4EuyA1PTPovX7oQo8ISAU37D7L926CEd5
wVnDokkNTqi0LhvWJZCJTs0nOhPpI/aUobG64HOV/1mt+Xrll2vZK+2xNTRWXXyD2FpGygIKR9dn
8msk0e6uDtBgqqa3CePuh2EbKC5HvwCdgnPWqoFeTR5B61ErfLRJTiYmGjXrcYKJl9QXBz2wsEZw
6sXALhcjTlH1I60h2/aSMHvtwFcifbdZR2gemYvF5fuFz8rLtJYgiQIcYBYm4zhUvvb81S/FQ/f1
CLb3I+N8qboo1xFcLpXOnZ4jIWLbeEgEF19FB7C4ySGOZXlmRfLnWSdaMR9+N/NkPckdBsR5xQkn
rBzSob2iSR2C8diaJsr6mm5nGtjfcQIcS94U3xOyL+fvtP9AQjWLGMoGNl/YZFVQJqwigoULRFem
Z2yaeXT7MNciYkjdZeQSKIKWX1X64mFAtE4FbxzdWRloyswBWfGzUJGFrMsNKOnZL61MVZJIO6Td
xqmngqcQdxldeOJfdbu97OWJK0NV/sIEgtvBL/LP+HzThAmKVpgHg6bS0Uo4ksdvK9ELBuydgR7I
llmIAXG2GZ3siMLApfYqPWHvLKa9LxHMt4/aBExfknD9mFmn+Rzfn5oFai5BfZsg/Cc7K/pJRPMV
UmvDBnJXAw0o/kZp9jJaUVmOE2OBwA6k8RT5XHcbpFUQ2V/Kz++a5S33Vt2gcPg3iBjDyifpKZmd
hwtx7vnFcOjPH4Ji2bXUeF5jqUVdBCU9xPz+SNm8j49ggKB3mBa2DbK8I17KRXeHNJGEwZ8OiBEK
fNboz3W7CcFgW1X9eg6FQSgNWaKtdZwVkljX2la/hbVqnUq3EHNYg3vj9HOi2LLc8ChvbuLXWsae
vwZ1d1jJZsFp7Jdj6/g4YhbzJ6hHMQv3WG+gthtUftJLq02PvpqJreelGfJEen+WdNIYQxNlU8Jj
X4bKB2khEWsK6B7BIOZ35bAew0EfokwCZFb9XJ8eNeoKvfVEq/HlT5zWfTvIBsupbcvkyRX033xl
sPUq8R8gK4ryUtqPExED3Bw9FChWknEUkiQGPLcz605dqa2PcN5hOI7fG4mEgfu/PxqhMLpn2REo
9fYaQWTwrd4VE5KoolIRtMiEk/0wBaSigkae9bKrsybP5aJcxMOdtcAhz5gbJVpHJryapTId0GPl
ycRAAltMKuGEWYWTMsQP7+ahU4ezGJRBcmeeuCVrA9MJXFln7SEaD/gA/CAIihO1SBAfoOYJumbe
i3vOuqw1InptrUIfc8Rji6cUcYvU9g53GmrrCN6q1K3PqyTcroHY+cdoq4wx0lIbCF0RoNzDuYcl
PrvU1Km9z0aXJTr8ekJjUWf8IXy4IJPLEvJtFoCZMxXREM7dOZSZehqo3YizIK8oQ0Kba1N3YipA
uuwOrpjA63d0Ea4Ku+/MXZYszgy8H2xnBf737blCvyh2rt8zBFVBN/EdG2hq/Pi8xbWNEAa1CqRn
Rs2mQq1YThkAok/i5KKkehv74mc/XUzaUpShAbNZSLkQZWmHf/QBpokfXftjRNJIr8STPFd0P1O9
csYI2Ted3C5fC8WPU6fh3DXNj2XAD8FnDCpgcFebvLrc6gXOB/iaCD9fh1JAW0TU3JIJGcFBR+H4
tbgFELyxPhWeWsWynyuc3ZnUf+td0JR9ldMiUAm/OG4V4uujfJlC/OPgpbm9APWaw4M84WmTfDsB
hWwgDU5klCJuHa9DZy+R8AFw7HwUDB68G+I9IXIRjHYS7FPBtHd7Jr4T/vHTt8Q1bholYnkl/Oxv
ryS5km/3zgOTMR0igz5LdRUDfa7+tb8VhB1R28h7jFhMc77SoWRu5D+a5LTVGF/AO3PAgS5NyWvV
SudPYsf8CGpB9c3OiAu54Uu0bcpgZEioak6LA/FUeRdl834IjT2CJBtL+nSnl6Gxe4G9vdlHMYMO
N62yIcyRp1MKeFNJYFtrmLeV+veJpXc022xkrvp0QnjznXOJgzAkC7q7ssJwJxxAMYINeX3AzanJ
9ZE2Q+P5vrDlPQrEWHA4O6hvZGGSO145Vh9cTV8+7UnonnTpOXuaTJjh/8pntS97RhncRojUwaGK
p9T5VhK/3MOprysSVdocsYpq7Mj1oWbVvwM11vrSXLfTHe5TKOp2P83Lvr2iZdrKQIrAmp7Su52F
uMJG6iVgME0kqh1AZfjNWQXkhQoc19Rx0LKu07Hu6bGFY05hpul/FA0TO3N6ivoJctEPIyY4LEhu
Sn4LYFCyKTADc+byioSn55ALmI/0SaPG2k1d5KzeM2F59mrxeokxvlESbxR2JsYSswIia8bI+lYq
XI1Ie7YF8T/Xudq98nZPXBFHN26ypf+5Ha+tTaY+a08VIQp+hckKgMtktAK7MFJZMt68cPnlQFnJ
C9wET+xiZ19WzIRicyIF8hKxwxgfnOYudNBbAfvkT7jrO9Pr9gbrQiYpR03RPhOIIXwa81T/Ze9m
EQjknDUwyl16LC3fQSiw6jUIU0AdsbkGOH0UvUdGMyXa6jRvE/yzQL4pSexYHWbtxENEZIh8IUUO
i8RMHXnd2qNsqUBX1ZKPmb4fc9T1uX90ehVS0b7ieGZ/G+7Yp1l/xJYkT5YTkxiNFdau69ypLbYx
80zdsR7DQhW/jniaNRZntKVfwag1vLhY9WUBVWa5QDQEyJmGxHHXeFiWL0+Up4OP9Tp2dhVBF6/o
3v2/AuUBBQXP2wFq17DSFE8lmNukh13OnHM4aJIsKMpSrJY5H0QskBWi1d7sucYHOQRmQDZqO4Pd
JisYhSUxZ89rWXBzt70vJDDirI4BrZZFEciDZFyefQY/fG0KYijDM/F2mJWL+lL7bHnDcMigNnQ5
RWxl/FcVgcc1uNcGJq951x2CwVV3loGhqmI0I1MSIHPeV9RPzLPlDXfnnA4RjxHyY8anchIYCX5Z
bseAMEahQz7NlF9m4mRVrpfSQhzzIWuSja9JvRmNkOPq64ycFE0XRqHTeXoxOrQQEoimmz9w48yq
3VrOuanfekY3H1pQcHdL/BPBqSeKEYkZWAhKPQ06X1aR8+c3HW2LJhXLSq290pIEdrQFnZ742Gw1
fl6XlEs9yJAqAld/nc0itJPvSFn1xUCKVHbsqx0siwxL92PqnI730CcqMk+WsqWiwYSQw/JyGhji
11eYR6ep90S6qs9yR/lvWncKP2Hx5tU87juXHDY74WFq5eJI7dU0rZ4KT+9/qxY4Cz0r4sSKzV0a
Ku+HiPYbwKvhQlKRgJf5Ha+Ci//hDJWSdPiHpVToDlifzM2DRBLYTJ+BiHNJkUCw8c1YeCPqgK6T
S3z2sMhMlNN/A9tyMbwSgJkV2KKzl9xSOCk878X1JYVp9Ix6F8VkBzRX4ddt1mDECcikBm1mqltx
+v9JKb0IYNhdVrV4LY9k89bxMW1PnV0xufxqIOM0CwWjDkESHk/l7SbJUicsQx4P8xWDCz973pMC
LNjGGiJIOMAglhxzmltI0b/hnlVyvaQE7gqSQO7sNeLVRbfAwgdIor8jDytxw4DUkaYLm0Mtg/Th
AHTHZhajw5mdY/djFSz0VXXJjIaZV6l8DMQO2mIcRgVG2Oa1DIviMeXBhIpUQ6W3lrSU2pHnobZx
Cu0OPBnNilEuaAkjXvLJY/ZEBXUfdplZR6lf789iJ/Hp7RXl42KqvVDNszWIb7epYvBDFVjYw96u
UIwrHldn6I5rEOwvqg1Osi6EHCZv6Wuvv/v0nz+7MamjXZB1TqKra2ROHUrfxW3afXMmk+mNq8L1
cbKU7vZDPASTkvzrKO73qeFiCk67gJe/M+BPVIVaeTs872Y79Q8KWKvnTK43bCYUPseVJukEi44J
WG3F6aKj1gPeojIAJ6TPhbAZu7O/r0VTm+IegBBFjRCdgvp+JaS5ATbKFNOLmsz64wNwo5/2X/Cr
xlN+o/OakrK3mQmhMtTjE5fJn97s5ksr/EMmIRlp+42RgBSG8/5LXdJM/G5Vi9vXnDDsetvT+U2L
VfrGhHKCLpjsrlHJM8ln+fRczAlwCLTv0zNqSZG2lHtdNhGginkMOtA4HaF9Mo8yBLEv4YMJWjfD
7SBmqUckDvyA3bQdbjwqH6gEQs4jFgVb0w2OecQVX8f3N/1G0WavMiyvc3s+lBoKyOEXWpnWBGod
2bOKeeqUPijiAgjEi3gBcuhBMJ7DFrCsRLDLvoHnHUGOXsWbrde6MMJmTn8srQobYnq3c33tAcDj
O5eGXt1mYcl3BS0IYfTulO9MOAFfnrH2OD2T6Jb1fvjShTMsSmIo0zk/vQf8gwsjULUvfno1lelf
ZFWmscEDCCPMN+8tYSqdDB2lQnO1q+vCFug/FQ7Ss+gr0l4V3DE4Hv+hTLzTetnnpqWxuQqAeGa5
LP496YIdu2gt08ltNdbxf9roVk61Gk8Hz30rsP+H4mW/flzL/H5P6nZbFsBux4exwKLGgF4ZAiKD
kSXTbcpNhqSuKIuXeVhK8Cw84NffdW7olFLPfArRdmX5GNIwEqPdhKiW1wlMR3sYShV/RQxoHAo+
bWTE2hAMyN7ZVWsAGwoDe++gVQ6qAI/N+BIGyhMJL04jPR4TPISil10tNUj8L6R/BGWhXYw3M2K+
fO6nPPu2SrM3Dn1nRRSC+luBVF+2/qYYt7e7JDTs7an4SflSISSUnCl5H8sgXSsPH6k4MiGaBN8W
xR+T7g+Ffmsr/8aho+wIrDknszZV1B6xHo6cIu/RYHjVfIQUind8NIzs+v63EeO4B3mdc/x7kAvj
PI2X94BCb6b92ur3OyIR6NJbouFo/kYZ7Z9OjoMuyiOMEYRsXyvmF2AUYdGZ6JXku5oakGcuEO3j
66snAAvDXs8s0LCFLgbx124cFg/ceV6xbPnmwV3d7fQ04DtRtQSpXRyVHU1nTpzzw36A4EnnZTlv
KzHDnAuEehzM9TwcqfZbVq5LkkLXx3W8fHBxAgxL01qHywrPEY2MQQiqI3GfBmCTpHXocnZWZZ4N
Y69NucqHyVLx1aSh5vm2PXR68fnCZ1cZ7ZCfqZx8B3RcwhWE9dlPhyZEhW4FNHQxYuVJRRkAevII
dmueczPET1eN0369IAnOADgKGLGgbMN1lERlPFn/gxg6yUL1QKHEww9R2mXQi5lIjMCQ3Ss6HtMW
VXJ7OLysx0iXpsVfjhsD+V/EE/Nt1XIlYqlyZUb29ePQuKEmwOO+XQIZOgYkJ91HVaaEH7jBzT+d
JGZv+qqEPXwOiwWlcOoCts01M22hqiQjUCInmpanb1sub1CgcXlIQMaC+6Cz9duwa4+YNAx4qTuU
k+eiyw7ka2LxvYdrsTxujOp7bEZxp2Qn28SMeo3bDoDk0NaUITnODOsQ1V1AS86AfcFlhBQXOb+y
sqHYDa6pgsprsXrl0G2yYS+TJwAVAz3FKzhy6/C+6XeZ4QqE5AKt/Odt7X75y7rlAgyYCkfL9nA6
6DM8avf7rgU3xO4vQN7C1McCBr84XiwUHP29BhapjhHDFV9vpAh406HHzJvJa501VZ2FPepk93nT
mN47ihzi3+eQ3C6OVxV8eaIl89/m+qXWK5GN0+2KOyDwWp4/Fmtvipmx7I56nLnyMKB93m/esWxL
P8v/Av+BzOndc9PyXp16sS8Vm3BRvYtlgeWiE/Qw5OQZHAug9BKmOfEZJMYX6BDCBzHJrSNsVtHB
XHLqlNa5Y9gDkJ74Rd5m2PzmUsjERj0h1GkblShdjBwErx5nt2F35ZFr8WXzsTSc4DCqu2qNCYxO
/J40HBpksX6c2xsVLJ9j+KqmaPQCkGIQjRfCYLvKTS36QjjkwBKqUaJ9fhsIeciiM5XyV1tL7G3v
4frm0r1eoY1daoJoCWymRi0YyJLyU5OKjlwglgALHfwjxq5/tBOLLcuSsx4+LCuyn1ikJKKBcOWH
csWGr8EpWN9kg/k8lAjr/x2jmZA+jwBCEwkRnmoFpe01LJ5xxUcPXsSkoNpwFqe7Ulwiedgw8WSm
CiXe+aK9JhiZYk9d6S8ZcpaouzRJT3OhYnSOEJLrsNd2Ri2ES8xyJXkNuI7ySbdN9YNcWKz/f34q
eShUKnAzHCBxY+cnOSZzAIXTZbZTg3S5uORSwbtaZFc20wX+cItWq64jX+5DD/SH8o9lFJbscenD
Vz6HOx7ekmQxJzRl/S4DjLbo+qxiILG7qN+jSRAyiZhR76hnJ/58YVOCG+8NRv0a2WSjO4sxLmIc
8Izrhx+bwqvQ0yC+UmtRHsOkCcQZd2M8YJtjYFsZ4mqZzMHI/x1nbs5o8eCpkCRDdP3r4onJFPfZ
3NlxBAhUxLTJlzU+fTrkCkMVbx2D3RopeO3x8kTtNDzQefztV6Hryw3+kyjVw07kcrZ3lFrKhXKM
m3P95WJLrX+BLLFT0wy+coCNx4/qRTRrdGPV0zdS3whjVf6ydJLbm1bbTNVmMnAXZcLt+eNB6h/p
aTG6CMnNArLz4VepxiifX4aSxGvajSXF1bs1BARjqMok7WA5As1ZZD781ay+FxxCk7IdDVKkQdaR
sNJO0qzCVViWqNilefRhUoSBoLAkLaRMqlcmvAPuN4dLwzSuBZf5XXVRXZp9wshcABIfF5IDtyEw
btnKU/kGkzAphj6OzjVEHUNja3nwPVPgxfPwVH8qLHc7j9jSdNsFNYvpqeOLgluBGhdei9WwW9vz
I0g8wrKCszH9WPo0/jOdDnytJaLOWWygNASIbToYM+/6eD5f1rgFHpyuBryMTYROMEJo75eq/CrW
R56pgxlDIOiAxXD+DgfVB2JAQtYEbhRRAW0CxKfcT+l3DUkbErKkr50f3tZUxQSahtWqgam/CS22
jCNxSPC7LgCovjEQ3WrghcU7tZPuWC7+dmTLu4BZ0vzOwPbjHQcPW350m3YDZ6+SD37D/X2371I4
9vxjWASf4KyF0SRXFcCTDM04FVObUIVoEvGQEhFRFUIUrQWFUQ/aPwcemyPq6moMUCaCf0g4hfk9
5WXl7WZ+dEzn2w8ZrwbsF5TbxDkFSpjeSxfkthVMGHbSJv2dLyIsjpWHbI4IKG/OO/0w6mtbnbCZ
jsSMSqxV/VYH0+x5TjjuA7PkIsqq2NPAOCfiSlO4mVYmSOwUgN/jEE+VqlcJtsp9PcZccII/6Vr2
gJAmFIllGFpupJ6oOODoJsXqJqgomiBcNhX3pKlD2J26k/ZwtRFeGHUyUvbWEaHQNVYgKyFRcXLQ
CKHL1dx6vAb7jmUAtnHTZaUkZnaxFPFrbP5msiOBeKfdQ4mz5l4COWd7AI9WAeKvBv9JWzDIzuMH
x2IRsjaSzZX6opaK6FQJrf7mhYflX1YqeeJ5MSsYVW+GYngDilAXcmseQWWoM37K7gAPqzjyPwsM
Jg6HbQEjPDBhkZJCn7ZRmLPkWOkot3b6LwXqtOWWQANOQsopGbWo87qIfhVCRjkhNF8emkWXUqu4
tqhMwYjc+BBNnk9+T89L1vOtQIZeHj4DKOO1dlDgtH9PTH13EBVdSmN/n5xS9FOXaBl5mC0YsMFE
zJvWyfY4/yaWnevYvg7df+q2APz3LRyaPsgbyr/Ax8qUXDcz2VIZRTGveCPpFREa6XTPqDKrI55H
wLeOkVR+tKjiLrVf0j2EByV/zfAfk55yKGxfS10iFPX9ist3koxkRv2sbJqIbJiz4h2Dvh6SSnxT
APwOxbK9Jy7G3z+xPwnOMXfpE1S7xUhGK6eKN15BB7zrlzU1RcyO930nI+dIE0zeKBdWpXqLSi8r
ncEo45pRU22uh56yFjgoLecvQR/1jnr+7fjuCu0SX+3DZnuWOxLYSmm4emqV6oxPVmRPtp2RDJxt
5ibzxz/IyIWzeNUZOiWiUWOVT8NMj117dcmK4stMYmrrLMEInrsBQ/zRo/gEm3nBvH/R39VfZhLe
eiojWhyOt9ziIHIOJrgX9UGW9nRdCXKm0SbppkqyRRCULpx2SGLMANymnVZdjhizRW/xLT+CEnpV
VQHhlNdwfdKwoOmL9uqYC2NLbtyCJ0ym2TaawNVFKNZjvxEAIEAvl9F8yuCfx1FzD0eLbunKvJBS
KCnXCHlCzdhBqUXyqjzplkMx52hexySnMGRYBfBYML1PMhO9KkEKiNGlCABY0ZDXrRVHabB6WEpa
lORwgRyTkqzJvDFoua8+Wxcfj0nL2AWFW1xvuAfswrcyTBS8gLkfmMHyUTe/HOOd6lgQzgQ5cT5E
RCoo4oMnP/zq5vSc+bDvWxZQjcScHF92IuDRW7+U4sj6tTt62RHHx032T1LE8O0hfLABvv4fJaMj
UtM/fqcvS5+ji/AX2h8rR5i2Lr/uMFZw0jGMCg8OjG2VgzxVu18RoSRYM8fp9CylkHUexwqvJGtv
dZ5EEZSoFpdfoCCm9+yy0pDths+mXPUdnMYZMSuQBliqVttUeCc86T0TFH1AZcmK6z6xceGTtilb
Iop+hC57kbv3dTvGu+ODvdWmyC+RJhrT07KgQP0L0BcXOs6godoYQwqu0wY5rG2zj0ZpM89VpV+g
Aq7MbhRIcdYJgqHa+cOLOwKa/aDYDcxVW43xiQp8RpBDi9NdjaFNng+aoMsODUB9DWhen9/Vjm1Y
oelsI/keHlW/jmqOVQHUVDJmVNHX6KMI4koYZjm9IDP7NrcQ/PIMxaCkT9W0tPg1hoh25DNIxLbO
Gr5D8Kj3envV7lR3kd8LwT6GZK1WHavTXXA/OXJH6er0iuOhZNTsLF2wvUW+/Mk8yv81CiEgPLDO
cILQxqy9hgqHSbCniq53iewHuIhYQAjyIiloftOSC07ApuzAQpBHZXhV17c2P0r8C5Gq0ReLxBQW
IY7VHj5WHtrN0Sb3JQeriGVFfZ/0SSbVej1+VsFkira02FJfCBWuqY7obWL/fCxs5zdd3D6FEVij
xXsE6DMaGiuNu3WZnp+V/fpJBFsApEMhiFa19oiGnhFUDficmp3XH0mnfyvXEoSdvFcrNUh+xt6S
d4qOTol52NhuluKF7mwT1ouyd1bdeLbOgHip/iIlgPuAaHVQLrilXh0KDzyqO9le2IAd08uWr7e9
8Xu+uMjwER859pWKu6H7lo6YyC1SvdtxpABNCncqsdICeqFHpVNSGIEBV5L3vIOE6/092yRFB7aC
WW1y6+rDBoPsO4eF/tQx0Go9TDtrd97cpyLeWqevAzpmGzEQHvzMqH7AxAmeACGQYiwwQdAxKF5D
zWWaFGKccnZSk1OcP+OYW9Djhk5QG2GHYGJC7z1Is1H3M6CGGYJwpao7K0dURcVNBcLeTL3fGUBc
ZUtRtvvdhU6aDEZb0Z3IR4bCC2mcrofOtjoObMEifUt6OQFbFD1P0xtJK8XdfC2VyC60TrER8tqP
FBHKM9Mq0kfLf41Br3KQqSmQ93yCsOBdkl2c+CnpfFWx/LK9BkjzKWTe/u4NXYNpcjHsQAIus4Wa
3jRciOspdO5qsNlhLvodTOtslpJtjyAW1JjP0fMVJbkkn0l9B0OWjqlE9SIjmfieqy8O2fT5YGEk
Q0kXqeJngEvJReiyX2vVvPGmEZ4XeownAizHED8gdLX+FqbZtonaSxEPEf6wyhIASqd3oryE8SVG
QdE9ANKLsmE+tto9SurrngPsdR7n+WUMZGxIOHuHxZ5IYNxrtzhDIWLrkBe8R9DZ7T16wx/yoO6r
fOnG2c/IjVmn9FG58VKN7voQLUHascG41N4mZDRCO31NrXyErV2Vh+0OKdEjqDzWbaHVmF16ZjFJ
meXD7dXB4HHHBQqJbyox5sWOpKEvoqjdae/s4CrpedeLfbCT1+59LulHZC2UlfcMvq5LRljdhSW2
pPprU9cxvKlyofxWwQk43RQtPor25uMW6eccZFvSM7iO/TikpSLtDBQVzu/czt1YYSqFOIh5co7s
BUwGR3/8S6Qg/GPg6es60aYFnLuQ03k+ciXH9ifdlTpUEYdB63LmQUUsfOavJfi7QAFSe7bP5mEt
awiqJynD9qZZWgcdzbUSTBonxguA3+3a32VDxUY8/yXBztB2M52W98XEQaCoh4kX+W4C3sBZsREv
rGty399RhkaFlaFzYMNgjyNDDj64jjpd7GuEg29++3D27a88wbhBOm2vciBCZBq6yU61/xb6kYel
5URLxQQ46HjtDDdeYQoAwP4ktSG3dk3I6wT9NZP0tlTqeQ45N9H4qpXIrD6VRUuV2VBSZStCIK8/
5MwlkvdKSDRIB/xXfoi56ES7tbRg4XP6Dn0I7gFk9lZP4B4kl9uYju6Kb/ywcv7LoO2lePsGd7UM
wAag7Syq0JalVyf7onYhwryyjY48EhK0Na1gVYv5s30Zlz0gDoqDEYVPjK5c3QpZqSAdW1BMB70y
mfQgzR/eCUx7x/SF+FlH7G3dKGTn3eAJqsVwyN2NeCna/8HHRZqkgt/dtT8tCi1RQNLr4Vzriie9
WnYq6tyIli47jqhKhmoOOSlAe8Qq0rtLjodjTM0CQDTvuiCJdu8nBAOxvbNnQL0xT0+6xsifcm3c
qkWqyfy3SY5XVPqtKLQQiUxPVKiWIUofn49AiHOm12Bei37TjFB75fIvrI/FwiomikymA3fw32pM
Q6TgBQ6/MUs6MMW+WdHdFwbiUETTlYqZDTxABBWDnmUf/ZfMnEGNKY1RoQrmEcZ67cI7Zuxi0/K8
5I3U5/7C3n8dreCNg3kgNac9lya7mAvOTrdpyCkcp1B4XAllPCRIHiCni0BFodrj0e0/SsKziHHl
wa0GWf6azQ8zyOAZbijdFc2IuAWiqy20XnIqcEv35E4O/OpISugqgmm+y3pcYA4oBHPozy4nhPvG
C2U94zfJimAkF5/w3CYV1tupwHk/71If9PHq9aHhebgIrVK9p/1SRJoyNs2gN2SusWDDqPJY2YFF
rHmoKigNy5FNoM/0VZ7fJ37+og6Wbest4CA0ZiiX63YTeA8laJozAlmr1bn8ytOkkh4anuT7tawI
C4NCyckU4qXovQSpoURNadS1GZJBQ1G8OTzD1REESPuPtbAWM8b9CZCPXgH79doWSZfTsC3mqZ/x
b7aSWA2nXIik30zSYIdDIDAo28x2K8fD8Mg5VqkVJAF51Z6SKrRJtAZb8eFNjtKqEWE3vrMQwJS4
5nM+o2WUGtTeZt+7F7E3uxuaW2uGoAwmftSQODT9bRydI1+k/g6jIVuXbkFt/KiYtPuQZJFdvqnf
Y3mDAgN3lbuE4E5yCCiTe8VrdkZMEgcNRtrOEeBXHTjgl+j7f6+LlcV3oy8QVAre6Lc0UCrqTYiw
NoRY74LMcDZBxYgEkt8VYvbvUpo4jDC2kfV4jhfcnkabRV0WGkeL/02BZmyvjKY+00OkgiUhKHtn
dulvl7waNW2dDnn1q3ECHaSRj1m8HicL/8a5w5MmybPjDhBE+jOOndlNjTPgQybin1/5BG20mK1x
sD18bK4b+UACzISH2edmby3yZ6Sh8OdDpz1gshh1Dp5HOm8vt01/s8MTzTeL28pllOWePfLQzJUF
SXCBYrlIJnTp4jGvJedQtha9hllJQ59p08IeVBLPWNLZTvfuAVBuMXg6bmh14hWfRqVAhTFU8yaf
dnX5YtADQ4LOx4hrNyk72kOY/qmPLSxhGtgFGoebEPdQIwhk1rX+vPfNaI8j4OwcZ73QW7FoqsQX
IqF1dmWe+i9LhTeXQM42w8WNKs9vNyl6RtrP/p+MeCSpLp7sZJAUYqccu57Ssh3HaRT5fpJRg3Qa
xbphpXdZLP/uXX9q3In0sn4uMU+8TH4/1DPGl6triZo0C2LB0Aiq6d1tT1yMU7RoT3lsbb0d2V1d
7t6utxmveqAwFBoZ9sfzDs0T62qWsdQC0k7i0MZqSFFkqinKrsmRcqoOpwV8eLkwTs6Nb3U/eLo5
YuOJOOBr/hYEIG6XfPIrgDOnlMhys8pd1uv4tfJyn/xtnMWMQ2x5AweBQK4Bg0DoFUgCajtMqWxY
OPpFmNtzeKdxfdNyp389TBGPh9K9HCZOa6S1NFAOaq0rb8ZWL+nANTumLF+xYfZ7EXFWKYmSXHAy
pHCjJakSijU38fRs+snUkf7BaOmwidgulNz1N4cYDuMQRk5T+iyJ3cagDyxSo6YYZC467bdhDLuf
cYqJGRaNtN8WPX17LDDt8oVZIQ/A95piY2wlpSRePVrvc6dKIXpEfZVl081bunhEEF9E+JmETt5b
YbalDM5a2F2nWNqXHrhwl/x5AO023yMISylYAcm8czYgAdwB+PA1Telfmx+6oQUuntYZJUObCirE
uvDXRfau8sPJLIx1DpvJzj8yT/oU+V4gl4dNMcZxzKNqMtDY5pR8vUe0sAIGYPpEjdh8Soa+3sfy
6mEb3SXFAiImSwuoAq8CYeXD2+AH/+J+W6sebs3bgfGdezbzzc4SeIsAP/b1MXJkr14phXAk2qod
F+E6+jZ7bWKEfa6cv+C9b1dFPSCts19Y2pb+c2ufFx4inqdbv3ypGAwXL995ZHQpsYuaE+oDZVjy
HcvLQmKmd2pkfqK7xHsXzJIEFMzzpHuHZ3++ssskmTcvSZfd/oZTeCg+BVJE6R47b+AKaMfmW9GR
ogFrSyziGlss4F9rdZFc5xSyPiSVTkbM6EC5fhGM7Ey4k9TTE93Bs1cXC5Fl6wdlpRpt8Gu+zKSl
BE459KPbHZEXIxO/giTS0+m+BT4rDywBq5o7VOsMl+I2pY26IB2LT60q113MNfPw/3xR6mIbvDcY
pHRdIUswtxEJXxZREMpQ+NxVXSOeXhtHXtDmzcaYOS+T5eZIyCpLBKuJcZv7QDy72z5/86VFZRQG
hWItbxM5tFMh/F2REH3RtNt9h8yggS0PQ6k1GpXh25JHWbmP41PpkpB9B034u6RND6doCN+YHGHb
78C5wf7ffbwUMYx3E1624NH/ZjivyBj0l7pGjGwsZ4QHRLiMFiHYmixqMB70gE/EpzXcrCJ5KhU5
GFIelTR10xA4XcXR2fCrCpO1iqn99hMd2gCKYiDKmajiNj4TDGcEwGpHX8sEHFw0hvt0ia8Vw+4O
OFdXZuxeMlTa9VCImf0wo0bwkw9IaWJ3flnAUP9GH9Md7P2I1dBxJcC/PU8IQdHDXuIvboFyvNwa
/mFQHiz9SKdCv5f8NNGJMvhO4ITYSAdF146fYssi+zr0sI6Lo8A81aPryzUtC2cYW2B+zeWYgzYP
Nur0vAypkKOvM17Ef4MlIsQgSpXHUXNp0+PIOk9czY6QBNDGNsaLEUAUet+z5lztT6ioAzCAo4Ku
ZEezxEzo68y17qBhVAB4zmYfmTrCW+LJHQeeDRVlBICtISeE7xUQ6lscLN8NGM8C5n1PdVRY5WVr
uaDkU64KAEmb7Wo7qwRrSzGqad8abVT/z31e2VIdtDY7WA+iX1lyIpwvpfGOcHZd8wQo1wPnZeh/
nHRvI4/APE/tXBIay1itEGVUX7S/0fTslrckH3M71jHBFy4LGYahJuZ8txAmHVqqNMaciTwMjdwB
lFPJUeI9uG9Sge9pHAv5yNzucHSoMs9N0Y4IEuk1oY909yU6djPreUjGWCW+1V6b6yMR+SiPAsrO
oZIuA84HTe7C7FmUM+7VoI19+ufcelA3C33oZP//XFg7mbO0f7IYBG0TMEgF03zzYBjrePcWS0gJ
5ipNY5GmNAACrgrXL+8aM7nmdbuB4zv1lTdeNcaoqetKPBvVvN8snZhaAL+LPuW21wOtM4hJFWoK
R8+UuK3D3ChOhEO1ymGOfmAKlfkeaLg23dEdmM/8P6IOI0IAZM4NAeZxRzNMYUC9yr8zFdJMjPcn
mYJTDowNE4ZMwgrlYd3hc2zes4u4q7NmStP9ZF08Bw9RS4Pw+vkwuAgRCtRkS9Jlz/OiA+3LEAnA
ffJJCe1CVFjV1yt1I70VwJRzyxDlOC5H5sj+q3kyErPyFiVznhShtHRcuw/qn4zw1lNllJcIK1BF
NTzo7TolMLQ2g90NE66YcsTgKmRLOkEXrlPYMe6Vbe87dj7+zy63SEaxyd+QeIFie3I2YcJdV0XP
sZT/kECIDhGBU/Dg2YTKd7K2inS3ivJ1d2SUJpEyrX25K4IDEiLcZgfZKSxjHJ7331aCxblnqQKq
0p2aL5MNgUdSETfpv9Zvwsn5YWDGN/LqRNxs59/DeSDRh12p3shKPLwuZf4hh0oCFCp/K8KRVd+i
N8zk8jdahb9HFhvG9yQPcjttggi7yCwtvf2YAK8JJEw174AVhxPyQKnqa4pYRtx4vJXHepbsKMxT
xUfgY7YdNI0B7/pFHX+YHxZZo3YoK0+mGl53dqDLJz2MU+V0f5/N4ZgG4t7awFOvUJoex3OKH73O
NlUK/xNBBh8HY+e8FgnadhQmzogqm5ST6Mxqyr/AQjOHEcTIMXj7yMudP3gzuBnqdi0zR9mm4aYC
eJSDCDf+jWD7xGKChbaTbD1LB8vwr8aNpfKYLEgq6bPBxo/FLrmc/wK6gcJOZwYRdlSygucp/mwJ
QqZ1nVWgVC0Zv4VMilGYxezy9F3rDSnLQXDy7EwNckhff1Lee+QwpGv/MZNMzyQ8JOWv23SjiIsn
WRQl+W021ZHwnlffrCYoWgsZt6UxdyNGGs6PW91lFmGNM5eZJIWUMk3qMZzw00sg9o2q6LmQUiat
glJ1Ca1g2i3kESzYyEvVHkVNKusL4FILoJbYtIL0Jhm/wOdFGlkhkwJh7pgtvdB5+flhApNC0Kan
exuisMKmzG6+dMYxqu3rNNICYmSmE84XllnvfuirSWVoR8270xFLWOFynwjlYFLGYaLT4HscgqD5
Q6rGL3zKVDX2u5T7sEc2V60k2ciEJE/gIjwdja3PpOGWjwAeTJ/hKaF+5BUgV92mz55L5+L0QYAt
j/x/e4zwzbIaAng67CUxJd6S22FihOcAuMkxtte6xfX3vtB2tmMxbiQdugcnDwfRV+wLM0DARXBh
AVwbfODpWLCGd9Ep9enhG/HFJpO/1oDVIbqZoGpU87tWbOhR1PnE4fuUhoqpDyannuvAw44u74VX
GFHBai2JaUKnk0NMiirlN+zG7kr4LWKWNNuG2G3fxZHB3M3xCwQD1EcQFwtBjcnT+JcHYewGszZx
YJ0nJHtPUcSHsBQcAhOmZ3lsh00jLlAvOrl259j9aYprt/UgQU+fEOhXvobkcqHi55LLs24URmPw
R2HHx10fFERYaP0mC8D5SIQAKIrvVO9vtlXOvZfHSFWUc5oTFCz+4QFC/uGZGTx3DiyaWSj0+eG7
p8/9OqmV+A9SlHpAvGxUH/WnhERLNGtwMCHXfN/T4RW5l2/YUr+5Yjw56wOuRlJZJuTwyZwogzx/
PCE+vI/NQ12MDlG9rq3CyTTZTHbRJ7o3vY9SETlC/2vl9i3rG49LtXQzQmjngbjxHO85qruLuO/o
WoUQ3/k4Eh8CcnYTASEYzAy2mwJNv0W7LDVPmpHmNf+iS5lcbsfyfUD4sDcPBtOmRqs6/doroppO
zfHM+UkD7+KPLIxAVAFCMVI/JcZd10YYeb9cgyIXLGE6mmSlb4MXBauoMQ0mAZdoaK02UCami27o
0Od/+R3fZVVHHOfmCqf+PW2u2bC8aJlt4RfVYa6NT3GHkf11qAdd742mo5zDcEaCWt2BEIT9V1VN
4qiE0FfMqJwyurFe9/jnbhvA2s0gI8Y2PHDIZVTzvD/HcMZRLeaIaNfZSr/sq0llr2vbbSBgWgQ3
oBJ31tSBoczrhnYZBhKfkboyK7ejDaXRq4l0PXI0lUyyBvOsRydRuzbeQNaBEJyYVSQIvu1H11/A
fjbmpi0xhPpecv5QQ0RiYWdGQ5LbidiNp4LJeySO2oV0IyLIoGBxmzsyRfaDBQJS2MHTF1iCGRJk
/7+0oAmXHz8sLpIRGDpblor8tpUfLpuErFFvEaxdhdobwVd4dbuk6EyY+HIJekkAICb+eFqxisuM
SJ1UYkH8pHbFfAdZ+j5YHSvhcf+zNrsG2DFCdc0hpuQYZMjsSh2H7d3+mcIUT5QgDpugWYdmZZCf
ovZNFS92jEinD2KtQfojw3Do/q+6N9AnzgJn1RMomWfA+oXzz/42cl6VEjH6EpxDYE+Q0CwrN543
m7dNA2XkpI0yzNKXQYotZiIbb7LikHWzrBBf1/L3DtfXVGr4ye99OOUBSQ9tCc/Alo41tzqNzxHd
bd8XA9tq8RqfoizO31rU/d8esd9VBbam8k/4TrP0fHd22lIqmDmvKDVJ2czva9hCJ2mTSF+P5ONu
Kp/ur10poB3buc8h199AlGo7rbNRlB3qdid+kyfaYAyw5bFMRdOl37uH9x7f+eRnnH1vLI8c2uZt
l+27dStTczM7/9QMmzhd8Pskg8yeCnU2ch5qEThpsn/ycgAcmavvh1/mWuH8A83rfpqDsHBdCA/N
BajwV0THhOWQ+Ee5DDj7McU48RqhnVfABs97UYz4GMVN3E1Z+4LBYczQpusMGRWqyeCns2H+sR1G
s1EHV1YcI9RkX9jBiwvwuef6INuByxu9ipwxk/f/Ysgc5DCt1CnrySbgGDbXiTdLaS4ToaEPiwLs
o/Qy8el5hzzuNzyirzLMcy1Jj07nVQkY1sYBqPHkH2cx9/fsCP76t+xwg6sZqcLeYgA5dl9L0tnY
Lo0VR4N4UNcx0v1fKDQq/gqxSMBs4glh5zBnNCKIKBoYQu3rDbSiowAvyrABwPO211ZQC93YMjIS
iCCcErK7f2RKxFeh0Sflj0x/S7NrKkRGSZ9X1HwE9obusAqOlfkygiVdvktZGGt7TIif6pEO9G6g
v/WVp6tmsI6H0KApdbakdCZNsreETnWwhQRb3/YzSSe/K4L4dhjw/EVQ2YwtGcDeuN+CQUU39rsb
cjLkZyTPmiWMXQkQrs5J3F0k3vahogGCGkv8+vpDBCG4gfxsHyrOBSbKdmXl62ZmOZOyrq0IHAJq
Cxsnf5AhUidmLUeeV7kPkWkdFejtY3an57uhYAe3T48FDIXAYtKJIAZT45+wwkBAowZBQVQeRHDf
QFeVQNAYNkW2ZkOemkSugBcvyvxDvSuDFjW+N8cLeF5bK0PcaK1TpO/+TZXPM82NNqbAX0u/gmzO
QlqM7e86B6tt4ehL+RThKhabuDOOW6FZNcKWJkbYG95ikI2IFJspGZ6h0W+gdsa2r0fXCQfY/+mq
0/wa8IND4mxJDMPAWuMgiFF4JU99UIpqF4TZIzaE6xAbgGu0SaJhFXQE07x5IVvoD4Z0tUfT8mfA
VbMkeMjGnKybifPAwC8H+3XRRWwQ5hgmInT2WT0bSKoiccEOCzkbB7YKsGJMGlA8N42jwDY267LC
pGO6dV+Vv8q11/TdE36uSNKiJggnVsMdFSChhz8jkSJGbDyV40i3KwhjVxQ9cJ+FSdCb7YVe/jL6
0qut5l6fHMBOCC9dJYYrE6yQMQzelyyBm/ePm6MLhP1Abga5DVj+4MbHGRRlqLMnVEj4Im58SY6H
huVzXxGSx2TbkufUD//EsR4i85SfmCXL0aKLKIYBit/q0zkYf7Hm5Wb4zmXd3B9Oa7wZ3XSHIq7m
O1oniIlRbDJcOIgwcAwlPqtwDyhdrfxcOVQHrTOmOBOxh4sM7DVXMni5wA0rdNSQ20/FQG39SI9J
ciQxbDYAVr1Y08vUb2YIEAHbAFns5ylsWpNueV9vWPWv/+mkBIZoAKdYxlbtW4+4pZuIcWLCnA4I
uk1OWdoix/bD3QC9swj0o/5e1thhN1nIMMOgpaT56vLwoDydbW6e2g4SWZ4sRjS71p6pXIn1TaEY
2BodDQnf8so6AG33KdCzkzFyNX98mXlOlAfXPq+h4Oit20XXRDij29sO62pzs+lu7uQ45exe75zB
XeLwoLbB+b7h3G3Bopu3KKzVnS88pUknQUZUTxoyCHO+AfBJwN31nLpjI3ES8AZNgbJfCwfSI2KX
vktb5yNkbtxoSGbNwIQux+TAuKQYjgSK2V5PwUwM+LWUZqKYcSDJPLIBMdgi1bqKzRyORfa0qw3l
2mFhS/mOqXiyZXVOwavrSQBJ9Xe8FhD21ki1Z6Yiw8G8Q1/8Ud6jRINttMqps2mm0PQkOv4JYtOC
ZrDnIU+jDQtRTHveuEpUYXW49JWDwepAQSE9osW+aRrFNYzqR4KrJZGkSSqRPaL8PPUewGyOvB8R
/j3vyhT1EqHAHjrz53rKQtdozZiIrJY7Q6/3Eq7WRv8iSiGB7c/jns6yTk1ALP6xj3mueD7dIOiq
D87x5DhhWwXfq2hHNDz8/2rwr6ZP7XvnYGAHFA/tlztpCpKyTGQ4/62H6QkeiWZs9LppcxcjUzcc
w/nsBCMB2Rwyr7wzmWSBjy8cLIOj2WJB8s2iU/oCk3D9A7+6m1DXH4ao+RNiXx7zxBrAhtqJedMA
T6glxI/Qh17raINJFA4UD0It7Bnm5TBEJjclfeP8ROSlIeBfPlwea4W4pUEQYWC3xAWPh+PSMC4Q
HillRGXNFqejJsA4jgYkkMJUkYsMfUvqhchoBfkjiAKuy98U6xx6M22RNG5w4lvOLU8kpwdlI6yz
4JFqSNQnI2cSHxUZir5V7R/IAvQm3LSjSlPyOMiivLUayUV9xxnk2VhAhNWoczYMlymdcN3CEeUr
KkgCg9Ro2uJhXNBHQgDPJRjzFrlYoJctblryxopwvy5efva7XV3Ee4XG6BM/vRfhQxXaEbfOabu0
858ow8rhSI5gAwIMEL4342XNsIlsJDIKQwCLOIhuWx/fA0jUb7oPE1t2z40Q6vDGnCE+hkUbPFIp
XL32EOH9zmJuHYmKX+QA0WRF5mu0jIvMDBNEDb5ipfn9z/PjxOu22/NGz2rENGz2EGV77CPsN2j3
zT7UjWfLxX2yEiWihr3WUnAFiDbRdgdGPmwQHSpwNMTLXOh6aImm+xFAXcmCJYGntkqeGjx/Mya6
OkO1t9mUHmFm/f8Nj+xWybxVlr0xWsCa58xE1SZzDFyV5t7PUnKRYo40/rnv+ytO6g2am0x3J0jl
b1rASy/tDMQa4N6cpbWGdpgQ//vLYqe0BfcLgoFqKkgcObLXTUoLjglt1X5wIHZNrGTpqIMIcos6
MN5Rz+QF7YdhDQ4g2fBeLgWFSuDknpcJ+DJ9/tbor31w4SkMrvUSbtSap5adhPOXrIHGpSDlxhWa
JC76jYL7j1RoNnZe6totSAQDHT7nq00/dpG4fHVmJkN9aFPJv+exYTdcR0pl7DTdn5aAsMkaYxqs
8jg7HlSzGt9dbFazbidpzXJD/sRp/KF0c1q4xyzVgy4D6M4a06ISzPe5uRXrRG8TQIPyxQd8WDWk
5ZQFqem1QaSE8QUZHemXS/1S+moiaor757LNWqcf/BYLtp70SVuUQB7X4+irHR/VzJcrmJY9TqIe
Uxw8B8v5NN14l4i3Z/UKjJiTldzgC+ewc0+y/sfYm/JhijHe+0TP6aHTaB5jWIHxDHlmhNvNi+Yu
BsHyBcdDq9A8HO3ULFGCoA67fuubSlkSBQPBJ1JVHS9ZaeeYwVae8ruZV/Zsx/OKzoVj5jYgNIdi
Cr+Ef6TUihy2WXSlcpuxtDbtceaKncA3Qc2qRzetyhPCeX1xhclvTCBUqfm5kRKqSVmCu5UHXByz
/uBvq2N1E0ztPrUojW6YSMaOGjIZHLT4z+szkAdDPEynFuHegFiEFdCAG7k1wpLWRdFJWPDvhlKL
TIedbob5F8Fcyvc3tgmK+W7DblMlwjuSnm2WvWSTIpfJ3+sFFt0U2m3WjbAULqhb2sVbWGV/B052
LAMynk2YU5oGF/r6IEO2X5iE22cBgXsuwBYvvxQBDb5u1yHwRS2ntcNUPn2ROURLTODnZ0bOToKz
qqKiwGc2f4FgnT9IBph+XLXzf0K0rjsFXPuu7O1mUOfmSfyLivBAoqBOhWW80eWk15rUxrC+g9HN
c6638hkTeNAl1piOM9HMWSmMfHEA0PRiATtiOzBN5+yv9rzFRJhc2h58WlKd7m9y97ClMbRXKB9Z
DAmU6M54nXmUQYIp8QBmvnkV9haioFzi4CNJ+/rpLfbB0Vx6ZYkyxelGhJVPMIQMmtopUe7YTWuv
yyEFRoO4hytN8bGNvJ8tDe+3quRG/Mc2VuFyX8+CgvuKtNWaIluwzGRzKWCfHwj8+erbsoe420eS
4ukX44BJXtRpd0bDjPNxw2mtQaF6ZIPH7A+ieUouSWB2xt0KFAx3a7VhsEoXWDVBn68Xa/x9WXrJ
FDQOEFn71X5ZknwugVBOwZXmazKCcWcIXYBVmRHt5JbFWEJ8qBR1ljH+QqZMM+ajGxUO8//kMwfk
w7pJAwCjn9295mugmZ3C5WfvOUxvr8iTOjTUY89ig9ZK2aE+/PaOFxW+I5RsaWC2Zn2ph6Awa4pR
qcMnyNX7l3FHYjlXHWWIkJwRVYeCWXetAKRm9YvJGUYUw2fZtJCCALW8z4ad3icxSnUTRicYy5yT
TET/yY5/uKoCeJ2fi5oYCYRvc7ZppzT9Q1HZt7gK7JNBAAqTmUpzzRLKfbKywSeTatvcE1bKE9AE
ZsBvrm8ydOlmC4hOYEm3HIlI2uvQiYsYlunYkOogD+fPm2xgnqSSKOTGRl5kZnXGMNvsEd6mZQUc
XOUy5nvb3ZpksMnYg2H+RC3/1pqQ4y71G9AcxSJBWgYBy/vqBd90fdYy0Ry4VC2swzN8elzb+RZ6
SN/FTqzsPGZzfJ1elcr5PxFRzAc4I2YaGEQxs9qP7/S9M+h9UprQDs3d2eoB3ovwl4p9+VzfdLZW
E7/LMfH4OJIrhUYt35CxtR+2ZI2jKIzOw9N4njjcDA5akh2SC1p0yDbzHp+yX5Xu9qOFhtDn6tBe
VPDPlOY51myrevpgs/EFN8Z3fa8qmaX7yEPz2eHccraSDhtnjdOwMaiaaqHAa/G6iyU3Ls33Ib+L
b2qpjJxuGcnLvgLIzFWjDEBB2Oh9iSu5Rti2hexbFmRVIllDn1z1DtSalZ6zJCGGGlk18C4st6x/
pBu5SBqhLbbdECiPLxjwQHEXnH/4AAKp+PG0cF+FpHlX6LX28w6X/6Fmt7NzH7Bgk6DhvTRCvmi6
4mrgFAhmLN31F+UionpAzlx7Hdx6ejGK3s9Tz0yIDITDqTANL87lLPU6DC2Ynbm74CZkOxeIU5kJ
0rU6JnzdsjPhXkRdP0NkvnOQj01Q8K+7zE6GtdOP8CJMLs760w2yUYthsygIF2uppcHnsBV/5FTT
LNUuMbLYcwXIb7VsXGnBWPA5f88KSoeKWzP5WDcQRfb4PrX1K0RJOhzsFpFjOORlYEHng0HwI0UW
MiPY2XKfjIDdnpD6N5HCcLzXIKYkyIrXlk4Bh5E052UuvPUV1os4QEPFjEr6eCPxjR7UMdl2VA0Q
QvTeAQ9MV7iFAnB215hzyDLfJVU7lcMgQXg4j+FwHVnMUsmx2UkFv8GXOU8thfqtwjrw0/owOclU
VDNAKm+w8+rKrw/4WGD/aHWqZegdEmY2/FyfFlu3tKatd2N+zaKZGMJfdMvuTBGyZARCmCgjMoXQ
8k8XisE580UUuBJcUtfiTD8s92D/YBm/5rr4Sa6p/d/6D8jEW6UqCDs8JcnijXnZMnDSXSN4iEiQ
jjvtOnBGToj33c17fX7A+PLoQIjk6K3rNPq0bEqPnX1wsFtYZudNAcAgDfg/us68xxOEL4xhXTD/
ZfMZIoqk+SGmFT7Lv3p/MwU2YRjcjFBPQP5RDFVz3Soq/WnfYCRHzmhKRXlVhtbc7xIfhSJhhyxo
ShIfr0iG/7tmi4hxw9B4Q/M+DIr5fmjGbBk/DDFEeGg+M9KvL87H2ZmAB7vixjc4mLsQYhHhmhWf
AofRxnqb3kaj77n61paq/WaGlvUR0sosljiUZvoQAVGGeisYPL8XnwZ+sNFh5UWGRrWEtr7TL/jW
HPvi4tdfpQViLoYlD7fRiqf1OtJrwlTvAEJjkmhTYd/k+oA6HIlXhys9/GsW0amxUu8XaZPaj5oQ
OO1WMD4NW+3L7ssmTRyVlob6BXAhaEa27BXEekrPwxiS4tJGRxkcMDRrDV8bU7//rgbX9VL3C+qy
OPmVwt2/a6L1oUBhrkseTqpLGD/e8TQ240kIkikwb51mjqQuTA+NSkEhdtUUfvwPmSIKM+MyvM+/
//eA4YNrfd5I+p3Asn+fmjPFFbRvT7u6ZqyVj6YNffxVTz1GbOJWjxgQ4ond8YGGbYxel0bfxOKQ
/9glDEykdc+X/lmMYAMs367/KzWe1rzkAgqtnJJQubVGUmNycdKNdljClAex9xSsaQjip3h79MUR
B2ncEWMHyx6/HOSOWyXZBF7evFkk/VogqL5ZI8WHqSBKllmX9NzlBY7qT5WTR65ukFTU3k36Bfui
qCqERe34/ZfeiPnyJ4JxvQW7M1GPmrPQohKy/ycliCzC1q1Wh+OeLcdMMuU8ebdHq2adl6F88yW4
b33cGS8k2pyPch9k9MT3PofmLjiThrbHJD2UtTsbUmDfjM5AhkTr8+qzZB7BtmwA1oR8N6lIkYTx
/53x7URn/Znjwubf/B8tQHclV6JKvCNy5hRItVEZYn1b6VX5+60JN5YGK56din4q/mM7aKTPjTXh
QEWQPC4P2K9/4c7P1Np4oYUS61Za7Fg8Ic0b1zslI/+qi6QHVQY6eixXFiUj54vLHx1jXvKezl6P
edSxgiu46pc+3oEiMjLwzzOwsLRulejEmkrdK1SFzPnlfJf7zNBILFY9tNtrT2dcpExe9wHxYIfl
TB6jevBrez4wA7N1/ANt+RH9x4qGh8wMYEokgdEAtUFf5ESYZnVyHHmxxW9+g6A2YCzHYFz6pO7j
KxVMx0gppR+SkmUYzUeCbM3EJg+lKdw+ikFh4x9F4b5lrkZviq+JAMUS+4GnnzzCWrIXwI8HjP/5
AODTCTDUPUIyJudFKtwnF4XuTgh+ogpszzWpadZEAAy+cXRVYe9XfCtCxC5BpzodMGHZty/Ujm8N
YYlDmtq3hALBadzCN9wkeLgaL0QzWbR11xUo52JktIkQr4praHmERlcoeHUkTHPK9sSQIUIpNvHh
jpT6ijCtIUItV1eG3/LRiZyQYAOon0UiGagiVcUlV2msHZcLas3xdyNjvWyi6i5+O6seb2K4h4as
99NdUJj/Dg2qUXnGg6gp9Kb0QcIRjHfthPWrJoo8doK2SoXK0z+3mO32rNwArxHe2ZQPut/FfxEZ
+cZlN5UiCCeI7yRxqWYXv8iSQNSUdeRpg2xd2NfrNto3ZE3CWnCaZUxs7S1btZpo2dxSeGbDpmdV
dsPfKZrSedAov6mRubwD283+uWiRvX1QKvJBkVRJSiLL/SpgPpQpwNBQI9MXOgHy7nzWSfiZQ4ul
IQACwGz4bua09dWSB12WFZawav68kda4fpiWlFkHxnOyxZZfH4PcjKq2WsjP+Bn5HeJh1isAziYu
d40WRHf/SavMcQQOVa49PaJ5Q7l9zFxxpN5dM5K9ezzcFRPUdOYaIs1D3I95qiPVM11amPEsDkC6
U6JQ2zvLV7QJ0x1gTs8hpdrchb+RhEcyH/EUdduR911Kb0eIZvzhZIR5xj3Kxg6MXFeijuq9hiaq
BZCKy9zk5F8KL54HfucEryJmXywLv4Mc3/G0jdORWoPXS9Wci9JYxuHLkevFJRX28Jzi/6lQwKl3
KV22rGPWY2MxOoTVa2ahG9FebIfjtJZWg2V6ytPCIS652EnWq0dCrmFWuQ7+GziEalnaIeX5cZUQ
Lwv1qZb+ohRjK6D6eonASdWrDFj4dA40kBVjwtHL3VgN2wFzbfgh3uh5TNU/joEiMjsIpfUdwllk
6wB//r0+dYujN1lwNJIN5M4Hnd8PlO8vjP1dyowLldv3WCX+HJJd5nlRBAbdwL+0Mfu7vvejvz2V
dZy07nL7SVEMrhYFRHPCu8EFpHEys32zbpe9OsmMu6iGi9wY0XTljQZ4wsYeZYvfqFX4Sg1g2Jxq
5czrPHDxh1N1NtX9A4a/Ind9FMCbIk0Wiv4jDG/lHPLOe6r2C0P14JtrKqLA7nEBoTK/inz7EOTR
6Xt8JBWtewQPEjFwnxc5a4w9tmf2q5KpoNJCO/XKHXP7bTKAm/uwS3oShDbj1dPCoine5vfmjCvd
MUNxMQAHqdr8CjBRv8Zx2aC4rwefiSZLoTtP8quY9QtfHUv4kzbimWfaT7rb+49hM2G1/El+u0Fb
Hc06bQzH9sExN7I56vAI90U6QcLzXiCrcv6Ved0juLKKsUtAR2aF6MEWs5J2RFozCNSKHS/Hxph+
umoSp09HgHEd31cZuFsjFg/nC2rHFhIaySZhk7h/x9CocWAPaRvQtN+iZW+yk2CfI8BtqAZ5KmdE
TUQJiiuyUOCl3n5HI8jJ6VZvup144h1obs2+aBVOCE93CkNhT1vvNDLJFBtY6IfajXdZ10dKYB3t
WDdTogyqgJMt5oE6W6LQNYkU0K/MpGaDwqazRF7ui3EcV+7NqOyhXSbQIsfgH+a2Ybq5lTg2cfC5
Px6GnapQIoeQ1tUzA88qjKsmu2c+cvkx74pQ6KO4OEFa8bi4T6PvfBHVlI3Tj93zLIEX+t1sRPoO
WnfcitC9cvqG6oHYhfYDjRaCVZUw63tOWSaKDWyYyxxC76EYHcTHavoHZlMPv19SSAhYzLMKfQB3
dENNmsHH1y3L51dDBv2MbinMRwf2ssRPlYvHauas0Y+jufcyak7YSkwHhowVYkvqCUwJlFawmcai
HjRrrU9bgDoWhfiyLWBiYdrBqBuS0Ov+KcU2fEA8QXyowK5Kl85rlRqZxSlbC5QWMBC73pMiihIn
QFM/Bcx+Sl/aN8VNXMBoeKkzCVDmEOPwrd4Aj/oX1NFRXQHKiDvAbvF9PBh9wm8sAbeV7gjN8WfF
dlQOHjHGvOQ6k6fE7Rwb+FN+U4nSzALQVzIGPS10wNYatupVI78PFqSqhKYpWErNDLAzRxSGBOeq
/Sw8QoAK+utDxVc4DAfx2R/76zF8sLLvGl5739JtMEN71KUGNuS1+hawofEGPAsH2zCSVMDxHHmT
8AxpqkbAeMoGb6G4LnKgoUXhLgji/qgnmwQMOGikRB49ncP/CaYJLMPSycGnpphB8TpaPT+eIM7a
S6uMhi1v4o3qd01ZnfkBbb84yiijxSm6YsxEueTq4QM/50RX9+o+8Gc2nCX8e/R6qAxfWhYlvlX+
zIvP5T+Pcd8NTeizX6y47HdjRLlufS45OqegDPRr2EeBchq2nrELeYQH2dktEhAh6dmrQTMfjJbY
ZFhOUznpmqSq0fZ9zUrlqv6O8ikf74H0iGe13OA7Ktno/Ud3hXsmVPIgpMOnqlbmMQtYpHcHbWqZ
rNpuxykAvfGWwZQnjpuwAo6pYzPEPeIIgK96WzRhj4nB+zBPsMYgZXsgFTTCFRIyrW9ihZ087GM1
zQoF5z3sBtfhGh4LOS4gx/KCEku1cnmfPQ2KnLdvnBvrYtof1R7mc/mVwthS/80QYeeeDIEyShEd
OIneHK13nlrBKXJzQfjb+AUSGggK68y0L0dq3982IKpbH/yQ59vUuNloYLtXCz3jxC8ixe9/HeZ8
5/yrNl2HrYUVnZUzv9ahp1VtxLzRKAAtqE6weoUOTkHEPB1lACrq8iRJ3DzdNzwgOzqZknX5NSK2
59wWUI7zb+ez7+sd+WYvPu30IaxpLEeiVPiRbzBA1AUtUQF+oYifXlF6J3zJAygpXsjiy2B63/GU
ThZ6qyJoeKAs+WOH1Q7juy1soJ61Av+7cCII+dXF4HI2tsxzT2jx8HHb+OkJS+y82tHkqdaghsDb
nuGm41Rvj5Zzp5iSxyJM2Eh6x/ZjwXs0yYH47ZolgZrcLsMoqe8qHsju+hQZWg7XyJKyH49LCyI2
Vh7etBCxh8kH1VCvkeZTc5oSwoS9tCXke7MlS8FCGgmBhbW3yLHQrtnlcRR5Y5v5k1oXf4eH/UG5
oCAfUPWnhRwmgFQDIo5jVgBzYJuioeESk2SpFczaLjshwWKkMsMWxq3vNmcN4TCZwksNG5We2ro0
IAECprrEctapHQkcG1UEfukI3Y8rRWPxy72Q3yXQED7CWDd5sxjswvwnpx68bD5EAkAUxfaor2gC
xTe4uiFJ1+FdDhch7/41iQ+53kS3QWi8SIzlB44CJOHPhJ7u8FL6BoCeQDFrtO3LHuHI+8mr16Na
1cOZdhB0xFBbcDdG1R2unkozdiWDbhBDbkNig2d7wMmWB4nGZ/dE0OP/X6eWCE6bZKshn8WNvxJZ
eKV3ie2yEc4QjQr1KXNTAxN+kb2Jr6Pl/b4nA347PnggyNrDz31AaN58O41NmVf9TK+Z2i54lgmT
QvctDHM7sfG4lhWRPg6BgDbCREIA6JZ9a/Nu4Z1MMuMk5S3A0tCavijECQAY2J0i15rZEapu/Ryl
yasUvqZEG53ZRNRmrhkjt7mPYC9gbVGb6jlFWNUOVTNc6Ra2P6J1YSdd6nzbj5KaVG65tmJ3WdKF
6bDGiMqzbR7KfHJrEpleG4FCTEXvWO1qmgr65ZsD9ds1XACdpZqIbaVq2vZT70+548JOvQe5Yv0K
oOdpMjyrQi4X04NRxaXlyk8RdVliZypQqiffP9BMqvJ8VWfKKEKYUrXx4W32ebmHYjCNTJEkFdOu
3tjSLHRNwmHzVWbdPdho4fco3d7lrjOgh0SHypy6Ug5Q3g1Cn5uJI81KcyMlj35g0J81eJ0DWxQN
aJqgWjMZQkHMAAiskkfaIfzyYDRJJh3hdP4xaGRvNbCodghqvC/0XIzaWYlUJhG75W0yt0ePj5JF
dChn4SrFyH8wF2q/9pgYwj3YztDu9bIZQ20EVfP3hRV7lNzWso9JYnt72PfpKTKqH5DLD1jCNmhS
Cjt0XhVxLxTWoYS8FCXm+0EKiiOUrI3f43Lu7lPhLIr8h8+cGEjcf9wkfwBxkwSFKPvhJPXrXmqC
BRkPWKu6a7rl7Uuxh89dSj8JM3Y+9Aj2cy9onduGNrP6V0LQpKvU6qbcElzHlwri1PCMpYyWt2SC
Qfpl72aNxAYT2wAV01mQAGzBLuFAyW355CC8ih/7j6p8ZM/3VPoOikd3FuG6l2Z0Jt8VAl4Sr9lM
ZDu+58SM5fqHNtOWoQmQ1PQ/nZ94IzEN8MQNkm1xOrP4HJJdfmOQ5MxDjLd+Wdrp2Tc8ILvG3+3G
GPdBeN6jDQnvUvsJXlOEw1ePjfyzDOsHyp1OgQS3qSotUAyLU4ODJXhWrR7aMPEKu779gyxdeBlZ
24mv7QYDIMdwe6sh0uL/OClamveNe8TibzxysYvJGwYbKIlvCzaWp5MaA4EBUy6OA+2A0tFt0Eus
LKN+fe8kMemqb0dp1LmVxoapkymd/+zJ5Aju8stBF141guLbwljm1qkUrNnqPWdu2xZQrDNZH8fZ
1ATGts4YaE1Fir68IRBYgt1fJKarI/dZzFxjjdCLvzEf8L2TVyYMGi1KGftmCV+Ux+SfC6HAEx9D
MVHHJC7p9SYKCA0BZxVN9AXnIsqJ0bq92BuFNcjODb9A5rQXDcCHGMmvPlS8H+cCBiy1yxdhfHtZ
IeA8YJDeyA/iddiH6AL2TsagVMpWRwVGagJQ8eS3eKafFcfoBSmgT+jYWAXxCuB6l04Qkxv2oYmT
MO4qMk1AzJnmQMcifIqR2TlmmMAaYw++cSu4K2AE/ion6Jt5Am0GU2cNJO2M5vxzznE8LxBXsEqV
UEssf0D06wqJsS0y3brk6sdF4XtKu5px+kxWRnfaWqtznrA4gAG2wnnv3sSLmQ5tDIkhzDVs8Ocr
VTjrCJQKF1UMDdXjEzsLWL08qI+TWH5WrOztkramh/TwZU+cimW0iUcqNY44uapHwTkBPcHOi4C6
nPXhj5qp3NZqhSYWwbxLtexcyj4WJeX+FGwhippiI3prnborMKvesf0hlvf5ofKhd6h1lsgGgQtV
IXQGDbR2MbPmLTcxTmL+U4h5VrMMTMaTf0ZrH65wpb2XG3M7hNGu96SnPQfJJX1ZofKfunflYPIF
E+YM3U8bskLePMNMuJdZ8LGflICAx6+LqZunqz73W2aO3gpkgFnwOVUmXxGV/Al/vGxourwOlUHP
hRp+689Rqcjlq6PFr8XAlj4CRQaDjFtrExPn41shscdbi2qrBZIQXg+LriMW/1nkF+vHcQJ59I3V
DZcWe2KNyzw2uHeYXVvtAajU02jzBDrwmo8fwfoyuSzsncFEW19+0llWR2sZatW5jAzQqdB3Fps1
OdZGcY4cedvj5Ffh/YVdwH8Wt4xtr2K6sTdq5DESQ06n5bjFxHDHQ1GB/wYroZS9bAkDv1doJzv2
7BSd+b8vm8w7MvmFB0bYAZMM3PP0gxPF5dl2xV9WLrZ47fajiCUmviV2bmCNb76tbKP0hnDjVnWr
adtfkt1BaGEiq2XgzrC3kRIdq+HV+ags6y+BQN02MH7SZDLIuwlv+zlwUHHiGig4x0a5vf1zMme/
tT1WAJ7TVlOoLwBoV8CHXKkH6ZzbBI/7YxxsjiLNf9k5m0ig+wllH2QfzUeeSx3Fqgqi2/+qLzpP
F5db9464IGv+Zp03+wzpHPkXd+DstkUYbGDQQ0ZS7DizqJYyEkdfSSgbfi+6g1mPdvrHMxVTbCD6
VZ+xlTvjjo0U6rI5qrEfMvGifYzUwbpXkq9LGKecefkaDOHYupeV3D4Z2pm0kJmuzkT9EVV9X4Q+
xKnv4g95T+afouBULdMZ4IOJLMhVtiz7OY4DjVoFqPVrrgQRqJ52K6l2aMAoGnwdaq8Iz52zpDN+
FwFNFOoANCIxzMlmiGkVfd042s/wshMjYsnGzOhSzq2+
`protect end_protected
