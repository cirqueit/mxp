`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12176)
`protect data_block
sXYm3pHOo5KvXIQ6qKRDK3zEASr556jSdZPWXo5Kl3TwArKvR38O2yLrayP+icUShCypT4xi0RYM
Zu27RWOvlp23Ywc/Q4EWMpkgwNu5vYl6KXSH/zLuqcxEZBRhKS2LJvI3oq58m/fi7ImqcCO7d1lq
6icRctqBfXEaEaN4YFHQcAGGGYVx5rMFLrMqP2YjnkZB4k9BxSAq8yq5iRVfK314OLeODmulQWJF
Ebkzee1TyP3Hz6H5dbnoqeJ8DM0NB7WLUwvp1x+nMTS1aZaf7GVFMEb+qODwVhp9HWchulUGobbz
mmWyFexRMJQ7hDxrY6C7BHvcq5Unxht/AS4rgBOCk6jHW1HMRVwy5ZoxPmXVhImFi8GZvqoZvUBF
H1CYXnt0nKevJrwKe5zIXxmfl7SmDnxB7eQLbgpCxXsFWo9p7j8t+qGvEQlQuPmkepjm5rSndI19
VL3xeXOh36oazWB0k2O167nxDAAgrt1HKYCpHhWiryvwbDV4cl7iDZYLxO98xEplytMrBZIZzI+p
InMBfmHuBbWKq3lNHUnTUYtRAyibLZA9WQpRqXd+LHSnU9bBVESdn9MNONpGroA+ikv/oTfMJN5f
WpbMSvZLPoYt6cBRX7FmutE1f6GQB/VHXU4I/Xq+Gvl6IMZwlZDfprbc4o0TR6WtnBevyXcZrf71
6zbZCc6FU//Ny1Y6yooaSVPRW3JIDTdMzz+LJy4vpFB2HGfrmYXJOzA+xrxWSQ+GIeTXGYYRob/x
+9UoGwtX8/8Pwt0Be9+jA/g/eyEo2SNjKpKcfuqhCRuUPMalC9KURxHpk+AgC8RMJb21Duimesgb
GIaaOIa8j/uvMTYG2SYQgqlfucFgebjozNcHIbL6NQvYl7fgbD1QKMqtHSO68k1j8Xl8M3RY2VN8
W1caEPPLNTf8+ZcHiSVeMy7Vya21eCfzSIXKpe6qNy7tIkVlXGhtl6EZe7qnV7PA9mGtzPzCIw6x
6iGZsSqB34TtTyJGboQhRbP6yJj2FBb6gSNUQyfPNVY3z/m/91j3cmHvj1eUCL7I6ANJjpvtky9d
eNe3zvpjgLw5TZjx5ohLIEYmA8mzwOYgkUjLQkqFVNzKgpKsBWKFG3pJsrCVAO9SgHHSigvgXzB5
VapkLKAwFf3PJeddfR4xh7T/XjT+5ZLNtinWynrTeQLvcJqxS7P6aBi111+DUgHtBmPg9ZotxYsC
rZKMYrx3CnLVb5E7g/lAhLjdU18+m5T+OPrv6EKGtj2+lmdGrLvhq+rLpNRBlMCSn+C/585wzh38
GfjyNtgMhqsdY9VE1ErJ2QHkUv4XowTYvhBBUkafEYVCLUcHwQV2XU2Oe4o5OAvrGgakLI/ycQVA
US/er3rdvkjJ2FphS7OUKaL28+feKMJNcWTIBwVUEQ4ZQmHF79HRAzC6eKCdhAL9/xdQYW5BMqV9
1olWHXsb2ls19o82mjyGSR1UtxOcOnp5YAJ21D4JJy1EN0Q/51E2iG9ZI+tLaG6oVO6PIPofUsda
50ejQaRIr+rQAG2jDWXQfmjqjIrpVWURkEnz19sLr7ctRqIAL4UjKimd4XOzAxXhl7k+v3OD+d+6
3u0YUo+g+Zul6yDdzdumb4S5rrImTNzlDAeodBbfUvkyYOnLvbuEQMUcsT7HtJLkubhU6UuM3fdL
vm2sQW4UZVAkLqnAxvhlYStQPOIZin4HQb4lRbRLAg+cjBgkt6NtEuBliZ7RUxbEcjiPUn80VM0i
B76M2R9R4t59b5YAvCbYz6TQE4qUPipRc1/oEVgIeXOwSqfj/26EOqy54yLYy0k/w9as0m/3xR67
8reqcQj+LaPpsCSysOYqAac14908p/9YA0jidSjcHIuN7rNJFu3kQ6eqO3DEbd7MJjcLy/QecEqa
5aNPPK4f4lwC3b7NhugKipObexnii0nxH1wPV2LmJ1V3382muCzeV4T81NH3Hgtwpmr4z1RWY2Cf
x4Rd5cHo9hNqYt9981bn/pUzIYVWL6HkJXnyJ8BlP/qBcLVWPyr+qja1g0d+OGFV8EEvlyGKvA1/
m/6y72d0EdTrFmbxjk4/z2TdgElXm3ioMu3sbdhrhmlIFzGFaTj2udPp/o1OxhmYVYrba159/alH
SVu0/guOhTgLPfOHYaQRprLKdiKf39Iq4dpz77/yfE7Af9ghNpsxoGUdk7o+4UWtnptMtf14Xpjo
85VdqD8ppnkvgScc5C7uA++otPmmC4b29LvzFLeNwMkl0bPfurLRiDOyJYl1V/5OYVduX3my5R0A
8+FoLTEftSnvu94NBR6CgKdZQPs+5hRNwBajaJwzPBh3i6CoDBBfM2ESwz2xN44x0CyKXPWC518P
UMyTulafcW2ghbtHPPSrddYuowexGYGSxZgsPXFtKHwZTxuzt4nnJTiqsKykumBmayQMuEhjBN/+
EsScnwzWoP3KNlPAtOq7Qp7es1rToGh5BHkn6SWnaVY1bDM4lYAnqghcD+glujiui8m3+48+ain0
wT5TDdwlXGKr4h0//Hrm3Vxf9MPCS5Se1cIUAGlbIh0VqBQfXZ6SmSfiq0dOAu2DpcQ3l8POzgnw
sYii8dFHbn+uVtNamVSd4ztPr1uBk4JBa94wutPnHs8WEDQFG4aS+Mt3R1MhBieZPUyh6ZoyZvPF
V6uYKMgRljTYdcBUg4vjmBO4x4Ddq2A33cLb8X+NEIrgGG7AYRlFbRO1jkG+5VuGng1EoogJhyjw
NsHegBIOcErirygSgIaTnTXnH8zRX9h8F26DXa/UU5Fwm0W5d7TP9hzkx+w/m/W8tW5sAAQunA+O
OA9yHMKrd2BaX5DmZYU03sQoRmMmzLyZH0vNoEXyqHsYRodKyMY+J9NMWhexPDJFTjig8c0NmtCD
3srQUztKn4JrI9kKwDLnCyI5KwNyrTDPhzbCYirWC+k9f9WDJyG7g0SrmQiEgyZ9oYKhrU3j8kxe
JmR4tAKcspI+fsidBALHlBgDnZr1bY52FalUukRXzw3RIyqk7obCy1ESw4ra9ndo/mfqTd2l8CmZ
7b0U5VK8hE9HPrbvvxH5rFpoAqWD1kgm28PiFWbQuUd0b3vw5Ob0Ew5oCvDbPOP2VrzDSBqdC84D
uHpJ9ZocFwfUTKXFO48YVgYxTeRbkUBdCbdnn2WEq1PHJG0i0mvW5LoYwqYsxMo1rdb03TXPtOWF
dCKGupxlzIbfAr2YGASz/GKaGX5g0M39b1n1g5wNDsmd7hSxuueVHgp2UdogBePNlp7znKoZNFp1
01mvQjtKz+HXvbI3mOuJZ3xjwa9G53cLjRJPH2X0Kyr2TkTCYAhSO76qV1sFfOrpwlqTRlzbiFrF
zj2HLVWvJv1Wqc/93j5PycpBaKvZyUAMkqkGmUw+KlJJbIacTc+MlDlOBLI5Hb7EIH04kP6AEeE8
biLrR6nArLk74wYaHhoDuLN7emBuTVE710QH/mx6SCGvEmzxj/PVjCHCRqNeeP5uL7ZY5wkiOQ1t
CtwQtOqG3agrHJ8NwwdnUQYedCn//sEzTGWrCN3bUMut30wxEIa9+//jfMvq0c906AujhUC1KyLR
wZq332ov/oTxmIYstonhHnehN2/ie3C6Ko0YO9pvyZyjbnDuLz7Jq04dGZShArAdzFc89m/9E7GV
a3KKmc7rOURV1/qKBrBpylBuWa0mXbuOcbYuLxVcFT5cr8VO2d1/ww12cr9Fgs4ioccz3DNf3j3l
QBEi5eYRE41CGFldGm2JzAKftlEqlFSWhpLWSVSHsKt10qo3/g11hpMxDTEbAwougP91gwLdH0Sf
XMdJjp8v8LA0YjkwnB5h+O2fdjYihhKhhWstDv8xBIFQkKV54XUW/Ui5x8eoG2K5NXoFszyIvvHU
0IACyClnyuBrdHkSOFWJ2K2Xwy/Wit0oeFFVU7DWrzJJs1U5tgsG5TSC3KCOw+PgJFw2ARShkaq5
I8wyqhsrkvXDqK7dkMtHIc28silatppY3hhmCUEXXVp/DYeua5Vs87rsU2wzjViv+ui5B2v+/4mG
BMLToIoprW4LCLdEXxRFpqpLpvMRe7D4J1VnMvsvLEYlXfogKjfH2R8QEz6IJ0AATU73MeAO25JJ
RPUaJYSraMMxKe1iWk/oA8ocwGksRlpaE/H45XBbsafWlljzzSeuw6lf+bKNAzrjKj7KmR/X3oYY
g/ZoE/mhBNCDG7JTIqSuBtuwIqPJHlP8ub3gJ2NzEYRpdfMo1FzStY51Oug8+2DHQL7bkxA6sxEX
7H94xBesXaiigmc75SsVaAmJ3/iTO3YfWtaxVkZTpo5iolMGWTgFNA6KzUAzSNgamwDQrPKBKdJY
zglzx5BKm/YPwP5WZ6Sjtxmw+pnNGdSIEAnXMJblaOi0uo5eB2G5PlsgfA9rferTFqwrvC6N3OUk
3WvEBhQFFWKzyvEOOaW3zjG89vOhT0epWrD7chxKHYBGbQDSPoZVrI963WF9ls2O7H09W8bIguSM
QU6Zjg9wY6vsiByTNCphAaotug1Qjpigd9Vj3jDKUFAC+1obMwisKOA4FI6lA3mbEeGxAHCaznT7
Jpn1jS1susN6sPBP6orAWpTmoC87gQQjbdt8DOZeBk2qwaPSJ7DF4Fx6sm5LFDQigCrMhap8x3F6
xGZeVeDZToArb9bN6eBN99KBXyalMw62uKX4s9UTeK/lKRM4z/0og36XxDGOp2tThMZYmSMn5AWK
9AL+rMN2/ylod9dCKMvilRmDSTv9lGp1QADe2/axUjl5HopR6rGdZfr06zXFak9QtR47g/sI5P7i
Mb5ybbMsRrrT3f7a2BgTRUHG9GwG469WY+m376hfMI1w0LpEb7Lvk5iMQGtmAHjinFqA3j9x4lat
EBpfcGzNDYhTFspWyywsx5DygdjTvMJD3Wn373Fy5+QAGwMCLVPJ28GBe9ebPMPjaqwBxB4doyHj
oWEXTuwPhgGrp6sjm7+2vNlh+nYHEJRVBHCj6blr0xC5URGEPyWfpHBQzpwGfv1sWWjhcNcHcR50
DwMncIXTNvi3YR1oT5xXMFPpNJ6166GiDEgSm7BFSms3i7E3siVob0LvrBELBMgrcOssTuQuTVIr
cz9P7C7axcmQMhEr5WVTNx/OlzfxqJOynXCvKtRFORtzxnpvjcT+Nql1j0iXu4rU3xrdQjGZpEwy
/FhtGrbsgeEI9WedTe0HRL+Xu3V7ww7IA1urJSQpWI7qWhcPF71Iy5qDmudv3r2/T1ujbVJ4pY8Q
rTH69VOg/dbWZQRTkWJO+aiCtx5cOLl7L+rb1rb9IkgbY8ugeSfOe5OLGdvG/4f9wdvsCuGLz5A/
KZ+9rWHtfkHud1Lnf43DwJ4wYd38MF+IwhqLHj6ghz/rR1wFqmd8XIpvP9fTjdDdBmZ8AVX3PzEe
DMPf7zhrSA68J3aFooGL26f5tLwL3dsy79lRTyRz4VXtGp+8YGoA47VGg5cLQffydd+91brxSlWC
3Me+e0Wv+XRQeIyZC4x94NW7zjJ7tQcKy2N8nbxqLnk6OsV5eNuS2Z+2d8/seWIuNDVneyQo4qd5
CK+VZgGvGc9LR/KnM+yengLehdKrqNwKJAy0g7mOfkjP+/90LV1Bs0Fnt/jwjekbEAiU8mv/XPQo
jO8Q12NxlvckT8WamRwaC5pKey781o/7nn1gTDeiwsYWycl+yvOrO1/GCsHUO59wqVrCYjS/6pFA
sj33SA4tkRmAEB5wsNMdmv7Hw+mK+H1oNo5FU48qStVX/I4SHOgEPKfx313Ne8flQcbFIG8JyW8r
yF219A9I3akD0kXqHeLx5WdNgIUa7/xLVYh7jUkW5P5+WYIZPJK9Y60y70yI/rT7TlonLw89gZr2
a2KC21old+7YikZwges0Wugz0KJVHMoicmjpP0bOAZJi9gglA+OWc9nX5hMKv4HoTJrZLVaUpVWs
6GYFECg3lrnKlDQHNQrZm17T0PQIPSZlpm50vdyQ6OddOJBzeC7yHYUxEzpDmEXClbYCE8xh50NS
BJCWdESy0Vdr7q248lzkHibM53haKe+zUngkTtc0vdZ0ESq5YuEutEsXwQ2b+CMc/3wKRHXxkurn
ikwGEjPxKCk1tu2yglJDjO9nn+Vp+0MbyDwn0bt+RpokRdzCtK7Ref3apA3wqJYi5Hk82bG8ZcZW
v+pDMZnT7AwYC9yHsA69ekhkmQNm3ZgLAm00Vo4X+b0l7XIJDlqTUndRrm3YL2Q6KWNpjDdA58xK
UcYr7pwrgT2MQRMH+npPxf60ebBPznez79iH0NTVtHbiU06X1F6VC2Gr2oCjmYabU5PJLgt0WQBn
eDEakpTgowNENPTMsga0Kn5itij2rxITyP/Wu+BGaMRHWQijcc5uhMk/44aA8o8kgy5X9nwIzwR0
Kc9aHkjTHzTnIdqng1zHQaZb5AMnwxJwacVUhS1QpHHjDLX+KlN890RrlwnFbZo9E4LlR5bJu9FL
JdQNm4mTpu0vCDnOISqkjgqiv8jYUavsDI1e77ovz1nkZfuHmKH+nk3CI7C/l4uVtJaq5SCdlkWP
u06ODDD1ceRHVV9ECoiwAvSUIpyy2GcX3LhuCYcortBQ9o0NNclKc5IrX3HhO2eSUgwSblXCeYh4
xsniPT4kfMERSRqmPZio2JMI24THP/Bz96uLYbhsC0l2MH40AwPrujcAEIxDFQPaj4FgPDVd2ayY
gKmnJB45m9PwKTOZm4wZibwZO/BfCj1VjLK1P0tJIQxgoiGQS6keSuNvjElOVdpGyEthoTrv1NKy
a3ilTpAPI/X0oaWKL9vhNzcuFVOs033HxRntWOSoSN0n06oP3Y/zpHzz8kKemo2r1VViRQPDM9QG
iMCrufRXaTBPuUgy0c++B7gsB0skQ7NF8IQobQYseijsgmXqaRFkwkoixPHapOFV9Fyv50PfrkxT
1diOD8aK95hlYY3oM06tUgME7gxbRXzFYxjGeExKCUTnft0ubU7oRs1z98QeGQpHaStej8UjNPoq
3MeWBqcU/hxEkL3Z//gG4uZtz/ZNYEcm3O9QyNGCItj8pn07pOM6hf5m4QDMyzL/dXjKYNF/7//Q
jeK1IMaTuHf23jjC7GVhWmQ4d0+kGrHm3fK40agHgX3jIDHNON5xex2YzI8FWvn1im+00fdPpIlh
W3fChthAHix51tqhmm99ocp5QEaxwyR6Pj9XVCb5Fv+LHhzB2Nrn2aSZsLuEhnMkSvfWCTxf2HQj
2uuUlArNqy/TiTiK5e95/Dwd2mxPZ545oUtG8YHUx4laBHZbWnNZKF4SIKe9IWU3uzzSn3DfwlII
MQdaZrq19NDDK3X8AIafLUM2MNg6DK9bjAA/En0HaBdWRXWxXYjzNXdrBNh4UQW9OlJzOxHl1rAI
Lo8Wq3a9BI1SyegBngTEIBFBUWCSi+0KcAtg82zwFmG7K3oW68tIYwzHQ9qApYiMd2G1ldw1ebKx
7xBPpv6R1vPEQVfmHbzDdy0zgUwxL6XNNb6FqvENnNdLTAnxKtiNzoVBRuAtlC0M2oS2qk9wOGhH
Zs3LMmXbudQ+u7kHqg/KoN138yhhlQsAk0V+AZpuJA30LDkE7y56+3Iw9tQwcEszgIRtt9am5RB4
NnkrHAIggVvY1PXv7xmP49aptLvjhACWbnGQY1tSKeOA7kEEe8KvtSO46DkwBnJsh1j5KZIDOsoE
urGhf+6qdiebvSAT1ojE5o6W3LT4U4n9ibYGcbmOyB7KjhC7lA1+8CQNV3R2p+s6KKsp2WHWtSFQ
x8kaGKq6oGuUCn3pvKVisQ+tUF43ZkI82oXxYdzuiREk8UCCJphC7zAfjcO+vdZR6DXGUAQk2U+2
ZWbHcErFFgmL0YB6ou/XAr+t4AzMnhM93ynjco9lsqducO5RHcRW80OTJ3nw/9qMUo1HgJ6uqAWe
4uXYP9EnwSzw+qAz5gM0KOJA3bpr5iZNdszmnee0DuRo+Kxc3u1f0zIXYXLrn8C0EgLCUB8J8OQr
vuXAmoiZBplsHK51XEQiK9CAaz4LoH/cwgrDrE5TYFKgr9pBAW6BRsXI2WaTFhhkjUF7ed8gIBh5
yliIcav+nZ/9OZd5wbBo3hzeAIU2JwHXq2ewiFiu19BVlSZSoOKQXaWS4pAy2qkoFkT+Zi9n91UD
BzAMm0U6Xu/0U4vAoDebj3GRZmIaV5GM0+nKXwmCilb0cH5bsd2V3Me6uAThRnt2mVhHgTXXh+Ux
Vg/pUdOnGaVbafYtqw9wQ18MX6K/p8UuL+1TX0/49WWu+8h0nYhIzBdkXri4m1A3dP6J/gCa+MYQ
9Cmyp8tC47NCncrCPBSotEOCaNpPF4Q9HIQ1vOkpzYSxfuOeCVckfq7qcV5T/dVbKYsNaCaXNBNx
R9WWRROR35VOblqdylqwDm5BaTf4qXzXP3dsd+rwqHL088M0vpuWsM7Yc/sKt/G2ZJLeQoDfcN0W
KgsgikmrjyiOrc9br08MswbRVNL+aZwpD6k2DBC8c5x5LOV9YNaZ8cucjz0GkQ/XxrdyBJ9cylRc
KkQOxmjJzId3So8kV5bhizO8p3stXW5zPOl8XKoYU5JmufaY2unPxHaMpTMw5VyiwHDs2Q7thDiG
Ud/OAWvWsuZ8XByDGFvfWmlI8vxj4u/cr/sEVzKtKwoWJKB4sgICOUzqI3B5xYsysx4uykg9IDHG
ITwObN1HxnlHwAuqpxPi/kgLds2/ARIZbj3CS9iqR1nfE6dgNoBZbHWBOyY3RJAunzzNQAdy4+Fo
ilOyvupyaRTJHXUexvHO3OGUi21PsKLGb7xfgVRDqG5yJQzo8Lwre1IkJ6kBp8EWeQqKG4tGDufJ
ur5xvGIY9U5qE9FviHd95XM+cSGZyKiHvwlBp2tItoQofTyxEMHaaYK6BFZ/YYI1qg1FyTXdpk7B
Zzj+UN3pNyv6Kcfj1RdeYg0YKFQVIgp8lzh2IGjH0NFJM8sVWtmasZMBzX5OBZTfGzct+GJkQdjU
TZanXKqHhzNNrxScrpHtwszP2gPVKa31iAOQ4IXyjxBgSZo3ti10mBuyZBHxzMuAv4HeoJOKw546
EqCXI0UKu3zXgde4I+wjMHnHwmmAWiXwfd+Skzme51Cpo3sBuUvxGSYfg273E+QNppTnMbZ1Z23v
DqELKq4bk1v5kst0+dGF96Foynp1pntH8uubV6go5K9mol8p9voYyUa0GAGSW6c7q8DLjcCUBvD8
uThcRMiZl6uczw2qC9qPXCgzvL4wp5oiE0QpXknNvRqwUF+FVUVo01EucgvputxA2pOMOgEZEI7O
nqOnsWO6iRnXQ3lFitSKbQthLq1J0nXuPfbtMGS2BlOguzZM5iKWiXzF6fx7WtpF8EPCYIgr/JQf
zduEogLRGZrIGG5d72yI/p3egMogUZftV2y547Ab1LB0TQ8CEyaONOmNDovB/2tb7dCvH1SPk3JP
idP1M+oHt06gbuTeblAyvwwDR6sGxqs0Z7MJckXBosuQF+XZIglChWIT8QdXSbRImTTpRghLr830
1NPP2sJ2KWJu72L27AX9nrVQSH+R4cUaYjdAT4oc2bb6LAXZNRqQukA633tu5J6EEhrnsHjtxdKg
Me8w3mHz4+IFJc6inmYKSnceTCKsJ4od5j3Xg7hbPk5C90iJ0kw9cafWtF8aufE59dZHGlnEiTmK
n/qB7UhpkZsxzvzkNDZC/sb/o6MwmVcxBCUJqmqP+d3j+RHymFH6VoAQ3PXBYSbPyqOxD6k/hBjH
UrSMxwqWX/g5CiVBhWYV7H7bLs2huDwnVL9HMSTGcdPd9AHKnAY4keLieWqOUkbQHPiH2Txgxobu
5mg4l/aO6f3xeLmDM3Des3Apktc6O9DySwD+GBi1YMgGtUa50dNXPwto7C9KcXmfzVPtUnZVpZ0P
ItJx2n/An0nus5RplQ+zH8M0RWiV8lCH+pea+99yQDaqoghqzDlUvES/mcrtMZxgU+4Ggn7/o1SJ
LJimE034oE7v2kcBQRTsG0+MgKQth5+N7gWv8o+fZi0l0J4pA31FNrL3F8epN2DD6vPl1Oq7HUlY
BIsBb/ImDRNLwpm9QuKPTLCkjWbFU+phogUAGvcOXrNcDCdJthPREX+YvcEtgs58Yi7AsisF9To1
3fHmSybu8kl8gEYx3BBJIzHLie6UZTmyPcLj88CqTohH61v5e/Jwhj1l7tB1JXMLgk/qgH6Lmd2n
6xAllC65LCF+y+xCoVH8FrTTffB0mIfGKockQP/QcdXsZh9MHIcQj/SSVUIQKHCcVi7U11Dq1RAB
lj7rqdh0yxRMhNJr+oc4l9Z/ZFQwQYYSkxK7UUjtlnNGp/NIwIxQypg148kH5zo0Djs2HjtyqOyo
uZwUnvnmr9O0spzNAO34c9XWKD9zK66Fvgq0+sAjzFgrkfgfxdVKLfnhGg6RRBBI3oe1C68YL6Vk
Obhe0pgsxMD0MxbNYnF/zHYUVM9BwS4ryq0BCOdJcs3mZeYK5nw8FQd8gl56wGdDmFWvGlGNUlZe
jNlWAlHJp0/hdCQXJckKYP0zhMtoQztQ+SrwE0yPh30nAUCrP/tQ1FWb/PLBrup4j/xrudxfcFik
DwPgmGp9b7c35SZcl6Limtj2h8Fsn5Leotx9F9d4/vAwWBvN2oTXlZSWNp7a3TCK37fZaRs6Vj0O
GUA8a+RCq63ieOf6fw1hhzuM2iGADLvjMpwmjVnPYGsSE/jfboCNi793vGbSm0Ic9qgcZBcpGU0K
SX+08sihtrAiY2ruNZHAn8xSvUJzc7f+vobBL09lOpDuvv58PB6oHu85wlzbGyKq8Xr73MzJsKsZ
6uthIIXvlphqsuvi9af6SZtmrNFZrBp/HO/P1+aRqqQs60v0qChdFVPjCY5TmJbIFHCTplIIoYlN
t/jlqNiDw1LHeMYsbtGu15eXnU/2NWXDgW+6lsQC11AxiN1t8NEt1UIwAF4AlKZ7vNOLL2+MopSi
rq64EVE0jcsbhJ422zFSWwzwnRYgdm7k2qBZ7Bc6bzhQ4OzKTJ83IjNMs7Co4m2TBLFt6ih+22TY
IIkD3lg+0l4aba3nuL9fWQebgp5PAwBfVxpH4RW10IrzXi3tjTQjCmqP7EVWcvoJ+1dmC6PeTYDa
0t7OqazaQBeYKcE1YrhgcSkg/tgf0rE3GnAIFWPMvWhukXtidbpiBzs2cQPsBCrCH3XlZGn3N2Yi
0zS66wVXOsyBpp3kqpHRuCEgD9XYH7r+ermLC5RUJCpd53M6DNtm6LWA89pdAzQqsbuRfi4kOGZf
YlGuH/inzpyC4qi0kvJdFSxGphD3rIT69dD7B4k0XcaOmCwwLRF62wUskYSOIkfEYd/yKlR4hVef
bTxW53RQsOevdnB2Jhm6MXCtAORPr5QZm2qDx7ooUrPpzdqyfUkjOAghWBxxAgPko4m57TwWSFDn
Kt9k1QinAcSXH5i/+YihTeVhcrxrh0RuwVD/YuQHalaNWrVK/1CjmbEesZK20UhL8WwUZqOZOPRf
0wxseduNv6eZ5r3EQMunDMXvQuEfOOzDe1oE9rPYRuhdI4irQr6IJ+KNliXMi2wVDCCndHAraDn1
0oHUHUR1tshG9IEMHwekcJntYyZLj9U9RbUXb21+IDnt+RU7452/rs/SN1GVqixkI2oNNdjQ4yCD
TwaQDPZbZ0SSgTiq1FBzhVtj6+w183ysbqlNewVgh7xzC+ShtO9j9frKFlKaLtkNyeLsJesVTOb6
9QY6X2N8YL88OD49wmvAJiJQj89+6QtzDfEoRTFfz8t56SgBhTabdaGJCybZMKru6QqytDnFucui
EojOZmWsMsCDy0aFyZvC3qz4M40uH05gNc1Gy+0NR/YyJlZX8SLa0TLmou3GSEwHQ7eJFmoJgq6f
PZz5Dqj+uoEtYdLaYHgVc37B0fv7ZhRghUynFcsbTo7P/aY2mBGoWZkVKNwIau06pCJdgLzDfKpz
VvFT2CClMHG9tVgJW6SdzV5JhmFvJgIrcl18rIGLYAFcAxNS/H6cG+Go2lmysrxEtspkWIkisnbp
X2RPEL9gt1mmku/RhXuPodaazqcypm/HiCwWFq2g05jbIyEMwvaLzoCkj/55572crl2SmsKrALZy
EW4DFKeKoKl+s0RkBY4qYhiJF/avNU3YPpD/x6iPDxOxqNSILzotLfsEf1gK9LtiwxrTm9eRZyX1
ZzLtCXX5or2F/0PLqBsJGLH+GTDJLZDzbqOftrUohdb2vYovVlqCh4dHvSpZPoG6U4j+kNZ3H9XN
uYEDvuvfTLUgGdSCnBO95Bix8DHyZeC97lyE0a8HLNc63OtJcAgXff9SfAG330GqU4InvCmWRx89
1nlG/HIpEsQmltndOWdx0Q00met5wscVzbJvu/s7jPhzXEHq9V+BaA1Zt84ePp2IfT1TpWLBgocL
Ymq8UbG90l6JImTYKymsYpauvHYxZrYHuXdWWPB+Mq/XYUYIrLAFY7PV0NoBQALdtb/NJmMySaNa
EZrVKo3wE6dtwqpeUYeFm2vZZ7U4fGR3BZAP9MA8szxT8kuCW7JlB2VMIChq/zd7DYfAxt27XtNW
Tf8FlQaaYMs1/qlSHrkbjuoTFGEflMPkeC1KkGvV/CajoeyIgiGSnkgD+zglJ7PpdXnFtX9z8Fow
idl9TuUFrrS+StLvy0CH+P4pYR7dHIEjc1VPPEr5hmQ0u2qf1KnX/ec3sdd59bRTg1+P8+CmZahS
hdmW/sJBpNHtLGkr5iLJx4qcOILK/fZ0mo7oNv6oYpvWUHCW4JCPeF9nX2wcuLUGtjrmIY0vntmn
zVBecVGZVdAnzRVLTpCHY+2EdnZVcaujFog0XNZzzCtrmBhmyfx/GvO0BU0RUIDX/tnqKki6aL7E
pPez+fWs5pFNGyb3r8wmUyXCzW0iI2trernp2aqrQ4CEzoPCGvjDKhbUVK7Z/7TEmf9T2eqRlRt3
6aDv8PlgBYLiRCy+XVcyztkVsvZrzfc4+EDc8wBlp4JWLZ7MfFYAF0uPJGQq5pZr62q6HKQ281Cn
1undoc77J3F5LQgqPHYpXVIJG45zmGbRqDIvDk+E/SVpX2+FLiIHglIVJxuc3sebu0ms4Bsr7Qc6
f4QcBzqTB7efsh7HRetS0DdfDF/BNKUTZ9xFfrhKlEl0d+bWfbBklKaxatAjYDv8GGkQ6T8lO0td
2gxI7FF3uz3QGJFcyHzDuzY87msRiL8vgQGRfAxf6n0y7Oz5FjQrPJ6h7RMRDm4FFoN3cty68uB6
Z/2AWUh/V4pljH08L1eD9AnOHTDs1/EZuDx2pIWHNv7btsNtqi677GY0IgXwaVuNY2l86s4EazDm
PgxRj8d5PlIQP3M7f0Z9FNRPuD01jIayyg59Y4dzf572EIkz3+db5V/Ac3FNIFCe/aMNKZ0HICpU
q+ytG5fNo2kYDPNSbxnI5TVwvmFA/fg2XJGyCZckCbXzEVjemSPx4W3G0+/os9AUyI4BBJJgdJpy
uW3K3sMmhC9sj3DC89HeYbSwWHwKCrRYsE9iUiMkWBABDWflMqik1oCSwGHBXKxMkgYkdVgLifDD
KW00r0Tr7fjUMSpadLBrxoPn0LzCz3Iq5/9P7Gw3OyKyPNHhKFgh/EgLXafuLAwvp9SHRAuYunz9
b2jdNFKUT0jLPc0DCSDVKm4D4lv+juRwkEF6qBk0PIQkebJ2/e5D5hAP3QZSM9VSg9TuksDtk4PY
wKmm8/Ue3JrRwVGObCl5ZX0+9TgbDlwumHQbi6j+J9zDLW7CKORLd1PH37B7B8H0mukrGokPojP7
3cVwMwb2zcC2xzVSZhf+sjY24B7QK1e4wyLKGHccig3mr5cNgpJDheJdQ3cpHD/zPy6EWyscTr16
YCguSd6i/cHnnV8ZLLcbBVxWwBK4TAtET79xPKEf4v35QHQMNQe0N8ou7ANYd7kUhiKZjLGC04uj
0MN2iBnXOd+x9mQ4u6kcVc5eoOOOuGZxixozGH1I5IKiCItAyWXx41Hcg6DZGztrYlzszkeUjnVu
gvMtxdBUuGbMRm+9W/Upb6C0J0G8sY4XlGsNxb6R/TjyD1rpoaJTKlrBTpVXSLsjLhLQA74CmLgt
NXLE1JKgY6cpiqgxmK8RwOF1FXfQMcn4b1dd40V/LXt1ayyoo2u8a5d1UjEMfq1RvnQk964wNg3a
MUbtsP2m/KEZnpMy6+J1qY+1FEyPNjODFl3/TbjCkUy1o/qJNz8jZTxmBNyuGe6zK6tg8DlizOzp
NV/jfjUFoFGlOWjSHNIGRb6G1iV0EnM/llkhljzHHpk6nXw6GTuU4fRX2SA+i6BELuQAdPSl52nz
x1O/oJXiSYWr9cuOcy2SG59riZtEDgGy8HvUPf48CRJZXbkxk4L21ZfhlRujSkcTgjbBHJA1JaX2
wEs5yFYU3wptTy9Wxfofxa3oK3BRb7UagH6ZKlVzpaNS0aqpq5BoUzJmXggGHjzb2g3IPIi0wPD4
f+RM30O/u3Te0HtvMh8u+kloA3micdtnQXp1IH9JLS4xI4xi6QBigwUxV0wSXPoqqY3IoE4rhFUF
4Ul4TdWRmxW39I/5T11hj7XNyi+wBxuytk86lTKKSV5dGis/NtjxxZtQsRe3LQv461fDF9pUBnKv
RHcrNYCYpHSVT+/AulaPwa1LseH3hGc5+DvHVJx/PUdo/y4GXDCobboApf600tlQmm+XEjMYpM7z
zNu5UAdtgLdQnQDwITuThAwWFgQErvOWpvt37sjcXviOlzX92UpeOAG1+Np2fAs1GUBp2E8k+W6d
gIWPyy01QXcn0IzcdqCtdUs7xoiH6Oc6yuBhna1/y7y0lRg0dtAzP80Rx/trd36B8uueNtfTyaIy
xH1Rnl7rhEF807S2Rc/IMymYsQvapvC9CkLtpTCozOGpEsevvEVk/L0md0qWi3F29/SdXlTiQP0L
awVpqHGCBzVaOAX1hbFlS/Yc8LD50pmb0v96JpmsPYXyIjqI6JYGJHBEwcUhNu1/MDw3diYlTX6i
kfR+/CSdAdYsQ3GEGgQ4l87+bsCZdeOj9ZCqS5mv5VjldBNjy9R7BNp8MN+iwOY8/cvIfLEbeAeE
B9Z1PNtFrq72a5IIEYxtCehLowhSzBtCB4lONCw9CMoNh2uWAl5MZDotYs4LC1byWzuEeFOe+1Vl
ZGRzZAijKs4lr5fLTghcRimUyAoxl0di8AMxtcnwEG4AjGBNxLMrWpDPR2EzgSNu8PDaapmzneDh
yAXgMFlWzHmVsd6+NGFytVYljmnKykVh8LWKtEyvstSYGFBS6EZaWANAfsVp3AOsx7NZeZ59lU9f
XVQ2s2bVAx7T7Bs3acZJ/nMiMvqm0a3bYmAW2p5TK9MvDXlJK1+MU6g/gESMunV8QPkvbxQ0ZawC
Ss7sGktNw4JfYIt4P4dmQO8rRJ+N34r8fvwwOxhJMx4iZkCcDi9ESzqnp/HzEVoH2+X6c1moXDjC
/razgzVprgHpfw7fhMuIQw7U51NwkP5ssyL+lwq7ouMPR44DKBVDPysDKCaOC4q0WYq+EfqMfz91
RxDZ+BoxHONW4xGR25ff2qM4zfqXnDWqditp6z+PShUxln/NAzfTEdBbyNMyy4AJuRq4SpTZW68Y
dlYVCmnsolJ8J22okiiodiU4lbREpRW9XnvajKt2rXbzTCzIdvH07Eje4wnJJX/4VCUzjJoJdQY6
IC6Uv7snOKiaWRtrdYs2tNjQuyeeIwgEpT6ahEuAMKNFZrpp0Wl1fcJRnACHKb4BwpOIl+0nACum
uNBs9lQt/H3z9MGwtFGoW7vmBHnrIUg/Gm7UHwh/jqJFrqgkktEh6TtKFlHSVW+hZhXFl6/s3Cct
nIy1S5Gg8vk8qzipXjCYG/do8h5Dycd/mgGfjrbsOnjFUJuyyf+bcdsq49ljuAeNWQx4t+9HYFFl
qCASkfuI7lZ8PLGs+/ETQ70aCpQ74K2yAureGt5uFTJHdr+vYUE8SXiEp+kjXJsLcM+Zk1adnJb2
UFJQkBtbQP0YvRY0O4enpjEoxhV0LURN/ucfH9VWX1Sg2NZWPuaoiDpUCxKnkv6Xf3LM5cr3jlww
tV3kFcVp5MevgKF/ChHLYbEyj0tkOIMqhgL8q552eHv0WFECEykT6QkT1HSuiNKitYHeUReFcGaC
m9aBuEGRRgcxlm6JND5ZC1Vx3aoVmCSqSy9HiAq6O/z6waqFn2XRF/DZoCipB7CPL584iFweo9OY
npAD+DgYgDIk0tBjAY5YVQnZUSFX50hJNy4gM9qTsCghJFw=
`protect end_protected
