XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����1e���z�ڴ��@�th ��>G�DN��!xH1?sEj���n�&�l�}�&3(�'���Ϙ�y�J��̈́���5�H�fI�<De��L$�f�d��uwkRvV_?+��-Ġ�5����Y�)?��+/��N®�P��a	�t�R�$m�d-�{~p���`sŅ�C�ŋOL>�EQ##�*ŭ�J�g�ΘGI��S���,�����x�W���^�	�1�����s�߭�6��ž���臃J]�&,j��9�d_�!�$&"�[�Å�dO��Y�Ku�JNNd���^O����[o�#l+����V�@�;�x����+9����Q+0e�9�&e�zѶy���]����@�K#N{�ve���tCn����\�����
�K���s6���d�L�[K�4��鼦cfrC�E�;I�=��������$H�Ɂ����,�kr��P���d�k��y=14���c����1�m�{�{���C��_ø����`�G��4r��-v��`�h!���Pi����o
�/��A0a�`fkg^���d4�?�vW���u�*��Kܧ�x��t7�)d�:�m��S��X��y3/�XN���S�l���H�Iā����1s<�>c  ���O��(c�-�� (����9��.00��u��u�ۃM����k\�����ƿ����+�N��c�1�2w�1��ٽ���S*�5�5Q���t�tڼ�t=:`n��HO�E�HFs|{ѷ�<kb��|�!��M�XlxVHYEB     400     1c0X�gB&۩A��'��D����c�]�EԆj��9~�7ηpB�W�w%�d�V{&c�[�2,�].Y7xy--l��LH?��$
:�%833�M�����!k�������K�f��� ^#LbQ��zE	2�t�v�ԙ�����*A�r�0B�bJ߾M,��F�0q�]cL�`m�X�^'.��.�L�X�SI����\wd��p��[���2�^��'��!�MlfT�c� �H�<��qk3՛J1��k��D�3����[:��Q_h�[�҂�,�
��+���Y7K��`�M;���V���b�1��՚x���"�����	�G�ѥ�\�J��,t)e�ۯQ[�:���(@p[p�ʮ����|� '����;�W\�����uF��)�yb"�*ӞD~�2��XE9~�Çs��B@��숼!g�	"�`XlxVHYEB     400     150�6��k��"���V 7��^~��lk7�F��qJ^����;ʓ;�Q���2èLd�m���\X��ݢ����a�~vgD��Ke>���\�Ԙ5��M)2���+�Y#*�<�5\A�\.Z�l���9e�_xxgƩs_r�u"�hՂ�G���:o��q(�����3}�7� $�����	Y���k��II�<ʨ�l���ݥ:l0t� ]���П<��C󯆙?�:T�ԍ۩��t .��A�	{�߲Y���v�Ӣj�I����I�]:+
6�z�4h)�=|i��H�����wЄD��&�y�S��;��W��q$y$��^ն���&XlxVHYEB     400     130��C��M&��]�{"�Qޕc9�׍D%�aS�c��B�bZ������>e�p�{.�w����[.T�G&�7��+�����ia���~��ԇP�o� ��!��h�^0�"��U����#��gː&�l��2b���׋V��p�+zp}̒+Mƣ�C�n�R��э���x�ǃ���H
9�xK��������pYJ��9�DO�@~�my9��~u�g%8�.Y�Z#��׮�d:�^����+��| �k�J�̚a# Ĭ�!|���0������� �Z�������V�3ԗ}�i9;XlxVHYEB     400     160A
t��h\j��&�E ���ꤠ�{�H�����O�WbDM,r�����P*�k5iDJjI���h�k6�� ���'�aN���?8��"��n��h�Ge�%�н�[���=D���l��ʶ�~n'[�0�.�|���k-c��'�w>,�?Mu����'=N���[�{+/������,��7vՀ�R�J6�Գ�$��al�cz�>ǉ���Y�}![T�xQ$,����̨��P�8�n'��'���K�@y���(,0N@���B�"�y�2P����~��/�)����Q� ǐ�0��'h�M718m/vv�I�>��H�8��C�m�s��g�ʱ�C#6��;��˲���eth��t�eXlxVHYEB     400     1e0��WG싅��(�Y=�Y�~��b2�V�$�
����K�+��j`Y���f�$�z�QBp�$�\��l�Qڂ:E��@���Uz��w��n���u�|n��qп�~��<�9�W�<�U�]�A����L;N�cǚ�da�m�t��J��7�EGC�?��]��Z�Ym��$����s��&=���dXA������%A�~k�ch�O2�U�v�ӅR�-n��W��a�#0vM���J���MdwHNU#����,T�!o6�QS��3��PySѾ�>
�lR��x�P����z��C��J�V;���;�g���8��q��{��9�o�|g�8Ӎ��E��9���>::���X��s�#�I�kr��*8#��U�ێ���~��b&P�{����)��+b�2�/r-T����>��]2�,���U�nL�No�	�6�X��R�&6aD�A�}>i�@�
�3�prXlxVHYEB     400      f0)��6�p��3��o2p
�lOt��E,Q��<����[�[��v 7�c�+Lq�Eɗ.鄴��5�8N)~|}KkLƲ{ ڊ,�+P7	-�~��6��\�ѸuO��:�m0����6j���[��lp~>m���N����bB4%�x�8����?H���b�>�t��F�7��.��,R�TW�lFc�9�h��/f,�.\��Tt�2+�D'�d<�s��*�@�؋�Ǐ�3��H��XlxVHYEB     400     150��6�S�(�=V�t
�5C(��z�
�v�.��e�66�ٽy]'I�*yn�Zw�~�*�������t�sΣh��(�11���]���a���q&y��#�=���gJ�]�Z`��9"� �Y���<e��F_�-fg���t����2Z��Ei��htj��(/ZA����Y*a��-O ��nD]0���6��O�7�JR�s67�ur=L�O�+}0��"]1�k#�X�i�k���u���0 6?P��u��m�H
47��_{�t�6Hg(T��Z���	�Ȭ�R2�x���C1L|ЋRhm����㑝}^�B 7ͮs9V��v��XlxVHYEB     400     170�������Ų���w������)��9� k�J-�>��E��xR���r�<���Yʬ19�eƾ�����g�b�r�\��	ah��1�A.J��V^�^*�^u�T�<��졯:�)���(�a�X|:f2q��ؚ0��/���3!s��M��
�ì0���D���pp�iu�D(�t�t���K�ժ�Rf�5��E��P�?uWX��_E2�fa�������ԪLJ3���0I��^(�k��O��h�����<UD��]�{;��q�N��+L�΁�oR�v�Ŀ�;�<�Yf��Q�T�d}
��Ԙ9�ޏ�t�iW�ҋ�=
*6)� W�e�j�O[`�����,R�ԏ�H��XlxVHYEB     400     160��ݨ�`��K�$�	������"�|N>71�F�,�r�0�u4�=�����/T���>��8;��B���;l���x=�Q$�\���K{1�>��6�s*L�H��d���B��V�
߇9�O�Ψ�l��֖�k,�[)d�A���
�wӚR�0��'�<��!�l�_W]ק��f���|���q�J�Ml3�PxvF,�Py>h|~1��vgG�8'r�sN�L��=�ޫ��sm��Ԓ�M��,�;��g���b1VnOsdi�e:Z�p� -�CZt����Zt'���'2B����!�o&�V�o��Whњ��s�Er��e���dY�y
<O�j�Z��Đ�XlxVHYEB     400     180���ð�vk��h��I�>.#��Sߞ��� ����TE�	Y�iZ�[�ЅԾ�u�R~q�H��U'�GL����^�/�¶ϼ�&~HKO��f�Ea̿i��:�l���=u�
%��#'�34�'Pf��l@q�A��(:3�ડ���
׏yu�y��x�r���y�C;_2�����=��5q�Yt�dh>(s�G�����ԏrbMD���b�6D�-Y��eYYa{�\���^Wz-}�N�A�3��z�k�[�g�pԴ�S��&D3����0�b@Ǫ=ig�XK���5`q�P��IiwE�5�#l��_!
��/��r�}�T�؎w�i۔�$R"^h4�miQ?���O1��g�^���A�=G2uB)ѡJo3��XlxVHYEB     369     180r�Z�ӿ�� �(���_I���/�ws�^�ɿ��KTR�(�	
�u#��h����0*�@%f�G��7C[����W�L+a�0��4m�����(�ϚK7>�)~�I�o6�J�^lB������<2��g�[�0PU���/��tih�h���n�r�r�	6��%0q�f���`��e�ow�ۓ������X P��C��<�ȔS{/�ѥ�������&�I��������a��)7%�T-}Ŷ�)�9�#�ʒBs�|�	=.�뗠���i:�GY�����Y+��P%in�56#�n�ɷ���i��/[����R ���Mt�!3;
��������~<f�lR8���z���w��*����B�Vx�i-F� �h��(�c���T