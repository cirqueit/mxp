XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l0Y6׻)��B��x���첫�#��ts�t�=��F
ۼ����Í��D�E�7�2����)�����}��Xy��_.B��L�H��U�6�ƌ��ݺ��] 9��+����h���/?]��.�k��+ٚ����M9y�ϺrƛJA�Ʀ���5P�SAm��6�n��V��S�TNv������>�t  �4î�)eB�hs�?p�Lڦ�ǖb�R��Mqg�k�4]~�]b���=�*-��oV�4���4;"g���iK BV�
� �^�m�������=E-v��\�;Y�5!�g�Znh����srV�)���3N뮻0�n�-��|�q1^���6+��,���LP�6h�\��K:@��L�7�9'.K�*sj�0�[dYg7�E��)�{!b�g�!����壃Q��]�7���.�|�Z�l	�Pz^�$\����<R��N��KM�,J@�^� �	b$c��Nm��D4~� ~�"*�����U.���^`�gAc�ہ�{	t�xOLp�㧉q�Xk0�*-Z�B�Q���a^�Aa#�AҤs��1��j]�C� ]��.����|B�cp������M���p>�U�Un@m���J�^��G�7�e���8 ���k��L��sYy2~v[� 	ċt�N���.�␚���Μl��I�7�1�L�y�U�7|$�����!������I�눜�'8i��,Ţ�"��i����j�!.�O�����U/H����M;lHSdEIj�#�wRgXlxVHYEB     400     1a0uД��}�!�/���ہac7Ώ�y���������f$w��Y��`���j��`^��t���+��{Ө�Un
r�p:m�;A܇@�C��#���Nm%i����I���|ny��*��A�"��`+�m�C��ٹ�P�mX��ቾJX]��s�aM�Hi�y��5Ҋ�m�I��|p�/Wei�IfDY�Q�4��[����n͠oנu_�n�'_��a�|3���v:�|w����s�u���x 8��5D��e��=���30�Յf�ק��c-f��eg��_~�S4�	y��S�g�ww6��4��ή�S{��9G��(�X�F
!�&lDs�͔��""iE��٤�T��ͣZj��T���
��7	};�U9�}�<�����^�3�"��~�����r�K��p�6jv�����A�}�F�QXlxVHYEB     400      f0xN��@���NՄ����^ٹ��Q�\�0w=FI�4v����l��[�t[����C|�P�-����2tں����w��Ć����<%3ݾSW��F���E{����y�}��5."V����'�.ޙ�0D���T���􁈣�3�����Ѵ�^6�Oo�neB&�4APg)�C9�b�J_h��/�%��GM�;�4��3%8�t��i�~���Hx["����7�r	����8�ρ�q񙍤�"h�����XlxVHYEB     400     180~���G������h6耸heAYޕ�� 	�D�lT}	��{�5�}�r[4�d�o�·a/U��$;�m�}�@��q���p&��t_T@Q�#�6�����ۢ��ҭ�=H��F������jzZE�f!��-)?�ks�ݨ��n�%�L�Ev�T��G=��-8�\D�B`�aʤG�n,;66�������a8��~���*ۏvz�	��.5���d�^��fk�kZ6Oǣ(�;k�\[�y�eB1By���q8�ݛuP�cpx������좶bDi@{���0�	d\0�`7����'%��I�u�R|������Z��Jݢ�N��щ6>
;��׭7a���uB�����'�ц-�|(�iN����^��#LW58�:��hXlxVHYEB     400     230bL[�Av��BE�P�?xh��S�� z ��9&�C�4Il)'ԠPm!1�#�{�a��9�]MA��H"XTd��IY��j�*4�L��~��]ѣ��	�ixU�#�4�;��`k�QP?�a���0[�+��i��B���T���v�C�^�����2^(��8�B�2��~���W������=�4idS�a�)��B��h��-	C}����W[��;ac��Eb��Y
��o��t���+���Et(=�}��Ѓ|2	��:Q���DH�����Z������Ј�6:�=��=R����]bJϦ��<1�K?2>p��KLg�=W�����KЂ&�h��W>�	�ٌ!�����8��;�E\�='�tv�K��Ő�S��K��<F64��_�b-N4�!`� N\��V��E.-r�<�7��5Ue�޺��Q��7k�jiM���.,XJ��n�U V���3a�f�S�	��&�F�+b����Q9�z=��<�?�t���ܯ�;i���i*YqŴ�oD����(������	]9�݆^ٌ���Ts�\�IT����-�pXlxVHYEB     400     1c055�Zr҆�k�%ᛥ�"�rD���)�?��#Y=%�yuM��DƉd�J0�{����r�A/ٴ��w�)�bdSȑ׊f���v�	m�8��#�_����ׯz|�)y

��պ@�iP�"��� )p�7��E��\[�J���/�T�@��:����	��Bǿ��I�!�Z��RN�9�>f�/L��7'J#P���1�`�٫���4��Չ�:P��YX*{F��ҟB~`�'���lt��W{a��\�=#��j�LE��z"~-f��.s��~	���y�v��pt���˽b��KL���Gs�2�]��k��C����t%��:�7"J��r#>�@�&ݠv \_�K��#b^	Yi�m��};c���/��VD���� D˺�� ��y�r�A�v�9��q��
:��zq��q��� 4��	}��XlxVHYEB     400     1a0�7�iX���
���dGz�MF�5M0���j7F~B�p	�Ɲ�5*+�����X�k�����
&����H.ɰ�%���(�-���Q��2
�n� �+-Z5��}����p/�"t���J�[m������,��Z�f�R�s�"P0��8|��Ns����m)�hK���q�eR�^DoӞ ��f�0��#�����3L�mcgᄄTt|�y��$~�G]�k}�ml�rC*+�F�n�T1���.�X#�G@�����K��qU^�2#Q������t�`�o��|V^)HE�@�CY+��������=���S���_@�^�ɌQ锈�Ph�m��rc�4æRh?[k�=k����8���	��#y��V	ߔq��h�����;8�>��Z]v���>H�ay����̌aXlxVHYEB     400     1a0��М�j\I&B�R�C�"��"z����+��2|V�U�������-#@R�$���f�7�!w��v��K[�ώA�xZ@G����rDN& R�|�A, N�"	&Y��wپ�H���9M���eW��˫sÈ[�)�i�u«��� F:hI���a!�qK�~𕸥�Ø�E��&҅�y��x�P��@ !s'T���\�v��Ş��L��Xz���QI�RK6�p�L<SQl2� 9�D����%� ���Ȩ��B2�����X��T����0�Iq)8����u�0�f��;����wEZ�[��*���F�P��� �QޢPmHI����v�ȼ 1��E
��EB�H�m\����n��K��V U�vvV�(�?��a�F��3��.�'"�V���G�XlxVHYEB     400     1b0�Im[Fq?UE3Vd*ǳDɭ#�Vڇ޽�b�U�F3F�~��8q/����T�p��:�4�l�$�p�)�t6�9��� �I�I�w�y��:�]a�Q@;��0���z��!!���M��aFƎ���Ϻ�����x.	pڗ
}H�"/����[`7��ёPTvx��$����6fŕ� E�_(x�B�z��R�!ڳ���f�r��ۓFX����<�X���D�4b�o��#
�r�����3܋��Y�>gԯd[?ߣ|����sq����{��N ���H���d��mwż�b���(j�u"0Y(�>ܧ�( �l����,����U�M��U�?_�1y�c��Hq��V��Vq�F�yӢ��X�[�͋�T_�J8I�uռM�E1<��`�,;���.w���F�L�3.OXlxVHYEB     400     1e0�)+���Ե��K���` q�Ͷglp�o�3҉�7�i�@_����`'� D�`X��ca��(�y�m�����V����Y���
���Cq�>^֭BO� ŧ�)�(�24{�#��b��� �J/��ԕ�(�� ]�gZ]eD�A+ouDA�]��h�Ų����� �r�҇�TFg����j0;Gj����T���j~a$Z�+3���	�)������n�(�
Ѵ��,3���/�"vAJE��I�� Д��H��U��_~�A�W�ܪL����.�u��80C�e�Q�Rq�����W���Mwzc��T�G�׉F���_��~����f�ͯ��i��D�;��v�MT����5�$�\V4�J��߱)�,���`֥�'�r=�]ÿE���,^�_Ö����-�Ȭ ~�w�� �������,��	�R�ސm\f|/'�!����I����HI���q�)��w�fXlxVHYEB     400     170�&�À<�����)فt�"�<�p�2ר��YP9�Ң_���T�k�~��#/-�{�~j,�-oF.NN�����"]����
�W��P��f�L�ـz�:���ZN�\z��]#;�:�
mw^�Iͷ�����R�����ڭ�+#����b��3,G�"$(���m!�>85�^�"�����[�ynkk-N����EO^�h6z�Jj&��Ӎn�[ N�Sy�R8�}��,1���Ql"�ȣ���1"ε�7�Ȕ�� �N�9��jY]���RS�+)�p�%�J����Hb�6@q�5�P��o[c��eg��z�k�u
f��L�#�K%/n�D+���?����}�����0{��XlxVHYEB     400     140�kK8F�_p۽��ڭ�n�6�2rؾ�q���������u��#	�+#���q�L�~P���1x �-��gw�2��C��:;�2C��tDt� �#���Xjl��y!&�3H)��9�F���_�><c'"�"��X5���+m�3�a�oZ��Z:@����9��"2��b��xd�h6O�9��٧�� a��1:�g�gR�������=6u;�
�E�ψ=�N��CM�ng&�7S��7�%�e9}?WCmЫ;B�P�B�����<�WT#ׇF{)1��a�k��N�q��s8�ZQ�L�ꥸevoT69�^6Z�Ow���w[Df�XlxVHYEB     400     140"�j}S��*���l��S��䖳�@�}ϯ@5��������Q'r� ��6O����G=��̥{B�� n\s�y�yv��Fe�in>
l���i����4�}g���P��P6w#A�Oڑ�R����1�6=2�����G�=�U���t_�g^���u�7ە���4�Yʢ4v��C�?���U$X�B��sx�1'�N.�ͳ�l
�j����h�%t��Z��y��DD����/���nǵI�WǬ�M���� �ˍ}� ����ٜ���z7�>�6UBS($�b��f����LW�8������de 
�%XlxVHYEB     400     180;�#��6U�O���P>�C��T�b�L����>羢ވ��	�xh=�3ݻ�9�;I�v"�����C����R�lFfkd3d�VFQ�T�x�a����e�_�{��F^��m���Ȼ�[�'���;��B(azi��-ƶq� hH�9/L{���J(�Y��gz�9I�Wvg���H�%���dD9�~�]�Į�j���6�x̝B�����b�d�������N�{�K���ʲ��9��;�-VSbV���{�����b�Ӄ��)փ S������b��-_-B٥B�Z���"$�z�F�C��C{5�l�e�i-}��c��0� R�u{�!���Ȕ�%}��q�����E��I;~��l�v����T%I���XlxVHYEB     400     180��Lm�}���B{���-HcC;Gv:I�"�}e��EO6��v�|p�d�_�1�
9������;�ͬ!�+��E�~��}�$������1��/&�/�������'q����>#0��������t�?Zbڢ���;·�����#?|03)+�q��*>Mj��k~ע�a�M�f��YBR?WW��(l�u�@��|-�3��dÇ�.G�O��0/����-�
����4��7����zSj~� ��2=���]��-�/�:���W�T��S�d)L�w���-Q���~��7<@�1����04�8����	��#S�X�k���}�7��ci%,�7��f�  >'̏��4�J�Jwu�R�
?�`��XlxVHYEB     400     180c@������A����Oh%2���d/7�d�?�9�C>.�2_���%(D�B��������;t����d��9lIA���{�en�41o������U����
��'�'����[���%GT�/t�N(�:����cHa� �i�v�]:�֫d�}����{��J�Р�+đ���=^�h��13�Ǽ�Źz
/ ���~C]��X`c��|�<Tw�)蠏�����2�x;����Y仝x������`�mo��uyW�\�R�dZ�4¶�v[�*���n3�R-�1�ؖ�Q�������*f�.�Ĺ�ii�	N UTC���XLtRx�#��yAܯ�Y
O�ꪟ׳=@�Y�`\�q�	]����/XlxVHYEB     400     1a0"ck��O�H��O@G�o:YV��xb�:P�Rג-g��^��y0g:�C���W��n�,0yw��s\`e|�-���YbGLiPC��ꁲ��t��Z��ŤZ0�%6)l�Tc-ſy�J1��v�*v?�p�϶�����6����1�	j���/qK�DH�h���+�CD��;�K_Z�ԱL��IY�G�Ucw���?3w�����A(�0<;T6[�e�����Wu�cY{��I�C��a�=�w���>W+�#�X)����w�0����㫢L�5�� ?
�u�~����ĺ��@��4l1Da.B���Kwl���ݟ�l��hŃ��Fz���<��7���!��\=#[y���!q1�����:bϡ��}�S\Y��C����m1�]�Hh
(��?e����q�4�D�	����<z��4l�XlxVHYEB     400     1a0��a��ǫZ�3ƒM��C�h�'7�3|�f�te�$2��b�󷊏�2b���T	��zł9P��P�
�Z�9,nt�cE?M�Ӊ�Eó"V��6'������qZ��iG�҄����\b�;��5�5���@d�7���t-��Gp?3��$�Ӱ;?}EK@QFn:��!-n�����}�"D\���ܢG�7Ho,3�K6�b��ܸ�������FF>�[~��Ǫ/�a'X+�\������x�LU���+�6a�a�T���V�"N��q>W����6.T&�~cg�J��k8�Qϣ���:�I5�+2�jXxY�:�9�kx�5]ƚTǨX6Cx2�k�n��B{E5�������'Ĕ"�9N�أZ�s|Q4 �pD�%����@._Ԏ���b��5��H=� 3�XlxVHYEB     22d     110��^�081���,���X�HH��.y ��e���W������90a[w�%�v�����_�n��������4���Nѥ',07������a��.�Q���8�b��H���Y��q�qB���hF=��,�e�ٻ{Q*�1��ǝۨ3*�<�x�r��ԯf��_�w��o�7%�k?��o�5��{�^��<���	���
�-y�QR����M�R�K�g� ���zE!~�x�c�x�Qs�b��������QVt앾����^