XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��AE��C ����6�) b���uSeMi�>U�>�Б&���wp��z�A$�qG3���}\��	�q��Òb�0�Y�y��ʾ����~��u~�|)�WZ��|���t�����`1����%l�}���vu~f����i��c��z[>�!�pD\x��u��w^����*O�^c���Q�W���1����_��H�G_nQ�^;����2k��PeY�n�Pғ���PaX��!�"��0en�y]bi�O[6�R�&�Ct�2[=_�!�p��S ��=��s�^'��~ֱ27:�駯��1H��&�#�v�ۓ���ȑ��������`s̮��i�U[Iޡ𼦂�(V���&��e��zc�gS�t06�,~����Q�fĀbՑ� �6;=:{�D������\�+�,o������"Vk.�A�]#�]|�����h#��]`G��A9�o�x���|��g*@9j�0�S���xԜ4�̈�]��Iyр�MGo�J�ߤ���r�sp^P���#�vv�J#i����_
ڇ`Ps�b�A;��Z�]�]Y��O�%W(I�����P�c��-���Q��3��Wn�$'S�(��D�-�ɟ3|yW�Z�8��)�����*:鋅����o��i�(/e��u6u�U؛j@��~v/�A�=y�T.�����,��0�>S
� ؞�v@ƞ�Д��2�Ea���!!��2�~��N%�\FMV���]�����N��#	�b��1�y���,�]����@	_&�Dn�H�9XlxVHYEB     400     1c0�H4D�bV�qb?�z&G옃�<Z5���?����{9	��vdG�TѼ���,{G�;��K V�g���1���U���z�*-���O���tm����9����A�E��qh���}��P�D��>�j/N��T��i��C�?!��F�Z��	b� ��Y���Zw܁S�p���Lb
�U5EY��YS��������^�z����#r�ju�⥓��,����Ǘ{�_�Qʳьt����3���Խ�S��0�7�� ��w�zi����U��z[������0Ť���٠<U�m�޹�]���o�ZX»G��յ�]71�^7*S�䀎N!�R9�������~�6��G����G�51f�@$�|��UϴsQ1���F���T`�=nX�c�u>��2C��قe'�m>���cO�>f��1e�Ԑ��*�y�]�^������+jXlxVHYEB     400     150L+*��2�d �4䝪�7�8{��߈,���tߞ|��?)ѷL�/�3�)s�����j���t΢� ]H�ù���N;�g�<��,�c�B	���sK ����=���1^XEKn[}֮0�����g�R���N�R���kFZlx���8��%��p?T���>A՟���*(Q�ϼ�`k�8��|�o�Q�n#�g��y�e�y8��LB]�;EO�p�^�g�K�T������y�Z����?l�<��YD�v
�;6E�K<��ˢ�bؖ?lwm�'���2XL���kmc�d߶�r��捉Ax>�\G8^�����߂U��XlxVHYEB     400     130範��6P�sIM�vB����JK�W�,d������� ����Qi27*��߀�M '�u�W"e�ȝykױ�ދi�>t �7���Q��	��ۍ
��);���IX�?g����g\����4�-�v���L\3�g�B��x�\��ī�P�䛆���C\�Ýn�(�~�[�~΁�eMƌ��A�6�IR.t�������c�\��@Wو�'|�Z�;����c�1��e�;�<�m(BI�Ok��>�°���0���|��O�޾�L��=�����,�J��0AT�t	�"��XlxVHYEB     400     160���ل�2���t�ɲ� ��~/��ަ��M�Z�ڛ5o�� c�컻�ɂI�+즪
�r�]�s���j7�8�l6��,Y����2�z!v�a>Cc
� �o$B���ݱ�X���
%fA�&����Y&5�%�;?�]?O�}Z����� �{�+̈Ԥ��"SU���muʹ���U�A2�TjB�����.2��3�pX_�G�hA����,�8�o	��b>L�kT}K���!��Jzհ28I��<��H��<�p]�=@#��ԁz)L�ݐ}y�ʑ�ۖ\&���n���Z#V�Ӕv��4��5��N�"ƹq+�%�P/��A�3��нs}X���~w:sj�̢XlxVHYEB     400     1e0��n��[��1��l����Z����䘰l" 5�����d�:9T�����Vj�bp��{ ��U��Na.V��[�9���r9(iQ��(Y�&��3�A�>W��f�?������	@�,g�$C�"m�,[��f񋾶yK$���v�]�nB����ۈ����+��0�b��� Gd�P�^P���-@�&�*������A�y�t�z�fn�v�R�2���a&r0���v��]6�:iߎ=�L��K�2ƫ��~b��Z4Ö�1䃻%פ{�:��s8tѼL_��>��林���K�^*���P�[�����8��1��W��=��v/�c�)h���0�rX�&vI��{p���O�#ໃ|j�A�q����Z�5����IF4�w��@N��,���̦p�Ŧ���H�G��i�]0(V��絎�^��q�1^�a����MFu��ȴ�<�SQ�N�#��F�$,�2�����.XlxVHYEB     400      f0�?�����P:�\����)sT<�s��a�f��~���I���,��a#	��"�}A�f���u+���4r@FR/o
��gb�)!P�Z�-�N/��,��>�kgK�~T���4��=�N�F�=>�"L��t11l��Ԅ�B�iF)��>e��_���8`"sU^��|�x�&�U0��s�zQ8A�0����[�Ix�3R���x�2�Ъ��թ��Չ�J��$fڀ^��m8XlxVHYEB     400     150��
K *��E�?`��(NH�%ǥ0[t^��X�6���c2�FF�q��jk_l�h6PF,}�)aw1\*
�����K
��%���eĥ�&�z��b��~c����S�d��46�}�a3�V ]ѕ&�׉N:��Rw�{�<	aY�ZA7�����U����}�~����ś4r�)KI�Q�����L��v��N�*�p�!�B��6��s�/,\�y��'����X6U����Vf��oT��� �_��5�����7Ek�����,7���z<B�Er���O�R69�UD���kdU�0��0�^bI�B�(3��u��ߎ�o�٥XlxVHYEB     400     1707}S �J�y!��e��)S����=lk�
�{:*�
��Rk{��h�'�5mAE��أiQ��S�dn�|o�&2ć��ݤl�v<?H4u�]$�aJn��)�t���,%��4�+�If��m�X��e^��z��f�9��	���a�K�WӴ���)���(�v��m�Y��g��Mp<$�s�D�k]��q��@M[e���0�a�
mD��8&\]m�(kP�7>�Wsh<��ff�:��nab~�f{)����(P�g�t��%�����_��_Og���Q��u��B�*�|�ގ��5�A!�M/�dE�M��hT"7V�i1�~;"���]��n�$��F�m웻^|>�L"��ܞ1��{�C?ޚh �J04XlxVHYEB     400     160���i|ֳ�Ң^A��8��l�V���D|\iI=�(�yY�{�\�
k��[���l�&'Ĳ^�<�7��j�3�s��֎L�r��y���	4�ur&[/��1���o���»Y��$�g��/��2DO���`�����A�*����JWbHq%�vj�N���Y[�0����w�Jvڹ �t�^��D�h�u�������u�����
	lE���� ɨ4PK��YYx(��)��~��@�F�U|�g
`Qє��ɛB^*E�/�BH���<3X��#6`�CW��J���u�n���׍Mv��[�5[������r
��x�}�}�����k�$��v��y	�1<�XlxVHYEB     400     180�؀�^�V��9} ���d=�q��뮷�gA��矬�Ē��U�͔qj���tfd��EB�c
D��Wo�H���8�0�mVQ�<��k��f{����H��`���*��t7Y
��.�]�*�f7\�/�o5����~�sc�:��-[�����ێ/N"�y�[a�ϝ���O�a�'�/Ѝ�W��V��n,BP���.�s'<����*.�F��M<D���Mo+�>��{�c��^��h�.OnQW}��~�MI-�e�9�	�onfk%U��/
~�?�1-��ƺ���95JT�iׅ�vG�l,F�j��m�����J����ˍ��wW��9�t���_E[P��`�АU�6���ʉ�jnt��7�+j�2ão�XlxVHYEB     369     180n�^��,"C���y�S4%v��AR! �i}��Y'?�=4��9�j�P!i��b|�\�s������o���(fp`�a�Og}��n�Ho=�{���?(Q���o6'��H�鿉�f��Fb��H0UR����1S�] se���i�`��@Ylz��+b�{��U�Y��I�6Ī��_t� ��=�O;"I������U�6�\�U��-y[��ۏb����q�G����\ʤ�~��H���!�inx�U�v�p�|����w0��)G���CW�ǃ�����L��>�'ft��5B��ߐ��Y	���"B�d8��'Y�>;z�����if���ޖq���-X�v2B�2��%;'�~��(.