XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>��Y|�xv�|��RU��bA�[�s�,�ݪ�Ru�ê4ij��h������E����.8 ��3�q��#�̆�ܔ�#^�?��&�qxs�V��x��*Zxb�-�u�g�D4��j{�O���c�i�I=��U��q�{��.\|��á�4bgc(��D�w\�T�J��[`��9eB�y:������Q�S��q
�?�q�8kL$	
!�p��4H�3.F2�lU�]vuA�A��3�n���W�<y&���J��d�{�~{�+U`ՄO��F���Y���[�H
��_ɬ΃�a8�����C]�(�c�#t��?A��"����K��[��sب:7�$ا��@�L2� ��R��=a�>S�˨��e�h�4��on�����i����F�5�/|��tU��*�v�-:!|��K[�E��p3Ð[4���t4�S ��#����d�4��P<�����R������:O��1':�2�G�B�C�����Z}�V�:S�m�$�q���~	��C��v5?2w��[qs;_gw��AN:������bm�m��6�;��
�طs�yz��D���O�M"N�o��� �
�@������Q�c���j�ſ�����NIz}u����S1���6fw�����'�[�� �q�#��x[���p�pYP �pgX�,��!5�"�&�x�|X0�y-���!���P�-^Vqƌ���^���@R�^�V�l
��0���L֓w��� ��8lW�9�vHvF��O�XlxVHYEB     400     190�{�e������Rgi�q�pgkc*N�ӹU=���oaB����}������t�hD���
�!��c�l7���+/�Z8I�|_�Ia��ڿ�'g^G����r�����:[�k�пF�{i"@�|��a�Q�N��q#�:mS �d��`ȩ��M` �D�ɓ��3T�գCRH�=��SB$�@X�8Ai	�]�6�U�A����N�해%� c=ʺ"�S��xJ�+�m4�m�*��)\zH��R��x08�^y�_��"���<�=G���,�B�R��z��zdi��g�1�^k�la�j}ۦ���'�钢LR�ѷ��'߮?���}����8�H;��|�~͇ɨ1K���$|�ێ�i���ř��iG���W ��NC��-3XlxVHYEB     400     1a0�K�F��5y/%�m5�ԗ���iV1�{(����g�w�L��|�;!#!x�V�A#�3]���)��eB���r���V#o������u��܆����<�xF$�*����8�HU/j6��7������|9!��A%���ކ -δl�;Aiy%�i��}��b����-=��������?�� ��t�P9A���9v��Z��I�~Өh>�R�e�A�j '~g@r�"�;W��.��6*�$z^�@SU��}H,�>x�'|���3��`Mw7�%բ-���p� n�nmۼ5g�:��>�3��|u[D�ޝ��ӹ ?�+����2�1��͙�Q��u8kr��eS,tq�:���+:*���f���Y���Ԑ�Y�E"��ð�U���f&�����)�(D���]����.XlxVHYEB     400     130�����Oģ7�ri��1���g��w*�YN���GA�^"j%1H�C����=�ٖ�RgA��*䬉�1�C��D�[@���S����+��w���S5y�gO�B��߅x��f�0huŐ9�OȈ�D��f@X�E	��n����6߼�\����`de{����qU[�fPW]��#(�J��o�/��5�ƍ��.���ܡ�ΥR(@M�;�kR�2>�3�Q���O���b��ҋ;S�l�����6�۳��l�+nmGj�ŉO�m�M�8e�zg�\�B��=��4��_��ڬ��,gXlxVHYEB     400     160�f�l��A���� ���t�.��c3Έ�&�U�A����- X�;n2�A
G��[�z^�ϱ���2~%�o��_�܃If��m)�=ˡ��$(��uM����K���N�-��c3N��ꂝA���zvC�a�&\_�AL�XJR80Ԇ��ҍ�N�U�I*��zV��_��I1��nx3̨�n�p�G8��T��G�h��b���	����Ru����o ��rxM
��%xȶ���M�jQ�w`�p>#�2@�>�5~���	�ޜp�&3,x�L�'υBCϗG!���0y�<�������\X/����~�ak�B�Λ�d:Y��8�H�=XlxVHYEB      3a      408�
���<���J+�����mO9j�׳�yI�5��#0�F�֣��4��Atq�ڄ&3�i��I7