`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
U0jtpFPxDzgLDzmBY+R/+TLbCK3RtO2PTUDsiAC7NDk8UaJhJIgCacyGUozypGYSHP3tZLnwevNa
uL+jpypc5SBbdgAc3M/Pig/i9qnWRG0MPgb80jVQ1YptInpAZnvDvEXX4feY9kzqFE/v29Ykv8z9
2jEzcXeY8S7gLJfJNZCiOHYwqSDJIAgV/A59hlj0s083SHLcWq08WiXcH89ZIxRNEtbJZHg124i+
xbUOdR2tuoUN5/m/33LL2ippL/GSdq57T9HxpEDtlya+QaUiuuLsPvuF9dve0SN2aSuQUkLHt8i/
/LZBekOH7n5SQ2gwT/F/A0lz7KObmKSapmjuCxdrdCh9orWMe8tQsSQoPcNWPRSbBI27jII1k+yN
W2S4ObL0QIGViwgLhNdMqpkeXL59d68iPz2j5GLBWFTZ6XuBFz8nkhJ02421zIKGHlCY5NGBMOXa
loYO4kk+JZvSRuPFgrwfAUS2UNSIL1Z7I+AVxZCuPVxI+fxmZeLQ0YHO6QRnHclnqy4qXowqN14/
TZ8OlGuE+kKYunqtoEsm7dcvbjCWOzglAM8keBsAx1d2futiIGkxe8fA0QgytcEe2O2LdEAcipEA
Y3OuF6p79ahp7KZEI9V8+r4Mm2WjQfSvdKZPCb0BQUT1iudIU1BSBAvH820u46GMLBislnUNGugp
WrVVOGA+brK1Nmt9XkA6wLyU635TMQiBN8yI0WPiV71p7ntEwDlYDgsKhQ5CVBPRAkbu1h18OFYg
pP/tJUna/jFIdZodKCf/UljAN0gssKx5+ZNrepQk/5SHhJrsNXUDay+X2HA02ruJOmzcHGkOjWMp
mwK+ZS8ObS8EyDHQajyVHgW21Xuzagf4P0lUp58BJB1r3SMkdOSVe8igrNSk/8GhOj5wwOjF4IXw
nshldYPw4MTKrhTemyIv7Mzl7ndvO21cTuqfokSQmCdUhDiMIzR7YZC/mUyOcDK2b2q3pFxLh0tf
IBpglU8hCYu0bCYQgMXJWuVnjTaB0IhU8W8ByzJcunhAAuZO7E/NJcAI+10WtbH4e98c30d5JojT
6hKSh0iR9BL6uq7LjLn6z33WbChsHfW2k9qbH7bwNzI0KZhMKt437LZgPZfM55ndCfXb6M8k24S/
JwoWpn+CoorQKzXWeLOCD22bqZDgvHaJDMCzJllnW0OPCyaPtiAqCj1iXQjt3iQ2yicdQTsA8YqC
QNUN11S3gbgmal8M9Zmn5YgZ8ToAbGnTd5ywoU/+1LyDamTxOolpdGUmRWN1lUf7fOtoGPBknZ/2
duQcFMdYJra26Y1x0bw3xPzqows+Gv1UqSES3gx/v8eU7CTRMLPfaQ6K+wbpA2QLh3jt+uK60t7h
IcqKQQBeCvX30VzIPnPAF38eni/vEP89sxcO5HJ9TGL1a1cZwvV6eTo58SvTK38syHtiHOSw8pvI
yL1MqCtxzDEO7M894ir8G5MOllKLots79lCSuNF+EZWZu8jFepLIl/b3SaC8G0BY6DpI0itwOaJn
M3USVl/5DitjOo/gWZ35ub68ap9loQ+CSc0UnwxXpsMEczMRaJl1xyKFmeegTRKzo05vnernyRv5
+V2ieFFncp1lcT6qatYtZHBOIhWn82WpwloZUg2QizuDAbCV4fdzwTVhQTY1FCptfkrOyZYcmL2T
q+whPofH9lqiLLkP5j/Dev6cm4I/JeTFjtt/GN43QQN4QOU/wPBRpeSrkYy6AXkAMlWs/u5e0ADe
ki6J7c7EzbgxzW3d5iu5ppxbu6zjOYdwcIiu6xGvmGPbQLaUhtSutbfoN3ioRwaATLSTvl/stCZb
AE5CVkJ+ekiUWIIW6e3vUWiMYuJasIJNmv5vKRFeSb1kjjHCwtiezPQ8Prdj3JI+3/2fhsWQuyoz
N05mH3QApxNe84nK/DBrYQNJlon52ujAid7vGouZeuKjc3J4cxrJwj3MW9Q2pCnRVPv6nGYSN09J
w5RhGliAzOc+Fcxy9wAcpfKe1puIUzr7dCOn/1mrYlLyuI3kXZ1ANvILgAdNZ9O+1t/XcLssyApo
mOKZhwKrWXuFIN3B6iJ/VujtsGfIgcgPDWqxWlltD+usewmWA2d4ddc8bCIoVHh3wOOR0OXOhsFB
m2+IRpvAVFR5wB8nQMmbP/bZtzkrFxUxcORK856cS3atQ6Z1dXbTQb96JrQHMymVJqk5mELc072Y
u8/wP0Q4JQbWT1RVGOM9r7+8mq8Rm3eewsAYGDxGxkYyagll0cicDGZHiax2yuZX7aj2Rct0+4b0
LU5lXGQo4UX401JCGAGJ8Te+u6Y36ftmkWhId+AY1NxPvjVbUWUALNnqgbQ/+poD75YblrlqRWRL
qNsHud7URegXej1IR6mDXO+Xfj+wetl4u2KWM7jc+tCLd5uZA9B8RUNpb/QWlGFxW/DT6nkb50FE
7SG6s2Ejc57AYQww8w4MzYrZR/XmldsU+f0Y9zyboS00DREP4QNu0aXPUhd2kmLIvvpCvVtzb+ws
d4p/sZ2rJ6/K+2Y3sOd7y+sNXSZusLqR0HXIK0ru9zKlKUSwxVgxT63zpdwaqZ70Bir1R/6wJqMy
998frKOudh4O/zw4T44IcO2/asplpO6PurwGOJ1poRSEywnGIcpCYr+FBNNPSKWyZ9GtYo3unj2B
UDI3X6UE91G2ZlQIPlfV75m/ykSUaowlA7eCVwMv/Oo1/fNALVEbnV32Ictg8Eqz5kT9koR6Am8p
sGZ/odX5m+91p4kgTS9dhoiFCcMyigtrUNpvTUBAjQj3LO9VAGMwrKBkH14hzt7gBWXSMmnHPPNy
CgpdbcBdYvsg0Og6/NYUHXr73fcxZpol5m3FtlDhY89b20yFLhAPmGaEohz7WDU9sP2dNEEX9+WZ
8lGMCzfmhBX8347MzfSMTIAOClpgiPfPI0MBb5NTtKjlxHietfcZucx/hYPcoNt/5Jdf4CFVfOf/
mZtuqXdLZa1WRh0bjnr5FhxTpyisFA4K6gYeVCgPvcuCkWEsVxmt7FBXS+vsoksJ5Whb4Cuf7gPK
o4Msku5VefBruj+Ud1Ejo5XZkmBSsWnfL9QkwD/C8id7hpeFbyryeVNKoaenv1b5FRyroEri+7N8
I27sv4V2yW4Ne8tfo8gXMJbpomrRv12SR4gFlEIMBcnnXNbwWUo+DAuwpnyv0AJ+tSe7qAZoek6E
NawMeVJ9QmRdKGb4t4f+XpT0iRUDUXrstJA1PAh1n9K7IogS5z5oCq/lcAo/xGcfNsMd6g6scl3F
JZJQt8x+V4+X4kSWfWFwrKynpOHkG3fMxVht4/2tz2l7u4cDs/ipN2wktf4ojBhWOSE3UFS7t5DM
B27Afki2B2VvYrRRjcuwSZCO02lRNqlxzG0Kdx1SfbhgIemqCDYr0408Q1kCml5+0V9/vC0SJA/F
2NwEMg3kCn3e99x4ghOiFxHgwVXl4bJ7DNZExbytwMP2EOmyY6ciLjXc5hslbLuG0ML+e2cXL8HO
nlfnIGuO4jIzpVXu3iySMhwjNcxGQ34ehiPfDspgxs2KPZikzf03hSxpk2aUZOmqPKIlom5zIL+u
3TYf089fitWbeArpZHvpqbdL+C1E0LSiyO9Lv7hA0oR0JZTwCGW6auYy3MvkrwYwpbIbIlD4wqEL
YipfODlL6t81jgzSxzsYE1LPz6w2IwLPXtnOYda7VDsrY1W2JU3acB8MHrcd3DyTNbRIjgm9ehOj
Iyk9cYl9b5HJks+g5m6rvCv2k0T3VGBQ+YZrJLKyEO/H8+cXLwMfRCmFO8ULWwCoLJjbP12Im6ZE
rFhUem1w1nyf47deywKEISG3lRNaJV5jZbBMM/EYoBMEpAafsR1aUCriwD00j5iXmSJj9xnbLEp/
y9KiU2WgTYoEeAS3EyVzQuYhVdBUoU+qyq9RsTXUzANwkFlJv15AP7UW+jGJYt2CrjyKF4ilOi3w
q4YZn+ZTbj8IjwT3NfC+4Qs/9TQL7wwSCVOB5S8uzBmYS234fp1g6Pm80MK5LITo185kNX96doPY
OD2JEjTWEPhkWzbFKtfFTDHAKDxfyn9k1hEPLBuQagRmMlIeOSNHjH2e69uP8bfbfJE/EaGJA5tl
KpqPbFCbo9xEXhcvSVjk2XSSwWVqLlvutUt55mwc6c7LSh7+s9vQYthOOqpjLbCQ8p/yjjlDTtrw
Lzjc1KOHGOLMQoaUM6uTn/8MHkKRp3Dgm7rknzWjvviCGcDcP2KlkfCzK20ehHwoNFFKBIsMZ8Dw
+RSbJjek0PNLn3ChPKNs/e/w+YAgPbdIqpNKmcyGvC3UZk+LqVx/u4ZHzQ3DF7MjHPKk53X1QBJY
uB30GBdLwn14RPKyM16XO2HlNXCoi6v96ivFlZoOBWlM2xrPnaSbSIAY65UNlJaW6gKFVvWM2649
pPImWbGYqY7OaOl6Ac0ewJ9jH7WYZR6Q0MFTnnMkyawrcAtnObdtuJSzVxaL1hsOAakdHcQZndO/
mDqHy2jwTFWusJFGewZN85pfomM3Yvge0vb65u5SBDCQ74l3n+MFBUBv8ocTovggDHHC2e9zwu2v
bCwGIdWKf8QOdSMY1LZ2bdNwjMggimIfqdXsPIHRjYg4FrtIR/OSrcpHaTSb4xyVKSkszT1IO+Tt
cniq2wNJk9gB/eKJjbAhglG+DpGGmqQq8f+X
`protect end_protected
