`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17472)
`protect data_block
qV40GFwMLlkladyjp+hCnYFAV2kKk9JUnmoYFu76aPFETozIQimxgfpqUKsj/7BOl7MkobgMYHcE
1wILKqNJZunLUHloAJQNln4h8X67uplC0GiTv7BEBQW4YuuW7031zid+Cfosfltkldi9JW9RCdSy
aONWDQAkbci1ZlLWq9ziWlOrglfHbHnJSYLVbHLeGhLCkG6qJVMRzW5vSv+QH8Uq/6BufL4H4IXa
4O1vZFFBIlrNBpO9JkFMWsQqv2rMz55xZFxEvVs0Cv3Itema/Ad/CJRUqbYswaNbqlK6nydxSKVK
B8rpNZNgBYY7jPp5ANeT/nq2bCcWwtVnaajwnra8hdgGLjsEHJtKHgfa7icg12nRXoL9fDVwyIwH
+TlRGotTzlO8MY0u1/TOmV/izMxAg5dtRje5Msy1F2lJ7fbxjH9Q+M8IB1Ifo1DHxBaU9uKLCk9m
6LwkZ8udi87hlGh2x/VM4/UAcseM2lLxeYsB3TKKFS5C+mC0cQuk21DWjgo3b6kTTAMRec68VJHx
GRMnWEC7K3s7v9koZMkO4Nkod+gtqimK5f5KbF3RL+hbFv2NVJBmMtBaym6hOz4k8kewqsCHqwc2
36BNXvE0FSPu8FYCTbKok/KqibfO5pe6VQtEUixvYSiTldbjVshSnkwah363R6u3AVPVfUpZpq40
6fyNTaTxxIjLl44r+yPXNzYPxtSdcqJdGsRA1B0iY5FqciL556zwBzG5hfD1RbGJEMwKYuIpeZMO
7mUM7l4l3H8Jw6nwpeKRpuRxmFEWaVDp4KnsLkOPQwowngOJaqDxl3+3GwpmgTOuA9VkZBP9kN/s
T0sx8vjnzgB4I6H/rSOOGcf7l06baXDZO5JpTg7GrMuUBOaWuK9NdFHFGIaBcgddFp/hZS2Dh0km
0rXFnE1aVmbmonQ1h6TwVaID0+rXTGzYAdo5wDHd+DlOb3vpjcN7UGkMWCpvGjEpmrl8Ixxi2oTR
XBhtBHic04irUMdlCmcIFKaIMWMHAiy7jMV+MSC+vzJ3SdqhI8KsmXvwXzTjAKRjB+RfCNBfFjlb
b/P0Hc43EhgQSr39LW/S7SpI4B04DsbZKqfX9PiE0ngEuuzML9FMi5A0pWB/M7vBEJbVix9LwQoe
+xJyRwacX6U/Jz84OBqKJuLbrCY+kQIhE72FV3WDL5y17h2RBNZ4puP/dXSUI4SCh4BB6/DiVSgu
eFPWlXOBNxfsBRtOahQbQ/5P3jtC2+9oQd415/xSlwDQ7nXiaIS8LbCl1Rkc3RlWwkwUo6hm/A3e
7f/El8P3t6zWjxaEwrlcZeV+RWvPeWyaMGuYaWGDNX1plGM7UAUcKpeMGTg5NsSc013jlwyIjd1Z
FGnEGkjLTyAELYi5l5HgBhgu/1Tut05I+A4B2uX0h6AEeBciABcKfaScwgS3xMj6ZfJKEGU1Jsv4
+UIxeT58+9UmpY5pKUeQerhaJLnhaq6jMFgQS3MSiz4ja2aUi45a2LUH5HcjhUfl7mzgVnwZfbcB
X+EpADt0AA0lGYEqEYNah8g2sRK3A9m7jK5DRD0zidN5Z/yBQvO1buxDcjSZ9fZPYdM52UEYdrSi
ZV4Mo7zxmIhSoosAKwWQiXMkKLRZlIyOzgOkwPeqDYdZVxmHoM/KFOpsHU+OtmU5/8peA6Ba1DEh
UX/6Mqn4GL01mMjQVlGTlLgJcg5e21k0Li3dlVFED2cUvM2M480EHi9aAeiAdOTuzDcFez9YFRnL
c2kx6zHqla06PkVClZ9ZZQpQcwJOIqWoC9LKUSy/qGesiVXAP9ybLh4iTyZwukOBNTWOQByYWvum
c52/gxwXGv+tmWYtvMCAjoPUVmXfik8A3cZO5K02rNqylvZJtUl7n+wsZO1BkBp+oe1IKXu+Oe6H
HAwSlA0edMizBx/RCcEduRg5uv4GFSwjir6d71dOslwmRxYD0KW9lVFtk34Z4Q5GngRyjbUebBYl
tuH2i53uXeB4Js0TeNAZj+zWatC/GAw+jtlY+qtWqr/KIoGJ3Q0n3gdIBCPP2aaFBqXhuhZpCVSN
15gQBGi1TlRO2gLuXBBlbb00TZyIbB3Xzu6WSim6Af4mjCvhj8ErNqa7AE8eP2MGCvn30zQ32Jda
zwGbzqQ9simjrr2SWg85T80rqpbstD5Hyyk1pQEMadiWCpHQp33AaI05X/j84hbks+fpRHiTnDVH
xpeFXA8yy5ep1ceFtzY0bMmeVhWP6MJCOhNwNJhBPSSaGjuPYsCsCFtfdn83kFqZTmXr7atGpo+J
7k9om54idocv3HhPvUs+1s5zt9+gTGJy+pmoE8ptzUvI7Hxm5GV0ASTaPSmUIiE3n5GuSJTP/mK1
JGOpz8BJZvnQlOTH6qSHjqFBymuI5YaRXDrATcqGHdR0pGu69dvwZsZ6FilSbX/7Qr52xFahAUjP
jCYtjwhdN2i1FfwPnwKM36D7Eb5vzeN5KQW7buxrDfK7+kgA/DgM5mDMnZje4C1ecP7dDrzzF0Kd
15FxEmO02394q/CImZjw6//5mll2W59C/s5Qw5MtjzF2t6OCFkHrLx2Qf/ku26Ae+Sa+mJz1l5Jb
RIQYEFfINWaCzHDI5ZpXt1wnjqCBKBPtymvTTygMtKkECkJjsBatC/kb+AnNbCkslut0E0LTprNX
/0AcmGP3uzmXHp8f/gWq6eIBKRUFTmElfvMIg/o1dIaPCp0WxiMagMVo0Jv0tJNklM5sdPhtpV6h
bM8UquphkuXWedaSdX03XdqjJh8M08vD0lkLRuHfVsXEncUymLKp43+CvJ6Ly4TU6skKxjLTkETt
oz4+EQZlrmEPBPWubN3Ssa7/nA80+6aLT6ZZaoBGWDwv6dbuqwTY/oJMyrdaBPople4kKouVpXxK
hMLut+2HkeBGwLcZsyZ4KYvG1WnbXi/xneipGsBSfWNs+8aNYq67Co2aGmadNAO2TKaVilSjX4jV
FGLtnp6MtTbNoBUpoVBawazK9FXs7tlPi28eyJVwcticwj+UtVflEL4m1dBgANgGgzOtl5tI85c1
zBE1FvJddYErnUHYrnqZhLH8nMDy+RonWC4Z0I3hpaj50TinbVgZiYmJmUq7xUg+lSm6dddI1etn
IGXi+iTph7lTlfTEpUuitE/aQcQrm/a7kkMn6SH+XJvEFToBTltcaZ+nBPTJr2p3xoRKsCDFOyvF
fS9kCFhBxPzxoyKRQG+q7/NpHHKsiSx5Jinl9ujg69QbEztgcFsAtGeeFoBvXmVB5wZ12U/IubEy
IMsfp8LgHRVGTMQqcNGY9Rt4DZIze2nEiiJidBrYpFWXQ4pwXxx1jrZObonThRKm0vNc9R70MhUZ
7fyTccKyg/ofvYFlr/zwgFxvzChiWrMOqL/O2IO8my9xcuZI1qmbW76ufVUHPKgQ96Z9kmpMQYft
IJxSpi4zSGMa5YOmx1AQ5sVXXiKtRlQm0v3R0nnhrus06fkwT+14Snd2WesM5yMGzgsdM12lQ9gt
U3UCYa60cmGezixiS6QcoPJPzr4pKbl3WKmMbxTEjLsI2dqm1o2xegnxgCYwzzlt2j0+rWxOhSjd
VRb4dLJW3InPY6+vxr+cCIk1StBWGDN8pTxfdr84R32xpkvcK0ce7Y92u5HlycFw6YkTUk1swamJ
BmkjNus2s7entZFxkCzwsqxlBvT3QUNnKZPKP4rpUd/b/bJxxAZQrHQX1RJ77Ws7dwDJEaGCYOhG
7HH7pYIQj9XXfiWqMEA3TnuTPxj9FXX29Df8CAJNsfKq/YNA04hdvqLqXhaKFpQ48U52YvVvYhHH
7YYIEF95T/eWz4ztrLCfA2fiM5svu4olXWvn5Csvjo3TFcEtIE6GjofAVgRjgF+V9bqjGSSPvpV8
41LEjQ+NN4mXjqPtJvltXbKwb3NGT0trs9Wg7JXTldAnbdmeV7RlNUpjrAG3+tgWprFQQzyfMvcE
PYxhsaA+dSQV0/r05XSGV1n0htjRhOXQfxrAeUiwKCf7hLqZdQQE9tOeb2UA9sRFuFkQY4DSORLc
1wXFktbjjUkbsxSWOfApkHWKDPPU1Jm2H+QVjMGlcqFAsY+LoO5RtdnASr0QQCEbvJQSFbtXsj0Z
PeRe7xIFnxh4hZnxmZCh0cWjd9L5oAo6UqAsYTslNvCkKaA6MLoKEBQqOI5ecMbKGXkH6EfmsDjl
LWqXnWcd046okZmiFMwzcv0DoC3osY1LZSbpjE++m9xRHKGIje07DqKeI7uh/GYidUEpXgPJgWIZ
jTkcB0BqjPKlJIMdlQoAgnXXvXAEwcZ6ea4lIOFchTPfqdvhz8PeRF0AFDKXGk9vI7E4YUb2Kk/t
65Tgcyd72N5f7uZJqqUosmYrYz/nCnE2SupSymhxvlPi9NTaepyYLHdYbD4UZG2XDSfOldYLf3hs
lw1An2bG3bgA94CtdvFHohJrByma72XKygjqlFo708g10DR55VNmeZoTAOyr4thH6Hc2jCx4H8Pd
brNIADAYH+1eFmmpoZqN/p8cbUV4q1vaBzrd44Xq0VrqProAgeB2gggaO9OJUszk2EiGOq2RMs/k
Y/iiM8q0jV3K8DmjxwYx95g8BzGa/ExSuuNlltgvmM22+zPIH3N55C4UxTNUhgetCMYzNtlXEwN5
Nglfb2envsk3tTT5TUPxKScwmU31tqq/HMd73gX2L/dCcRN1/o4ZPYNbEoWYafHtqL/WrdNwi09g
HZji42QlroUg4XixPQ6tChh9MrGcaxcYl4m0U96QSlWLDCU2IzanFxSid9yyIh2bk7HQSxZMi17Q
NCGV0ohXKYZcA/TP1UktoJgtrq2Yn/54S2EJ3IdPAl3Cg+ETXdgnCpvdsYkWbROXAIbJ7pY9coMM
/66BeyRX/7L1ULFpVn53FQWGHJMmrI4Qh7wqdnc6aUIqlhY2AOaNuay7Vvwhbs61+VeaVdSFY5JJ
TRjM9Du3KLzwdaWIVj9r8M6sYxtYLCgPF1p6oWcG2gz7grZC41TrwKDyGSZqy43Ad7/KJJrdfDSJ
VPQ/7xe6/PmLj1KiU0PUXIRnxnwMX/toolssC6jsoPg54P+j3v0f8l1atpcv2TLW891S5tgRRLdx
ftd/l8nuQohQ0a7jcd/Z9WAj+1b24DpRyEQ9eWmRtOCW7g6xgBj24KZW+/EjHLHKWzjAH1sPfiW4
lWuHt4KhrGEsABx3h22nnQDQkfEcJ/hfmlMqnu7q2U3+yxT8Su46lFj+b7pabuGRmu1VFvh34DZk
gcCBSSrfvNQmVuxoVFAtKQ6teTS6xqtSWlZ/RJDmJeZynJB7wjbsKCBQUJSga69XunBf7On79kAy
AqZ/aWqyOPNtn6sqB5uieo20xuot0UYeynKICpuC2uA1SvxzcAAsGZfG97pObZfwC6ykzL0olaZ/
V1QU+yNDtXsQ0uoaZKoSDP+2jUHX4+Bk37IfwIp7FvhR/m0BQ2XU74piXlGS1svQ7eadBqhoFaC6
HKOq7en3Py0q/g45JlYpSeZCcOcoK9yxd3yorVZro1gdMGOIBkM9s3+Rn1Xrne8PBsvgxpDVhjZf
NtWKrXb7zbQlwo89KyIHYO+Ec7NMf/+8bYVNLnthKHAruRWy9cOimgyNJvzVUPrynq/PFYZgI8l9
L0/KNZlMWKmW9CNUC4F05GfUBXI9lIFhbNyGPBXnHYE1MYz4q60zGVe/ouxYt3DID2P549+jQ3el
lwRI50IPqBJyeBs5aSsv5WPcYms+bX0KIOLwyL6mOij9CApV7n4lk0khThpwe2N2evkUdfGyatfx
jwO67iIOxYrD8FU5Ckxhip+LbfF7uIWyyAxVhSbR0ay2xW76+9fMPUmIH9eGiDNOoCFjqjpyNJ31
okladdOahM8nfZswCpE766pDkjge8hBSIuriL0MjGWVp0Y4GPSflEOs70AFuCrJFA9hB9B3PmLCg
+mR5d4c2HMdFi/CtlcSsRJKBXB5Y9ysNfQ1tizGUYl3NDOGXAbvXvpYlltz+B5WbGLehIGIzqJXB
CWI5f0OmNDbowqy0YR9Xyodnx//5EtYZq2PyntU9JpL2NvOySqRvR4D3POtqWcN7ebDj79EufXrN
sJ6+zV+O0ldsh5cXkpZQxtQX5mgsuxqZHhH/9rtFKnMMduGEHGtgLM7XSUmhXUVAcn7Ge1U6iFLa
mzUgonhMbaJgRW1oZAkDxwkYiPm7WDF8goFaYgj3ypgVO1xcBQA34KwGazMOH701NXDTySVCA6pm
8WUBvn40d9iWpYqP5mFcctnQ8xt9P5hjWEUMpwwzvXJK2Y+EUe3m8q6HUM4vuoZHFgsI7lY8tUhh
snuu8oZv+Z3T6jGRpvUifB3e1XCsmqsy9Lu3RkYAWp0wzYu5xqapKqPhMuIGJ+m2KkKm05kxva8Q
XPLIFqeqKPRA2a5smjUvYwE/pUQ9K9Hk0dqVdYtWp2apE2gQH6PjyegAQ5EhvWYlu0XmhJRQcRsb
pBsCy921PofAxEn32i0Wq+gpFAYDpqMZRK8lgZeVlL/8y4gP4d2XCXUCJRwXq1BvnMkwf1Eanwnb
aLLMKVYNB2vpVYpm7Ir5v2YbUUF5ARv2os5AAjqlD1YpZynVPSKT1RUoURL6eK8rO2SqNyVJnd3g
u2uyZbAMomlA3BwO2QWGF56XohA3XyhPXRyE2O8fai8RZtZT6Qw9RbEwuaQulkTj0zfjzFSs+lgm
kXKGmKGfOQ+CDYEoAu7Oc/SOPPVoP4eaJVUap8we7VgyIiakIv7lluTAB7yJBOQCE3JGLRlnK8fA
PWyBXoUv/Em8x2bpZ6mnU97xkQC8GadJJ4qUk47sT2f6K+8QRq5ORlpwhG0HtnAqm9YTXd6ZLiVt
IN1ByYNhFuVufD/Gt1qDJT5GlOIlYymLZ60OTYKrpnmX6e4Hwz6PTCZtY0zDicxk5q4y02pInlMQ
X+tpPVtSDCNlEgS40/9PdLHmDnvJeHKhF+45zm7Kfckvd0WMxbEUxHqcmQV1+Ssd3mPOpU4+EfbT
qP5nQifJwXEwmoOsuLOdrRqSO2f2PePILkvqNgdQB2EI7gQfeu4XxsyBab1ylR7qWTi1OGxrRrx1
ZZyXu4sx50ce6gNcO7cPc/VS73AC1mTmA8PeMLoDw1s1hPkjNpMgsyMiiv1Pm51icRFlDT1VlBIE
hpdbYpJziok9ql2pGcgmd6fS0wywPSdIarI1lEYldf7nMeEVGTe4dMNJFl5ODCJ9ln5bnMm/iwlc
1FkHkYy1mWTe5+8dOoQYQ1hpyvwe+CWJvHKvuYSpdRLxAe47to7iP8t4tH/CN080Vjzwkq+fMlwS
U6leQoMtmLesac3b+RjdEs1fyJlshDmizLVf1UEM3GuYCxJKa46EoJ8VN9xbYOewND6ooF0DcNP7
EL6i93EaNolDCGfUKUkMBvUYF7TuDVwnRSAxqTxknpaN5RvTl32nOxIw5ETtwlGN79c5LLkecPMd
7sYPFw14pK31jS1d4iWn8ZGGVI+urfkbMG6IPQrh6ZP6nIc1AdqYBnS/lVy5U8avG1KEb03/iMuD
3eToGukr4haamUJdl7zYVXydjnoAbDnhOPHVXQ4G0BNaW617+tc2XqFx07CYz4Yt84UwgrHQbYI7
yKtE/P+HO5HrvJgvT+YI0aPW2bVGs+tj3LOcLFwgDWY0Yqgg5P+xUBTRz69E1n01xNOMytlZNPoN
K+lam84xWGV5Y/oPyTwq6Uy2k5Zg1ZCI32yFNoLWjdK0Pe5TKvLIE+NZCdHvSQJ7VkHu7Y/uaDR1
VD8cunlrobqtrLEbx+Rj3ynl0ONZQCYFJ5ZDuDqkNl+bIkuJNWZtaaVntAui2p86mYahdoAqp778
55CtXz/zyML0OrTy6AZfvtMJpbIcc3UlWZSdOEbIaqEE/fejaEWXWgFhGoqTrT386dsLIong4oWL
kCF37p71XY9m5AtRYUgTTW9MCJOzQv4f1PCv/EsLypPDuco8EZWZCkjwIlWtmb42qzUvR5Ndb0F+
Cxwzyn0fWksNfaGJwt8DrV/RtHDPJcMCxzP8cftU8LbRp2OxiGBYSgHgEgCRdlvnAGmVTxV3dDYt
htjZ9TJbEGgZ1erWl6Y3ULAfj47eMNTp+D79XlvaXfQhEyg5Ocrag632Jy/q8miFaeisfnHvwVsr
r09Co8usjbODewpJW3NKohxYVR8LQv1L5IxONO8N19U/rSErJwDcVT2k5xe7yunvOQKv4CVq5lyV
IBm/9ra4PfR7gyckAm8KEMrlrHogLpuNGvGFhse8w2oPLrp0Tcy8/CGEAYjyNy9geijuz2b2kEhS
NV6NAJ3nsmiPMFzmIe1klVU2rmfA+ddIIzXDHxH5l1Dj2wHBoh3p0g9l6rtRitkIYHzYVQnzr0yn
+sCVHBdCcWOFF+p3H7ZzLeqVZGEWTEJaMe2xrrhZtD8SYVywXVYiwkuDdlE+p8+l4y3XMvnjT093
fk4jsExfDlF+Yw/ewzkOd0HRmjuV9BhAPQK4GNEEcUupYLLSyeQ9LT/sU4f+1KNnBAJqOj3gwEkO
gaKlKTA8q9m+xuYCV/WtGGIWbGWoWMWZxuqME8za+HtjQ2sf48A938Te6yksk/uVyoybJkiXGuE7
9oap3vFDf6fgj3JOwC9Ys8/qyXl3vMhrLRQxZvKY/TIHA0WKAjGlj9QmBpBq4HhgHYkcwsgM6/4B
Pe0yFt+527Z8RQJdVxcPdN/b77wO8SIBIaexg/Cy9eB/8PFnUbNxaXegj1WcA813zLAehArImsyu
stBD4JbW9h462T/tkiX3HTNOJxrPNctV8Tmx6LqauBFCkDg5HyoLpS+IbC4qfW4Hb/zyUe1lQ3vL
CYvpazvh2USf6A+hEXJNbE2f3S1ufFS6u06RUCb8+RgYuGkWwMo8oSQOnJK/9jv4KWaMzrhu6X+x
jW1uSyRFB2V9viPpUluoE6v4S9JW5jVRfm6pzoFAXqs6FKnmwoAklg00okvIKMqyEYNmQT4d3h9g
GixhDogSPmOUwNBjvAiPu2m5UZCpAowlWgeTmQpPD1vNsMKHt9qZMwX5NfkbOHe56ftNnUvehqOJ
CTyQaFmnwGzviGK2gWkgj7pUbd8mW8CgYIIVROFpsoWGdNAEK0Nhtzpq2pxw2J8u4xeyK1bNR53b
cTks7lH4BjI6rQUc+Udind1kU3MyRn8h0nUxcGbD0m+uTHytLHdRL4v8cVG+DqGPGYg+F/CyrF70
zkq4CMSg+tpp30t+CfGwClkM99dEstf8xqbWI9D3cVltIc8w1bwTGf1O1wYgVcL1HbxtOAwILMgp
0u/5EciCxOEfpj+pSGb1zitcLxvobByeRjT7esANOFqdclv+gLEUtwMkh4nb39VX90V60/FUg80F
Aghh+MbywQOdj+DIy9NM0QHRori+5jss9/XkY/JQdCWrk5lAbwHN7t+c5Q30UidWUxISmhVgKPxA
zvQ/foJrEBc2LmD/ZrIouNhLRdQ6G6n469+0Ir7Ry2fy5sbKshK0r93p4yCBZDZzqx2pKuXhtiBM
ZwdfnFHHf1cAIYsbkAHOlcBbTQ5BSDBnxFlowbVewdokHpkovWbLdOCrECc9UZVOAPUvk6pDUEa7
M9NV5SeIB+Sif5N3V7Zku1+ql6bjdboCL/6ERVN+eFF5e1J+aEeGEo5SU/tm7KM3sbqcNnvtQmOm
JjwBJsDj6i+6LrqTDCloIyPBLsD1ERGq/yyO8/E3IRJnnTPC7YbjtJajQGmHwjk0DCGEEBIM49Oa
SIQVC5mSXxlO/NfTFYGyaEjz8J3yCNPuf2YwcHKeRF/QXwbViylJ0PqtsOAD5ENV9oeiDHkuLW04
KoLUsHwNrmXrGwckHc3EspbyqIH+dQ3m0mrfAN1Tv4GlySMcq7poEFPF5k05IdE/FEU50KgUMgaa
5b0RHq3t8fhHIZ2BSbZZkOCpcyH1F8xjlYXGJCiyn1nU1u7PsC1CXNDTXjmu5xy37PBtzgD/91FR
NchqhrJWsdYlUyDxpoe8AyaHV7WlrODAhxvC+1r5vgya415Pi6czz067nELJo2ekEQZMKbvXwS4a
v0iqu75/HeBdNqAeAStYFoRsAJVfyKXyaIER5mrPIERS0AT931GEUqlbhWtYgohscba4FKz7Ot4t
/mJiP//V8Jy2j3jYOK5rDJ1Q2/3XbPUmwBJbo9uYYYquvWK+d4h0IESSb3RV1XnsBiMp6MrPCkuD
aMXdeUVc4xaLIwojWwoSR7h6IJcJTiP+mIYzOf+6meYFNqrGiuhf4b1nvyXDIdGhJX1F2w55679a
VBnP1yqzX+DMi3FGdX4noyvn/qkBKZCzG2DjCzjl4LPcJA7D8aC+fbTdCLwDTswip/otzAs4k17E
KLfAMwJvp3zczML/oXeGYD+FZrLVYETfZxVVjoo3e2ToGx11D8mS6scstTYnsLF4iNltqTsoA9KM
nKK1/Oh4wlWcwleY23PtggN9MHN3LZLrnm7xgPHcjLgu9FL5UZPAHjRf1FcMNjEZrsbMq09XOEzX
bCZOIvshzVKm7CV9NpPiFn4kGckxkW/5woACRFb7TCugKyP9Zhu1FQRR4CQIfFa5jQsNeE7UJ7Na
mGozu0TFW6pplDQ1TqNbGqHhPOjSKO5KNoZIvNyQxkkLwvaU9FfrwCdEDgj1V+xzSwYp13YlAXrY
peqTbaVuoMz3DuKYdhCflrlbDXNzMF5W9vWYmHgGtEDlQHqhVnrEQYF0zOlAmmuIwCGfuRcKEiUx
RUVPm0rSiZvokuFb2G84aAPd7N7dqrPsF/i+NtrlWZhu0Sg6IiTxIRCd7mn58scctDzlQopE+19K
DmT7fk2MBl+VkamzpRPIbZ5pI+eIMcLStyfkBMpAaPBmdvAfhwlrAJ4qqvw+1ipdOv2IrK2sP8fH
Px52ijC/CZH3VrcVKgG/tpl64NH6CuhRuTFCU4OMFsFHTAlsb1mrqukuD7N2703Db8ji7jbW4Fj3
xvIdhmXJkywNC2PIrP6zJgpAljosDE2gJkAHccMga6CjsRIVaAEbd8V1Aq3C54Y7PMmz/Ofe5uRA
pMTTlsn3iS83DbHbloA5WdxWVFMY6HNxVJpmwKIwc98Xaycj6b47mpGfYsa8gOlAtGjdT810yUNv
ehcK8cOY1PPRWmDdJ+IW62cOuMmhejQMHdxtgpN2eJPOUjYh0OcQsUm1T4DhX1wb+6tOKJ5fcIag
40YDVjhz1JnG9YNI1oE59k8BWEsp14ZTQkRUj1kO8FBZVO+WZUGzf+rkOuePIp/CT0mGF6RILKnX
X2sOLsGKfsf/HJxrYHo7Y3ng4jEUEAgM3bN0iwmgIZkksWyvx+uGMo/VJ/ienlnqKfTIAirYih+V
N41UnYU6goOil8bO62g5muqEMJy3PwkTWh4UVziagHYVuaYLJvj03myttU5vHHt+WhU4r/KLlMbB
5xVYC5kmSQvDLuiKZgqDlV6IgcKefuXOSKfdT5Nq4ahgvDVEN+XsE7T+LfPsl8HFPfoeVSwHUnel
Aa6kvHo6QFJwmBYJviBbRR9JsbScu7r1uV+DawmOxJwFca/A+zfCBAlYE+/PI5GQEt2cMjROKvaE
/qPgfPKmuwZrJA1MF3Obg8TCHSOCph1pP3g8vyN4ycJd75qSADyOFcUP1PhWYOA2xyJxDz1fefeJ
fkuQN+kZZw6U0jYbAQ9pv0jhQ+Ndu9kY5KzEKr6KOmiQ2cztFIOSa6lyPXO/VBba/JECizA/tnOC
CoTLmnvmRY2hEeoNHt1+w/hR3JOq22I8BYXmruzpJKhK8Rha7DF0FAlwMHMKUV7vpo8o/OR0BhIr
bSdeiqKd5yvjTDh7b9QUHD+sCaTZHwU4yi/9aPv9TZ9iN1tNoU/eKblKVrc671AFxyiAX/RHai6j
+6bTw8S9tcVEyYgejQRm8HoeRPcYrxndHagSkx09z5rKfJs3+5STghRydQ7lP93N5qjYsBqXqY2Z
EwXVebSZ5Baofj2flZ3z2s7d/O+diCf82+VfFPBNaX6F8heTlbKaaHBVpcvBIL/zgyvMXuZJFrkg
7dRQfe8UZRnsA7TqXFoZToQniuIdx4IGGWeRbPELlHksk2R1odT+rlBh6HvKl3rajtUdAr+NUq/E
5mtvildgRRHaL7jZAoOYY0TiRKUCIHHCDcgW3XjucvrZi/9f+08GEAfxzYnljOAFt0RL7cNV48KU
EVYLhEdLRhrsG1xaQC/cBDI/kOfqEK5gVj07cWTclIXi6uGvmcP76OJj1l2Vn/vCTzd4wdWPnGfK
axyBWCgguVMiJmMNBgu3jwcwV4JYXBTxFL3lUJVpIcIGg7gJzLsETgUKDmvxN5xwARoQSIOCf7LU
ccc7hyYjkgGNirpltkZGh9kEd355KOrciOeg3bvnJNfQHWUNz0xczDXQGlRhkulwy3kh5Z1PV4fa
ntXynDnxrzUehIZYvKFs27ERTPLYumWFTjIk6qtIuOZ+Db6P30nE9wnKq9LEcf5SeOiti8zkLBef
XBh++Gb6/oSJrJ4l3Xf6EuSi/7qM4bW5al0lBACWcg2B29DgAvI5r3OVMG+90OJLCrEQnIgQa6ev
O+8/2aA404oO53UpW+GLQHF5PJgOJIBP7dVaGa3/216gHsS2H7AWCvoCNcEHKDXP1cNEKsfLNhfU
VmI+kAkNoDvkI9iwkRYqWfoYRKeer+Yqc+CEVlUoI648cNVGnScsFL2f4XLnIefRe+dJDz7ofgu/
MnOOXS66sq0q8qiRyvhKL02dtZWPDbX919xGHjpQG5cbwhU2Pu99u7ag9GQfuK/QMRfrrf3ldoLQ
exLPD+oQx4Ozppm1JxGIp1upIZKYFQyXZQKE4OIMoSGbRkoqW2tanzPgN6PWyv4F26GDU0+l/cW+
K5pua9LI6sA/Rnrk5Az7cN9VhbGlMAyqfnm2triCIDYarYNFH2bq4CzBKvAKapJT5BDKd1IvKSCB
FdORYULP9bY9lmG4h4o70PbSGAHEzWct3sridM6OEK2ynHyi8Mj8MsdpZte983A3Lo5uO2J6eQkv
0ppfJUslsaURiSDi2xm39u7fD2PrEv6NUikDi75NXVHkhMzETOB+F1xji29hWfkFloXHQhOQGAeU
5th2YfPBNQMG9GzSpwcvXQ7gAE+0S/n91b9qv3RfpIdAGsIp33/JchbfyFsu5hAOTcWwCk3D/rT6
TpDFt58InW2oNCb0WAGKBXjVPIatWhyBseXA3uNpVUV19k7zF0jQbg/14giLFdtvMLyU518jjxNF
gukzjotGfFwYhcnpLB3Og+kvBUvSH0qfATL9UmRj6/c4bsaupO2ZVEpQZNtofnsJiQVBWD82ZxvU
QJ0d1dXznaSv0PlKhLL5kShCl8DZR+z7MmDH8aNdvF2mchn2zyFc+jp/36YsYF6INPo5hk03sIir
GL0ZwaJHs5Y9WusoGwqQ8yrVuIlgNuZ7Bs/VsdbIFBPubVTuSKw8GZIawUS5A2Nlw+Pi/IPcFU36
FcTNeKvPTR2qmuIcexaMvEFxRhSo/dyGNWEHkgTh8fC2Ny5QSsSTmklPmJrToAirzMAuzZ6OTcl/
DDc9aky2dPbSqXcwxoosEdVW8qEXhLzvyzvcBRj+xaRv+VP3BGOcXEV/F/e0emQtIifaH/BarPc0
FDzdR6/P1+FG85nvOQiC/ha4e5z/Vg7D9wCgom7htVBT4iGesUG8kEzf56BfCE71QN3iHSpAYenW
LNpw67cGoGRgzS+AqU58Y+VXPoSBhjodnZuoqemUw4HCW7n2NU74ZlQHc6OK0LsD/ddkg5+o7Z37
aZvEhwSpKs5hk+StjUCNz0hrCafHf71g6V3Wb2Fv1aHYVTrSfBNZl+aaeJqes7I+aLwkJwk8k/5/
aE7iktfmdkIzuc7mBbMRAujokdtqccp39bajm0OxP/pRY6A9SOMFlS9c60w/cixG2EdS4gUH+VP6
Zx+0vcYQW6iyp29TJyjSWMg1Sx0/UwP+LfJgMC7nYmswgR3vNBAs9CsssnasEnmdA/lp0XRO8Wl1
Ds1nxWHVYcqc1FTyCYtwvcSAojRcXP+CWQzyvzQNWv7aksEX2zLtVARvQT8vr0wJSbFRfQ1O0WNr
cKq1QMJqrQxU8tC0VewidosXO/rgICgfdkxbcew7vboRMRwSCU93QVk74mHdC2xDcrCLBDuuhz8U
w17e1AcePcACxXnHwZJogQYKNQ+bPEWoPHj0M9xJM97Cgx8SprGr2A3DsMLacHS3U6Zau4IFDJMg
B1o7LvtJPzuZADf86JoMyzczTG7b698RP2FvT0ubhr1FVilqWT/orB4tswCX4SOaockJS6FV7//3
GAqFymy/0r3CEdb1g50bC2JojRthR6bvdyyGV7QXzAGHINj0EZZxItixPicGMzI1EKIkmDZQh23k
Lyq8UIbJiPKtXJEQ8uk4tV69UExSSinwZ1uuFLJfSGiCanzWCw6dVuxuqwp0/07UBTLKtJF2H99a
mrG1nVdI5avjbM4wnk/oxTiQ/vEruHp4KLDF1KWImZ+Mw+VuvqFdVOTxdAxI1hSb5prGUPWGh85X
XFNY2ztyQNFntX5dXv9fA5E5812GFKWn73b08pid2bfgc/Np4iXPFjJWBNGE8q/lZ0mATrSSefGo
ywiw5tUrOxuUQmD4HqzeQJ7xKY62Ivrymg9GmqMAf/ltlepgyD8iJzDTCf/VymGAxiwcEBHXvbdb
+wdJjRCvM76XzV24oXvb2Uzg6Myeg9UvdjYz0FZNlnkV+NlOytqAUm5tRzDH9J77cL8Avk08rMUy
qb7ycgQDpWreW3TX/SYlR9ZrlqnCBmQ7j3THU2AThpq5yHxrSCuIiBPDdWK54Ux0REiwmix1U/zx
ccQkLUP5GtFCdyZyaZKmlv5QP2dLKM1EkzP1X9eA4mh5xNUCc+PD0xrlnyXlH+uPWjzfHeYzlPS2
SisxFyYJcHrMYBa8qp1VRL9IniCMUvYq1tNFGmOriBVQJtNlHXFB1idTjR0d6w9OWJ4IvUBKO0Bx
d7xIudfZoyKlUSDKX9hF3WMm3KoPK3zWkexZ87e1y26cKK8Dp2gAym2LaEoHQf+JqLWPzkz9ebp/
8gWYy9ArbHiRLDb26xcBxOPdmP8MKBvUBCfAJ/d63Y2vYVNZByMe2FcnUDnRXIgjyKROberXo7nS
ItwNWMYY5VucnXJc+Mlsunu6tl7O8fK233ShHUlSQLTqmKtC7EZHz++5dAZ0qVoHh9BJAmpdMPhH
eGaw8pxJ6G7v8Yg8syPYmQbirMJvhnu/KE4ljXkGsJZfMwqYo6NJ1AXiRUc/awwUqVaLh2WTlE20
WjGg2HRpqWkGjfyeOyeLaXy655oxq6OIxRqy0G0F/HSOB04AlgKWCYd2ouSdzdjydAMULlUxmV8I
ooM3nzJyarW/Wz255BSvB6NiMZshGwJ8Nr6e2602kvtT06bZJ55Jmqx+/nsplb78lrpf/DOw1Kxo
7pwSjPQp67QxX6mW7mJL3nSeOkQ9XFcAwezQjuo78c63jSZEwPZxUYLrY1P/Rc0yYHTTE1Pkemlj
9dgQI+5iRskV+uNhWpLhCLcB4TbPjQ0zapEX+Tt1XQJ9h9VWcZeDSsuzDB+7qfAtuduDPw5wcx1O
eVRolS3N+A9Y3OM7yRw7OiqEdTCrNm1lsmqrrut+vpug0JEMueX/fBPvjSK2n/iL1KcWgzaxIXJ+
Jklr/hM1Ok+OhufERCC4ozSFb+TMv9QQhiEpQdvMMbUq4kgp7RfwSAnrymYXzHujnmQpjlZt/uwl
wqrNSKHbvLeSWgDWUnzgvy58g1XUPRC18v73xBb5TtcgbuNndc8k48QKdVS8rV0w/hNcjKJqF2sn
mBFA7XQnjUqxFsQD75f+pX/dnN7J1GM987Yb0fKLjR8MrzaoAeD2VH3x2pDTO0CuzZiuuaX2QMgM
Osh1yZQsxZ7GmIttQuEIPhlRTKMc0duwafk4QKM4kyRsFtGOly7RCc8Fll3IXhN5an1G6l3b8nS/
JeuKHA7+tHTA6TuNhcpFhi32p+ROXtM8RnUYE6akRwkC6bb31WKuk47FHutyoE9HAMUgwxcNPiHk
Pk4xbepGL9dRrffmhgB323KE3KTnIjQp28UzbAK2dIVJU/bzjxeI7xpF56PCZf8ysKYOzC/rNyjn
KWkZeVurDiMSkNE/5epXy8byvV4XSgW0IK+LnOhVWxc/pvc8N4sRClNzPbgQesq//Txp9ttZ26Ge
8jD/A3+p0wm4gx2GpLTz0Wng8Ad9LAvCtooqV4jo7uPoQPXKRgikbb74E6KH/ljXDnTZSh+PyD8Y
q8gFIZD00rglPhKkmzpOpkupUaxbl8Y/spjaKoFZR+TKgcXbTtwtxgZeGysqAzRckVnVtCzA5db3
UP0cWrq54GvY9Yp3NBA1dH4WKOx49I5Tml7fHXV1XQDXxiNTFyHQfz7VKneH6RwZ0+nKoW8+EUdf
5ZxZ1SzJRFxd3kxCOzOkyAs9K+T3pxpwS81NO0/3QMkoG8HuhoGPBZkpbnNnPond98Hk/x09Hjy5
7zSGYSKXUU0af2u358L9avHQdMjZvfx/5i1MiW38kR4ZZt6kLszFIlhXnOZ8QO1/xE9rYqmsPHNi
GZmW2Ftmxe4zU2gkWm6cmJTLkgALm7BdBVBGcd2jyVsEWhhWJIvkQMU8M0Iag1G6vVrmvxuvM38q
pyIRA7QaWwubAeaZdAwGLBzdQat+nomw2KL0uUmgObuaRqTuhnAKpBmefNZJJAvjFZd6q/6gQTeO
acEkjlAB37Y0Pz6ccLrMSbF2vBPiijdz9lYfQ6qRBhRIM67HF954zJWMz3GNQBpsDB+lBhAsPYSG
aRnup/42bGYz6ZArdJYk3zfHyxWfdgsDZByJnhpwPZzH162Gi+dFh2JkA9I58JKTps+4wq4BK5IG
I3Vt04BR4+vQosyTvTV0Vj5CvRVuGXu/v8tbir8z+zzt8GiEafE9yzTU3HqpvrQAAEM3pBZeOpYq
r6U+v5mKLDopdn9MnUYvUNeNmaiEUHezmvmUOVv81952W4w6bRtnJpwUXgh3w0NB2CMv3vgOL97I
OG6JzBa9xlB5gRwKkmSV5sTzRbpeT2F+Lvq1slmeEyDbjBrVpRtiMGeV6EbQLN6iIWpaiZg7ZmOb
axSSKAdfWIvsVlQgeG5PevSwJSWthGd/a3To2edFwhZMeIebXn+9KvUpBEJmViQ/q/mZAX02D0KJ
8PuUtUhawjGJ5mGTRt7eyNsPcy51c7BBFeQmpU2QmClMvzCO5cvwmOHgYxe5LRiEqqFPY1x/GWH9
igHukx7CK3kv4Dnm50ZYM7DCgb1vOB6TG6Ey+B6GBuUcwHrxxwq0Q7JATs1T9XYbW2PWrxKr223r
o39LicKevGNwJSAoURtt6daE6YbVOMnXEa1aRhpB4R5+ixg5ewb8KnPoIaS9Oe4Mxuu/0ngh/7UU
VhhT5xNNLBn0xofJzXfs8kLjGwkNJ83yenYtGC0ZeDASlHNzZlgrYOk2M+o6gYKWxyvUpsiEY75T
zdGcxJPFBbNHedElCq8t34PfOCWeZODt8h3zyy0o/7Wl22V3AOxdqcbjAHQbMGxe2+0PQekJcj7v
Fk7LgtH3jCaIKYQRdmT6ArkkYJLNFTkK8tiZs7OvZUQQXA57pDdALjQk2/fQl2BqRr8EFsD8p3kv
eTKoRsYjwB11A2LNIy/yCOdiNg3l6j2b44xADP85TMbVOJ+GVzyJ6nEGkBivovCf85Df5/6yv4gx
0FVZSnNbrvqjpQplHDGEsbLPLhzBhoS6nh6qT56XfVzJQAYW8wEIQW5XNXdXTloDshcSbgxdSi+W
Oejg1cJlMY7RyQK3Kw3nFK1aMhsp9Cs0TStIElTbTe5TZnzUQyRTBcguDk2zV0DpBTQxy4B5AiYB
eIjKFjT1/ZXv9Ni4F6UE7M/8c4bvofo2dApXD4v+mRsqCe4TDp90zo4hnqP9SdGtFhOs6h+HuVY8
+9Vf1DxjOqeKFUyrAHHLgwSGd4tAYMkKgiqhnM6qZrqvltVu8pjGGM6sQHVGo7KahGSP4ZCn8665
O6uoWDnTBX5yKLmFAmWziHNxA+HJx1nAHI2PmfBVY1dyEQ4V0UH+znXHvin86ZdUQslbn5uydxOI
x37HE4wzTUz30rk0a/U26MNYmqoHiewrTJx6rY8wI+KBoDUM6kjiMTc4d5r2bcHvw2J2FkCh6a4O
2nSKX+6qh/9+m1OSDUOMi1mc7DvAjJoHyZXAdt8ioCbLSLD3CMlPqVTnCcQ/S2eSLeVC1TiSIGcM
+/1+XH9qBp2O/1RTeApN77AVp+a39UHsKp1itjQakQsYXte8FT2He5k3wtV+0ZcHY0zvVL4BCRzE
MlN41mVa7q26WAO8YhzoGosBDLK77ZOEAXIqmf/+zniRxD46PQNKjLGb8N5h76aWcRh74Du2QIog
qzFFCLXCVytRzTZnzt1TaTx2cRG9VrUO1dIs48y7bUGxU/m5DTShL5XL69RFT4R/ozIr1W88lcfc
/hqqRDMW9CzPGwLzobo81XLvGxrxSjpnnRPVtMI/tjzekyLwFCiIjMmg5IwrystfXCzkDhxejVyx
2H093ltJLuWnt22reX0HRHh9Rk1gGiwws9L7EwdRJ5QMO2JxAafb5Wi9FrOhhpcIwXqL7NYLiqnW
sT+at5XsAxEI42GEvtATjuXZA57fi8OIRUc8S4RR7ffjCM5v31bHRn6MbdAOq4mGcxvVyK589uZg
+csrRSTNystnfVJ+IkSGQX+Wh0m2HZrqFNptl4Xvu0M248cHG9OKQsjayBRPtkymCd1zOTHSf2BG
PODGex4hj5NWKIjti3bu6fxk98DbyMU1mp7PYmIVY3NV+co8wcFXUnp43xKK2UPuBSOKMYqTZWnU
NLe8b5uOuJAWeYCff8hIg7NZvjY5zZZEAK1VFrM3bFdupm2P3Qqm0kOZwfCiYiPAqCDbEFPcJB2z
fPrSZQPFv4Z7OBhWa/S0Z7vhp5Auv6iDgGASwV0nlZjuMHygQNeACjDG7Xn021TMnUn+j/qh/v6t
PwFJA5ChmQo9z8atslf8WDNSJRMuk8LPkFQ6ViJsO0OHFBLv2rvbKqDlRim3avhHrs70QwaEZoBd
TyUYM1+xnnNgDoemnMUmzlz/pHdJSot53YWHh76+u06fyot/UQtVIOQECmne2bRvNu222wgVGyvO
iE8XDM5rthNJGVLrOAUk4ksu+RfAYBZJH0Ky6JEa79mtA04R/Z3nq0SjN12dHwbULuPvCUQwR/QM
AiN+fJ8uhgRdukQ+fEhZ8Sv7LWkEbOBDbeAd3NQQzNc+I4K/0B0jptI2ywDOXt5E79S2BlZ4ovhg
4kPoz4ul9QoDrvsDcrlf59VnnDYLT7hVgNgERydiFImt4vy6kPP4ipYcbGpvpRuv42h7M4iV9Mcj
ENqELQmzmzHolWXuPNohvKU7d5YGiXaTfoQRcGgCTvaTBZHxwb7c3/LqJck8SI4qdM8rYL+KmcPo
Kxoo2m8IB3uaIya0DSSuvJOb9NM4kWZmWKIV/yxaIM1sgxx5TYYfu3HgdMa552iuXdO9PXPDN4Tn
4rZfkPIYUZy1PsxFX7lyYMx2wukydrMOA4MS4BG+OuRkelLyhhtaRWTID2uLjmcT68v+2WKx61U5
b7rEv+jyh7TZVqws13cK+n/jgdeaHwMHjEd+C7mxpbknOxqJBTpkO4Okyx+adevpe2qKmTLuOSlV
spTO8Mlr7HsLz5T6JsNJk3pdgCjepoK3elJkPr6im1zErDexcPnmbwJdLaO9NcWSONjQxG1blxRK
/uwdvIZIJoLLDutoM/Nc4L3uL+TeKego3rYU4Vs0LZGzVScAYJJUepVUlxhZEtg2T1XNvE1bNFDn
ZT2XFeXVdaU6vXjITAkX7fn9HHAc5WEg/WMKmPFWEB+a2iRnna0SUXKCsgcPkRdmScahlvk3q3Nb
NAz0wFMHsPJJScC1BoAF8GXJJTRewDao68nrppcXmfh+zc0LhZqQ5aCijeQjN3UFOJHkjT0Dlk0/
RjeXrMKAezlrUpNli8bDVGKtJp8ectEVl2lgRixiPQb+Nif0Pi+wtetTDZbfQT3wA6BzZL/Wc9W9
pXBGQ+AVconOUMRQ4OM5r0DGsw7hRba0sO+oyZ1UgDBY7pUaYuJy5VLP1YaP7ouBUlhSMgLpXzSA
mfogrWFfjWl48LprvjQQ3XnUrrJCsuqOqehWiJ0O59dWp4B7MsoercgltWND0GanjJTCfVPwd+nj
j7k3IJtm1NIsh6uGTJNSro4bdKFBL7yroEtSb1d6HWjnpJ4IUgka4VkO6VLJ9FolwM05IssmXkm3
vr2PhPHtLEGI6abB4urPEgpQcVM/v6aHe/H5m6VwNXPVEQ0fDZJZjVmPU3/8y8QRvFn1vcFXK5EE
KUrfBMBs7wsMub1hxTFgzJbc00e1I6usYHB901Q7nZiNLVDrqglpBLzgp5pTieNoG7m2ZhFs/XA/
KJz2YRNRsAnbo3Q5zOkSiXAyVRXSlvDfy5noziIWcLklDdp/7BXZnHhFcoL9DBFr7UTD3smGSCrg
toFaVe6EOEl0SO+dFDmRmK3I8BIAW9/HInEzEgmM/HF1xRVzIeJd/oikXgmV7eB/O8Eb2G4/HxDK
scxLO1fNLsf8tQ6T1xOjOcXx86eoQt2EcBMEgL2uvajFKOXfM8XhHWNYtRuMZ3IfuxV3y+rAB71H
jBVwwlSnnbkoQH1Od+moPedBXT4AXOFYMLl2BL8MGlli3PfmRCagFEX+X4ATiAStvR3EMHeJWOPV
gP6aziR4zTMu/samZ7qTHNTqMUjia8XFO88gfjm0OI7ql6BNRUPV2kuBm71P6AKDlmacjAQn6aMZ
XgzIKsftJks7+qWooBIFMZLfVkH6uGFCdR9NS7slcSvt/lgPhWXBeUMULs++ZeqSHilRENMDJvsu
9kwnHMHU3GBEQ/4oww4CfZN2iKo9HtvHPjI3ncHTgEQ64Ae3e4Ju9vib9BhZfX66A0G8ja/P9BUw
qQn3aEI8nmfxh7Z0PaOUFUvua0Az1xgPtXfQJ5OCjSpUsEjiMgasw0OKBV98Ku6/GiynAfKzWde8
ceh0LUKc6LVe+4lhGq0/06bKZU6bSaI5F/CNxs1wNBh/pdexv/onrPwqubBV6wxi2hHSTB7VuPQ9
9Um39Z0EizYSOV+6+bkPghz5ZfbFI6c0ca4VTnNfdRujqgESfD5qXz//YbFtl2Pj+kYTVFQbikPx
+KWo+UNULQ1JE5dOwhSECrMk6BGy7ZxwPhZh7fBytkpqAzxs9za4F78ME5+C0Gz6+bua3NCTWAFy
XMrTJCIIAeTiyojcOJ/Ej1R7mTPSxU+7zYYVAF3lGZNSAtzfSiA/t3AAPkGUICe2r3vGp5tAuHoC
8ss1+V8ABUCrTs9OzLYQb+haH/kOJejIgDiGU14Bktkwr5bC8b4bdvNdRYuYupigzQ1qM5NivVjX
Ug/RpWhZ+iAhc2EaWP7OAHDufQAwTNxsL17Zvsy41c4Vw5eVqQprCsPoIW3s8pikO7De9C8SnDbo
sd7zEYdDJIZBGU8YaNKwfT2hGqJBoReX2QrUniRSfdBjCo/MQJcolLbRB9XrA0Z4ntCIOllPN9w+
IPU4JLHmaNHw++G+AaHZ5nNrVenJJMxniHbsS+nEr725bmBmU9tLVstx2UDhVKQSb/Lc6k/eP07q
HikPLDLFeQcuGfBkpSMQDA3R8wtMkMdxer0+TU9ZPYx/4bVvBnyw3GVZFTZvb1vwFxx3vdOyQDvw
ikBWKf/axknw7KNLUJkBYS8cjya4w7j/vz8l53g+xO5MXH+H1WPV9FtCKPfsREB2vU9cIQhWKeOP
AtU+OkgsNNaal9pAUPxmVFvtNR8crtJ+IZJOkBz1LXJGsy51z44uZ044/TQHjytpVVx96q13uLwU
jgRvsYjr0h468VoNqubI3FIoN078xSc6EelbUv1ss3pGH4upTd8k1lGylq2FXl5W5JM7clCiragv
9hAhomc9M/OWlZkrfItActEgGm/KvMKWzArse8ppmUxsCVJOYjYijG3ZcdeAl55nR5nL2J4W6x/H
VAo+YOtQsPcp60ABzxh/fsyr/gMOHIY3oIy+8fhLsj4zlUGXHGTWTjuCi3QcjAnQn5jZqsNE76dG
syDRGmZgMaHRhkfr6hAH08zfy+8O2k/kNAfJrqErZEd25UyL9WZ8ZuLvLrXTQhEFMT84x0QYFUYt
zbHqHroLjCLh3j1S3h+nHS45LhuyggyEjOuqDED+3t8jzc6x7JBDJaX5SWuMAMXi0ap1x9l9H4AG
Q+NTdWco0T7jcFHcOvrYwWplepXYEYBo2omPKOU7dUqaMKRyBY+O4l0k8SqJTEhdU9L6JRcJ2HFw
KKKhM06N6YVbqUdLSaDPIzxQvElyK4rkmvBhs0zToq0mpZiqDD0YO/EJf/+Q2o/NsAHiOOK29Ctv
wbTZfdhdE4y57S1B7SNsjQIqLtrIQd8kKJmg1blEJkVFjg8SSUQMHC4dBq8sBZ9TFgy1oiiJK/we
ExH97oNQYn89KgP+GFSxRsqZfke9DAtgRAViSqG5+Oqqt9GMaHRiQ9Lj+DymWsMxaPvIo4UsKGCr
3Fr3NHQjawe2LSb8dSNo4yMVofxYzkop/Z1fuNxxTwsdJVLN9NaQbAadNA0Xs9cAS8yXq/VD8aOO
1aqV20daAppuw98DoqwiQO9yw84Fe10LkC7+LchgnMSeiQME7M3m6ryLrRrHZlCCpjfAd3FQI0Ay
do2jeS3svF+f1aBR6n+yzwnRNV5ZJy4/4PoqNMAD4G628cJr8qpZAw6AeQFPV40JMPdDdMmXUcPh
9am4aoI13GfCJwOBTO454DXnX/MUTxtJYSghhPcLVD5TymvFB4vKreLiJGawd5VKsnDHXwi0egxg
OggoJ8z8flN8lJlDwberebZDsfxzUoqHZ1cjAKeKkIt1vcgewKtt4BWAeVW6U2H1F+7hs51NN2LN
b4yza8RiKeaYlsRjX6LkXwOZnO8LgLOI3ZHqKs+otdZ2uOXdoht9xC3roHb1Sz7qOPDH0GSjzptp
Agp1nEejupBaU/pdHrHPII6tosDkZohjcVsarnK1c046Po8ztrrP11hEf1k9XHMydk7fhcoxd8Z1
92CiGydvrFUyRmQlH9n/X5hPyHwlNuzVevJyefq92e2xpb/ogjZqR6z9j6kn6B5RYusGojn95q7i
jlXjwZwJhG86W5dXJz7EBDp1UQPH5YqxIOVaPyzrwrBbYNSTfUjEvG1ZEpyO8xjVKDM+FEDJY7O6
IW+yWmLfBjdsy1IXr6OItBckn4731YdwRhlvBQ92
`protect end_protected
