`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7472)
`protect data_block
OxGj7egbtg7zRd7++3Ec3JjYj0qSSQJGf4bw2YFL3zyoIPQvMLBUCf6vQv5JQdWflnrTxgg/6eWG
W8LbxRCL43cIf4uSrQmM1uVDRJiH5oZ57hnq+nPif2eXJGTjkfJz+E/qefwnGfTnRcRUIwRU87Sa
2+0N8ELQjZy1GPJP9h0UVF++sODdJTInfKkEhsqsC+vuT9B8MHQkLGBdCjJsr0k21j1fVFgiFGXx
JnIhpIjhWNLVodsnEAdW3y2A2u5pMLt5x/CnQaW1yCtBg9cXcIBUCIx4pSoiXqXuBtkV0403yNmO
MHzSFTDc0jXaH+SJ5ofgWJZyLuAf/CloQxFwJDG44udc4cfEhBTAfdcG37LeuNfAdbARGiZIT0Dn
O3yv8x5XjAjN5FWF2Tk+8jpQV6OuVynKRSn+JcV+dgWbKTsffaZTozVysf4mmZC5ugvxx8OAma1I
vLBndt9k3b+pCfMTQ+1rJpKEsEba+V+MoUsz0dpll6E3S1MPbEpMIlKFFXvHt/4rFvl1xC7HLxXs
rvzU7bBH7sH6dM3/YiGkmVPsttqMIGpf+Q8tIDWMM1FWN9MvFW8doBdFbB+G+X4o6loOtZjaheZp
B2PZ+4OPkKCu6DB+JQfkuy1ZTVyBPyzaKbG7WVJUzQVsfm4Ns5hw1Z9kJBai4dRKX3qtg9UVWnyD
UakUooG1L1i0lsCfIagkqq9XXeSufPRWjAlNSgmtCUlyc+/z2khbK1AOmC0x+EN73Uou/ZYYOfwT
P3eFGrKIJdi+G5a6ndZYrqSmDaE8uq4C0F8bnARQNTqyuI1GDRCe5IaZ3R0gQtHvYYTPkne0ndbm
wKXPABve5ZpWSaP2ipz2bQqMklmD+t5dqtyXadPIUJ6jo/ZlApGgZVIc7Tt4WGsv4B/gHG5A+DJZ
sD2ZYNSuVIWw+f6se4CR/DSpylNESGYWPWxJJQemDlgYLr+JzNI99H3AQJQeQR1FO8Oc7NE/9jGR
2lGFdHJB0CXamtbYilAWSzNe7sZ9eIVLeKXR68jRHJoZqCeyD9PWJd2HkwhOePt81GWohXi9YsWf
gVvLXaVh0V0mxnugnqMNdL9vieLRwESFv78uWKiESSvkNSL4P7GesQQR4tf9V4tlR2+IGv8Piqt7
SPhIAybMYA5K3NJpK5Kzjksxw8mVIX47hY5GKeI+f0ICZpIbtQEkHQm3zFZkJnU2FOsTU89s7CQ9
vQlGe6J+z7mmPYRXghnz32mQ4zr6rQld+xoDVVnyIFbPkbSkm3Bh+8tz3ik4dlOjWhyD40hMQH2o
p/AFnuxEPvFjMT2AouwFS4Fb88Nz/zzdzu2f3JRbH9hwmhff8pJCeVu4gtwYH9Oa8TIMDslY2now
oNlJHyvcdBWwq1RpriiAT4mOY/pVbt16od0GCVees/vhh32q1VJIDMZ80xztM6XdKocfTbHiro3o
EAsA3jNNhFxm4ghUJuq7f3nzR0W4Coi1GXOxDICzz4INCu+ZtcZreeunVf1Ec6IEjuK/q1qpSaL3
x5vz/z2JXo0hU+0cGA8dvVpsfWHvQYAzFd0gqpdc6qeZ25gwf4i44oY3IrWoQTFLtfkJXxx5iJfp
KwurqnqgMzxDbg+Y0Cd8FqZJy4NJO/gG/P67mm+N0Q0nI9LlEyQRDM3BhZPzxB3KO3LZgyhzw+RD
7xS/TyaVpyeMtAaM3IzpPcYKgV3KYI9ZO0d6n6Pr+DCaq8wPVotepug4YsrdhccDAp9KrX8YmAFr
cZGPH3wm/XbUeAC4/OZJ1BEeS4GYkXVXj1eSvcpFqDeNJeDn7HaCVZboY3s2t22wmlPzXnJFxOA0
60q6RRXBW1cEt4gpc5Rq15o0EmBSmrZCHSSgaoG5R1qFwoM0xPheIvlthKdZcb8RRS9HMlSfEik2
qZr5TKy45wewy7tdAwllrs9dkBj+W9Ve8JJR3qqXi3U8r5NHXsmm3WgqcjHcTGfgnkA/H+zbDiLi
rAUI41a3ZAT4B0lX9cZeDyggoMj8YtZwK0toZ3/zwxiow5Z+28zLnogmcwwapkdotk8xz/zpTIzO
wED7pZGKhsET0g1ru+vVDcwuTPSiTXL6HrXm3IC0DMZLqKZ4GDigEvY2bRSiJYEYTis0KcCGtJOK
Xv0TUuQHTbBET4+ds3ZhNe7ukcuU8zXhyG7TGxWE7hAkLWEZcW3NtvEnikwcpUu94E0oc0AQkZRf
3FTfZS/1obmPkl3/q0T/6Z//RxfttlXs7ViRhipJSmhSC8nIHBfV7xJXetckje/j5nQvPfvvIhvU
UgJ4GAZ37CHZOyZDlZZoXzD4eWciN2uE4HckvrDxKuqmTTai53TASdvzt3+h59mpCo2vW8i4ghTI
KssDOqSweMadOuR1uAd4djCgyeZqQofBDtG8aH7Mw7ZYyASoeiwozaI8YpiPLy5RCjLmq0wdhIe4
kjDkdaDhJhA/ZFC/TIKYJsYaovEm57nmKxA+uGoukRhcivcNAd9Rq11xqmIX9WqaiTjLA7O2x/jj
gzEwzu4LU3SUpEsWMneYkRxQ35Ly2kEAmZ/K+hXnr8kecxcLsr/K/kNSGWq49z35YpWQVARk6OwD
bo/g74FQJHTGyNOh6xWm6JS6c568lb0agkZrHo4WWrNoJKk7S6fqBKw8P2+RsTpjPg7cuXCWaD37
rGQv9pw6TdFSU0sHbgdPmXBajbOLBARgzHVU+3QpNZ0tLvgjh8KnehlWPA6uILmtyGogQBM1mzmC
UTm0IAsGKjT21nqFpB9JtNqlHTiNG834GgxiMGCZdTEb+Qfz6ZhH3TU9TA0EqJATsPFxCKTzd6bA
r7/cfyg63X9uBREs2tkMH0mpVSDfeaNH084aJUK/tQaRSMkcAkYwraz0JyEhlbMLr8bSundFxYc2
B+YlOhA2QMFyjfXJMdqd8Y5d3eLxr64YYNkcdO0SqCxwmUFsrXptBptPawA8bWyjptcSPqJ/dfS5
dxaFStV54c7fHgWM01peGwhsehdQpZgI7sJO477OW1z/FQSzb0WH710CY9sqnp+5tTnXnSA8CWkl
TdV/hjZcY8tDIm+TFaXQ+/tWgOupP+csHcTLldgYdsGNmRkCmynVCSnQo97sYrvR7MfIPA2nDun3
gxBh9Yri5+HO2h6ATQ8whHvZW2d8jE2IEGxfENK3GjJxu8hRjfPkp2WxAIAZmyOiZ9UbVH2KYOvW
7tOHOjTDUpmW+tHGoT/OP1AQVNNbXVUvNnBuwGusHrBMBMQggkw62eoqYPVPjCmJlqwM9NaBwMA9
y2I8lK5vJ0X+ldrEull8FyuBKv2zCLpy2x/0U7aBP5m6rQQt6X22lzj2Cl5m4s1t1zaK2G1XXHdW
EN6A3OpOGaesA3zRJ9VkuEu+gqrvL2SXWFzA5tgHzJd50zFZvS5wUpB9WCX6joGdOg0GZVX4n4jV
rRv9IKk8JPYqrb/CvSUrHhvY40OOjEfsrvW0Qli6Ds+k84/17cXnDGPEZhg1Jdm7nljcWCsx2E6E
N88KNX7L9j84AFLdNnUKJVmltuWucCue/2E4EPzWpbNWfTTDrdk5YyTNeISfJmHp6Q9irnYBtQPX
pBXPJDoT5peK0QPGSWhUijqgmkOrCqenKFtrpeiPZdkv1+obRAZwCfxsit309GjinKUo0nBJjDRf
7808hiNXirX30PQ2xStiejc3kBvBP1MdNRVvu+Le0GXEjNVGAXvnlh9za9cZiY9frhdtG1xnaJ5O
9tupxNMj2V/kkt19PEI3Ch2GXb2ACFos/lwe5fHqtnfmAQOAMMWId0lbTRd3KtwWYnC9d0O6RisR
pX5XyTZ5f6qWu2VMOFgCKcx0uzkY5iFxxFOK93KNoPJVpbfkj4bKPaCxeCLZSOfGUw9tSP2sO0N3
EWGvxM9ejlmU28Jd5QJ9mL2apK4w6N1cUjJICoJHD2y7UF6H9whDSh3GZA/Ohdr4varnZG5kMJjZ
FFLZnP9NE7ADqSxDplUuBTQCvfg7FStpfMOzCNwSncLC9bTfhDHhj5F4JY8WVS/7c2pak4GWpQEe
eT8nGJiGfpVrV9ZFX+R+TH1w9lmGnLA3ow5eNtHyHysmkZtgHIFSo/fUKt1a1CO04nVDnqU76tDp
2zb2cFzBOvevpCy42Mtlva1JUCsk7WgKGNua3I+u6S5KUa9aYeVPSN+YRu4aiOENDLNe0uM8kIop
e0HW/hwEzB8S/HykZskV9uaeg+pp11itkQOhBlVBIGIKUcj57Bi6Aq2TJzZS6k+wpLO/wu4obGBJ
9gcGA1gEKr6DCZGFat9xafFIpwL2/XqS+UmJt8DBciZUJUuxLztgcRjXolTtmoQO0Zk9www6Artr
K2BC1YJvubd9uVnBJnYjgcdEZvXOn+t/ziflTnz4cFHyEvzoL7csyrqH39WtOlL3E9JOZp40pucL
tACItkAPzzyh5qWoIb/nAmR+udlBSoxydY81+BHReybkIcvd7r+asdpqsfG8d+CyLWiWrxsk197o
znQ7Z4x9kqGwaRLcX4jDgMyLwAihpiM22ECfEMj6xNG7A9X5NQaCSsu0laidkNw3kMdPdkuJvIMH
i4FTXhAT7WBzobMqc8SCZHRhb7dzeZsCGnLQq6POEHPClKb90RvKGlMWcljO8gT2NwLu2pPEW7sn
p90gCTz3PSc3hTdnzz6g6IgGq2Hs9iGg/U9H7JKfVwAKsV/GMzR9HwDHynFx4vxQZJlUqejmjPuc
SpH9CJcXc/htJlA+0XtmI8haSCkdfEjIPlTP4kZDwlzoiX0wlSqU/oovaOYggkE7qxui/mPib0W3
Pv9wG04sX9RCDuSKv7oZpzSveKvwxCgkZsHZ3aSWTAs0mknt8J7VJMiDbONkQ2P13h22uRTz1mKD
xka9CnS4c7KhYsDnK4xPZLcauS9+fZnSWGJjZk6tQeVKb41MV/cR/8Flf7R1RywSyy/fnCzsW00e
qMUqvPygd5JXdQjWWLTwJmnwh3zym2cnqFARCGq9ZE2yz5VTXeptf9RRx8z5XjZ16AWyypF2wdC7
a2TD7hZSIX5Ylo8jTLedAVRxDHCy9PwCIBYwLTHcIlQHiUR1tN5ZC7C/yn8/D0kSyVHQKu/y1jzT
6HMqIAZdlVptauM1ryAVgfJUvIG2U39Ixx63tBoFU1+QAPIoxsXclsONHcsuuuR1G7Lw7y6s7C2d
EUAjxaJa87E3AaNw1nkGgl23xiRv5JwESj/oLu+x1HDkzsh0IqKPCuxPyYhgDWnHD8hl6volZW8W
4oTdPyP8XagegZRQSwBBWNEDX0B3t1FqglUZaNO5VZhjVZenCsVpv//8jw6f0dy2fe5iaIypGBKH
RC+sZt2otsMy4aOrLdXrZFBXro5glpTsxmT2wVKvURBLvAFvreCfrdRlBUvYK6KuGZvck02Hibmo
L2qHqbPXvlQRfeIJpyHKL2MFYIT5bQD9Xb7wmbtwQrWX2L1BhY3ZDcMrmbUj3h3OYz/pBekqO9Lf
a0M1KeGF/lK+EW1pVRArpIuyNQMbfqFPcI0aESb1yA5ZyGjp5+Sx8L4TnFyiUU8+UXEQSQ+/zaaL
DFX3V+cHN7dXqOjho4DshT6LWnI5Je4yEIqYEbEtmyo9RkHWvlOusWSiEvE96vytXUUI2QmWqppv
0BxBxLk39PHO91DMVXxU5EV4hkYVYSeA4w53LoKSRQgtxZlZ+K+ZIanB+m0OotqMstrp5rNN2Wdj
PNTasFTmXeE3v1In+0w9XeTAR94dUjHgtFWSKJ1ELimEWhjUzEDDgdUur6xWG3PvHCBd05RS75dW
Ckuu3+OUkaRqzoutAWd5j6JwS+baMrvYcf04sF2T0iNXW2T+4A2dcTTYkrzKXmX9Nry/Yu1iW/8y
xhiIC5GyzCICpv+l/Hlgw8ZoMGIsV/8zlRxI+wYIRrU8sRvmCff2/XDFPqdCc4lVZhSioubTjhQg
Tlx5el3LZYyhdQek53tZ2PGrXIRtS1tsttq+Sm4grrPFofrU1e2ymz1zm/GEegsFTtskOqmQXi1V
A6tCW2UFOOVsUUs9xPdz20MLMvqwDSL4pwZlTHrhSqYq3Z6nZZFRc+ufoE2O9OV4uYRS6iuIMysN
C4x71RlHpY1FJA3XTOrduijuQ1uWYCHO/R5BA6fC/OgyMzl/P5Y7rvhSoeJ+hQDdO+hXiGE2DrIN
hBg834tWM5RWdoy4e8RrfGgWRtfcZ1cVfj3kwirzwYWUoGMXpj+FfDXbD/dO2nttZoIExMMCaseQ
CzkUkRHIvQo8QehKgsVYM+noVzNzh2q9e+htqKwgl+B3f/B3qfTWiEsCKq3u7KWo0izECn2kuTt7
x42rFW5gUpS3hvewksU6+Whj/fSPrZE7h1v9nQ2ak1e24u4cPjaQOGJ5ygGfjtxXqif3RLG7BRvc
RysqsEpLmM9N9x9mSNR15LB+EBzT84jsI2BZmQFjUBfXao36YbdTKLrFMWsSdGtst8+johNGe/c1
DPzHnitIiD9eNMR3Kzs0wix1aMHOAuZtY4gMbU8/LqvQJYaDyr+/JOng+QpVT0zPQswvYu5tZh0N
mcD9i5EDBGV0NPDMhWwPke+JAPYbb7/iv8iWTrBUF12hTQqMQ54AlQpiXeYxZ3jrwM4uV3C6TCXA
whGG+jnL9Wo74rsgZxMW6hfv+yg7uwVf6XpX4NCSVqEcS5eweLmBpxgz3uDtLBTr3LmT6GgvyQxs
3UY8rfqZrD8wPlD4HOiM9jYBQJL+mdr9250NE/pkA53cP6VUgd++x7Iw6MGpngd9ZXHx1s/kcE8L
k2IsJHmNAmagDnBANYnUGryTTFS1EjOD4biT6TF5gmGFJdNbHUnmNZWe3sI7wsmlgFhCsKSFpbEl
gblhbMr3EON0PPl8UMnRP649+0LZKv5WJzwWYCOQVXm4bBvzObgF0GSjH8gqd1zAq0Zq7Mf2wZmr
Nnvf4zNGqT1L3fbQ6HnPGmHH2c89VJ/DVmcyqNVpW7zXxg3yecDSnr47Gv/WmKncjaA7S2qa0sth
rQ/Y77MW5rWmt7heT7pM6AcCzYan3xBeZtYxcsHYrLKYdf9+WydV0mPKBbXL49ra57guvNjgQmE+
NXHQYDlGPinyjO0QL2ijbrgc6Odf3s93ejUAuEIKkphdC+tOjtPo/8pBCyKk+MPpXs+KrfjeUtPB
2obI7XKG49IgNocgGpUtrroUKWj64AtYqMfdeMp0EuJYYOaVgA8rnsjWAiu9hZslsjD8mFztk7Qb
DJblZHXSSYmQxGJ/2/SvHEgQzWxqL6YXfy9eyk9KAbgvBncjuRNv2W/BmWk9CSloNcprkrXghtjq
AYNSNWTGfVI1qmor5swlVP8HNxMPFxCWv8Wi1xd4vqSfLWuPS5qPq2iH6tzqV5TNKAhhPmoFuzgs
KgWsPGco/Bp20ySrN8A495YNNDwuNWgb/MA8Inrd+lluhvB3InTGCodSxQYY4JCYIPKtDsp6oUG+
AMT54HHcg4IjQztG1kC5l1RrJVuK5nSwS4FAlK6JGkspRV5Ynvwa+ZrPP8c9rX335YWVy2sbxy+U
Bb+9cflODEMWDsBrZ5xQZnP3NTj965YspCWein7PVhFgsRpapVpoJL5xJk6G+QJ2iVmRZTIPddrY
W3lwJaGOTf06PL8mWQi2h8+9peouhHJ02imbg0Bi4ncFeohi1Zu7szCZLQVFV2tY4M/Ue6/OwcaR
ndVz3ttNhArPizwLA49sO9b/7app4f0eZ0IujKWYvBjuyayzrIKIuBBH6NKkKi/h9G3/TcehVswG
98pwJU1s8cwsyFsPBWnO5UPs3y2kmiTXRLvpfYXQW71W+ctHNRr1/OtEsAwZBsL+4yT8XSqVbw0o
DXPycpI6WgQVC8/K+z77CDr4U3Np4iSgvBqvVuSIbutAClqlzjiFZ9evE7cTsM4AzkQ4/Mu25uAV
MbcOMC+xudMB5A/FilcSm7PS3ppNVTio4vJ7ik4GTDHG23PUfaFy5Ghz3suH84uOwhhhW4p8hinm
g5NI2N6dafJ8HFCjHAbxOJCXHuMTMOyoMfVmcmVe3Ave3zbugeIhEVp10gxsaZ/50/CNAUrbOXNn
wrSxjKgiZlLUuHUNnqsF8IyGdKN6rds5+W6ACLcthOoqaDEfsKZqi06K2FZ36N9djInyDp58Rtm4
puXgaBhVMt0JAn3JEg/cp8T54w6ijbfnn4nnWZ4eMS8pLx7EUOmvYQCtU/bbnVaC175De4l55Geu
M4P6/PnLl2+mmQFa1CztrpPksGgFVnmvkrf4hwPnrK9naNUpfu/O7C62ddBBClPGa3J1g+H+UkzW
gvWQyQ1J7P6kadJepXvEaDmXrgzZsp1LNcQDwB6rSIeMNdWt9v61T1LPXHMHTB2t0UNEx/689rej
GcI6c6HNb/fA4L57RezKhlOIZ9K3Q8lgfPIbalK1K+YL22Fq4OVEJN6cS/z1Kz2wkTlidWQM97Cg
ee/ifR5Lde4Yy6RsQjnVYmW/m8v+5MDKWNqrxveAcNRb/3Wb/gFgffGAAyFlJ43SGBQF6XNPk9Z6
17zVEDeNHor6mfl9VzzxEWqHgiqafFb9YEdA8SnEomJRzX0REy3uzS21oxXsWom5xK341QPACH6v
yTO+RvDM7/Hup8qfIqr7YlWrMnYTUIqc3Mq9/owT3muEqfRjm5+RRGU/VVuWT0yrfjMFGmN53n1+
y66Fv8AKbBymIP4TCA7CHYHaAz97lK/ft/B6ZDckvSs8EydEthUlJf0rPXLqZkTh3XgreVSVqxca
xcpcvwOdFe3UXgl4iYZy7rKGbtRj+g8JLKhdxNb2cM/0xzpEOCsAfptkgRligE+mhxt4MtjendZp
AP4TFGqECyJKCP8qLRn0/ComUHtXQsWUf+45hhNKUnLGma9XrKSI2SFUpVMOBxxLJZbmqfJ7CxuT
h8MnvRmHGFC0sAw/FFSb8apvrCSb997cIbBNJbFpQkOn17jnayVLE2TFepkX361qU5AFe7xMhCHX
mF53ESENUae2Ln0dr3ukDg7dtoLPoTIu5N0cHMK4DiFvU74Ojdh3K5nFGmaPZ5OMY6zGMX4vCT8Y
ZmL+hF9FUyYtTCK9TA37sBsNVTETEJBSM9LXPvhKGNKcNfMEtFbFLgQdDZ71A2+RQu3d0QUM53ha
/0VSFADsSkL/+DWbjOXLYJRRc9YUPhnGGpMC3yRltDJ/FJp9p67J/+M17C8GyjWeAIctBBAm0ROo
In4M26+2MH1zo+khjZDapHj0Cz13QHwYE9Vj26wGAQX25C7C8BDHzi/Nhtt5FzIw5Zjee6vxTqSq
wdbkeoT5+z2ISiXJpgQY3lsjiv+PYbNOPgb/WBfchISOMbNSAu28O+P9sZF9ExSf7lwjFhuu1U4S
Huf/KKN361XpgOphn7m1/9qdQ/paPKkd8w3YJZektiKrQYPAEPg3dnrZ0yJhTjpE3Dui7ILC6Rbv
soD+cZCd2RN5QPyD1IXTG2JLwwFHeO9JZaCnFD8l8LBfr5vk3oJhmB/E5Ft+wC4PN/SS2Bbk4aFx
E5hXebcCCTFLo7TL0Dz8J1VGqcf+SrjWrB5AF55c1spW7QYPFHJ+gDpbAxFfTEiDZENROO/mQt4h
nTfDrkKuuQDSoRi9Ou6i+X4PZ2XumsYNQpiOiEAqVzQFEBe3epYzfsi+vd3YMlNZ47TdI+VIcKb1
mbAHy0K03R/ycLN/HiF7heUx6pSegvJIMQs8hUme7ruqu8I9rQvcqU8nG9H3ezafnnCKwfMlDPTL
Xs0oON3YaHZ8XaJbVhuJWIf/hsUYOWWD0Yg7lTTUhgMteGAEDBFZVMaffF6uooHAAqrG/OO+S2cs
LdXGyM6NHKOyZor6K5Qg4geodD4wBfU+aTR0UKT+UFwGaMznc1i4VNPF+sqrQvt9kGECn1y6GAPV
IuPC6IPyup0heKHtSVoGHv+NAyd4djgojBpj9SkogAgUB4TQIYqfIduqFIrA2yhfnDNyBhyPmVfC
7OAq2ms=
`protect end_protected
