XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Ã�4f��
��8��o#��w��0Ķ<8��3���f��!	|~�`e��0ǌj�\�ق��bޙ�����C�A�0E'�΅T�?���G�\j)���ն��ޓ#���iU�\���
�0	#Jb�u�B��vo���m��"�>�F�>��-�~�1����U�2���!��g�z��E�jNZ�M �o���4,�^:����O����=B53�����~�����<�������_~���v�� ���ǹ���:Aο�(���1�]o󁗺�6+
Q�Q����+
i���v��b�ϔ�HĤ���~KX!�^���B�憯&_��w��#7�U��(j�?G^%�BF6O(�q<@T�w��0`�!�)�!�/�_~�Q%rer�=D�F���F�w�p�W�%VQeΟ��0��L��h�j)�tJ��h�R��wСi�����xlQ���2�3���]$ �ӖhRfLUΪ�ݫy;GX�y#<ʖ�jp3��
|-��?�>�rr>S2]x�m����gk��b�1��4�����[�$�� cJ�.�@���(��=���5T����BcR1∲�::���R�j��3�8"���y�M��`u�Yy�*E.30	�-�Hg������l]UMe��]�F1�ZI�C��65�i�lWP�X��y5DyPK�h�\,�2׈9 �<�r��(�I���Pq$��~�uGd����c��G_���d{�_�'�F�yNԟq�XlxVHYEB     400     190k�3� ��ʟ�r�%���~%���)yW�D�T�nG��^D��v.a>�g>��;���5�����i���L�0(��0���tD"�d3�e�e����3��g{R͚�Dt�ߐD�np�O�S.��=C���Ф����b��Z���)�^�쮜)�;
c�wb�uz[.��)�-<�Y�1��V=
7~�7�ü
�dJ���	���1�_��!e
�J�#�*X�j&4�SQ*C��l �'�/�(m�ӻ����@��7���/qvǾ��J���Td&�>��Bfu*��� _ɏ��	W��r��{k�"��ן�ʴ����h�'���L���$�z������c�xG�XB,�r�9�[d�V�2[�0+l��&�H�ՠ�]K������B�:�*XlxVHYEB     400     140J�yp��hɩ��J�zP�νe	��$U)oϹaD�?^�W]\�U�;������pAI?n�n���H��!,bP��7���(sHY�k�'�����Y`� �0��wM1F|��(���}`��6� K_v7������e&?�5Ø�����I�ջ��@b�!�w�y4{�!�Q@/ >�O�@�oE�=�Hݎ�7aQs[�he�֬�T��a����vN�P��i�TJ]Lt�^���iZ�� Ŕ���wAK߂a�z�F7!'^�ș��'��S��[ƫ�A���ϙ4�yg��g��#��Q/�ÕA�@�B��� XlxVHYEB     400     130=��;��;����3��?Y��'�շ�Ct��)�d3js��äc���C7� �'�#��I�l���v6���`�2ߒY�s�h��!��	�5�G�ׁ�j��lCw�h�*a�r4�EK�<dd�=ǘ��QJu���j�i��~���;6����}�?~�q<�v����'8Ӈ�b�S�쑣�U�-uܣX�p%薸�a-���8�C\s��a ��0(�����/܍a�snbU$Pm���>	{�g��:a>X!���x�Źs�Q�p�1�eⵚ�r�\�6Fu�z�B!����XlxVHYEB     232     110s���Ƹ�H��h0�n���Z���*� T�j�0���Ss����"62�#��!bqk%E�Lة�v{J!���B�v ;�z��$e���.Ng>L����Ѫ�Uj���UF�z|�P�w�\�c��uI.�Rp�9�"�j��r��!<�����K��B���z�  ��L�|ǅ-�S@A��0�q$ZJ�1p�z�9$y sPV��p��G-�٦�1���'3���+��j�`챥��$�͌�ϴ������jG�Eu�'P����g$