XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v�z#�zp����GlW�]�Έ�.��`g��P�=�<ǡ��?��Y��g���lg�&�,=&���dPܰ�䦃�q���ý�}o�~ͽ��HT	i��L4N���p��t�Gn&����p�ȒՌO�.���w��/7r�hz�z�_�h����r-9|�|�����z����E���U��4����O� Y����6&��q�"�f`W[�qr�lA��x�+����[2�����>�K�$�/{�_����G�PP.
0x�8�[�Iۊ+���H<CC�ę^�y��Y�z��ҌG� ̎	���L�o6ʟ*��{���D���]%<��/.��$tE%̠�fN劈�U���t�4zҀ��Υ���Ca.T�m~��n��R3��&�����p�4Oc�2v���t�j)���E�>�nI�`j�]}o�-ό��g;p��8D��J]�����jH�m��� �p�T�,�8���/���#wuP�rWŠj~�w�����A�r�AY�i̙��_M��/��J�=�'e})��l# (�G�uO�1a�v��;P�19l�Gk�����?F,d�S<U�7�{� ���g�� ��\��%"ng�C�{Y	/d�1����Tf��)��@ރr���Y]���@��~����@��	��0U��T(i��pY���:c|C�t�{��UR��8�C@Y�ivL���'ԑDy0Z��ƴ�83|�0��A��\A�E#-��`��Z����XlxVHYEB     400     1b0��Ǣ�!�gF���m�ZɺjNeAc�&)��bN4�i�`n��F��%/t��7n|P�xW�L,_C�Ȋ�Ԋ�<�b��'� :�����N�7���y�y`mj������:<	�,�Zhg��ں.��y�D=VZgv�:���盿�G�O��+��RK
�x<�J��xnrK������j>bl#f0��\�	��iVv� !J�e��}�wE��?� �ax��d���zo�	�y���)���KB��9� rot2�ĝg3t&�=W��.��ML����H�F�ķ\�ߙ�N��L����h$y�����`��,�5���,2d��Q�Zd"�W��
�	�PBMӧO��]��I�I�J��g��e7/m��P�a�T>+CZ�/�'��S���)�p����Y���@W��N��D���?XlxVHYEB     400     1b0��X���|���X�@�����4�M�k7Vf4m�
����A&�v�Z��(4j��b]�x�*����E�{?��%]}�"D�`N�׃�Hq��Aī��.��(�=�՗���O���]���y�����cC�u���)�`���Ep�%Y�i5-�9�H�	�y��? ���Y��m�_^���_���K�ͥ�a' q��ٗ*j�����l9q#o�+L���u���o�Zbo[�NQu���ɵ���NM?vU��,�`b��,8w������{��Ť�C�0-\W�!����1qA�Ic�?FT^��(#�Yu{����,2��C��U�g*h�D�4�w�B-ɹ��'y#�ڣ�[ vt�V����Sjy3����K>�����EI4��WÕd`���e����M9R�iqoC���A�XԗO[�yXlxVHYEB     400     130[��0����vxO�ou[:������H(�
�Fִ�����\gf����R!���`��m�>��z���O2\z��'��B�o��Z��lF�a����)Nf*P0W}�����0�V�D�>��I"�=$���-W��_�0-��%�Eo����	L��g`�[����v�r�?O��)V���)�<��9�jD�C�e�3�esW	�Z�y� (Ѹ蚔�F3;�k(������O��;N#ю�_�2v�6rcӈ>UE�L�x������}vg�l���Z{WF�Fh����l�L�tra 
ͧ�ݕ��EDXlxVHYEB     400     190�䢙F�x��8�?��&n� ɠ��k��R'K	y�Cʅ��֊Z�C9��]��Rd���3,����d�1��Tke@��,z���#�p�����:�m7��+�����[�㠽��}���������<�Jz����S���S%�$=N�(X�,Kpa�y��s�x'U3&��2G8�>5V|�g�p��P��j̛(P��|�_F��ܼ(�C����,��iV	,VD�Ͱ:<�55�a��������-{����LQ������SY�1�7{�9�`�\RKU�Ӆ$n�J{�L��ݔ7���<�w���ܲ�C����<��Sl \6U��dL�����0���+����~�k���B��ؙ&���;�*0�sE�����B��l�-=XlxVHYEB     400     160;ކ���t�Ҵ��]���Xz �u�,��	�/���ʹ��$����K��v��U+>��tJ��GSR���ūἊ��'
�����+�Զ�	��R��)?K��{#7Ζ���� ��)�?���V�u2��`j3���{FGY����te�ziaUN���T���/��_`��<�?{1]6�M �\�����:[����S��`p�����E(���e-�5�IS� ���>��4*�䙿P�*:��#!ˢ$�v��h;G�Ѧ�@��֬[d�2J���Va��,K��("Ux,~����u$���$�˜{%^����cf5K.�O�
�D���N������dXlxVHYEB     400     1b05�"��Y�d���fz�9�������l 渰"(�ފ����݁�<$�K�3�4���D(K^���q1A�Z�=���2���j	�gX
�5���7^fOZ��Ƴ5�W;�:(wB'H��:����(i���Wr-q��E��m�
Ϣn�r,g}K��n|��Ȅ-�2��U-��Ֆm����O�R�Ace%���/-�%&�� n�<����<�r~���s�d�i��aQ�*���u:ks"�I����Sx=:�=�FBtژ�iJ�ϋ:Vb�욁�݂�>�3��/�5�L�r�\ܿA
�/s�7l��粷�°G�`�U8+���8/�^��R!E2�MB��女+�
sL�q �O��?108�� +���n�����{�䱘�/u~t����[t1�5 �}7��f���XlxVHYEB     400     160���4��`|In�.����ﱻyp�(dE��7���hs�`aIa7��	�7�����Fl��@��Wp�_R�y�;���O��/�6���R�$��X14��C86�	�䉚�h� ��r�U��;	��^�)�Ou�#��8�'TOAR��u�"Q���X���2�����I�6S��J�.�a�b�x����|��̏��/"���~���`Dk��	۳&�A�r�RP���O��20����~�2�_%�2�Q�DDh�nF��a/�[;�!Հ��I����]��x�ӸP��%4F�	~ݒ�f&GŁֳ��s7"T����m������T�z��-߂�8��XlxVHYEB     400     120_�5-Og�C8I��'�AbA��I�>4�O�U�G���/�� �$�w��<d;��?�B8�/�!��h�T�����8q���%����qg Gf"gC�q/F��V�M��7$���أB>w -a����$���BЈn��ߔ���<����.D�v�𴈨�W��&HHA����"(26�H���^G!��,������4�ϮTO�-i�-2�(;�zr�"�U�؝O��^�$B�B;�Q�S�.�4�\7D�r�D�Wy��Ύ[��d��z�^��S��xA�Q�c��XlxVHYEB     400     190uK�fhH��M��$2��T���[��M�#@JO��%��������jY(ʔ�Fq��J. �Jͼ�|�}Y�t�˔��,B���V�����2�YGV�a�O��/*=]7�U�k��M�/��Q�۝v{�^�{����F<(E�$�X��J60k�To.��"ˤ�C{|vqX���pIl��y�" Cy >2�	N
��:�{�pr���������!��-A�77�<8��{��5R�4i?PR��]׼Q�;�W��o(�D�w/o���W`9����]<F&�v������Nrd���#���`�t�PY�i���I�$a)�y�N��19r��z�gH�Jb
ԍy�-KH��+�7$d�@�Z��ȭ�ut�Ҡ_8YP�(�W�w7��~�k"XlxVHYEB     400     140r�ńm�3������+��hP�@M����Ũ�8��V}%����;�L�#��b��������I�1��5�|<�	�#��m-���k$��
u�j��I��=�?.�1m��(�g���V��}.���8-�r��Sy��S�7G��lpT�3ȝ������7�g~bjc�"���.�].�x)M��'�j.���K��xz�+�~c
<GB5^`�ЂB.��g��I1��p�9݁�s}mV�Dc�<G4��2�A���t���?���	�U��`�
)�9�'��7 R�� ��r'2�WR!��XlxVHYEB     400     160l���i�/�ۍ�����v��h���7����1�N	��Et���~輓x�ǀ�F�9B�:k�#p|E���ӡ�[o�~%("�W����G��hQ�)d��J[���� �<���T�(g�[s�u'���y;�`VaD�r�z�T�C��%k��e����Al��C~�y@�:d%
'�+�IǇ�Qi��A@w�b��A����h� ���pX�o�XNi3FR�E�4����t_M���M�U+;���N���U�S�,r��N_=��N5a��?Sv��~�;�'��	�ߌ�MN��
��RX��7μ���Zw����?���bZo/ �Z|n!��hzXlxVHYEB     21a     100o���Vt��X`łR�\�����夦P05y��"�Zߕن]J���#[��^|���X�rSU�������>�ߺB�ϛ��vƾ�BXez�̐u���e2(�C�43�P}L�����m'֭E�FHw�9�,�8/��:��)������{���F2���Jf��?����t�<�Wl��=�+��h�����̻�v�E�aFA�yտ.�6�̲9�H{s�*�e{z1T�}�������B�>�CDR~�;�n��3�ҭ��