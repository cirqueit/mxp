��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���?f��?_v8����g�a��!�9��>��u�}��-}u�Yv#>BQGzwv�v���;�Zp�鵻1L�t��{��XP֪2�D�p�x\X�wbBi:6t�����o2��&^�	�M*���Nt�.�C�4�W�W����H΃+���rz���{��[s U[
г~�#<����ġ-*!h���X��>�;��{P�����th� 7��s��ܱ'gJ���ȔϦޑ��b�>�=
���]	��vT�8�µa���#���DL�S�S���8�����ɸ�zZ�u��cCj?P�{
��|�%ꎒ��u-n����{��A0tt!NOk47����{���^膓U;���vj����ŀ�^����N>�N�@�9���-� �y0�tw���:0���ޭ��<�Ne埀H<4�el�6�|Oé�r($^h�����������=�N�z]dB���va%*�!ٌd��݁!�)����[��Os�M'Y���,8&L��j��1��Z8�?��A��V�/:���`��Z<-�E��� .�M�Ve;��я�L|�)����ج��Я�����J1y��$[(.���o'\��)�l��l�(�߁�
go)�j����!ݤh��}w��ET�j�UBZ�9��S���[f�+5O�ǅJi@3���6��@Q,�q4�5�%��X�g獍��F�ߢ#�T߯���R����`$Jތ�ΊH����b��p����s��E�B[<8/�'�O#,����gbtϫ�r����3�� �DZ���1]��������e�K���v�ԙl���x��&O��&�vI0��T����̫�\����i���+�b��$0$i��;d��k�w�S��T�n�_�]�=qo8���k���V������|b�����oh[U`g�����<�P�M�4�9��$��e��� K���+!ڟ� �"6YyQ��:$�a�f+�MDױ�Oe}�'��!��S?��(ż���jסȀ;X������a���o��Y�����+�N3�_� *�9Ds���B�m��A'�7%�/мd�o7ZܠCP�n��+��Đ&B���K=+�:���nj�k��6��f(�8��<�#�%{Suׄ��Y]z��R�﷌�~ .s�Ķ�N�� ����4�����W��B}�l�4T0́zJ�ӮG��,>��Y�QN:���.G�F8qeF|�����U0`�@�S,)�IP�31Z��ρ���ƪ}�q���u�� ��'J%����װFc�TfP<�D���^���~�sP��9�����]��V����cI3�ʧŉ����Ɋ���:�H=O�,���]0;�����j��_�,Qu��4Խz����ܞg��j�v��DtU��_g�ڗ