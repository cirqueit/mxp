XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���L� D2��*�����'�^�W�5�:ۗ�O�3��p!e�	UDɠr+f[7��桊�"ѽȏ�O-��h˽q�1"�̒Þ\�{<�|Ho
�5Z��k����ޖ��>��ӃTk�Ц��X
Y4qu@����o6�:�5�7K�޲��}���K���{�ʆ���zA6��V9ے1�e�vN�
z��l�g	��Rsԅ��`�rN���
Xj��d?��1�/�:��J޼b�^x;��9�~�'���O�BM�&�s�� ����!;�Yل��H��zW��Ą2
xi�� GGa3�Q��j*lL�wu�xt�:B��N��[XJ �:��f�bS�HUB��ң�AY3��z,��xnʝt�ޕK땀�l��s�&��rp�P7���ZJ��q�!�@
n�@��rRz��������o�v������	��z�Z;q�]i�o#Ɯ;$$��P���
��	���6/9����;�n_��va?��pLBՋI		i$Hj�`�z�jnc
��X�A҉G��!BD-RV�8�L-0{�ZW׾=���mX��ԱEKD;�1�Ǣu"I�c�|��m�8��޶�2e+��_��4��3�#������E�Pә ����_{mNo�b�w�#��#_�H����8G]��iK��/cmTy����D��7A �%��K:�W �,�� ���Z"���N��n��Q�aW��*�D�ó_���I%e����������y��0*�.�(l�XlxVHYEB     400     1e0�?�4dmsx�aC��
�R�G��nSĝ�'�A���(gqP?�P�k[^�i��%���xmըU��K�3�@+�ul����e�q9N \����2��g�C��2U�ذ�.�S%��!%y�)��k�R"���萳��_��9e�A:�d�!CQ<s6��r(z8��s=�r�ԅ��ea)f��͆�Сh�Kx{?ᑁ��n��b3u�@��v��A����_(�Gi�������ݱ�]�F��XI`@?+5^�Gs	�϶�,����r�<6�V��A���{)�f�Ld�!@4̈:*��IϔJ�B%OJ����Z\˕���[i�cq�mЮ�=��jG�o��eD���y�H�H' [8���b*�M8�H���Zl��(bA�h��(�R���
��7j�I�]��r��"3Ě�b0�Sq��9'�xi%]3��!T�H������Jy���y+��嵷��ºl����?ɝ�ț�(XlxVHYEB     213      b0��z����+l�E�����%�N&_���c�.�&Y�ܼ�`f�c��8�a�ЃJ���=��;�
�h@�� x��nvIia&�b)ǻ���u�=#栐]o\B� }�!R[X��ߊw~ _DqsC���Fÿ���Bϵ����$�@��Ґ�Q����!r�R�
sԫ��9����