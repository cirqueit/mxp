XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X�O{��B�hqc�ڝ�������H��1���\XMZiN�>�46���,QO��[���9���LI��u˙����ݖ�a۴�'�X�M&�;�$#�p�GQ]^C��O���8G���K!�Ax������L���z
Ҏ�a�i�Y�V�N}f�q��x1b���B)��ϧv���nEy{�^��#�Br;q��*���9���ߦsJ�W�7�Tb���#0���F�UPA{�Ljmxn��y�F��WXY���`���H�Pk�^]���_�8E�}�B�����d��<�,OC|�o�F��^������z� �y�>m|E!��8V��\ղ&��mNCTj����RV	��^_2>V�ͣ�&w�y ���覀���D�*��;<�a�,��K���q�����V�I�v���-,mCF��W�+����0(T�TD$���N���Z8�xv�?��H�]^�<;�!���+U�';I��F_�ϰm�q�GD�Ra���ޟ�Ɨh ���֝ɳ��Jv;�����{�4�I\>�sa�^W&�~�3(0�%@��
@?7��	��+}�&���kl#s�P��$MO�C�$�]$�(��?wO2�awl�a
�H���[Z��Դ˦w�6��oo���w�
[Oj����b��� �:+8�ߏ�v����a���1���{��Q�������u ��ľH�ύ���1M�i�{;ږ���`��А<�s���7[JqD{�L�}4�A��3#Ù��:b��*XlxVHYEB     400     220�����'�G���Lx����p���[m)�
Ip����6Z 鲫:�~ ��9��mFi�d?�������W�-
����/�\:��6q�æ��Se����M8��^_jz�	�,��U��BD�X�"j@�%�	���w�9���=b`��R��kP�$e/��	z��3�:�{'9�5�q�����|����t/Z���H(,�	�]L��4����:��d�pt���H�Q:ۍ)��.Г�.��Cg1M�A$�s���5;�*�
H��n
�� �ד��43qPSSr�(�i��;�ūN�=a5z���7.N?r��ʬ��d"��	:\1m��YѨ�
��|�b�S�߇$F~�XR��Y0��q՘���I�����a���(Ze��o+E��;V�R���?5_�H�^72��6��1��3l��)���%_~��,I��<����ܒdL^D��q�v[(�A�0\�@B����^�����<B�fH�4RY(���QcBT�2�Q{eW")�`g�6h�$�ܼrO���XlxVHYEB     400      d0[l�j��}>�M� �<��ܙ�f�C#�1�,0�t3���ڽø�B��vKE�#N �'�����5@�n(o7��{jy��ޱ��+�O�$�-�V����"jL1�1Ŀ�W� �X��sBIk�+-݅���+�3𭓷}�#��e~�o�RN+�4���ب�25H�����i����	N;}�!��`ㆧK:��wӦ�W�PG�Ө�XlxVHYEB     400      c0p@xӣ���@I��1�[�o0(��=.a[��r�=#z�re�F`�����;����@���K�L�i�h2�eYo��uuo)�g�FOC;�f��ɭ6�aɀ\�˿�쥏h�f�t3*�Ioxސ��x˳),�j��١�=�6�\�h�	Y7�y�3�5��#�t�@��D�ǁ�U)��\Q�ZXlxVHYEB     400      c0�Mg�\��&�b#5�Y��{��5/�/���������}�Mྨ��<�5���`�i�"�?�H\W�(�����"qa�v��=�6��C�v����
�ʴX���o{'��cTiy
��j4���h�:LHt�ea���&��XL� O����05���u�TE5�*خ�Rs��j/>����XlxVHYEB     400      d0Q�>�Rg��r�$>lvN�i�ZKr�ڃ
�W��Gl�i-��P)�К|�4r.���a��X��(Ec�� 7g�k����MS�R�A8����z_�D\�4���S��\1�>gt�6�Y��絊�I� ];�mZ���Z �ɒ[,�6��] m�w�����yG~{23��@�jfY�}�S��9.>�#IT�N[0U����XlxVHYEB     400      d0��P�!7�ڠ�<����K�oF�Une\��q�l�L��HYj�'�r݁L[�������	qX��eX�̗�f#QM�_�;R_�f��LM��ڴQ2Ǳ̃���/a�>B�}3	��z��~G���"S|��*ȧ]���"�|��6��{a��y"!���$",��g`�M��c ���-ɵ#?)�z��$[_	�-����]��&�XlxVHYEB     400      d0��b!��W���,C����A7���@@�\=xC�����tHjV� ��p�5a�Pt ;L�5@ײl��.ш�$d�g��e5S���쑸U`?)�/�9��J��1̻�c�����	9�h@] �/t;�]�@7K����6\�<jR0m�j[���n��b�SV�o��$��+ 258�K��b��V��n�����roB�f�l�=B�XlxVHYEB     400     170��%9@�ܕ��>\�vuj����%��o��uK�4��P܋Ψ˳����rL-U8��mq�^�2!��U�Z�w�>Z�\ =�>����4]�TW.s����Z=��`��8�?�$RF�ӈN�����u��w�o5/dj �{G{[�[tj-�H3a!0��֬}U���k;T�u(���3)��s�O�����w�����2��L�L��  ��気%9��a$��$T~c,��C���𙷣T�2B`��K�F�g�+�G���܉a???9����'I��AL5C�귶��[��+8�b����m�Gc�s���_Ll��F��n�Q�U�O���v�k-��hT���(z^XlxVHYEB     400     140}5Yc�]5����c�jR��K"{�d{���ϣH7`�Q61�#Rc0�;~�>�%䀿6)r�+>)�#6B�X?�4B�	~��8�W�gL�<�lw\��+�<^^��xY[�ftj}b�e( 2)Cy���yY"���7�y�tk�5����U�#$�n�:d(�+z����%�@0ى��L\�q��{X���i8�o�|ݢ�jW�#7l̂d�1(�h�&B�M[#q����˄RT�:Lx���]+`��T�֞��(�^!��H�5��֛��^1� �xJ�u��':¤�	��u��,Ax�١��^A��c���C�ס��}v���7XlxVHYEB     400      f03E1(�{p��sWu8�Zo�l��jM���7"1�)O��H/���N��Ee�a+f��F�t�|nн�1C�y���2C�e,ca6�آi�1�0�f��g�߽�dIFd{u���S�:ٚ�X:d}=3�@2��mw��N��݌�Ү7_C�~�"���dMC�L���z���\!��BU-�"�y�S�ѤВM�q˩rX"n{�d!��]=���O͸��^������j&��XlxVHYEB     400     100&�W�U`����Su|��e`�\�$�Q���Z��ލ�h���v�8�e���������&a�˾�`������=VQ�o���:W���߈]ϭ3]VQ���#3b�o��*#�������V��ܿ� 0ĮQ��������]!���$�ǘ�F��p��4����eDZ9��T˛���6�7D����8j��C�QI]b�(�O�]��`��~t�%Y	�E�atAמ�.vLq����Tc(��7>�C���Q��XlxVHYEB     400     110	s�׋Ԁ�`691ٴlU�D��M�vZ�x8�eHY�<Q�]��[`�eo�e��(JF.H�6Z��]��ށ������b c���e�V��8�ye1xjB:�V��g����Od�%��Àǌ�\�?g�����|���9ݡ�c�ɇ�5�9�3��F| ���]ʍ�>���Y��o�����������D��vU]5�	���΍1��`Ym���h=�w�V0%>W-rŘ2Y4���<ju|�$�Np{]�<W8��XlxVHYEB     400     110ɷ�q�3��`a��R�K��1a��6�@x�PT8�[Mϡ�l��������D�a>�+G�[
�<*R�)cc�q�'�e�x'3��#�N�ϭ��BE s����u��n6u����ֻ�V�e���;�n?$.��=[��?ݨ�$5�\.��z�\�i�,V��XL�K8���$'�3%��0�����./����a�g���U������$v�Z"��'��O�.���|ȍX-���W+Gz�j"r�ٛ%+T^`�-��\�fs���XlxVHYEB     400     130��L���j���ƣ@]��?w|��^�+%�"	o�J�h���h7����z�NI�9�aZ�'�������%�C1z�I�ln��3�Q�(0���z;�B��;4s�.�aR�e�/����
���q�|	H'(k�Iz���1��4�s�-qM�F^�m�j�p4�l5a�����G�*�����l���ʣղk|) -�m��e���*�7�Y�6P�9����8�D��@� Ӣc�s������X��6�BS����:�h�2F �d���	l��Z�!�1����Z�8=ƿxfvҴx��XlxVHYEB     400     100\-�1��㲈<���-b���.�D/s-���9uI�����)�q@��E�׿Ԝ6���/����/B�&�ح�&Q�'�W#��	m�	�ʯ�CMr���ș��gq[�;�r�X��1�i�c-��~��3"N3\�L Y��i�q����M�n[Xp���D~�H8���C�)s)��'1�.h�EFaO� ��6G��cay��T��y��MQ�.���d�&�u,�(iy59,��:BZ�����}��x�5k�����X.9'�$4�uXlxVHYEB     400     1007%���*|�f�7dQ�e'E���/�oME���E�3�3�h����q	�/�G�Yp�'�x����tۈ���Y��;Ɨg��겉0�f`���B�Q�Q��xه��X"+���W�Ă�f�P~w����!"o_�wn7�A{[)��<\�O\U^�S�m�Hc�h��9B%�uD�����y���p�5?����e�'�Ӵ��N���'U~)g����:NlI���i���Y�P�q+�^=M||T!?u�XlxVHYEB     400     100����&犉�&WbY��H�7�����,�
iFZ�6��P�
+>½�xMr����F��b0z	|��*\p�s��⃀�@�/y����ϴ ��e/c�N����׷@A�w`���.��Е����)5:��6;��3���R�b�9�K{��m � �~F��ӭ���`ݹ�!Ӳq�|��?�Ma�S?�#vQe�C�s�����F�N}�����	���m �.|x/����6� �S..y�jf�|m�ݲS���~'XlxVHYEB     400     100}]�K��qj�|��]�%��1̇(��7�	k;FʭGK�[4rC�Z o�-� �	�&湬���(D��_?���=^�����/�ݒs���k{Y�l7�š���/<S�]�>��Õ�� ��5z���í�C,��ݐϑ@ʨ�� �������𷟒.���t�<���JCpÆ��#�	v;V��as���jt)�`�/��
Z��_��d�Ψ��lN�HS����_�U�zo}���(�VׅFª.~0�XlxVHYEB     400     100����]4��ݖG�[(c��(���[�
*o��@�~PT��4�r���:ay���BW���ETT\?�F���߷�$/*����ASoH�=!;e+�;A���U�#&s\�0�#����6�������B5f�o퀶bv�盟lO"u�_�~�ҝw�r�,���f.%�4o=�<�I��:��^��(8�����j/�·����
�m�_���d���I=;�/��^s��1|~�CͬG����XlxVHYEB     400     100�͌��Mѓ���9ێӉ�U?�B.u���]����-���W�b��I��p�6cEL���`{�Y�	��#�Ӏ�����PN�����~��)����A�Zh��la�Ҩ4c*`Ċ/���(I��85R�8"E.�Cw���9�v &g�y�a��������JG̩�K_'��H�2g�:{��
R��:�'8�f����nm>]9����J�d'-�d4|�y��OW�Oǈ~r��k'���b�Fm�XlxVHYEB     400     100�gs�f���"�����w���V������ �ڵ��v�%$ja_zC���7MH�ۓz���ZE��A`]G�2�ɟ���� �ȑ>3���1��}#�W��*��U�h?@�^�W*�a��g��O��h.�%�)�9�K���J茀�S3�ن[��(\�h�27���7髵���xG6]01�(�x0n~ r�2VT���q����65����L�#��<�?x�7K}Z��M`���Hv�mb,XlxVHYEB     400     100P�.D��$�8S9�lKP��şp'��.T�¥�g�iV�����҈��n�,5Ju4,x>�ݭK���fh%�=Y��� �ꇧ�	i�_	Z�z�;�z��Y�ȩ�?M�@?w�"}��^�����,�+�(}f\c�_�1�|�na�"�R4�~<D�� �U�_$'l�=���`5( 	�	����dg���p�2�	��e�{� 0gH�-�&�)�p~͡���/~"��w�l�Y�L�A�Y`�EYXlxVHYEB     400     100���=���p;˺��.�F�Nf�e���0c:�K��C�#���C_��4��gG�]#�{��/��f'�L�(�:�-�*�#�O�l����˄8X�XPԄ �N�֥<���#I�9����>%���� JE���)㩻��Ո�Q��B����h��ENűq�7��0��q�f��T'����A?ʎ۸�ut_PQ�m�;���ykGYko�ɩS�բ�5��4�J�hv�ҩ�X%E�����s��<MXlxVHYEB     400     100nn�? @�I+j<�C
�V[��`H�ʄ�vƻ�_0x�$#�qX��`�H�������
oɍDeM���ń��Kj#�EV�����W(�>�a�7j�o;drN��Il�k�6���<���͓P5Z��k��ǨEu4���w��<s�u6��휈�:����[[���\Rh��y�D�^ڴJKfS�:��&<�$��E�RF��ژ�^^X�"�E"���yw�_cE�	�Nw�<�ͦ����]�~x���XlxVHYEB     400     100��!�ˍ\b�9�(CѝD˾�m�F:`B[����I�G�Wg���h�f:���HuB ��@�st-n`�8!X���k���&a�B�{\H1��}W��0��+�0���*�_62ڋ��-Jg�i�w������%Z�ѯ�iQ[��Za���p�Iϻ9x(��;�XE���2�.cPTO��R| ����:�S�鋠�(4���2�E��(yKft@��������<�~¸:E���6��y[q�Ȟ-9u��#�*XlxVHYEB     400     100��;���_H��zD&/%����3�|v����\#���o�ƇM��cƆyn��m�K_>:"�s'/��k]s��x��@5у��G��a�"O�ǬsӶ� ���8���p�~�6N��%�����b�wօZ{A�~�RR wm�Bgez<�|�a�g~@�	���c̎�.���&��6�vC�}R4�hD��u:�W�,� ��"�Ǉ�����'��`j�gE^5�7�G��bL��2��g�C�3px��XlxVHYEB     400     100D<c�M!��d���KU�Ӕ�^�ܥ8���#��;��p7*1M�>��*��A6se�:������x�����CS�r�2�/���N�q]�N�HQ�����2\�C��FB�
��
��C;����fx_�!�0t�T�����ق�H?�l�tp��k�f�_�J5I���3����42���&[n�uz�����5w{<(�e�L���<|�>7�="9ݞh��8���9s]1�8�ݫYM�8{!���i�XlxVHYEB     400     100�Q.�:�9���L������)��r��sQ�i	����iC!b�_Z$_7���?���Sop��#�o��0�=���>���N/��͊E)�Q�h�#�K��'B���`�V���fF�:�1��sO�O�LF��������#W� �z��l��B�LW5A�Sַթy�M�� x��6�Q��{�(���M(���Y�zS���<�0w��6��eD��6��v1��s+V�ˌ�y	��t�Oi���cQ��XlxVHYEB     400     100��j�4�AQQ�
�k=�������?註��@���!�k�q�~����$�'�p������R[X	D
���h!3��4����I�9�08��.%ͼP�Iނ�y9����N�i�A�
�H��t �ƍ�O2��v��b
��* �w�?�5�y$�&�v+���iJ\�7G|�w��msEr�@P��r�*0 
v���Ǳ�)5N�NJ)ORc�(�hħ���Z�v2�AvǷc��s@�pZ/�xm<��%�w%XlxVHYEB     400     170������P��#F�������#��X;&8�MΪ����錹�#\��֓yS��Yg��ޘ������xwM���U"��9�kf=qj(i+qt�I�L˹L��ρf�\T�ݽ�Qy`�4�M��|ŗ���fN�d<|����S�Voaa/-�p���'��m��!��5d��j���m�^�+S �B���I��"��mMx�ⰗP�١�	&�
�%��D�>[(��@܏����8j����xX�	�sΠN��x@� 4�C3D��{d��^��6��))���IH����#]M0�_���$񗵺T"�e�/O��3��U'��|'ݛN���p�8t̻�g?�)��,��rO����+�XlxVHYEB     400     100��X���M�7���n%	�q1�w��� \C����B��tkx������܇�yQ8��9�EՕ���ˊ6�k ��Er��y�Am�����w��֙Gj�����	�X
���Q�����.֧��W�qxLUGu�+��Tk�6R��pw0դ5(�O�/��&Rk���`�j T���=G�O�
oǞ�"/@�~�A�	`�V��ؔE[��z�^r�UƠ�= �`8	8����Nʮ�̩M�%ᕚ�W�ڭ��.&�XlxVHYEB     400      c0�8vJ�&�Q��3�JW�{4�	�T�q�(i"b"�aOL=������N�eX%,��2�^?���f.���4o�̫�%ga^�GeSw)U.F������2�ҋ��;������]31��@:�dڸ2<�*R1a>��t��|�4��r.�R]�T�$n�3�%�I;n+1�`$�l>IM,��=r`���XlxVHYEB     400      b0����Z�k�xO�D�a�9F�k�����Ϥ7 =R�@6��E�Q>*�Qw.׬�j�z��d�4Fa���P�\rHx��.�|@<�C%��������(��h�r��s�}#�_��floewD+#�@��@T��s���.�/ 酐�|r;�]BzT|�����{��$���XlxVHYEB     400      90�������X�����au�G��C�Q��N���jð.��0��e�G��	�2��]ʲ��m�o]m�(Ə�_�n�^'So���W��N��E�P�L�f��hϵ
Ļh��|O�����Kf�N��۟�N��P��$qX)�eV���XlxVHYEB     400      90~!�t�0<n4�����g�Vw�
����}�h�q�^��p0�� B2����G"�r���z�����B����_�KBu_���š������a)xs��m���g_��L��bp����^���V�o4��6,�L���XlxVHYEB     400      90)��n&&��!7D�x�X��?OόK���
�d��ϒ+o�ya� �Q���荂���?w�Cm}A|����L�3+r	�eԳ<**��)�f�{���O�2�f����|�m�']L����h�S��OW��t���pG>L����'�XlxVHYEB     400      90jq�4L�d���"q>���u�@C梔b53G%�� �]��Mnj(pC��R��:�w&�=R.�����ol��118�
�z��Z��f�6©9�';-Q�c\�$Uz��������	�c����͆�B�*��B�:�������XlxVHYEB     400      90A�9��ja]R��K �e�����y��j�t'#�,e���B�~��H�DI���N�w�>�_�}SJ�� O�ѵ�9�����T��I��k�Gzs`t���6��G�[3l0����?s�%� Oo��I5i�Ɨ�*"1�[�XlxVHYEB     400      d0bS��&���F�5��Q��G=��W71;�LH�Zeu���;"��O!Bʍ3�ƨG`u(���5�ٹ�~�1IH���5f ����J�Jάv2�T�;dz�����#OjVD��0�e��:��
�˚��.K�u���)���ևIX�Jf��ֹ��~��1�}�ܼ����޺�ǀD���J�t�0��`C[�L4���EXlxVHYEB     400      e0u��g7�짾�oۢ+�t5=b?ڪ�O;�c���b�j�:A6�m��
��A9y�k���hiwNR_oۖ�2q��8V�l�o`�QNx41NE+G�(��bxC��54�U�S`�v��y�yM"���<��bB.�^@%K;�}x�Á��"�ƃ��H�=��00Ւ���aQ��_#F��z���l�+�ʤ=|�c;U�q�b���;LS@XlxVHYEB     400     100�VA��nd	��AL@�ً�ʪ�:�~�;�
0���zh�ȏ�X�/&�Kq�%- R ��##M�u�e��5�M��ކ@����j�<�x݃��v�'/�)�Hv�d����@���/ɿ���Kx��	51&֚Ux(�"��n~��I['{c���[]�,�C�P"�-��R�v+�����{��5m�
�A�S��McDSK=:9���ll숯pa��m�
�����;H����@�g��ɨ�ފە������XlxVHYEB     400     160�X0^�T�$:��xi��� �Sfd?ӫ��!q�Ɓ��I�Ñ���tX�6%�;u�/J8��$�h��n�:"��?��]Q>L�m�1[ؗ���|�$)�t��աS ��WHL���8�L���rI� �^N4�x�I<��"��j�uPp.�y�+����U<s�:�H=�sl�[�c��럌��z$���8�q�$qI���O�
[��a�B	�zʱk��߭`c�I!�Ll¿%'Z�Pr���"c`(չd��ng�|�3Ϛt�ݝu�9����֟���L��`�Q�~5_�P2�ˎ~cÆ�Fw�C}��@e��:d��C`��m��V�����XlxVHYEB     400     160v:1���㼞I�Ê/��=k�~H5�l���8���?2q�Bg�j��ZUjOM����y�bG��e+�c�)>A��P� ��Ov����8eB��������#���v�і�o	�+�u>�F~�(;e�O��;-��!��!���tK�#�9=��Q�����z�̝f���1#v�t��P9�Lӌ�9~�o��u�3�5�3�FM:!����iS{EN�̢M2ܬwy]&/�9n�w�$R1���ߟ*7B��}O��~������Cϻ~H�
��3�c�钋a�ui�S��݇�TW%�l�Ӷ�g�6�������fۛu|Q{q:��}�e�<�եXlxVHYEB     400     140���`=�?K'd0��D�K(ƀ\����S�X��S�@ĺㆫ᛭A��$g��y+T،�Ϛ������O�k�}'i!��Z)p-z�O�̊Z��ZR<rW�q$��u㿽n�D�����=�z6�iZ�$��~҂�"�+uF2Xߚ7������9K,b���N!o�rNz�IKkM���WxbX�k��|�؃y:�<���8S�J������)�{Kp���������	��:�5��:��j@�jz{GQ�x�B8��?5��r���zBƝ)�o�L�R@x�K�1��8�,	���r�j�꾙�t�<6XlxVHYEB     400     170mk,�f�ë!'p���E�m��huH�4c��"��a��ܦH��V�Q��6��<�b?�-I����9i��v�p%p��Q¡P����,�l��O��v�	��K9!�H�7l�;ɸ��&�E�Z6�;{M�#�������&�$�����1M�o������5oE���Gyz���bb5�'��;e�^A6��5l��h� P*wT:�g��(!3K��ACk��:c}�믿�c��ï��X�=Y'�8յ�V�~�k<,W�j�5�Bte�k	�$��X�7&������-��6vTdE�������vPnu �A���,�H�".�4�Hh�����~�&O��F�$�\b�B�-�=����!b4XlxVHYEB     400     150{���J1&��+���86
?��oM��L]�cv&��+*�R��7Uj�q�~�X;aq��*�1ܤ�m�g( !h��#�Fzqe��6�T�.1���)�>�7��^�@���4�"�/
v.�zxǓ0t'.�T�FK[+��� ���f��G7U�O�ǲq��:����
��#��#Mn"�<�Y{��]��9��F�Y����Ata�5
��/��5���S�P�`SkA�����J!Z�9L����o,C \,yEP8���G���a��s�E�����Ę4��>۱�z�=��ь�?<Ec�fhIds���� 2)�	ƛ������I�u��XlxVHYEB     400     190d���b�k»Ҷ�Q�aߴ�~�����)�;I˶W����Qcw�h8T�+4�A�zH���a���}a���=8�2X����rXҡ+�7� J� ����](u��sਲ਼J��%�����f�s[�^�!�������D�Y�'�Az">D/�X%B����d��!��P.Z�M���|�+s���Hz���%4�
[��v���,6�ZȨ�a/K�%N��L�[��̽�
0#��5H����;l�+#lЁAݲ5�y��o?�����*��@FU� �7VLc(W�>��H��+�Q	�?��H�dn�ٯ@-!��ѺA�蠭�-����o�ѧ�c���W����𥪖w��-S�bP&�sS���{�"!z;L��}�J]D/��6��Ϥ�@��\��mXlxVHYEB     400     150T�]��c';�eP4nP�����T-޾������{F���yè�����,%��V.�ke��U��ؽ�zv��5�}Dd} ��ky�F�,��H���������̮u�x1~�Vhu�DvVK���9C��&�5MD"�t��Ǹ
\^�A��ހ�\������4�A�e�H���$H�k���������}�r�)�V�dT{UOƆ�t%SL�~ �^�4�@�,�������lc�wɲqe����T^F��M�h�,�n�F�."[�*䪑zmqNG3����#e��l5<�b�������(���$�Zg�1�"Nt�|��x����CLX�t�,wXlxVHYEB     400     100�F}�Bo�4��ZՖ�(�@��؎���\����l�	Ή�#�r^��h�!�f�{d!��xfR�r�@h�x}+ߦ9��7`G��\�@G{z�Rq,�dB�Kb��_!�<�̠��_)0�q_}�s��D��=�jаZ��Q��諿27a��r=���m^��C�4�U�sE�ֽ�D�w� ��{R+JwC�6�4�t�5���tY�P��omb���ʇ��>�38���&������7��?%�烗���i�#m4�{XlxVHYEB     400     190��xV���*Υsp��{bW0��WC��8���@�jY�f���6�z4{����]Z�T�����p���	�R�-��9�(c�B�Gh`rN�\עǭY|h1_ݶ�;����z�����Lc[:����?,��EO"�av�RZ���[c�)*��oD�!�����>	t��2>̠p�xcvd{����A��*���t�5���63m��j`_b/� \�}�e���&��3�g�ժ��f�pF(���)�7#v���L �V�zJ�'>*�/��	ߐ����Z͔�Wx�ĺ��#���VJ�&x��I;��A�����H��>5��8O�a���� X�֍��+��W��Ux��7VI����C�^�Raj�L[}�2���|��&����XlxVHYEB     400     140��L*� �y~����Û��x,ݲ�2��*M�V�(%�ؿT����ņ|��z�wͪ����Թ��:�)�i�
��=��ϩ�ݸ(x�ͻ��(��,��rdہd����/��)Ù��!QrC+K7r�� >*��9{U��ŕ;V׮9� �]AF��nl�<�u5d�_2.�\.%|���b��,�s���f���vm2��2��1�ߘtk,�E��.��_I��0[���Z��_'��R�@�k�3�#���qF�����~z��� ��`_�dS(F<va�ey�,�r�8�l�#��ŶJ�XlxVHYEB     400     150��-�<��0@6�$&�g��r_�|����kWy����
�n�W%���	������:��;�5�$kc�=^�QNK�'f�qN��>��ʦ<g̞�-�=m�Ϯ~�^�- �3�fF�z��.c��g�,�y��,�V���!i�=��ɉq�$3޸o�3Pk��.�v�ۊ�^�m�eר��;�C���Ϛ�j���h�9��t0����A�JFa���g�Wyt�o��S���[C�,�ak��Os^�H��l����1۽QZ���l��x�L�\?���yjҿ_�q�|��Yh�fe��6�� >K�8��
OV&���-�)Ҁ~�"yŚתXlxVHYEB     400     110䳏���0^]``5��7��;�0���q�+b��y�,8���sHo\-��p9�"od�*�Q�����,�r)ݻ��ٝ6�P1Xvm[�2	C���Vߗo� �;i���!�������1(A6����?�����&����C�KZ���o�7]��a>�*8�m��X���o����B��^-]����*��;1v���|�����'
�e����9�����ܰ7�,ʩ����p4p����e�� O-R�VPi�� �М�}��Q,�XlxVHYEB     400     160;�v�|O��%W��ޫ�On�>�ˠ� �gz�����{��|:��m�V�?��:��#��F��t�i/n�ra�_̻�p[�N��5lұLQR����a��D�+F��Qyڸ��I��.˔����b�)��qO�j'"��5D2>W�3�ј%- Y������n�u���(lr;tö��E��� >%7I�@�'\a�G �V�Abt�����	�b���3I�d��X�<����2@���J�ζpo�8�؈c����p�4ۀR���\R=�__O)��Z��*"��Qv0h�������em��ȇS��j����ӝ��$)�`,����y{��Y�XlxVHYEB     400     160�&�26S����:��g�����k�[O�VȠ7������ڵ�0�S �x��@�J!vL����:u�O��l�j������X�ݧ��}�}���&Ϲ$i�	
��������~��r���.��fo�H��$�̃��@�D���gB�<J��mKC�!�JRt��2K�,4V�>j|��9g��)go&*~Vћ{�}V��,���t����a�� :E�C��ࡑ��� �!-�Ғ:a�ł��ݡ�8�G� p����P|�{���01s=�Ċu�vq��j�<xNGR!�vѸ���~P?~Q�L�����&����;+b�2��@�I�n�֌IB^���Eam�7� �hXlxVHYEB     400     150�з8A{Q�ea�k�n�	�?�I�Nt�{��#��B���ıwP�.�b��
���|NecqRn������s��eFF�O�f9&K�W�w���B���<d�^We��]��7���bq�l��Ǝ�������gr��-�T�l.H��7��.��Z�Eצ7�e�M�\�����2�=�_t��R�����<oz����{����b �$e)�r����JR�R�րi?0qV���l�o�H�4����V}��`�ݛ	��"�e��G!-^*�g��Kf~��d���Gc�|� }�e9jm�|b�N.����y��}��v��.<ﴂ]��9��&L޴XlxVHYEB     400     150�A�U�/@���b����%��Z����d��x�]�f�Z���mYs2S��Lr�h©:��K��zYu���T%�>G���V��{r]kH�[�E�Yr������{,��\���n���?.�O����}���k�I��ɟBawp�w����/8��J���(S�A��5N�kvd�t�|��H����pT?�XG4Si�JX6fV�7��V�@|�*�A'}'�\�b \�a �N6���7�W��ОGp���>�l6l)���ƈ��ێ�%":�©.�T��u��(�dNd6�a�$�hk"�SHf
ڶ�,�0�:a�������n� K�0@�)�����XlxVHYEB     400      d0����{�дh0�F��`ÚxK����h����V�M7�I\�G`��7Dk�E��#9�}#�-uqk��n$\��mJ75y��g��+J��(�5��b���a'���0w8��m��b.��7S����U+vDT��~�7H5'-4w���C'!z���%(�r��W����� ��l=uW�_^��[pM}�4 aqS)8P�\�b�XlxVHYEB     400      c0G~4�_#���;%��cz��� 	���L^�
ݠ&�z�u�0F��1%ݔ6��ׄw���M�2H�_�ؘ�j\Ÿ�چi�� g�̴�b��|g-���@��Z�l7]���:yHь|M���Y`Czs�c��J�H~����a�f`@xU��:o9�-v�Y���ln��*�r��*��GXlxVHYEB     400      c0�lIJMM���L����N�V�Y�<����� ӫ��vFa�YY@�1kl�6��s�	�q�!ݑu�oC�n@�c���.�G�'����[7���~�'�~s�(e7��`4�q��:J�)$��X�De�^�J�'!6���B�k9��V��!C��{5f�H�긗̽t���a!C�S�m?��vXlxVHYEB     400      c0�Ico��^�o��seoZ��sJ��Y���]Dz S*c<ȐPA��["�;���MӘ�$�#���=�f�fU�e����b�?"*W�H*q�zV��j�H������~�,����X�f���������t�����`i���q@��V<Ct��HF��=\�]�B�ߔ1~��Y:q��CġXlxVHYEB     400     100�.�2�U�54�c�4��p�]6�D[Z~6��v[yh��.qp���$�c�\���c��62��7�߽�����k�WY�I�U��IT�����b4a@�T1w�d�7�����u ���C�m�B��,ʾ���}r�� [-�ŕ�emZܸW�_��LP��l|H��$�P���C��j�U~��v�M�E)Ju��`��4������	pl��x��c;�d+��?���ˏ�j���$���"��t��XlxVHYEB     400      f0$�o�N>��#�sKCׁG��U�B�11����Yec��y�ua
�2���X.f�Tr������+Z(�o�d鸓�ć*�M��z)����̬�Ě���i�Q�\	&עW�)Tq���w�"�{�rT� mW�
�t��$׊D}���#g��02d�]��X����CS�7u���*��H��"��=`f��޿���5�H�%J�UPֱ��h�M[����\�FIK���<5O`���҂����XlxVHYEB     400      f0�nd�g+�IM8��Xwp���]�%�/v���YX�#��Yoʿ�v�g�%κ��ֳ���x������E	�lFQԥ�@1�f�pt,��^�&B�ftv0-\�!=[L+� ��ll9*�*A�-���T�r�)7ܬ*^�B`N��g�X�D�
����%H^��o��(�z��&/ pD���p6��\��e:�y[|��c:ɩVO����pa�t3�BB�>IVQ����[UXlxVHYEB     400      f0U�3`h>��u�*�a�*�J�n9�x�t�8�u'q��j�?�5���F�7�-��ɥVu$P�q��|+^��{��ܧ�G��bBf����Fs�)�ڧ>#��d53�,��.����Ո�.|�nN�y�
��Q��Q��l�:�υVWFMdȐ���4��NR�9�{kju�Ws.F�N��+�vp�
���ٌ��p#����v��(��gz0>�6�	��&�����g=Cէ�C�KXlxVHYEB     400      f0~���I��D����/��4�� :��Y����`���B >vRoc���n��Y,�t�^	%c]��4�z�ےx�wfDqِ:Y?ƺM��	�0�o���n��t+~�'bc��W�=Zd1�w9e?�4p*T� ���6{���!Oa���i�TR��g�(~����V8D��9��8c{��Zj���
�|����3�����jCѠi�Fh�dy3;����6ԝI]I�27A��=���XlxVHYEB     400      f0���\��N�NL��֒f��?���z5�C�2�c�X��P�Ф��E�\���@���h���b0���j~aO@��)	/m	a��9F̧�:��"�Y�们�[}�`G�X�g��g1�a�0�(x23���i$)�3��T�}m ;q�
�'e�W��|���0�����s����?e?���;aX�K�1���2sâ���a"�ʼG�pؕ\�6��Huf���U
�ژ��{)O�iTSJ�u�XlxVHYEB     400      e0�9�$"�f״����7v�`��)w�my5��Z�d6I����<��OA��m�.`"`%F�ǅ�A�*%F��D1]����9�w�0(��ū3ܘ��D�/��h.	؆�\�b�,���^�gX���q� ���#.`0�{����`�"��*:�);���A�����k���2h�`t���CC�m�u�W6R�o�I?��%�㬣�F�9�d,��:P�7XlxVHYEB     400      f0�ދH:/�O!�S�Ws-�{�AB��nB���k��A�}������U��0��c�d�s�h�>��܇���;����ꖔ�|1�l��H�V#��9"�]���i��5�����(Ld��+p{�E�[�^^}{М�L��ƈy�S.e���a�Ԉ�QjD*����}~�{������^]A�}r�V���Ǧ�N|��w��˕,:�J�`	�蓝�۴�2�-M���_�}qi�0V����5Z�)��#Ɏ�XlxVHYEB     400     150�P�'���! ��s3?��H4���B�,�76q��J*��/��VS�\�qeVB�U~�O+��Y���E���&�nU��}<��+v+��I Y_����5����r��K���q&�G�{)4�\�RGWߓ�,�=8b^��6Ytk�������c�,_KH��Ӯ߶͈б��w���HB��%�>HQU#�^�-�ڟV��i0����H�d=�������)g�͋���V�����b
��9O�\J��u��}��JGOӮQ�f�n���t��>� ��9�I�QJ\�M��ێ F0_��[�����}|�1G�#1LKEXlxVHYEB     400     1a0�׋U/7�n�x��*C)B���|I�8G�J��l8̪3G��p�����ͅ��e�Edd�]/�yo�1d�J�W���������f����.�*-�F����$<�7��.v�Zߜ(v�-���#]��^ǘo~
]p�*�Dk�@)��UƢ8�a����n�����b<LU?D�W�����)& �d�!T��kऑ��d���i�]���5�3�O|1kYO���8
��>;r��S�J[ϯ<	��q�^���y:j=�?�ft�����;���T��7�7_4Eg,_,�1YGTvL`�5����&�2�*W/��}���ώ׮�xkb9��vy/3�@�R� �%��6�rT�~)��S�X	xGRc38g{�Ԙ%A�Gkt��A�z�ޖ@� �`'&�M�B.G�pIE2���)&XlxVHYEB     400     150�R��@�xw��μ`їW8�����s�5m_[�j���jl�j�")��)W,�4�z�7�*�^���h��Ғr�*�/Y���2�~5���@���^�đ�4%k���䡋����t�#8���Γ�s�7��-΋�A���W�[�k3��.H��?�ɖ'߭�>g��bsGP�+|0v���N���5��w��"� �-U�!b�N� �DN������Վ�T ;�6��E+�_����G�i����Բ�����u����Q��Q|�s�-� �����L*��e�񫵭FQ|%Z�=�4d��)�vj��s��C8����R�����g���.�&�XlxVHYEB     227      f0���탔G_=���
�vc$���(����q�s�y��1B��HP����=Ӧ�iA~���.$��r�\�7��ѷ��#qm�ĳ���+��fv���� �y�`�xK��k���f!&�s��Z�t)7���׎�P�ww����4��h��|�}{�=�{�(\k"E�#��@UR%��|\�<1j	M��Ã��;,�l�R�\ʤh^@M3�]�r����@��e��ˡ����