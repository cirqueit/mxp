XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4��D�$�J��
o�26N����˃g���T�l����J�ūt��M}�G�7tO)g�����,N��`u�"��~m�`9��{�~E����jiyq��-MZ�"tE���n��&�He�v{��4�^5�(�b�.S��f �1ON�+J�V�N���䨤�V@����U���?*j��t� 2�|�f���,��Qx�B��:�����W~ZGW޷�JW��w���I�Zp���[�S;��I��n��h�`����qB�͉I������,�e`�۬��:v���Mo���/'Ud�T'~zp7|�,Sۭ�v���T�R�������m �ER����)��]"���٤��#����m�T�{�*�fV�u�A��Wl�F]��`*J,e��aKD�ͧZ�ń?�or�|��~�=@�$��t�o���q'||6F�7�"���S��I���V!=����p�w}9����A�3�վ6�gܯ�[�⻹|���{���-w�]J�*�}4��/����)/�>��$�_�}�b{(��7������F�ta>}���J|lEcs�Rj~/�!�!�/���n��! �x�Uh�\�MT,y�Y�,����6��_�dh$|o���XA��]��z��^p���}��y�h�lY޸�B��A����7
P�~Qޚ���|0`���CZ�"��@8\��W�a ��2�"㥗�Oq�q�ɱBe��<J;��Hе�~I`b�cc�e�w�yj�;�@�|r�!0�XlxVHYEB     400     190z���b87�|] ���ޫ�������4��,c&7�X� |����c�/��Q��	���A����h?aТxs�ٙ���u%Q��㠜d�CH��.ɍ����<�
j�v
�p�|ӕP��9:�����:�#pР�7u�jODJP�]}ryڅ���x�.�8$tv$�F�.��E�M�_�0/�-?A%|_K����U5Vr�ܳ�}ywa��j9e֢2!z��~�����o���^��t��#�69�P�hp��u��;�\. k"��P��#��|:n���a���������>�"_��V��͈f�t�h�O�|H��2�d���sq��t���̺N�;�����@m�6�u�#�r3�M���|��SKL��c��$���ʻ�8�PXlxVHYEB     400     1a0p�e����*6�E�]�9��&�F�DW��s��[��D25��fS��-��:�� пR�ExTܗj��h�	ƬJ'b�T̉��L��Dmʫs.�7c.���y��'(S�wR� ���-����C$؂��R��X��w��*3��aO4�/l�=�h���.\@����ZͶT���yG��гx�y���8f��M�\	����(�ݬ��nfs��7�v_�\�h�󋴩�j6
{X��?����S�Cdȇ�8��\���S`6K
X�#\�����kC��Fϰ�瀗��D�'�y�@vV ��0��ӌ.	��c�ؿ�ɍ��%ܑ�o�nt)R����{Xīܼ�u��_�	v�����{K��Ϳ@���P��4�V~�8ѿ�NA<����X~&��:d���XlxVHYEB     400     130u�"7q�H~�2s�g^�F���/5��1���d�N_�#'��{o�H���,�d,:�I-�G*��������Aq�jw��roNU�˜	[sP-���,�8�s=�20ݙfV���`i� ��b� y=�2��:�<��l$�O4�N���Hz�u���"߁-caZ��c2d�#>�@ F32�&����>t��r$��p�ę���0�|Grk��5�V�MsB��X�K&���6�mz��ҥasr���0�[v~������|ץ����-�@S6��  ��߹U�߮7dz�7�e�GF��V^�D�XlxVHYEB     400     160��\�<� f!94�$�c�;�v�yp��Ǵ�(��ķHy)%;-����8��F񈁛���ZE�$�,v��q��,�����:���މ��P��xT���ʲ����8��=ې[I��-�ށ�s��>���Kwt?�2�v�/�LJL�,���B�6~_B��b�I��Qf�4�o�j����x!����1�,����nw^���f�8i@uϬk���,������%��X��uԫ�T��c%�1� ��h���d�Ut�	�'�,��no�?���%�0!�P��M�����u<�;���Fo�ʥ|<d�Q�|s����z�N�;�)i\��s�'�bXlxVHYEB      3a      40Y�N�
��������k���[M3Ns�Y�&l$����mg��~>1�wK��NU��	�����f