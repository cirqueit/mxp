`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7104)
`protect data_block
zDnro7Wf7ipZMMZrEkbvfv6qhqUmBaa+iqWkK05vQU7QFYYTEVECke/cUqGSF+zqVAH0Dq4XsXfx
2XuvyYHGiZX3RDU2csj8X/h3HDDkMLt3gk+jJAKzYfU2r17d+N8OQINhOyOcwC8/yuo1lMKzlB1R
sekiqml3FuaERHZc3acipKovvQcVRKQ/AWxAldrgG8ZkfmQJZnWqA/wMOwNEP2bkF1GcC0chOtRa
xs5uhCxvQvpVarIZoO6GmkeMdYtL+Nz8ofCRXeaRQ7lNZ7zPcJzyzzzDqqeUWYH3aORmMvcWmVt0
D4FHcbN+kdcE2oK1EiCXmQhpW1SLLg2gQKUHhlzqRQ9kEzrQ1b7TbhXmQAjjzvqHq8WQ1pKEMwaO
jD3UUDvbq2V2ApCScwMJsaDRxtaBz3ElKEF3KMN671GkMKvmayzrwWaO+t67PkO4IWUkMrIJfHMW
HVp5c0k/50ot4yRcTGD8Mky1b9W44gm2MU3VA+r2h2y8jNUp2F38KOTO+0fI57pXJBEb/tPvOtgA
ms3YBj3q/mO+uDOk5FR0iTlM1ZqC9tMWFWAABwXQoGaLO8r1pEcQ875hzdXCjdlrn1MaoTtzDUWH
t1MLc6pho2ZR/5G4GS6cS/XnSjsqEvoY60AX//8uhZWQO56Qv86MzVWuHS66+hq9ZiglFBkUn4d+
lo/arSU8SH7XdX0eyS2sesvh+mzCqEfHKZbE2GYIRuNpBf9jzUavOIjYN0A5TLIlrv/vTkUkzxGX
W9F5QVd7LdxtP8QZ2xtJoem5mq4MSnFico2Y5KSfjyZdZB9/jjianK6zA3Y5329g/iObf+VO8Psl
jOWA8MbTtkVnd2BtxCI8CDscXpDYeT83C9JceRjeOGZaXVQ3B8vSTnG6x/L29Z6bjNZ8Nr8lUbo/
7IpWnA47PDFovS8G6LqhIHJ8vsWuIlgvGR5aoXpkOUJZHWy93cXbypoYYBTt4oj0LRsqYCkL9QdL
KwssRz5EczJduKyU7QYnK/C64fYsKDpr1DP5p/6b9/7wqzhFCgFpqWFGh79zsEz8/4nk1K1//XMk
pZ0/R1TOGkrqfYxUqCejudwDHqRyTasV/TuP4adv4eNtMBOC4f5YVBb0GpbYJoaq50FZhvFPYfMG
sNEddFiiEMqFosRDV82VDhX/yF9Ahmxk75y1un6bJhEGg/8RHbASaghdfZ5rf8ATlyUYvCHWuihN
Im5ZqR7tblVp4XYUis/Gta9gHxSCkPCx3DbOVaFmSc43bH27YEUr1saqp0sI3WCwidrxlM+Yljo2
itIhwtd7M23FnIxSrSOejhbxAYbQiE526RJlxLbXrM4fOI3jjxZBlKsVdPGSMEXadPTiRyDWamPg
E1F6seuPzCtTye9NSWjIatQVyc6waUHKnJjMmu2lOxpB/vm4vKpXC8bmC2gxbeDMUTu8AoveRCJU
iLW+R/aq0BfN6f4UsXwl8YmnDbxTm1goRB315hcDwoHXt4Bm8g/j6k5uiXSFsojpYcTV6PFD0rsM
ye3AhPO1/JtfqUM3NC4tKBzJtBAYAQiP+j33XC3kltYMX0SWuhfw0cdJtH3FcRlIz05HEgKoIlRI
9V6ujNjJOK7WWAGlzrAusqoH7STWSQE4sBbxPyioxt+0VZZS7d/ENeebCAdavhmisLa1ME5Hfirf
lt6rvkfkQRqfwbK/NND/uQ3WJS1ABWFyJ4QXUUMxLa0QcoUfPOf2Ed5Ggvbq0iE2fVe5dLcfPDVb
cutowj2eZ1dhJ5Cfw4Z1SPT8S3rLWinGG3KqHngV/bZ/rUQ78uKJznpUDLj0XepKxb0p/KP7DjqW
QLzx2h8J0+iqTj9PXiOFOUi/ApUgwsd14Hzt2hX56KCkCbfzRalhcUP7oKaMFHOwJSjUqjD5GSkK
liDGPCjKsmZ1fLP4JU5ZtITKLzrEAC0PHuiH1vd3Q7azVocl2+V3eBNrhewdWYEfExDwcJnI62N/
RjSMHvAEqBp1nZh8XQVqIN57DirUqe7GxP4C/ySCqliOXvzSZxEiPQ912d0BIbztlSwp6WpBMux6
YniG7cysg7g9+TlsbVU+WO3wTnOLhmEjtERnOtKmmSGsfN+IK2Pqe0G29wp213MYgnO2JxgikTNs
8YKzYf/LtVCETQiUvvmRk5IRLeRsHFpJVCZOOvxLksSuhWVaqxyLelur39ADM45IlumN0MTCDf5u
JTWFaGtnVma7F6xoHkNNn3eWzt1Y752A6w7YbxareFPzh53hXTH2pL6ETYtWwTcQ5QyoMOebEdl0
XlG3NLiOsLeDuBf+pFNEj2bMzntMO+KnkFwWjePeL3y/K89dRgljFmnEFHcV0vh79vAF62JPsiOG
HoUObJ4xeI++lIsdCCFey1uR/HvyBWXKYQ3UmqB4xJbKz+W6wOFocCr6xGzvwwed4vUrjSOnQEVD
5OEkUbg1M9JkIOZ6rnztfsGp3hwRvZLmWif41F/ajrafPsCYVHs4yzsQZbYsrdEjX3344kL+exTB
w3teCFM5sOYZEuLgsqBqfBCJIk3U1/2RlU/Ek+Aqy/MMeE9+uBaJh/0Sc/aFxvaIvg0i7B/T9R3O
QluEmwDUYbFeo0ZOHxX7Rjl9/9zSwsz5Zr/GGRhDmlcoVDEkKxj6sZj9efeOMLWIgE+RPHp+qmzb
hc59DVXVjW4RBntVZRkg3WRQUVif+lZgcmJ6oKij5ipnzLCDTXQMJiLq1ix2fMXnUjMh7mVksN8n
8hH06YIpZ0eSOxC5KzSgNC4gkjLpTCNjfGQ3hlHJDN8dXlsMshtZTHi64rpqOe0LrLXMQD9Ty+ac
pNjOzBkZI6CT1EJXzVVHsLTTuhWdz32+FzZJdvdH5OdWwjohEX/snT7fcnfYyfDOKfLUe11/zAON
pXiYxEe9oG32uIyQmL3DlXDLeAUmrClOHx2taRDm6DkXpn6JzWGpua0h9ncPKQ+OEl4A9YouX7XG
iLVlXC1KCjKbOzq/3Jej/srJi/t7y0IxfDOebMPiPBwoznicQzTgEFUkbOu2bzbFVj/HS8oDAOsv
NMEQg7Mda1rfDyCFLVHwwEDalmwLC1SGKtYLCG96COUXsnlV3nfIc3uNwvktRJbkVBm9Otp2c+mR
VvKMdWuBaIR8uqKc39RvL71tRvT6kJ6P93X+b23bHHSb4GSkkMUkCyk7xBsqcOT6nkSzXQG8QUbt
PI5gMHzmQQTOqga/+8IWFqxRIvIaFVukzgSIrDwSKGY2N9vK4jMxxicN6kRpVqGVM+YZXl4cApe0
gyuqouXbyXrzcaPI7F+YV2kb5sL+eFXOSrkDq/fpaiG4djm8IX7Mr4qZgK16UMfLNPYmUICNuzg6
6drDo3PDzdBzIrciXSrxN/ovQvkRSxChwNV92g76JF1Buj8orpuh9Qt7VM654ar5pX8GtTTqpTGt
x+gg45/QrTN1lVhwpCkUSzx/whEGyx689YHfFje5tM5yaFLqcN1U4DMPWrUked4+O3r33PURyprs
yN16KOYCqLEPGSbc77HO0sL21Zu9Ed9A8AWAH/tA3Fs4jp7DK/9OLxWpeKjq5xqN6Gvw3tBcvJnn
wC3j2W7QbzR6VsxItEDezql4n9frpmYc5eHozlwsDi4AdbAAIQIeVjLdIY4dp2mUF+J3BZ/zNikt
ao3+hqPPNC6POSjjuiQ1pBvqL4bkEQWziB8DVZuXxFdJBg1x7SyeSQ3E5C3QNLHAXz/QLIRAFCdu
qPER4jGa8uHx6dD8HLJjxq2hU68nkNRZa+2KJZfnsZt372qn3OwK9PWhMv0D18TjU/5bgidfiSnp
8sVJD+mWpG5rNTlf+PEn64HqrooLrBZMXyIWqBmoqMkdMKUxDKe2DyVhzhmhKbRRQRUHuzbHCwxG
rCjdOoptyWMTDwubsL7rr++/tejmIV248Ap5D4D6SkwEekt0IdJWP7A2sDQNu8wGRG5RzbnmE8FS
AUBmK4ztVhKvs3Fgeh3U+0l39X48XvY60ps8qPzQ5zSPNEVYJ4uLbP0tlidi39EfTd2/7i11nBjM
vIpXzwT91LCO6O1Gs+uI5gbMwmRXSw8ZGWpW7sS2Gj5oxo5+ctXsRVlOAVuoIYo3Cme0nJ0gk5pO
IXbIn8u3HlPitVTArQzDNwE9K/DSBVCidQs0vV0pA2JWu9xLrmOEc34XCs6wl/Sj4IhYT7TPUONx
5j/VB0C1aV/koRlQEzQDWvNds5RAnobVVOv8pw8Q4fMrqx9ENQ54vsbjGmSpkh0UR1rBlwdt5Ltk
0MXv7A/Dc21ZB7V2aezIHFjnbQWAXBmloC+nah1TXuQ1AT20s2/W3PuI890yWc9q1TVtpr0+xAAq
hII1HZF7mOoE8d5dr77Loznp8KY0BOmPHuo8m2fiVG8OsRZB/+UwWk0c+L7NrnvUl3G+DYN7q8e9
vr06MpFWzK0mo+ooH2El9GvdWooLwK74LYUqwJRxGayDixNDh3nhh7pU7Ckyi0Bgzqa/jNgwmJtJ
WxXwJHRHNC2eGjtT7yLfe949V45l+O3MhJC3ZDgelfwVeBTubSkh8jog3qMcsd4ytvH5Yop0mNhp
LB36o518aR3yuFiITXxmK1K++5jAJyULgTkmQ8x2p1BVW7Ag8Fgc9Lns0IURimtK0Ua9rW/aGl3Q
OjVjdzU36NPNLe5G76zESI5ydE6lhZngRjjcGoNHejr+yrAwH4BDSJrZpP3Abe2dHmOojog9TvCE
luW3dUemu/vOw7FZd01tFy0QT+tI6dxNnQ56zCgafpD0RGP8RcUmjEG2PMgwedR5vTehdVjM/Exl
r+0TFXysVtm29CmfVJFoROM8UV2RKUkY1zWHZZT9V+quMnCzaeqHE5ns9riLi2W/s+iVKjzBqVUG
bVAnMnlFcSHYz8XLh2FJI+q69WxwS16JWhRpq53dkH7SHgm6hztIec3irt9HkY4p854WGM8KU84d
lMU4aVNHRoXQhfDOzTxq0j1axW53thUF0tgRvkEY0chq3M6Bbfgdp7uuyqxFebVJATxuyEKhV2iL
n3r5CIfa0WHo1KGvsNgrfauLvSgCgC7fyarAUlCb4bSNP2BtcOEo+6dAcYAHxPLsgFJ1b/W1oZow
XAGUJ1FbzrzytZ4bCYf/tv5T2PsIvxJpMbk191/mdqhCIUPFX7LxsfoFfLLJVE1VNrb6/XCzFVPO
I6Kv8ahbGGKfgkV9SsJyxageA022Wnh94b2qe64tauqejYruSYeXc4ACzdvRymPfOjI6pkepIwUu
WbTeK4YJTwmFGdQkIHnqnI8TJLVXnKYYtqwFG2myG3tm58wjeaz2n2e/+3t1TztvuNllJX0zmNdC
VmgSzSgBwOZqosiegXwUrDjIldeMAfMAqGCEGlh+iAK1QEIVWjvc4Ebfndo57yy/qI02m9BYNe1D
NTHpWwtZeRzCda26J6p8Haql7WxHrUiXfTJYmSVwDLPIIkKrdHCDtbN5oIIHd9hovT6uTj9tBXXH
f9yYJbynilQCbxyv2z3KdUcHLZvAHmDjKwbrRFd6XJfLQIwqWCLNeH80r+wFkix2vSvUN2cC2TXs
95xK1iBhA50XMiO0iucAsqyEWiQ3KV1FYGEI64fpYBTgRIwbtw/kZo3MMz4xOIKWtgAAwlNlUm67
bNLlSPc6yUkOcRiglhdfVVoLoogMErdTsgDYTsVLiJsK0o0yC66FYoJSrrspiaKug9mOxnyGjcq3
U03R1v+f1zkRO9ksM9oCVdVgPaSR20iZgYGCNHMnS7aYRMj8rxIsMJ40W4BsegMxUh19ABGclMFF
Qqu3VvYVZOfoqesVIElh7URD9yLC5Tj2h1zlgvw6XO2zlaVeXNFvb1reE09mt/QIWXXeP28Jk6TT
5NzbJvoSLzy96unoz1T5h7pq6P7WprX24EHbUgI6pkipEsE+82i19yfEKNHlIDWCB1h2fXhS+ppk
Q1YPPrBHlplYvFaxb/O0r6f5Mqfv7w/tkPQgwmwbghcVIk3Zs3ooXsZhCDGMs4Ri+eBt92jcSljm
+mXArdrthUzGAzcFAHSYMw2vw4h2jvOcmYZNHNXyIhOsX1nAoyK0P06i32un6BSXTMll/GKEqLOG
rvmfJgUNm+94CXNQAjSe/OfEPbNAhBioXgzArs8gtSOg/UJ5v2v8vAolRqc48CHqh1VCxDhpi/Oj
NGhSqQkfqmhmlPdXEifaRfRq0LnGu2Gk07fpYsbzXoi6P2jlILDcjgEEhSYR1mkzpYWv8GqIbOFi
9A3JtSuJlzAYAn/YhTvOTqM3oDf+o1Bwxu2n8Q1rUq0X2Xg9425FfV3GeUG8Kr/miGqiuhErmwAD
zi3OFHL03Te8HuX39xaArQY4fIYxzkQzxz21t34gkxMsousgfDkMRP8aaw6p08XjIjnYEHFrrD+9
A50BjaKWgp9ahSGQD4cz6iZHifSxlbsjrXjGsqu9hYN+IQMbV6YV8Uag9jfR2niERLIbElvX1Iv/
NS+/4tb/7W4IGjFMf1mPjyedkt7VMpItAhcDYKnZddHzdhRbm5FqYll7GzONpd5hUpp0MdFtJjZ4
IljS1eshUMvVr/dJEPQZNJtxf495HyVSBnX8bznCs4pPdSRIZxqxxTp+GqLPyrwXILxU1AiHDaL/
PVioVvf38RNbGeWd9myujQ7zpUo4HTFPN+yTbfTnw6PuQA5BpSBhwIFw41wpBOUo6lUw6kq4HJWI
TMkq0HJ0r94xXyZAX8kHzKc0PMf+MnbrSg5P5E3BXS0oFyj0sRLzbiGO3pBMhaBEjRmyNTeCdmc1
MKu+gk/+zPuC+Y0K8W2hvVHVNloqeVwQAxYJ5qghCkzierykS075Uvgus6HoT17rpPb9IvmHZ1JX
iNaZU/hQXYphmeRDpNGKXxAEPJ7Mj4onXhGoR2FN1tSNeNfB8fQ9wVg7bPvQ3YtVJUabHtLI5pmJ
HjXBONN1KJ7rMmQhqLH3ti+WdIHO2UeHmSD1IdqA7xdWZxQkG8c5k6tNNFsFe5TDrd0QSDvMW+QD
dhID0w6aDXUwjDAtiKlRKpAy2NH/33nx5FoH9866CunJZsfoOgRaUtSvLMkqgxpMgfEGYOtx+1sN
4kzVlgmge9c3eRFD3/bqVK8Wp6hg5c3HAKz8gUqWLfAO8i86cikfJHG+gyMC/xTKXkQG6/dJZfoM
4UKj+JhThiRaw0XZKi+AWlzAYB/J1DBRKEhXSq8Y4Fo+LYx75A+R2vV63UYSihkfzqa1MlwhB9Bn
EuX4JhHn9VsTcsUiLlNLI0TceE6fxWwDGbZMmBPAjWiOBmJSk/U7Pe1cWJdAmAANXgQYZVP3lpNi
8AOy+YAp8r3V+7JJkpwKglzL9hiBUNX3a0FVmKqGjiXr0GFAUCqIFcXK85kqv7oJaH7gEdL6x7g3
Bo+chIQ4ZkYQDmknMwFdPAbhh2EXWKBa1eYM8ag4IbvImmzWx7Yw8tgyQyj2qWUrL/TOZhHRfu3S
i+7nBtt8qsKxwAdHOuySI7JePQLm+RTRH2NsShkEykNSN/N34QtsghsoakEa4W4SFFN5VoQ7/hEl
azAfzKUDdMn+jsKy42sjlJJwqqFfTSd3nKPiVjbVIzfnnUstruRseemjyw1gIVLmS5JWH3M9bPpf
bTt6GRUH6WErfLug6BFwJ7SIL4tlNgq4tGadqhjcEMH9DVp7xrYQyk1ZW/HSZggIyjcQoSIg7dbX
edHhzgEH38eRf/5Ys5EE7Kpw466XQ2W7vuF90zMuSunA2iV4RXR8RPxTXTrUYYfU48ch9lb0qOd1
1vX+Yc6qFQpyfjRgtNcuvqf2WA7rtg67bAuuiun1QlfZUwjBSzPjOT3QB5t8kT0U/QR/EIQOrsQy
UfEgPMzmPHrrWl38OP5Xfpgk//t3mgZuJ0YWBYENZnd4JAhNhu1E7DXfWSauMeUmJdj2xaJcpTnu
YSjcMj+IekhN1xLM02Vzw4seP47Q9jYr/NiPhCH4fmqkQb06UarRh+Gsu2JFPJmztUFcEv0nc616
nS7LmY8sjQ1p10ffglvIp8PZmOBEALmsLjw7mHpd6QDXoaMV7cIgZxUxj1An1rGsaSvjeKbrECNI
Fsli3ybrGJ2yb9mW/ZAJF66HR82VNQ8bMkBjM2VfY1NHpH0H5HqJMNHwQhsLTG/iIl+FIF2ro043
eEq2ZxulxlUeM1x7PMA0m8VYs9HAr8ZHDXt7xhcebTuRMVWWRyo4ObU+T+gHp545xrWXZfAICaDw
2OHA4dTt0QYuoZZOtc1rt6n9chvdbltCi5okHkRHjXfrapaAlgaJpnh3r+WHTr2eUs1xYynUomkf
+H2wLbhsQ2JLJBRwMg8KsSCcoz93Ns7Tt3AadPtpWMeMQ/5/86JPTWJVq4nObwEkf5pq1VCLgyCA
ba/FbygpKHerZwHQyB2FvFhYspVP1SIDK4jA62XerWAIgV933Z7ilhDO9gw9d8+YaB96n5jmRcPQ
TFjzK5qAV7h5ZFlsGuMrYFGYrilNFgEHRBIjt+geqcwLb9d8BfL7PeQbEsBYcWd0J4NZcXXUfB2A
t/hlBLHX9ZOFNOsTe5uSjpCMdIMQKLU17uvToTboIg1VrayhY7HcttaN6tpv/gXSpSzQ9DSUojus
yf/TN/XGXmuJ6J8nUKEOZghadabd1cG0IEP/R6PjJWYKl32jPsR5vUPbjxaqfgMlzwAPolCBcc0+
YH2/DXq2EHXDJBn/JuZ8J7PiHQWOs9/E8A1vEmVP8wfHLC9XNd/7PsdRTucCzpblktkix6TWaY4r
EOvHwO5NFRSxukXxycIxQnl9GOz/prNi7Kg6tWkKlQpVuB8j25KR3C7ADvDF7GgBAVH2zJkJ6JGj
fFYsUrL5iV2+glBrr6OSGRGxWZXgIXRPCuoTe/4EvT3QfmlPlwgLXykS4Wl3NEtENIwYpoard8ie
Lo3QhJdd9BBiSsTDLvNLIN/Y++0KReWKnryIjcQ0GOZn3rLbX3bxnzPpoz6MikZ9hPtipc/95LZe
2p49AKI9eIvCVp8NINOSehUI643Eiz0ECPBKkRf48yBUzPO0GtQ2dOClXb9gCyslRgygdcds7TMo
kSnfcG9TeEcHvk/gS+0FCsb/o/qDerEV/RxcpnQcJcrnZIDVFj0xbnmypq7R7IpVY0/IkiTIqfQI
fFdjKVBArd0W/7MQUnUjlKQOo3xGM77/n8b5Tqt9K9gkSUWWpWmkz2D10dcQTINEs0OGn+ZcdkX3
z0Hj/Tpu9SjrK27ojnFKWANAJkGg0WADEVe/9ofYtv460jxSWbXJGvnD0jVF/StgNQAzuENaA8o5
RQnGxWpr5LaNnv86X4s9+487M25UCkxh76haLaZq5NOV/ne3i5U00ixS8lvsznF8+Nh5NWXldV2o
INXwivRh9WtdWZlY+XJNzA1KgmHPf1+v5AvS/2n6zmMSB78IN5iS1vp2Fh/HR3FzGHrz22LQmIwG
97DRWTVHfnJqY8i+FZkDuG0Pc1lsedr4SdGSSA+K4+0KIbpT
`protect end_protected
