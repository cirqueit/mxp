��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����¦`���B�B��l�v��o|O�6nXWM4u�.ƶU<x�D1B�B�Ȝ���80�[a�T�����#���I��n�˘��/-��zۈ�<������R��`�?aG����D�\�h�G>�`5:��A�����ݷl`�ڕ���d�s_#�/:lTo��E�J�]]��7�v��a��_��ghq?�Dh�ɖz�6�厲�YG�|�?�F��<��Y�vP5q���(������w�I�U�Z�i�n��K��_2ڔ}�9=Iݚ��!��o�im��%���u%ٓl,�$�jQ���tPJ?�p������	�q+�i��f��������W��B*zE.ՏՁ�O"�:�3�50�C��T��N�x!^�9i�x��?��$bv�b�෧�AY�@tV������!���J�h��4F��ja�@�Jb���y�eM�h�}1�W8V��&��
(�h�U��F8>����`&�`�$�͞�0�<��l�aF)㑀i��sOT�is&>��:؈{�"f<G�i�渾'��Y>$�K�Ow�����ɂ�$Դ�m�����F#l�C��,=tx�l��J;��o��I���۶���)q[�!R��qǰ[6�&�y������
�5��Q������1�9]�T>����O1�k��弓Kt��r\�o �*��T�5�� l��c+y���f��Fw`ǭ4���Y�!w�jU�����c	
2��*`�@ޡ�L&�a���Q�L��A����E��gӈ�P�I��, E��A0V����2��\�Q�s$S���M�����vxaj�W���#٣%%���M׽i�PN�ⴡ�#�t���m�4љ��-��SW|�?�ʔ5�yc��*8!�h^�U
Y�bQ�r� 6��p��Xa!�҅��⼉ڮ=m�h`�S�;9:�X����wr$�DE�����
pP?߃}l�#n{,���j3ӫ����x�&�m���g��+� ��D�i!�&+�Jy��rE�'�c���̹~�v�\���S$c�(U���2$'��3��=�}����k��� �U��=2���&��)
?��&�/�5�x�|�~`������ �cO=e^�hd�]Ch��#
��?����Dt`���}� �{��OEZ����Օ��뺙��K[�������q����$�}~b+�g���.����Lk.���@ +G�����`"�]7=		ȗ7{�ॱ%n��X4��gٔQ���r=1��#w�:���>5iY+?md���EN���|��}�ƶ/���.�,�Y����Neҡ��!_��N��z��Q]��� b�<6����%�+�����1��wS�!���r3
���Y���f�zv���yVuO�Uo�V<�R�s�@��?���3��9�A��l�fm�0?rkI ��؏Q*,�����r=c�7� 6	ժR�i������`��\�C�[|Y����>�x�+,ӿ�G+�/猪,����Z�9V�U7m9U��q)QFN��Y��LzZ�W���S�W����IKcY3)�A�a��!k�ĉEu=D�-�N���^�����62Oizؒ�My���Xm!�lX��X9X�(dE���v���31X�p��PV�r�	��WM?�֖߉���ȗ�}_oby!�P!��F�&|� 0�N`p�F���7�o��I�!�̡䵆i�ޘ(�I6��S�&����k���ĭ5��r
,��e����[/���U�����	���" �ݷ�N��<w��eE��ܱ=�T�dю�V��*��q�?�< R͂���T#
�#J1Ѕ�B��6#�?[|����.��v��t�(�2�N��T�!�P�p������V�z� ܼ�h�����}�|RK�aTMn���P= liRR��d�s�n�y�y<�z؈�^	�1���ɾ�|�<?p�1f�(��y@L4h7a�xKK�1�]�~11�i�l���z�ȵ2_��l����lm�r��K�%�z�S�%�i� ��M��x����0U��\��ȣ�|)/�;��4!]�F����W�A�������c��$[�R������`$1"S����ub��#�e�w��b-n���h�Wؕ0�O���}d�^X^��6�'2f}J)����!ޢ�BUL�D�QJ�O�ⲏ�R��5rB��mG�����`K�"� /sYF�"����6�q�����L�MS)6R��p�$nO�{�����4DLY��XLkv��0��*:�{ �+���	,�Ġ�v�:������u�����u��CnR<����=b����t��ꥴY�=�uk�g��-)���f���*q�N�-8STE���o��F��V�C�+40MM�th�s��$�p��y�]i�L�7�`=��\������ؚ ���X]�04���t`�%P�TP�JBβJFB���m�O�]��oo�e

����Lr���+�jb�W.�<}㙁?�}")�쥢�1y��Hn(SU���H�'�����b���� ��A�ć�5RG@1[Јϼ���qV!�}Mg(��\��_	~ª��W�H��i� �
�z�z��e�����?�BIؤ>�*9)�Y'κ�"��^�b�i@��*ŷS\�����f�K�(N���_���H�5��P���Y��<�7������t�֯Vĥ/��ݤ�W�`�0���G�f���Z�Q�Y趱�<*�w���K7V�}f�Ϻ�H"��b
g!ui��wX�ZNZ$W�VE	Yy���h�˝8	�t*��!���U��ƺg���6բ��V��[
A)��,�a4�Y�!��w|� `y�k��FTrw5�4��S)-T�.��jC�������YAZCt�Y:��62,VV<P���� K,��F*hN����*v	�J��a�1���E�|'��6�V���������E�0M�\�R�����Nc`�;�CC����ͯ��?�A�y��_p2<�� ���F���.t���4���qv�O >��K�h�H+��͛����v�C� sn4RC�r��U�T�vF9$RY8jү����b�)0?R?'����n����%أ�ܘ7c�c)���F�ﴯ�����@s��<%𛎇��Eqt�А�!Q�X�G[�jk��(�Xe��J�x�Q������LeB��Zpk�Z�3�)\?�[{jc�NHg���u��1���<WkcF�3p�mb�O@���3�j��-7��I�0j��2�-�5�,���'��U�j�d�(9)��y������}EQ��5hY����,�1ٻ:����!x�_��U��ÜI��u[X�l.���{�$,H]�n"����2�|5z�MÒ��ƻػ5�)٣Y���W�R��Yi�Ϳ}���a�oZWq�J���F������OR Q�|�)ұ?�.��)��lNbX���)'@?@n1�|i
�<C6�0���\�5�S�.��C��������i��l���HoL��'a�~Y��D����Hb���U.a����[X��XĿz1���P��@B	�}Q�
!�ͽ�����]T���ͦ���ۀ����c�/b��(q�)������9�z�#�Ymi��D�Jj�յ�"BM�������[iʐ����(���Jz���y$�S�0X&�sL������,���J#4�;�m���Ǵ(��a%�����:"03����@dIN㜁����f�@pwep�ᨎ��#�F���~���c+[/I���8}%A۽\�v2�'�Oم�LT?�1�Ns)RC���iLmr`A%�PH��N�")!� ���\�[�-"Y��U|�T��{&ԭ��J.�I�X�?X�+��V7_�:�j+��T�V(�E�(��6w���/3zkp��.%'R둍�bJ��4/���8��z_q����qB������q ��[��$����	Շ.3\e��a���Ł�;�P6qbԩ�tt�]��^��kB[PY��g{�p�n�I�l�a��t&<�:#�X��v(�
�?<hJNC�O#!���ǡھė4�5����͔D��S��'S߻��u��)�,f�u�6�3�N�vo�e[&#�����o^ޣ;EӾ��Mi���c�ۤ��d�p�7ރ*�h`��>��MrZ�>��X�;�C&A�e�f�I�� �3/�	Y���_o��+�=��u������ݚ��{{,i����[�\�HuY!D� �|+rL���+Ա̶B��s�i����o��d�Rj�n8����8���[]��ㅘkya*\�Ϳ�+T+�ְ:x���!���)'S?LI���z"Δ���p*����cݥ%80��e`H���M����N`L��劼���z�k�xe���V�_�n�"��t�w<X>����ֺkx��ɴ�r'��2�R3@69��|ѳ��p���8�&��V��V��!��x�SF^�r"�Y� ,��ᵤJc��9�_�{��T*�d���)I�# ��Iȇy���0Q�������,c� �i��{�L)��0���sv*:�a �`����5�'n�	?�fa2�r��hQ�ji��+�*�Q��]%����+�.����a�߄��a~��O�?�ӵ�&8�۠�ʑXv,0&�.�����r�t��n���[�b6��}���b���m.¢��	߬�i�O�Q�����m7n�;���*'�	�2�m<�=c�!�i8�hv��?�<w�G ��A���B,������E"2�#jI�	�>9���༭��B~}G,�����7�p�,�9{EIa��;�͖'��v>N���0��?�1	(:"Q�uA��Q�̦�,=�a��W���޺�o+B>�sQ��'D����0ls��D��E�Ȧ�	�D��?�-��A\��Uojg~=����}߻��Aq3���m�^����)]B3���O�QS�@Ծ�]�*6w?A�w��ǡ ����iׄ���j���{���~��td�H������
#FU�K����D�7�}^Ҩ�~�cc[�����B%-k�ȅ+[l#��^�5��VP/� �������-6b�`����V��{���E�2���л��_^B @���`g�����t7���n�O�3۽v�Y��Cո��7�G��5@c���s�Q�t;��,;@���E�Z5E
�'7#)X�`�$g�9�}e�2a9#���1ޘ_�`��ǯ�LrO��*¿�Y6��Au�3���J�6��&�!���	�Y�&SX�XIn���VҔ߆��AMְ>S�
c(O~&C�zG����"2IZ��E
�-��;tg�Q2���М�s���9Ch���c�X�si
�iʐ�foC�
�݀�6 ���b�>�����uU��j|KB�˪4١�A�q)��f�n�DMyȶ�#/w���}���18.���Bi�wAܠe,���~3h/�eA�*W]v��>JTޖ�k�+g�
�A�h
��fA$c�r7u� u�"�B_��HӬ"3z��AL��R)J�Qp��n�ߐ��6���Нo�~�.C�n���Ώ��]L�v��[C�!l
7�<JHg���KUS��[dw�>��A�A������z�3�G,6�?�Y��R%���Y�+!`�#�pzɯz�D<�\O�1�^u�Xd|A�Hx%�UUsj��yڃ�t:+��~�&��W�`�i-wYd��'�mB�Iü�+k��;K��}�㦒f��
%]����PWp~	�;�|�8}�K�Y�-��f�:P�[��qUS����L�V�;g�[�=��^���<�	\f%]J���w�(�4Z�;Ak�p�>��?��m��b�>�-��%^,#1p9�
� v;fe�p�/y>*��a>�z	Z��l Г�dm}��ʫ�M{�>���	��f� �.<���Ʈ����(�tn��ay"�ڬ:èX,hA�����$�R眃EC�0P�Pģ�z����JmΉ���t"��<�q�si�3��0@�(�u���)5ө�5����ٖ�g�s�F_;��o
�&)��H(מb��#5l~vB�:��J�#�E	�[1�R�Ӹ�t��]k7��e��FLġ�'7��U��=u����P4��J˯�&��J��ο���r=)s�\�b�cD��*�E�X�Xx�4�A�&�R�Zh����s���zꕮ��(�*��HU�\��;�'L�0� BY���7����|��]�[gٹ�'(>v�����f�) x��֒�$ g��Ԝ�o^�g��S��q��C�QDV{g�����*�@˒͗<�|�46�j.yw��i�ep�e��,`����Hi﹢>�B>�ЪR7�v*�'�"ņ"�TtX�������Iv��HI:�6-�?ݛ�Zy�L#=?,Ӹ�y���w�Z�
�14+X\}�3�<�yV0F�S�.�8O�U���(r� ��I�Zn�:� �����C6����Ԇ3ޗv`��mA��犌�,��E����=��urN�a�R�*v�n(5��&3�8���f����5�6\���D��ư"cD:�
����ˁ)�P�k[��oBW�V�R��(��6ײC�Q1-�Les>�c�4����|�߻�=%#�9��3�Q�*����l����R]ىP
��XW7���&(���ɭ�{�@?K�#��M[�@AO�1����a|�qV��z��������Z�YA�Ŋ���JW�-�3��k�gg)�(8���ː？R��1R�1�V�b&��tI<
��f4��u`�g��'|
IP�y�]+ H0���e9G������=F�K>Ы�O��vo�c��7�5����@Ό�ohd�O���Z���I�����'
�kqT���S�X�@�oD����c;*��@�D姩fl"�Z�ؾ�/� �vT�݀S��2���^�Hp��`�Oy�'�KEUC�,�F��Eݯ)\�P��Q'kTXE,Ao��?r�񭏒�/�-�v�	�A;��NQnI�F�SZe/�J�d��Ŀ���U0�7����Q.1��۽^�U�("�m}5�lϞx��71���W���k���,�#O7�aK[�N����V^m�z2�1׌�P��f���qK�1��ӂ����d��!�{:���7�$�M��+��^F�1c���o�΀�}���ry�"�|��eϖ���5�b�AΚQ�A��b��!e�j����y�ƹ�J+����A�ޘǃvwhJ����L÷�q�������EQ�� nݘ�S���0[2n�� |����(U ���y�3�(dl
5`�wDK���X*�Yb��hn֕ ��-&��byD+���J%�J���o��-���c��t��T���O�D�e����V�}MM��wz�s���<��,�Z�� p�<ʜZM<`a>I�	���	�R�t$�~�8E�H:��9�^��:�����W�qw(j6Ÿe��C:<:�o����K� m@Χ(F�ӭ�j,
gc��Bo�B����$����cOV�D�;��ӈ[�=��m�����/FF I�0�Qw�P4���D���Y�)��3����|�@9nf�h{��b�|f}��$��|��C�[08�q�7
�¨�"����,�Q�U2^�X�j�(�_��Y.�B/��BZ}���,$��K[ź�[��C��,�TR����T�$O� �9V��F�"��FrF���ޑ������p��'��5@��L��RH\���7�w������DU� Ejz����F��rc/�	F��EC(n:O��g�8�p���se�����S��?����m�v/�G��.Sc�M�^Ym0�G�Fv� �rѸ��w~A�i��f|^�ǉ&���zw�ڀjI*n�� ����(i �)�u'Q����/f訄<O�ΗAPY[�-�.�l?�0�����*�|��;���Xʌ,|��!��  \xkoV+��6>�#�$@�xk�u(��F��kp��xy��ӥ��s�5=���|Q������|<�c�(nbb��=(��F`�� N^�8O��Z��l��t�&u�;�-U�ݪ��j�@�DKd�Yb�,l
Wj�ȧگfE]\檌vl"�M;!d�ϊ���	�@�8���V��G����KO��j��j�\��?�P&��BR��4��A��%R_�3�}��N���4��h\�ړ��m��������+�<���0I �����~f+ur�r���%�A�EF��I���B���i��-�~�jF}���.`��I�0�{�ɦ�vt;����&6Q���|�1ݧ��[�G���Y3͌�G%
CV�����\��H�L4��e�6�^����ID9�"KN��v�ב^��y�
�V�!��iW�T~�Z�E�1
��P��r����+���Qj��Y���7��eyA�#:�o�;��(�Pخ��^f�6�D+_?�ͣ����H��,��r��=�Zi�'r�jǁF0vĎ�'�!jt��i#�*Uz�ړ�{��zb,�C�C���rr�n���{X9+�H(ܮ'��m�c��[ycj�#��Ո�gǕ}��7nH�֓f�=�(}���~zo_�,n�Z����/����w�(�>bͨp�΋�E���~WVv��<��Wc�o����y��pB&�P��De�� u��M��f{LL#nl�e���&f�mvS�W�@£S�KʉsÝ
��KTnǾ���Pt�9�f�k�)6 �c�3�uH�.K-��vkW�6oz�׮]|/�Gk��#�f*q0�����k���h�vi��	�00���1ս����0����V��%+�&�薝o� ]sN�?`�9J�F��=�ڈ�_�s��;����*>�+I�Btݐ%��{{�Y��zjֹ-waH�,�R���N�0���օ;w6g�(�PJ�v��ń!�h�:�=;���*gS`�\�=�Û�g,4�8c����hQ��(٬���T���YJ� _	Ŧՠ3�7���ٮ�����_��_/�}����+�h-<)�(�j#�$�%�J�.o0G[��j��L�ؘ�����v�(�[#��]��ߚ6�Qw��9�w}����/ �_���±���[�z�\�m&��^�&t(i�+oU��&q�t�z�ۻ�-;q�m�x�d�")�Wo5�x9H�gH���g����Č�%0�DC���p%ɺ��if���W�L7{�(��9?t��7紶�y;���3�ȵz�}!�� �g�]�`W6�42����M���M��s��ilm3����#�����M!T�+�T74lM3������[7~�a�Թ�0�t�dψ2�Ƌ!^#[���������B�8��.A�p��}�8���v�N]/@��ЌG�<��i,RP�ƊA�K8�ȝ��\c���~tV*�
��SH^L+����x}�N�����ߠ�t3E!����
hN���k�p�	���>�.쀑��/�\;�q���|�̙H��N�@����1�����sWE��jY&�\�'UOsw>!������9X��X�_	��!����\�"�S���J��)���/5(�*��v@�v!y��)�e>�%B2��xOo�ŗ��Z��=���ц8qD�t��,���Ϛ�f���"��T_[8��oMt�Rm��Hx�ݤc�t��ACID��Y� ��x�g����r-R���y~T�K����v>�kM�ώ����G�Q>3����z�Y��G�H����`-{�PPp�G�r���Rq.�Ku�@�2Y��l�-�؊�¦r��Z�O��a9Q��j:��u�̜(���.
Y���<E#�1�>�&�Ά6�1��0���dA�c&L�ߊ�8�o��F�]{{�H)�ѐ�"u�B<���H���g�G��^�\J���,A	 m3��_w����Y�C�[�2Yg��Gch��u�~�wL����A��6���pR�T�V`��,�����Ԧ�GX��*�q�1*id<�x�"�@n(�.��^X�x"��4��%���Fy��+�J]G��vo��+y�,�B�_�8U���H�u�{�����$�<�o*��n�]@���k�;�9��f�X�S�brC�=�ݘ%�����Oq�ܘ��H6:^A�"-1ϫǒ*��+s}hS�|��9F��T�u�5]u۠(�WR'�Ba�����D����T���ʺ�e�7�+;���/�٘]��B�����9���,��i�g@���������5_�G}�yw_�B���s�V[�uh#ق8�/|~8:+,�'I�AK����Y*�њ�eM�$
��2c-+kk���'�=0��6�,C�cC�>�ZC�a`�)$�H�5�(u"�@`�^����!���q%���!Ĕl����U�b�8����p>��0�7ҹsɐ��;�����]����6���y����-��."����"x�4G'z�΂�a�n���ƣr��%6(M��ڛ'A��+7(��jԚ�f���M�u�<�՟$�C����D�!�@���	� �p��v��f�d�C -�Y�;�Y�� ���|�c*���vkh̨�h��G�G.�Kll��Zw�lCOt'aPX}y��8�92��d���Ky�jD�_�1��u��Wb�}���/�T�KI]�Y���!l�,���{'J(M���n<�g��#�<��-׳Z�d�\��9]T�!�$���/���z�e��9����]���)��ב��8�t>-�����C��*��K㔫���z+|�"���%dS�}�K�.�kY��l�!i��%u�!��Y��d����eH�V%�<`ԗ��L@�,
8�eiԁ �jr_hY��.�@����.>$�bK��R�>=k+���꿏_���y��ݴ�e	�����ޥiK]�-1&̽�F<-�- ��I�,�պ m������vj(����B�}��`Aɫ9q�Ŕ���ܹ��M��m*y糄�p�������X>�'����+J \��u�đ3,���l�H���bY�ɀ>o�(L���yŜ�f���D�
v�r���'�p\Z�aHV@�P+d�S�)��"�i�d*�J@C���EӐPY=�$K�UNˉ:�NÌL�4mU8:���ml���q��\�_�sq�؅DD�������3.�9���o�����q�ۮ����m�Ҧ j���q���=�R�:�ʛh�b']���@�m�W�����įdvد�$*���T�����¹0��.WQh Prx:�p�F���������ƀ,��ݫ���	�R�Lu~G*G���C�S����幜p)N�-�($&�})�yb&�ג�&2O=)} H�C�n��p��VC��K���V�.�	�sp��r�*��O�VM��#F�$\}�o��fAU�ԉ�R��}*?%_0�;�v�?�~��2�,s��Iz5�_r��gw�?����	r5�ݬ�o�m�[?ĺ�7g��3��	V�b�j|R'#�\]1��E�1���d��D��-@��B�g�=����i��X)m8�ۂ���JWm����2Nj�.�ʤ�`���\�z�%�5��UtGԋ(�+�c����p��n%������D��\������Wȟ�
H��gYc�nSL��M�k��s �����N��p��S�9����@�9_��+l��_s�����#:eMl*Y���H��"���T�M��0�e��Z��1����S���Џ�/��,���Q�MN*�ya|����4!���s�;�͏忋������S]��� �G�9��c�Wg�V/�11��ԪL8Ӳ���$��FW���Bl
ZbҖ8P=6)� �ˊL��3,���ӽ���1j���#��EI�g�|�_kf�;��}���n=�߷u��_�wR"�E�I�l5(~A����7��p$C�v�9Tu�#�1���!6�e��},�ޏ��N=-��٢���cӛ� ~Z?\Y�u���^�*Q��"Vuh�F�b{'9<��w��E��&�H��W0Yq*"�J��-F��k�E<NN�2�R�4-��5�~�C1l�{�"�0�l���S��"+i�k+�_�S��-5ђڿ�6��fT&
%�S���zNN��{��.�q�z)u��ނ��m�Mt��c<
��M���q�~e^��:���������c��5 B��p�����e`87fIw
�*2���BV�q`]JָI0\��R_���G}5<hϞSa���;272.��Fۃ_� J�Y�J�b�@���.�ǁӵ��Hah~�������tO�e(�L��䝸� Y�[n��~��[�e\����7=`��N��)��A�gYASa�g8QFC`Q���WdW�He@L�\�0}_B�cF�#f�Q=-�A�)��-�)�R� gg���"4��Tk1E�����l�_C֛9�Z(,%�0�)a��^6;ab�C�Bv���k����ϸ}1M�>	��v����(�'76M�ԧ�v�y	yMHw���3���'S�#ռm�o)&�Upӫ��:J�t�zxP�1�����"%��U�|t4��X���HW�9nX�סkh�Z�ҹ`�s���&�7�cA�n��� 	7��{�V`O�|�@о�kTƥ'�捯���?��R7�n��j4	��.����&�#��]�����6�7�B,IJ,�Dr�]ڟ#3�Dx�8�{�]��u)�]��r�ؑ7d�p�$L��/�Nq4j:���m���3J�~�������p{8f���Q��$�8�͌
	�1����i0!ˈϰ/��.�}:^��J�1/��^�47�����ַ�$�X
Iʇt��1�u��vN{F�<��!+k�RPY�cn��]-G4M�qh�j\��Q�e�l�{��5�K��C� ��H�p��@9:Aż����h�^c� �)��r�6L�k (��C)�~�$W��d!	���.[l���[^!�����p�r����"��u��ɖ$A�D����NB(�<��i��J�;�n3�E=\'�<���m�ͮ%m�!>�(�ɬ��>�tg#Y�1�L�D.t'5��C�'�4�*�F��p+`w���(�n�@���OS�����^��;g㕝�~�4��ݲ�F�<!܀ݥ6��}'�_�ؖU��EI ~N�i�ݡ��w���Q%)ѵ��O�p��P�iDؔ�^�ܴ�<�i�D�m��-��<��9l4�Uob�P�#H�!�A3�iw��y�<��bB�� D��)���'�R�y�w�8 �Qw��OP�a�v�{U���fo��6��kO��("�oJYr�+� d�9���ɮ�à撳��:H���Z���V�{��j���=�$��P��� ��(�1X�����&:V��%��)a�PdC���|#��h�^�hFp�e������M(r�������)��WYX��6�w��m�F���=:#�f����Ja�k[��d�S�_#-@B#f
�
ƺF�ƫ'K6��sH'm��e ������U� x���K�qw���N4������ܺM�~��a�4�~�r��MuSsE�������(c�+tP�B�g�3�|�/N�I˙�����=��ַ0�.�>a�Nk,qڲ)�"	�N�Zh}��+������<��Ѥw�:w�`jN+���ϸz����S�H���Z��h �v#_��b>����O իz$�0~�x�f�&�uً��8��R���<K�㤳_~^M�N��=��Ea���=�D�c��G�o�4�D���W��o�����9ьo/Ӿ0�o�(3U�����&��|�8�������7��<t·��s�w�2F�`z�2!jk}�߫�4�ԁ_����*Z�jѐ.F#�{0�|�DlF�4�ґ�	�w%ʞ���B<����G���X:v�+�����7bL�R+�E
y�K�i��ڴ�ԅ�`�	n��X��1^�b�n�'���nW���RA#����3��Df��(�\��ܖ|
Yb�n�Y���T���$�u�	3A%�²ҩ
�`ʞj���zw��OQ�V�cCܜ��+��.{L§ ���,���b�/��z�u��<Jy�*�2"��_˕��lݘ� :��ч��3�C�>���	M�ˬ%UCj�`U����E@@rx�Bb��0}�A�_<��je�T�q��oBM1���}'N�FE�J�O��(dK���[��^v��� ��i�8�G��p �����Y��A|]�]8���X��X(ļv�h�X˳�?������x���`6.+:�LcS���3w��j���a ��D�h<Fj[2�=���4I��,uU��e�A���񏿊EkK���xL�m��Е�Ky��q���9��	�(�ޓ(�9RUkf/^��b���7w