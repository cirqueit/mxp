`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 928)
`protect data_block
7MHkeO7lKo5NqZdD5MOFBW1vvvjNE/EHjXvvvD6tlbs6oJuiG6gaygb1O5Hk3uyoPs8jP7p+41OJ
kEutGGj1HWLc/tQEQk91QHD8M34W60LpLUh1TVymXfkxz3hBnpLioEAmMVwlCS6MaWwZpmwar/nv
6aNspla67H9vTwQC4wfqM6cI42TYkLRAHDYywov+sbJ2kn/Ay2DaKfl4GQjxHH9lOn6dk28lr1tV
7x0nRsw7ZnfHCvBiwg3HU8UJ86cDIURbfD3Hp7pNpIYucoNrYbuoREqotbczOI5D5nmVvH0YhTnr
mXyL/lAnGsCGQYH6NiJxJ9ZwM0gH5miYynzVe7sW3tFOQ57CPfPIQdE+0BkV2zbgKJVs1AycBtS0
3UY+oO1msN/tuW6OqeVuuXjVcmIo7S5vJmWODkw+Q5COiUkIf2W/WGNDQbGDU7arfoZTEwRmJaT8
s7poAqwwAAt9Qc1V0BS40xyOcPvaYdaoAOLjiArB4f29CsECAijryQ1+zUGnVg8jnA+jEUryoPpR
NaMZiMqSnBlT0u7VQJX/r0jiKOEtXyBuvdDaNeGh36j5rL8ueA3XfybbnXtpS5P/LalHlF3tFnFx
D2KYf60WOWEYBdUzfUmK2zke80DgVU/5GQvCjWZCXbWXX/uhFxSMtlo8av8X8jOh6uHAlEkCPKsy
V4sEqkFWD7Q1bnEwS6/tu9DGpkKYv4ILOraI8uqsxWyjncldODc8FIonvDqGb+XlRvElTW72EheA
CNocL8NoXYaQT0opC1q96Wz63CvzmQtrab8U66ofw8v2NK6sq6BjBa4KVRP5F1l+++2djAbIzxsl
wN5Dxgbs8YUIt8ssN/uS9qFHih2EuD5UnXMm8vjs0riNbO07ZZMQrVZ1dt6t629K+jYBmCoiDymu
rqC4iOzO0TwRwRFVk9HSfv+Qm5lDbSfdPr87NBJsVmmSwXg8Ns8TMNJX0EvH3Il7nwaT1k3/NkFU
czxZyt6jaxGhEyvo5/RB/ro3YKmW+sWof8vMChrnJy36/lCehrNyB+5uLTOqd4uLoSW+fbwgXZD6
a6Myxx9dGxqGUkfBGJhlv6XO+owWdBCguKLh7IcEjrF4YEylEhTsYun4Ls43Jzq0kU/Hjl3nSMp5
ZI8YP6l3zyBlw8sXsfUXa2bQjXEoU28x5unC1A/3aSOyyumjdUfOXzC9SnYTjF0g5i+0Dh5eW9LY
GVLDVFiWa8sjPsAPIQLmmg==
`protect end_protected
