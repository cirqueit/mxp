`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
1NFS6UKta2yY3axXz6O2VxQYWODi6u3p8HgycDp4CBCtghE/oySkq9jJPilwxALdX62WVV6AepI1
IIkUrjX1agj9YMnSN4G2ZL0ycRf692jQwwUcp/cPyv0EhinusnSV7JUUsjg5iS8uYtdTRqa6wr3y
NeD/WUFhtYiatbxp2nTsEUqu6haa+fLh48Nvw++d9wdBc7tRHWuLuyLvphrgD9wh3ztxm8MOC1MA
vpstnVO2Lb+mJZz2VyqMJ4oyURQ4EU1bmSd2DRAHUb6RVMCVSfM/WrhMOY/0CAFPNGmQ990CK5oi
TPIibb+8SHStqmtnHzNWZGyx9ZnV84GDFwOAf1FbW8Ahk0FIh4CblzQspuHdIEJQHpjQKo50K/8j
T2qvthKRq2aMpFctBpcvGijWVOZlUZjEVfZXISEoPuzhb7AFcIYelxydSJyF0ibpUzT/tHHouAU4
c3IRhqa4YRCzL07Cpb4goxefR+ZGadDWUYV7bWiyujYPgNjw8n2LCnjcKRnDVFcK7tsCq3UydbFO
nDbG6xShCW40v/dZqIy5HtTiznDUS4IinT3/kP1r0tDmusRJrOnWroHRhKlh3syeFUL5U5U8GWHE
Uzsl4L7UsYcM7FWfqVd+vYqdV0pn/NSsv50nfVCRewV8a8/kh99sFll8k6v8jLPogQeS47S1gwOT
p2oSfYV/CxziSyOB4FLGWma/0s3GgF/u3tcgvm/ih8mD9HDNgOrdJjNbaNJKN2OBMHqpb8iee95S
efXd5nevkLweVlgAgZev13ndVJBK3CdfJoowS2jmHtFz19WX7VGlI4lxGnmg19gOioCVkYCGh+U6
r/LSXCfMhutxUrACwDOdUCpuEzV7FqZwppfefw27DVi8mbwvLIQ7+2aXTHpE81ZPRaHty96Ra5D1
Qwf0xBu13mheaaNQuP0Hmz4OVGpX/Io+JhIh0ec/Ko8nUr7YrBjLrcCxx7N1SR5ixbXvvw5XozKp
z05B+Nleiwm3XxbycPSGghyDHnRNXqapP5TtVeY29CyNjHbRdeZed4RTf3jQu1aWpTlu7ekrAor7
Yo8+DWxIDDALCqPWRiubmCQafZucGuFV7UICSebCnjs92t2bCxP4dEUFCteekIHX/ugUFKejRx4W
s/vroSPqcPd6jIAybALbRs0dHsnY+0/LTFYT4ev0lilDlMLILdLfvgLTrv38njct9YwPyhVTweC5
tF+6hbvwvd/7TbbiQKUX0G4ix2/uf7crLVQFsT0hzYJ7hU/hcFcM/7/2sqBNiqyYmJ6lnPLBaaEm
aSOV32kySpJHzbucYWI+O0oju9Onbth10GK8Rtu39nfONGRJoXEv6rv2NY0IKM9ze1KThENwC2aZ
lLclVqHK6ikVXUb+TeOETVY9Z2ZLdXl79Ysr8AkZiGUGRpcqaKw7i9pH26dX3H8HW5dz+pq04Zz0
8dxFMT58C88L1uWYl1UFN7lrWDI7sboWr5o852CarzJKisLnhToQIa1Aj4Z3N6GOk4A/pHLGY0V+
kz0duRpwxqE0s0YRwd2Mti3zAGC2wbNS3RKwtiEHyEg5TvWDY3SFNbLZpRHPYUPdbWOYvxj7Serx
5pXaE9YgDCvIkW4/cl/nWUU+PlApH19yFgnXi0HBS6m4gZ4thLjGTv69LEvLxOgfTtDrTFzU6E5W
Kd2mZpukZ5X9I0gvaTUe+OVq734XlWY8ZHlybHjL5WMgUZMQArdX/iYlNI/zbpgSgNbQQ1D63/SR
WVtp0obhK0SWot3yWcOnlnTR0O2+azdPvipfOMjFLZ7OK2dfvvd0TTER3Vpbe1Qhzg98dVDQ0uVM
KtYUr5FcqL9nmxrUVf1GX+0A/dUigM58DEfCcIbJhot5PGn8fFsp4/Z0P5qnDB/ixA4HUnwKlSxn
Nnp1EjoZQOLqKWOoTjfuSH3t3NGwAw5Zb5hKFGbkIa1jZ/iBLYST6QOnqg5Bqg8svS6JMLJTuLjZ
7/WZBigkb0pWfMKL/nJr82agppbfSFm/TNPW+ZJC5S3gk1maE6HwpSUL0mCwU5fe2bgZ5Hk7ve5R
jKFKhQrHGbHQpf0FmDPPyo8TFpQI5FCOdSvw2PQchDtmQqa8e+Bm4TiRzGibmtSAi5qdXSOwsBFo
6iBOlBcscFbLJf50nWTM0rcPSw+2TtFcLt9xrcpOxVN8pQY3KSu/AKmxMVxhy8fIqDMX368+z0jU
aiVwOWHXUK3F4TroL3yzEESXQEi1B4DPRv4H0KeNf+5sjjGWt6Zp4bO4ojmNKBL00dMbzh1Eee4f
ERPs/KeF7kyYfIHegYe7kWEJ7oTR49V/svtWuKE6k8J6SqzbZ9Z55/pr98Fk92Mct708d+qsQfQw
8QpKgPemGDjiurKJKUU/KuGstyAImvkhcBohGGS4nOJQcU8zpBaQBDGD16u1niqKd3s9ketI4pcR
kQ5PVNdSkg6R2g90BVIeTr/jJPLAtAVIatwm1dPFTJ3dJckW0cR3m5nbYxeYnW8dKy+CTkQPJe7N
PhA7aVuraTeIBDFP5fQBjxo1N9ZEf72XWa6/qoIm5fIbOPJ/4iFSXiiWxP56LGhgTuGgp0ySDkQB
RjX5W0JM8h66GOKuBxGgrr8FJiufqSckUEENkv9lKmjXIg/+DeZHPTMZZ1c7Wva5vTCs+sz/x864
LX/w2WEBWjBLon5TANCZ+iS5Ls+bbji1xVjy6LIAxNBPbYUOxPHEOKWLKDUBs+Zque+pvfTIisUo
VK5k7kKs0dS3fEfINOwh/RqnZlhc+vMzjKCLpnW8iKuuHryTZX5EOfEEKJnCoe+JYu7jifN48dnS
MZ/fHwbZ8nCm4yMxzwR0g5zM6+2hW9WkQc3OxcdlhvbZem9nofErD2eL5vDHxZNjE2Ow48drVDui
8jMI5OjPzVarZl55YCSTo+oI2KkG9qj4aWkuUMcMCnGAOl7iyR945c7XyBE8b4F6sfa8WH/OdQ3I
v7dI2itRQFcdetqbSAaFavvCUQJWruPaN5iadJfWMKpkAKiQV4A5aDYTM6EK7o8jeG/9i2rfC/u7
mRTlgZur7Tw7kZ0B6/6VG7DAN+kgFYnwogaJ015WSYf/6qgP+rT7GBhEjKv0Rs90UbKLdTtONvmm
3fYXBfvicoknE3Ivq79wZDAqbLk1eSxZryngOoyraA==
`protect end_protected
