XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��M���\�[�+��No�;'�*"�ʄ�j��"���g<C��G��YX�f��s��Y)�)4��]7y��Fәx�O�U��6��l��e��6�.4EW��B�T��^#֤�_��͟o�a���}a�� u�vl��/gp���4O8v�$���]��}&��ǁt�3�K|�6/��q���
C�����)PߐT�9��m�-�<}y\�{UP���)Cq�t�T9�[��gF�0�5�E�oQ�⛾ ʸw��k�(�{?�*mo����$0�Z�~ݣʥC���}i��_���$����e��ⷼ��o�b9r��-����"���X��TI�ݙ�ے|��\�.�^Õ�6sƢ��Ԥƅ������a�̽e}.�r����	֗�|Ix�:��Mnk��F����4�[x�'{@գ[b����="�)�5!ٗ;y���2�r��]���l��G��i�c�z�©�P�Q���]cpl�aX����Y��~�m�
1��,�$����ٽ�ܷ�����q��a ��V�n����S��Ƙ�fH�֠lݤӴ�2��}t�4GZbM=1�Yj��F�@Tڊ��6���;E&��VWi"(��['�o��͸�� ���S�N��=����`�?����2Y�����hw!�	��[z|əT]'މ�8�9��;��<A�¦��x��*��x>e�`��ư��k�Yz.7�ߠ�����uHpdꢎ�^,��]2��Ȯ+}�[�XlxVHYEB     400     1b0��	�x0U�
�=��:��2���a�G���#�.��@z�<׀���l*���'R3,>4���]�K����-k�Q�B�����7��d.�w�����q�x����ɬ�=�����=��׆��Ù���\�b�~*$��Չt�Ȉ~���|��Dn��}P�\����c�.KX��!�5�GWT�F?Ϗ_^ԑ�_h���U'�wWV8�s0�D�{�]M��"rM��.O��~�&����d&	1�)�� �f�m*\0ꦼ�Tw���Z%v6k����#>���U$�LsS��Zy2 �뚃�o���� ��HuS6KiG���d�Ώ���R�m`�F�6ԥ	��@�g���I���S��$1K�%���zv�)�)�)WjϦ8)�EA�R�N��Y3��01)���N�jidj��	cn�'�XlxVHYEB     400     170;��/�d2b.#�F�n};xC7u���@�������}�R��f֙f������7���u�˚�#BGGC����R�~mV���_*�.~B���d�/mi%C���V�=��H��da�+���A�X(��◥0��+2���ۚ�V�z�qei���b��iw<e�/��j�ى7f�G0tihuW#�.x��?$ىTPrG�@}�~���͒٬>�����n�5!*s�w��IU!�B�(�D��*uȱ� %�	��x�d�D����'���p���F�a9���coA!��(1��Qm�LʁWe���(�l�Ȃ��&��p�OD��1��=ΜA1��G3v�m��T3�C�����\�����n�X�XlxVHYEB     17b      f0l���L�2GjP����iM�9�����N#�}�)����X��E�q�K��)�G̭k����vN;:6ݜ�����q��*�;/�:ҵ�~'��]#3����lm�x���G��9���#ȕ�KE�J��";�}G	��.��f�ez�Q`����vM���s��Q����9��l�8�8��b�UF��`�� �lȊ��N��U/_ȌC/��	�הӤW�u 3�+���!��<��