XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<ĩ��z̵��X�%�$l3���M򾄼M�g,3���x�}q���m9`5|s�m��|�&`�Β�T$��l:�9��*+p�xDW����~+p*V�_�s���6��gDn�V��:{:TA�Bh+9��
-}2��F��P5���T� �.Yc���k�I��*��q�_X4��$kkLrR���9v��rqv!���.�#Kv�G|�5�qs=c�v�4�M*M����2Z��;"(�C�^]	��0䘱��:�p=<�����HB����H{����r1��WS��Zqm}� 
�M�ٯ������4�}��Y�L*���-�x��ڛ�g���3K&���������&���!��#J�!	���!cYV���=�N����<��33'�ǈ���.��J6{O TPz�+:ϿʌU�<�KP.]�r:ů��\d�#L�WP��Ŏbr��������Gɰ;�*�}4w��?�vC�g��)`֬�^��E��������8��/�kdQ~�ZPfVn�d6�t&n�w��<�h�����X�D�PZ�4�wO�$x;�P5V�0*�Sw����bˆݍ-+��h�oV\�r��'�Ф>Bj�$`(R'	K�0i�e��w:�6�.A��II��*X���'�Ej�@0����x���ZDr�{�H�:_�D�ūA�ݩ�<\��i�s�~ڬw�����)䨗���^/�жaDH�����mj7��[�v����a2xf��Z�����6�m�J�|XlxVHYEB     400     1e0�#њrM�
��I��eƃ�R�Mގ|v[������&��rqT>AѩJk�U�>f����X�wUw��=��-g��� �����♝j�/V��x~u������<��la�?���
�+Ǥ&7N��RW�|�'U��2S7� �pd����B��~P�3�CRN�{���H�`��vV�<n1��i)��NJ2����}�Z�P3NJK�6(�4Ih�s�c=(�/ k��Al�/cd>b�����`�Z<p�4��.<1�aL��d���� 9a��8�zL%���W�Օ	�a�Ɩ���Y)���Di�P����X-�]%�1����aR�l�K���j�4zp#�F��,svF��*N�4�wꏣ�2?rB� ���E�DaɷU�k�io(-Q8�_�Lw�8O�o��rx/v��!�>Pv���ݮ�d�<��֣�uv���5B����̚.9���@V�'�W8b�l�U��:r���{�4l7f�&Χ��I�l�QXlxVHYEB     400     1f0qYXS��B"\|��A,'��:*�!޾@�	8�Uu���uf�Q{������Y��e�n�4>Q�䭓��.n�aƥ&\��œU�=��&f{N���),��V1ȳ�\� ���x'���t�p_�~CU�hޣ:�嶳�߼�B��oO�a��}�	*�?u�q���z�����H ���tZ�v�H#���i{����1�΋�nge�]�<M�Fޜ���R��m�([ȟ_�wx�1x���#�BY�W*�xv�d.w�&E��U(���L�������>+�����,�;��hD�;R���Ƙ��r�J�^�����x2(͡��"J/��<���yA�H��ťR��B�r�R��H;��=�@PhL��G.�f��F�{z��)l�!��(���ى��[���A#��FL��o�h����+��[���h�)Y,��ʴ�Xzܽ��dީ~���Ck[�!�ځp��=	�	~��8��O��XlxVHYEB     400     1c0���A��ɯ������W�V�A��'�WL1���@�5*�GRէ)⥲ �-��ʵKa�ϛ�̶\���u�:�����X��/f�h��<�Y��L�R�_��pTz}�훕I�����:�kF�������p����n����=�Ate��t�*ش�s���/w�{���t{M]xJԡ�b����鯒R�����	`C�§э-�i�a=wjB�gi�;�+����/�2K��E�ㆎ�ڰw֗��u;��c��������6�U���x��w ��,�ʎ�����I�x��VR��`�^�?��z*uCf���n�ؤ/���ej�n����d9�����Tq�6�3PR�����{�F?1����SP��+
�av����ɥ���c�ڸ��p��g�1���a���3���Z!^�H�I�;L��胸�`[P����^pɌ*��B�/{h�XlxVHYEB     400     1d0�rӠ����Ǌv�#w��qnz�J�������d�����A�W��X,N��ʊ`HZ��O�P�ݭ�B���vl�%��{�1Wo���|��V�{e�%�|��sk�	���:�V��7]��>�"Uw� E���&g��P�\���&�i���KFY���&$}ڣ�JS�w�D($��À�l\J�M�������.�"P��_Y&� {J=��@���z�'/#�ť�{q&R�q��¥�ot�;�x-cA��K������9T�~Yl��af��&G?��tG����ڍz^��Y 7K�MZ$�����ĸ��J�!�N�t��H�6��ɯ�y'!&����@�!C�}$�4��'��|��!����Yr�\O���,��G=��1���*Ħ{QfA#�~��%���0��W�[O��x�����Ylt�+���s�Cl�3��d'�;XlxVHYEB     400     200��p/�j�q����f�Ɛm�&����'=�M�� �$+Yr���G��@
��ތȿP[#q�:j���|�r���ʾ��!� ���aI9,Ԉ^v{���}��jK�M��YhX�ڴN���@�"9t����sx=�B�/\��� D%��Mלk�����/�/���ȍ�����Cs�!�!.�$MJ.K=���	�p�33�0��#7E�����˳v�vUU���<�}�ox�B�"i�Za6������$ �H��3��Y�=�?�03���)牰o��ɰ/��}z5[���T�4�d�%H���~��Tó��������7�@�LDQ	�%��ȼ��Xlo�e�DA(��C�c�SB����q4�hY��+�ޛ	h����#v���S~��@TI
�_�����_�71�o��/�P�X�14�7@$�i����F��CW zhlgs�`��ƣ���9ma1���>��D�`���E������Ĭ��jXlxVHYEB     400     150Uχӈ$�NR�E���G�!o�zez+��7�wcO��׊;S�U�ʼj���,���,���d�}�J3�h��\�a�y�C���B�NB?Vz]��Z
���3�&�`6�z  @TX�'*�dԡ�������/R��6�@�]��B�cƻ�3�.����mB���vh�_���p��0��������
p��Ԣ�W"�s
�O�KE�rgsk�&���_��ނj��g��I`q��K"Ey5�͈Y������C��#�C���;�\fbJ&�Avi]T�m���[��Ѐ �-t��#ʚ��`)
%�&n�$O?���b��4b�@�bl���X\ = ��7XlxVHYEB     400     170�5�)��`)_0˭Gr�Cj���J7�ڤ���*�L�6�Q!�w�%�g饻�W�����Ԋ�@� �P�|���~,3J�ݷA��[ι�����������l@u��af�������މׯ�6�/
򐰎�[.鷽�?uH����$�H�xn�&�%	��Y�k�W��gSi� �)7A�|�W����\��>\QW����`��!�{�Ϳ��DR��z���uS�'���EV�iҊ�����~?�]�1�go/q<7�Yl��k����EdJ�ͧ�Rq#�}�Q�2��9r��R�'�W��+���Qk�{S�h��B�)�'5sĕ_��,�a�vK�N�{���.���ν �u��3��XlxVHYEB     400     1d0�d�x��n^�B�9���?ܦ�����ؙ���5]�C%��@(�&�ĺ����l�nC��:Wyͱ�SݡAL�9�����{~{��{���"�T��xjeOυ��Zd\)+O?(vQ���0�]���B��f������% ������ag�.?D�� 4���ɂ,g�
�3�D��~��M/�N���J!��A��Z
A��%��f�S������e���襄�\�Ӕ���	���g4���Н���W���\�b��M.�Ҧ���#$;����݄�m����A~Ϗ0N�1�zͲ�G�I��NTun5Gϭ4���ڽZq��$oq�>����������q�C��⧊V���W4�CԞ*�ȸ��~�����Cj�9�)k�Vg��ҧ����E0U�?Yy�($NL�p�uF�|��~A�Щ��o�`I���&_��uh��w�:��ʅ2���]XlxVHYEB     400     190=��3�g__�F����%��aZ���6.ʹ�ϯX�9�0�&�8���657�Y�����k��$�Ψ �b�9:�p~ɑ��e"��*Z�:N��%�|w������HU��xV:�BCe�?V2 �zj��h(�!m��C���A�� �>\@��t�oW�����_�*�Tk.ܘ�r�A��ƅ��_);N�<�Wϵ���R@��c�J' <�
����\��m�cZ!C-�m�4jQ��.�,���v`(�X��f��)���Ip�����|�#�vr�7���"�X�G�-O�l@.����36
y���	M�8�G�&q/_ ��������vUܛ+R�+1��,�{ U�� V_
8N�Q5�t�n��pg��#��a�{c��({X�L�XlxVHYEB     400     190�?b
@��tx��$��y�"Q�/��_����Ϙ[޳�%g�*=K�6���jb����-b�^g��R?�2W�t��w�Iڬz2�qJ{�ER�L�>͚+Ҹ���©۬�ڃ��Y��	|���ӝ6ܟk�h�^���^j�~hs��\3�0n �N��B.ʔZD^;���a��Y�(�/55�A�85�V���`�I���=� ���u���.�ֱYK�OE>�B*�Hp�Ř-J��"��#���a~4ύ%���Ō�ͥR�d�N�zP�㨧ca�O&��y8z�� њ��K/ƍ+�hX8��MXE��n,8*��}��/p�p��&�Z(�kh�Xlw�뱷>XP �eh?�D���]䌍�R�G�=��<&�.�J��H��ߣ�y����m��XlxVHYEB     400     150��^�����������9mOŷE|'	�5}{�uy2�g0m��a�K8���&<�OJ�s�* �U(hƯ�f[��Ƶ�cC���۶�;���~T^��C���!Oa��UK�Z�KB��ڝ��JZ���⢙��1��=�&��z�lU�z�vI�3�OZ�n^�To�_��|}����i�,'�4�E@xxc<���f�IH�<����	=ތz�lX2U��w�V$�!��(C���+����a;�"'$@��o.�Bct ���m�Vb�ru&�Tx�G�nzꢷO�_.�ո2���ןR�>���U>��OfaT�x���?z!G�XlxVHYEB     400     150���/ָ,��4->C�o�`�z����%|���=[��yt���j*G`Ye�Qpo =3�D�h�HcW�s�2rQ���K�
�aqI-ǲ''���/�z�SZ������#��̤�WN�	;/|��&�6������y���r�٧v7��v�$��2��7+v��FFC�oh�XOI�2����������MVҴ�e��{�^�HH-��^��;j*���o���r!鎸Q�9�����L�]p��C���>���&�]���Wf7.��32c�f���5u�VR�ݕϸf�9F�~R��i��T�q&�S�_�Ĳ���1�Ku	�⃿���;��[��XlxVHYEB     400     1c0z��I�c	���@���?������,�����u���)�n(-��cN�D��ù t�`u��X޴X$��X7�"(~�._��Sd�J����!)�e��F[)�������<�_⯗j��"��I����� 4k�)W���,Q#J���6:*^�)�����.���������9�$�4t�kn���B���w��s�%)�'�a��?R�'s x/ߍ��_.$�N��)<���S��IS
bŪ��r3nQ��.�}�����zq���B��KM-~�,FV���۔j���rp��1�w{7*D]�竐�O�Hz�rШ:j�6�e���òi�ǔ����͇�� �{zܸ��&Jꗉ)����/Fb�=��F���ؑ���6Z����O��uU~~�N���LT����sE$;�x4�9E3��LdRP������)�T���XlxVHYEB     400     1c0�:��D�1"v8Y�����o�*�����U��P.E� \�M�Cs����O�����8{:�<�7���^��AN�����#��w"�LÊ\�2� ��y�&����4I�̕�.Zt���M�7Y�Iy���ss���P**Ҙ��ҽ�$(�-�6��������G{ۼN�l"@�r:`#܊y`�K��:�K<��3V��x�&�y��׈�ol�1ŗ�3>$tbB����d��Q	���i���)2��0)	�J����5 +Z &[���������+�$:ci��|S?j'����s��]Q��i�^c�etG��G���h�.���P�\��u՜z���G�(���#B����<M3���M�.Ɏ����a���?i�?�ٚZ/���ʗ�m f:�@�g/|�л�_o��v%�RO�K%��e�o��3����>�XlxVHYEB     400     170�0��Ó�N魧��ʢ�lg�����}���h�~��ߔ��Zml{sm���S�WM� ��zI���D@���n;�Q�%$6��iJ:��O!-f�<�s�d���=6��So�E��v��dDs+x�HTf��+�wt�7Y�ܓg��p��c����&Ď�w%�7mf�s�
1?f|@hVk�Gcb�܉��s�-�+x�y�Y�pgb�|�oJ�Æj�ƴFD+�,N�S�}t����G��E�O:�N�R\WC:��l��'��C䃀���r�Ƽ�q��{�3��	��D��_��~�(�<�� w	�k@�v�x=�
�˰^���؁iI8YTbړX�H��&�eW��Y�sk�b��'�����<d�XlxVHYEB     400     200wǦ'��R��(5�X\L~��-��0���n�b���M�	�q��ܳ�����7����H, ���B��iE���@�oБ<�������ջ�6�M�vD�his+�	|�0�syݽhR�T*C8.�h��D�@ehb��$�q��H���h7gf]��=s�)Q�(Z��䃪Հ�n����` L�|RRϦ`�9%���ʒ�3w��)���P�7k	�/��z�uZ=3����>�+a[R��B�V�Hi�N��w��HY-�����=�q��W|2V��r�.�/�:��G�N����սT�7����2Y�'�>}F?��s׀X̄v�f�X���7�{�;h��B�K��0m$Y�ץN��߈��Z��5�1��
�MX�#�4Kd��wD��_��I̙�+�}fr�߿<a~�tE���9���4w��P%b�Jl�E��h9�|��m�/��s9�����<3��@�������3���7�)�%-����:Z7���z���y�s��[�@<�y�;XlxVHYEB     400     210���������I�����>��"�?�Z�=VF�M�X�:�z��rUF�N8*����Y�b+�z�p7i{�n��C]V}1������+���Q�8����5�@Z�栛\uHO��6�*s(��^���J���P5��n�=Aad����QYLy��yCc����5h��gH(�b��/z����'G��O_�J����'əۜi�!͗�',�"a��
�(�*���떭Z�Ty�]G��7|���坓�����F����$�i=u*�[�} �����!�����"�:ʈ��+L۟�(}��/%��?)甛b�JR��4���աjY8B�Z�2����%��q���a Ur���y�ܞ�8�H� �r�}7��,�����<���p��To&�j�YP���&�^�8���5��^��O �M�3�t��Ε��^r�f����M��6�㇔y��A��޵@,e
W�p���;��O�� ��p�_HqC��W~w���A���u#S�����XlxVHYEB     400     1c0�3/���w�2(�W�wS�ٿǤ�X�E�Ȣ7��`K��3�6����,`k7G��o�:�����q�#jzP��W`z�0!��|���bO_g�P�S�8�<g��a-�5ˤ5����bV4�|�`�X�-�,ʈ�B�?���/�$wM�v�cY��}�-��O:d��x����h(�AJ�ʂ1���b���ÖC�R�Jb ��dYWS~*8���tߚ���h����!2j�3�*�h�h��i�,�\��͍t�UkUj�����M7���§@�E|�x����K���j�f�'��*��׵5�ū����u���O�=��Vv��?9\���)߇�����|Â���z�����JlH�H�?ϭ`��K��b���Z��7���0�Į��'���_����Q�,A��5u���#�j��e��[��wS�����XlxVHYEB     400     160���D����}+�0������u2sV̊����a $� J�
�Vؑ�@�l�@s�"0r��������F�_8��t������p�ȋ�}H%��D�Öw��1�f<�g*d��2t��@rR�y���`kz��dz���~����ב�7��2��3a�Qk}��q/4�:����.�,'��&�3�e���?=J��x�a���K��s4k�biБ~~���F��;�.vu��ii�m5z��ݲ���Ú�����w�����e� Xߗ�!�O�.��Q=Ң>O�IV���Ri�X��^ݯw���<WjF�,+��(��0x�;�w
V�-�Zn�sj��������/uM�03XlxVHYEB     400     120�#��'p���2Q�['��_�|���pB��|���S��b#�+�.)�n��B�E�V*lY���/�v���b/���un>8���r�ۅP�tY�._�ʑ���������� B���a!�cy?����Ke��7t�ka}��s��+��/��n�ٲ�{�����j��6Ӑ��Z�=����=q���b>1���O
|z�_L=�Lӆ��4�:p�7�r
Q��q�sA��Ɇٺ�PDM�P2MϱIR'꧚f8&n�;�����-��ǅ��m�m1�J�>����P�XlxVHYEB     400     160w��+.6�[���qۉ��[
�	sIm���?WRW�T����oI0�G8��+�`6cq$��a�@��P���}�L�,�2�#���u��t#��v�΅ڒ�7#��A�V��� ���.�[kf�P�*yZ�+�.���lXbp�kD�K�����}:�AO�'g�O�Ƿ��#��v��'�֭TQ��b�I�L�f%!C��^�:B/ԁ��&qꓡ Q�Խz&�fb9�u�OW��I���ym����-���ߛ}E�( k�@�_��j��e�Ȃ�����%A*�ڳ�q��.C�b��s���dZi4Ż�
*���=׽�����pH��ཀ��be���lCQ��XlxVHYEB     400     160�0�7,9�/aF��ޢ��՛�G0�ā�]���ۺv�4��R���a]l�n���+gK�_��RwF~K�e��pU;+�fx�&p�MX���Nb��\g���^�{�Yd����x��خ�- ��������i_�>W�������<��Rf&F�ޫ>���r��@9�*R󺆳���+M9��{x]��F�2������qP��+�6��B^���1Zݲ�5RށV�t��*�D�[��,F���녰���o�o�� 4JS���*z�8M]���j�����^�_u���/|�{Q>l�-M~��ۨK�T�h\�l��^��秇�)*�Ρ�+h�S�C����XlxVHYEB     400     200[!����lAE�e���uL),sH��!��usx|��S�cLT�N�2�L�6��ӂ"豼Z��o����/"f��<�>�3����Dh@����lٲ�E���]w��O����TC4��3]!�l>׽�_�+&���,|-3��{8;=�gL���3�AT�q]�J%1����� ���@��F�js_�����w�	� /���f��������.�ViG��s�/����.����G6g��jD���K�e���rk��ؤ<���_EÒ�ŋ��ީ|1*�Awr@e>dP$6
(��ڂ�s��q����`�N���[f�!x�yˌNq�N���!j�Zw��b��ݷ���KV�v�j���l� ���7~��q����7�0j
��O[�T���ґ��O$�v�.���W&Yd2gl�x8��O��5v��ن����@��X䰵�$@LǬYP0	
l�������Z��6�� ^|P��8(t��t�ױ��XlxVHYEB     400     1d03Tt,C�fj�w�X �G6o�2k3�����z^�t���4��Ζ�$ϳ���z�\D� '4��j��â�D��50��/;J`�W�T�$^i���BJ�Gֶ��O������uDʋ�8�Y �R'%ZtrV�]b�Z�S tNd��B���A,�߈�1�U���u�#	����х��y����`ʹ������qs�{��/��0o�Y!�Ό����#�#b�p������FW��	�2��!�IO��I���kUݕ�e1�-���#KA#��H��P~ݰ����r>E�,������[�X�ըo6Q�HD��hf�Tq�V��b�K��J�<�㌕��5�.&��w׮�nՂA>�*=��w��0�cX=M�=��8J����\-���ꉂ?��}���֙� FnL,�߬��7!n-�����o_c��MA�&�4~{���o\}T� �[XlxVHYEB     400     1c0[��,$�nۿkM�[*��MoQ���Ӷ(�	���'�l���7�]��W48�#�N��KNL�?��԰��.��*�{xm��ԙ��[J��f*&r���W*R_���<��6L���>i�;>��hQ_�u �7����
�.0��������xx	����B�.Oͳ?��ң{`d��Q��F��W�mV6"�f�ԧ->�x�-ߖ!!d��Oǘx/�,�!]��e���R���4���݀�MR$�՜��գV3�l�I�6A�'��<��3<biy�N	�0T5R"���8�u>wV��F�ѧ��K���tͶ����|�y�����poq�oE��
���Y^� ��e�%ENz<�:|����#P�m����`/@�1���ҥ�%�u#�L��ɛ���|��g��hF�@��s�!͐���[�Xt��ԡXlxVHYEB      42      50`]�^ᇪ�MҍWFu����H�jP��G���q���U$���qU-[�D�5(^�����-�a���*��-y��_��(