`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
hndNJQ4dIAT6hwiPoscBlw36Xjrg9SseyoP9Yt5HtE+KrDDLSIkoQDg8KJYHAt+2xAhksLoBqeZW
C9zuoK1V/PMLeS0hew9+CR8mIH4HUzAhGiorxhTmcOyar+2LB0PcmXY/IR+FwSrKto+VyKpR3qyO
34zYKD/F3oPG3uz9nvzjwzLNr0a0aajOMJQo1xniFemRdNKY2zWp2+PXal2oBXX0wJuPoIm2Xwzw
l/bPtuPKqNtdzzJVm7LfHf9BSpEtoU4UTzf3Kq5fJ236wbmKnFMH2PI41NFEhf8PqmtszZEAR3nv
BBh6vsUbv0WC2VNJpTBkADmgfeqYoob5cmR+xCumWXYei8XwwjkIHl7e6aHuselCeBUI8vCsnsU3
DXQ2TN2rAXljsz0FlOotIeTr7EZ4SyG3NaYql0A0NO4/EYxvlYkPON3RQZtM9fAMeO67XETjlpcD
28STmBvocaPPpTUpIIN0ymWkVjnWiSjJXGFuJks3IJSlfsgon7l9nwug5OfWsN8FxhzZE5B/ABUU
fGPCcZT1D8pWaIKPyWy0tvPQ/Dj5iJA6ncr+bq7vF4MHThtbBYewd63nIlVxqvazka68ZZDa+dLc
4QyMVwh1sWXkLYlZzWBl1rWrf/NigVxKfVUD+CZxeG8lW2zqwxGtuNm1oaNzZKNshlA00b769RPP
RmLMfvmgTapOxO3oLbdXAgT9EPTLCEXPjOiy52rYLEY3EwfMFuxnJXoBXLUrGCMlTkVgFzJ6v8Zh
/Z1P2I3OwoVPwQqRwBrJGWRuOkUxvgASIrXC0rnq1g0M8j9ziSRG8jXZss2encp2FTBp687tj5uq
6EBwzA1cQTDXVtzxn9VksucFL5eYCAc5Z5kJDbZHmiHkouuu3FU7RH28m/nqOq8GyQA9HQFGd1Fp
4PETpTBqzL5F8uQrx9IG7d7fM6hRGunzXJFQW3DWs9yfyoTBeicZ72EHHSZes9y0U84+5K8/abjQ
bRspxBl7ct6KPgM0HzIeR40HIpQ7n0/jX705LF76Jjgbc1q7FAfkGQ2GnGhxm5LOCA5/YX31Oy7/
igSpk7zNn22nXJQu2o2Bpc+if7QHuh3SlaTDsahjgjquiPTRT5NnxGDxEThfnIg4em9LVTO6RCmK
pqPxtunzRA2k7C/wo/HUGn4CTIPAIlRHHXQPDksfxq6zvFYaHB0gDJ/43gjoboH7qxWuOmKlBozp
u1GkFLLdlAC8SwfbKoQSRRQr6MVVtiTHQXC1VAMJ1U9YHt3gLvDJCKGKu/CJdLIWLt3oBQyEOSxE
0F7LjFwECYy0HQWHwSMi+91uqZRJyTMViwDA0GO39glYcWCVA2Mm2ZqZXXOk8yTXDZdHDZytOdnj
HRk9wS+4qydCbKoU+tA6pvtw1pub7+alATrpVRHxlbL3XiKqNqZyf32pgk4Jiil6NcppfZLTiFTk
QrdWrkMi2HYejmCGfcGDqyismiMi8Z7OF52aHCSCpKtr14vWaJbuLitVu4gak2BNK/XUNCZi1wh/
yv+AL+CVWobz1RpyQXJXQRALvURBVK4ZdM5TA4ykeZ0Eec4c4akOU1GHBFI3ZBNFXALoIqHiWbgV
iANtFiM1cYgTlloC1GRv8NNi8YDFT+ZdVXHtI8K0dE407fV3XmFs+hLEBOu+hPRRZM0BH8bifHvC
l+Hsx8PanhKBFE+bqdPzn/jVamGviGuGX2xGgsRa8kclb/44boOF9bvRaHKtZkEHeMPNslHdF/v2
3Q4wZzS274ybZHRPQPL55KmqCAIS5aIr3n41A5dnuU/dbqdBwr/EUVMo7Shl6mGkoEzA+5lDto3e
y1zK5wlGpFn2JS5Zuki2KVh7NHiMTAjLQWyEx+yFrIfJmYnyhWW7RLNAUWNQMM59vKztyABG8PhS
L/2+ZljBInsYChT8NmItTbamfJu3aa64OOZQl+66vGS9nEfqApLebWpE0XbwfHGhjiee/7ZTlnoo
Z06ga01evX+Vm33BQPQ0ieUq8TNGLTQgNE3BQhN2tAXVpPaYA29R9WR/PRzJsZQPFliZecSqrKwh
iJfbWGaTbbKRPvFqybIoYqk3NRaJJDJwU1cLyZTAP4MVBGsRD32wgjkVY5gpdzJ+3OpvSV0jBNi3
wKhPGbg4CeayMfB4dOEgIcLX1PDA6z+ip9NL+QNQiurvk/Qh+cCngUpnAmr9lKKKRIvRs9XUN71Z
cpUUH4oyTIxAiSw+e8uU+Z5I7ChkTNYIEfd2OSFsTrMqcUA4Ls4UyminUljI1BxqyTixIi7XMojp
9CaYCD/C/uVC5sPK6O4l5Pxmk6ED2Us62HphWrZpd5mZvYLzGeVgLqID2gE2TwFw8FDOhmLPovZT
yh7qTL7nY+TVlhcD4GutPoa3KNOR+bjeXRMg0rn+dNMPlBNmRVNQFPy3Nkgh6RS8vlCz13bwmR5f
SorCW5mFronUeYpRzDbyWH3o45BEFpKuDgskysqSNK7Ad07+KDqe1+m17Qu5cbM6Jh5utB3goiFE
gIpIaYyWKo/GdMqWtu0kBE4JYj4YUQjxsdVm1TxmmS3BEg1naeNyeiFqJqEVuLNhhPobsND7H1Wr
JLoXd676ixNbM2blFuJ8Gb9PrSlZyRgSkMM8xSV/kGuvkZoDWtW8XcaFKSLIcMfZVAHzzm4TNyYI
44R0SMGwXosDOEGYZJxoLYpkBVTblxGVnRUg6OT2rQOY0eX/ChduNXECqhW8vA6/buMK5w8ooReq
REQTPvTiehaUi2O54r4Wsm+WdohB9TnubTYvb40v85Lngt9ELjU5O4xzfYE4NmZTGZqPfKpJJx7d
cde6bg70qy1/Wn0RXCqsZ8pvd9JgpN3nNSbhBYUqpID3sE3yKRYnqwP/tnt7n2NwckUR+cH8091X
g+rqF6sezxpjPQxvxATHHv9ZaFWKIDY4hs9jjQ0J5RluqvD74IPE7cFN1UXuvSgxcpW95AbXg9T8
o87GXmb/WiVlolLn0bzp9z2yyPjtVKjsdjuFGWvAycdQ+eoyL4LQ8uK0MPeBZoCSs87MogGByzVA
SAYirFj9mQB4hPyoTNRATeb2CaFmgDyGH8hDlUK/oQczqAQrnC5Gl/KtQVibAwz+74yUnKc8nG42
DOvoQqeq5AxAnYXCGxKzp4IFNJ1SkhX0m1Xf7X5UWbrPVK0owIv1nT5lvT+4c4mkKNvIkLgQzW0m
Bo5HXabXIrtfGIa0l9XUbMmO/Y3VJ/0Xi2EfIZclcRhRrbM80PbHiZaOOXT8DLnWIx5HTQzaFK4l
qWVSdyZxiHRVdhL5arX/zA5TpK1wtWU4ZGUjeJnsxvVVgy7wGfCwFFVWudlmGRdJwJ7BK/sVjmGl
sotmJC81XSYg92zpnW9GTW9pVr7wiFCpLBgusDnuXs1dtlNe8JzuHXEE99Z69eyZOHpD8EFAAw3U
8AEwdv9MTNtHzvmJbF1ohcDrjFvBWoX+CqZuY63EOR5esZ5MCGK7VTG3JJWz5E346u5gXqR31vl1
1nzEP139Iiq0Vy3XCu1mbQvDsh2fC+IiVTxWXxht6PrtlY3U/Oe+kzUeo7imDXm9/l3AJCkCuLTK
3hNq812PSoq87d76KDK2nt/xgZ4Jli8s1KWunGUMt68dcOGHQYgxSIvFT148F0rnj+4vWixgpYse
/jsAsd7+6QoDMwwHUKSTKTMqI6Ev1f1fuPJ0+dNTXpdwJZEO8oxU+lynV8ieNXp533TeW+dQEZP/
V4VBOrXTlWURPsI/s/VK38M2Ix4AqWTZFfYCR9MFyrFj1ZNASYm0ZGScyNMVlie9LtHNyIwhgWOn
uimuAN4xo3vGmfnY+VR0GDeqklmlwSrPCMBZMJHFplrFtjQvtVG+AUo723sRDbZAQJyVwn+kokdg
o34DW9FMtDm7QunFYkXUbnTwXB8mZC/xIBZo/l7RkZzCE46TdsmDNEOvVZOWCAM2aJx+AwjHYnNa
sLvlbUJ6OlI1he2SrH3SMCMXwO4DfMjMTCqpq58omTl0kMkRO7zydxWF4jdBMacx6aLZtdnThErG
dtHLWnpgfX094eT4AmPLYJB4gbA2Rr+7jGG4+p3STmBpF/B9VRx2QS/nBckrfIwhekIBCa2E8mX6
3mD2ADw18b9+M2GAR3IBoauuApjxu8LojY3CowrdXClSVPU6gSsXvNjo76ffJdLB96eS5Gw+2F5M
ZfPp1gIJQKDd/rMmN5GKbV3iPo/Cl/p7bps6rhX3lsBmJnOnX6WRAvCdtnSpjhY/RjfDJBFM9ol4
XfguvoDn3FMjRdhQFYfgvrbjipi1U7a43VJ5DaZGEVbaybBSUqLqy/JW4KA5H8+Yo0k3gYLNQnEB
7RIt5wIJdnB6JRvlIpH6GSbkZKJZ/868v7rinMtfbPOjHY9JW69P/tpy4FDwv+nms3KQYZQ6TO9m
0iiSJeKaciGnHdQHf1EzeAm5Gjg8yq/ui4qg3BhKOmuPFFFAIwhF33ijUrHwhFWYTlpmEQ5wUJyO
ZdM0c66ACjyYqS6H+h9bB1GBqhCzvNc5TIK55gRdO657BROiIblUdG8VgBBzo8W8GoXY/QnV4NxE
1CCja4mli95X97q7DWOS5qfqaaWa09HSwJDmQoKhbg4s8E2LKVVV+W1KUnWPcuKMFb/dd3ntYev5
CRRJb+1R46tGkryCoaz9Ahztmedda0Ej85C7sjNPkoofHRheC3Y5fK1/IY/duK1QPY3Tj3tq+G7n
Fhi3DpjeUqK+HTqTGJp2Psv3flSrMQTPop4dTzWuPOguvpB6u9m8YZa+KUnNj629oWsBGfYzv5dG
TF5poCi5hsDk+hxMzidYbsHgMugyVrFImzdmZZ/1ijGC4b8vCKhRv05csWrvmESPS3UHQoehY/Qh
HKbEi2gnaz+7mIvT/HA91FETQzNhwSwM5L+7u4XAkL2QwSJkJWW6uzENhcF/mR869sYo1xSJb1NX
vlUnnh3l1o4epd3aTNqAjrlXhCQng1SmKQJW3bsTt/E2QOcLm5rZTBPIjCNxcqG0OlX0ZuAI3oSa
sfzaKLw6lJEC8UrQs328OBTtMWFOdiA1dpY82MFN0yrrwBHOWVI5EuJDh5ZCuoaUdCCAkGpUWpuQ
7A9b9QWnDG7Y+u/Gx1wEcrL7cTeQnGwff8v7RCq+K+/leLI8RmrasiLBI1BlMcaynD/nx2udQFwV
HvniErMfN56Y+HBG9RDbvxdNVYq0rSZetbte88W/eea48j/zTO1Js77c6aaTnjcCMIiJ6eUdHbN2
GqM5LptsQeeY5rizrvq08BCOlJZsMWySkUlLtOgWujt2plRiQM7mxY0dfPIlqezOSgLcN8ckPPtK
EW8wPqzPxIEi/IjPS0pgXgBjOvrrSQwShQtvbErF1EylCX9BLiyVmU31cefBOp+x8ZZtmwpIh5bF
diIYGD/qmhNH+Gf3ASzvFOdW4zOeq5kjZquvlQ66Fx1zApMgg1pnIl2RJR/TeGHdc5fn+p4XkAj4
7KqJxboYyuD7hkgd9E1fpVwYbIDg7q+IrgcHQ5OwHNN2N3LWFx2Ow+HSLPXBWm+YWIMxaKC2XKE6
ChESMsaVcQBUdx2V2WE7Da0SJ2r43D2tuWNmiRD7qfvLZRGWEJ4YOhP4MHbRlDWAsMrJLm2TsKdi
qmY+aoPn+FvT8UIf0ZWtkBjsM2WtRr3gtE+QOCA0+DBxfpS6w7qbwUXu35JMjPoYMx+oYyMWlu3L
VOvJVnkrc1nU6YQjpLxVKSc6LQ3QTRLMckR7U5Tx325bL8d7/MFdqt3fLWEcAm29xYLri1blCSS7
x7mqS4qtdwl23OfUMZo1zlQZNFVW+e/8T1BLhyZhGwxzyoeoxWbRzex+1gWvvQ/enGK7SlcI4ehM
8zhrkyHBuIQcUA58K6CnMgPY3j1EZtNa/++6Kh1iawNoTAPrGI6Cbtng3MgF4yZM0vwzrw93JD77
DWEdDlvhW71Q1a4DdrMVABEqnsFRjfX0Pr2D1XSigscBoxRi9m8jRlDAHG/vF5efcdgRZUR9N8fP
dcgIYeG6Bdi744wAMopJDAH68w6TdGVsuXYOkHhJpL6YOgEQJAnmG5+7Pn4c1T7nkZbQXhDZlYrq
WERq2IJlzC4NdX/gqHmRRCxVMp/qi01tDMrtKh0uEa4MshkXFK53o+UfsT9Nhv7Ou1PWIyGjzhQ4
1otNbr9L1DfaBWcx4uCOXTCs9XEcgH2r9Z0eXVse9c0q+A0eslHhJczRHRtwxChNF0J1fsIEuFEI
8K3xnSoVDgKZY937fFXkcJkDbOSX7KkbVlplVydAr4jw1ehd7BpI5lqXhEDETrWSStg0hoqm72RB
HH8jHl3u/Iq1eQ6b4V6Qgimg8BvMOCJKTPQa/DqmWFuT4AGSdkzxJLkJe6vxufqZ0ewXW+CcteFr
8sWxIuS/1OrbojY+XmNVPOFFGVjKT3oo/E8KGq8tZ5+zehZaH55xyzCbJSi9sik5dN4RMfkIAq4e
Ztczy3HnUhODNhoJx7DnzEXPTuDoYUj2skcLK5kJ0n3HKN48T+tds50wtv1VFeNTwC9wIqB0mfPV
dD0q8/V7TksFnjpREED9C1iwGPs8bZcpEs0MJz/6Din3nroJEqH6gr69+BAk24s2+y1pSiQkBRwg
86CgyqXr5vdHd4ym41acauUbiXXaxqDPJGq4TLhY1MyNoYnxhFohr5CvRBxai7nlECRq5Mq4FJGv
GKm7hyJsaHrIfU3HHBZCsmM9w64SPOiFzC1MNMyW3519o5zB42TXOXqcTykfgkXMcsfeH+FBzmsu
9UTG15SXOFconMsGB7t9YSI42NJIukG+gX8ylhSa8splrjakzFW8o9j2O2gtZobav4uC0HoMP+Sg
NnH+KZtd7g+53RS2vQ8h/4pN1VQfm5G6YENd7bg8XI4DsFmf0zm1PZi06XczGrS3CFOPOjIYofTP
U0Ap+GxMpCvuAuqNLi6QahpfZJTYukxM9YRAH2J0ORVtW69C07U2rd9Phtanjd0HGBrnhY4WkJZb
6l000jmtcASoN095ZfeqIRgb9nr+XzsrTuKitFQ0GQD42LcMom8n6h+7rjyNe/iEETGyFrttsUVh
tsgvol34x6aNyyCUc+2/PODPSw6nzhYYuR72WCGdk5pAcLrnVL1HXYSQCnQZGjklcbgh92M5ai7n
kNeYkOa25jiz91Lb0Z01mwyN/gJhaILg6bdpsur/pfncM7fTyzLCNVJaa8glPzDxftP6/MRfnP3L
7YHXpmhKxQ6/nHSAs2u/euUTV+5y3S6Sftid3RMNNEcxJXekjAK4fYD9+iozq+UYe/n/0t5kT6r1
mw1LTiMWxO3kfyv4WFGDGCJG/IscJKRWkMGI4Z5lGG0/hsXsURWsLkUs6eyU1lHJLpDK0ZoGjPao
w1Vp/6I8v2jysxJGOYboYAllm88GPrYao7rkb5VYAH5WaYg1BLFmMZrQpeFGgAG3EtfQaOwkmSJw
IWGXDG2nVyRJuAKuDvwG5Ry2skGd8Z3R2P0o81BHEf4y3vofB9Mn7pDKny7LvtoH/foyjh7e3evi
GgP+Qq8o1Gp99MtxCUmIfw+G/kR1fxCDpmSEj1BJwt2dQfKx2nFrsgaarUNZFMSwRPGSTRape9kb
66KhlyKCSq0gfHs7UpfAU5Vdr+g7KAvO8eQ3+kiKDSPmXvuAxMdN7L14LuifcO1XthvDX1AicWBI
3XeKX/X6Ib+1KK1IFDUByaiYL63yCN9qUsFEzp6TgKc1aGm2Eto/rbp17HZgFvl+SHpNrf8psUp+
34tHgR7+arNuVGimgchOmivYN1Qm3g2cgE/AW2t7gxrgwMuaRlaEFsDjUzWjCZwAKyuP6P0HCVfL
TNin1GO/cAAQa3PrmtPYY7YrYv0CKKpClMG03ykB774CDQ/mLlbZ0O9qAYwhg5IHw7sFTFQVsxVJ
ucoQFUDN6xdrLBnDs3CftPWBU3qhlSuvbwJJjPyOGX6E+ljLIIx09BN6d1uaLfg9dH6lFmslOen9
t/Nsbw6ZzSXuuPTJmL7OHQ/O01CgxL9AlgYHAzwS7fD8iUmb/hflWHpSKizHMgsYhREkgmgULX7G
Jr0itHxV5x9LjOjX4pf00gFY25msh/SG8lv1k+JS0LiCj2qShsDiWnbnAlVQdVCkqCLu8icU8ayZ
Jn8KGY24sfRsreqYja2okLZdBHpmf1b8+XhTLwuAfMZMv+/w4WBpWecD32oZ5qpXYXmelTbKy1gb
O9Kc3ESgMqgjhG52oJWRbHj39RJ2RPHU4iY2Yr4O4PrxDTB9cJsAkDoCYweY0QkLn9FrUSANiqs0
y/rww25PzZI/DEvAYD6VMPb+ExMN6TzypjQR0xoZs+ygNCOPOS0dHb98edwhdERnCX8OwIooR3n6
qWM1Mq2QR32zjQE1HMjZ69enATYF7gXII/zFV192r3FaSeA7oU4BiAHHJr5oBCc45vc1wtxxX5cq
RjV4cgc4McS/6eo3ywGxHiH6KPvNFIC7gmhprsesbQ/ymiwmw0SC3dj0eErFtS/gA0xYCBElKXg9
9IO9jxpKfO48f4v7Ao5pcT2h9qEBqUJdnnzCLogGRqS68C3mo+A2JQbWcrwcbal1kLfpcIAANnRW
vAvrIedlGjxH1UOwS6ESSPeKXBLG9a/jsKwKCQiHpEmOf95P+IeXchkgXEjpYSoBpoQEMzQ3UDWQ
S2bgb0SmS15wP/uym4fi2oQKG2ewb/97eMhLuG1wQgEVS7tNAVNpL50WY30ZxHlwvETShsjIlnXC
eO0VkKdfrB6EL/f5jnRKGeI2QFdzdYPQzx9GgLHyd7v6ZRoU62sXCeqtbYr77IjrKivwGF2D+cBG
gAeYcPvoSLD2/p59/O4EitZPDnwaev6GMl7swZqkqhQW6EC8vYXDpkcobpwFlXP9QvG6zKdjn38q
84S/qnzm6togImKDKkuU42X/ZcoZPk4XGlVEdhTyQR24BZqM62e3nEHGAZ7cKQyBYmy6Ew9X1AW3
ugc/WVDbteCni+z8jc9G4VEnVB8Ocju252DOwmkCvja1abnmZbpYVUHy4f66u9l07Mb9jKf04DkT
nU0C5dayG1MH4kbl23YWTjCMNfGVrbnmoq4WFIV9t3Kp+81/MNEa3VjVo9QY8ckKccOpgkiztTSh
fZVBZ3JFBvE3A7uu33A+ghBaQpL8b8Xa0R4SYwfG8jvPDRw6ByCHcoJYlemXnzvkD50xNwhXSXty
Tvvi1ICidR0lOXtD0/SPL0fq5fOAomfJWOfboYwKARMlLgcePwBlsMqLCCFP+Xe0j27fdFhIgc2H
rjGX39VD7YvHdhvOMGiYYh8No2OVZ0PZ4ve4XmjHM3Y4EWtC6JH0VFa6YYPeF81JSkcIHQhlkSwH
AiUihTi5kP5O9xWXg2l4THXL0N/bn4wJ3uKcgJCyr6AfkkycjOhPFH1jGkz1z49SP6GwYeBrA7ss
iFSDt5CS63k1fMkB9hTg5nvWYmv5Y1CXBvnHFVYwsKoLtEYDKWKV5RoxYRFfLPzs48adU3FRrQlx
IEynWvFNxdnZXLXnnNdna8po0SFmNZVYMLTE5DxNBF5Qr3VLLSfZnEQ+PLzXCM4VXjsuJmSTFPiZ
MZJCghtHzDvrn1kseFLqohD5kruevdl1mxPR2yFanGNhMj7dTjQ6PXmZOrz4WFj/IOzmyhON0iAO
kQQ5StPIQO3vUxDB2ZdSJoXz1UCRLBP9v0MiQvU09TlEk1fS8IZz3Hj4KTiPFhePRJ2TsAcF7m+B
rdt1jgssiouO3bEcChdAtdhVZwnzOgxnQxZDmJs84rIT/kPH7pOdaLiPfb0KFY+6bfi7u+114t8G
DXrPS+OEP7S0E6fxY9lWPzblKHsQjFTN0aPJliwvFLWKFm17I5YDZrpb236UySlG2jfAdz4bk4Aw
Vs40m3dmg5wqxZeJ31F87JwNDLfP4TjDzU2j71Tn111Ki/dpySl3ZxD4gxOSSQ4Zn8YAplGOBHr5
XcFDBILtN/fO1rdYQWwj9TNr4SU1nzXerpU2vv5qfMz8JqA1j8uvKkTdIyUpw5cVql1Yg8bqgLFB
XFWplBxYEVmroTVkTKBBxi9W3gACcsLJjSitk7D0Bm2n4CxTjlcUNE0KV+Gz4hlV9Dxa9lazWbje
sOY1D3SJgLS0EvMbFI6T1lmr9VgU4E2l0FAQozVdI6lpv2PCqe2oK9C0+VJ3XTky7ssLi/y2ifrx
6Y/AIyIVzsLBVVghkcwnAiXjEb7AaVqPudTlmOZhSeYW/fnzj78xt4K8XrhzbnVrIEn787TeSFj+
M/q++CBZ51CCc4b4bkUp8DQmBNX/4ozSZfJwn/Q5klHHZQ6V9UbUIzoXgdbWjJKXHD6PGW24T+nt
47f7Zi9+0Vb8xusawHm2Jo1JRa5RcdwSX5TUl3jlK0RiV7Tl3oq94rONgBSbSLYdB2X9TWeg5fyM
B7+sF4LTa5ca9h6EO4UFO1yE0RVO+ZQ3XJQPANbh7HqvurEwG0hWVCfFv3LBNBzL+LVv9oOXBU5m
5/qI3hcOQYLrVRgJHenLzYOGfrR9sDGsFq0OZhtfUTpHdXhboErXwi1/UgC6ASRkDzfAEicSxZFk
ZLiKxo2JCzkUaE61tgP1pbSNu+eWJFUlTBv8bp5CjK82P5P/CVq93m3XAGgVZTGgImHT6Gz8Xpk8
a+Y7Kupxk4v83I3QND2mQkipcCnlFFFHGrgNC6V0rp+XzBHeYf2S9tV9UKPmzH4KjJceWcw0njIo
aDqS1uXin1lSm+Z4ryC+WtHFymmI1wTCXJHDpra0cSkH410a2YLjuRdMBn85StjkcONRe9iPEo13
bAd33enqgS25MGf01ohR0YdOJ2mrwYcsYlCAfQgG5ne6BDr8ioRNXORcdcV9EOcG81/ZN1tyFZYI
ss65LGuvWkevFBpEE/ysjysqRxhWlAKBlHnAV8RpKuADYnlsmZZRaVBVuC/GClmdI4UG5AZnglUA
6wglIeXeUrA/NnR/G6lmShjquWweElvmEooJV0NVVJ+K1w/dQn92vSm9QaKPfHsVqT3HZuXWUmMJ
oxx8aXqnZdsnSULoKW8Bbr1rjAwy9mIGpQMrx2lS41CLnSCpD+wVKBehx/C17BXoWN0qBGZoz6Hq
zxbT0o8wZ4HhglcTgeIOnBpC2MgMzAtn061uR45H4k5acezVT0CxyHGlK4sCb7NeWNesaO8EEm0x
iqeXVbLnoUtt4E+L/e8f2b5rHYn1
`protect end_protected
