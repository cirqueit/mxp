XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������&I���rA/�s��t�2�E�f�E�D4u�ԁ�Td��V�	�V����,�QG6����ݯa���oXC0�Ŧ�*�E�~� 	���{*C�����ق<���'��6�x���3Z��0bX��I&�/�Saq��j����Д)��҄I�
��o�
O��M��ʑ��3��0E#Z�� _�$�6�+72��3>*����aXSؗ��F'n{ͬ���wI 4�F< g@�F�@�0%�k���Ċ�X`9�j�Q�9���'K�2h�ܜŠ+��(���K�G��I�EH�$�ow*���g?�B��&��βot����pv��}רSg����f�.�0I�����"OR@���kA'	�]��'q���FJ�C���BT��dKl�F+�����+���p��ٔD����ώ��=.1��o�|���%�)��'g�����bTDh�IB&U�O������'8�1�!�C��*sJ�Ү�Q=�=�����
^�aܰ?=����NW4GJȣ�M�T�>rCFЎ<@�#Y�z~C�t�	��3����%v��d�=-I�ze9ڵ��˖Ɣ��vi�.0!�D���'}�'˲���Xk+��az��f�!v�2����IB�/�!�o,�!i������oө�a�ӼI�P w-��Qg��3o�1S������Ue�n��Rb�i�,��B>&t���{O֠;�0��Q�4�;�Z����[`'�|N������ʏak�ѧXlxVHYEB     400     210�k��%����V����K��ɿ��0�}L�{l�l�^����E����,�"7�_��(JXx�y+@����+	��
�3~���-\�'���$W#�ǡRp\��13��5�X��Cw��q��$	���'5���c��=�y�?zT��4����h�����!��N���k�پm|�c�я�����[�u��Z�(3Q���x�]�x��i�Q��Q6�W�wh�|��hqH#^6����b���S���Gk�*��H�b�t��a�M�QOU����l0�b? p̺_�H3�!�[�Cz;�$v4�olȴԸ[n����F�Ĝ�]�J6u�>�I���YR�9��ᮥ�нt����r}�A�a,��Nr��3˴�D�/XJ-�K��O������+{Z6g���l�.y~#��O��ݫ1����;��3�Ī�O��KN3e�����(�d�	���|!�RI�ܣ�+y͈��t��4�HY�� &c�����i��Y��*�7��Ee�]�vB��d.U�:áXlxVHYEB     400     100��YT���h�'�"���Wr,=E5�g�C=�4O��{��n��rȵt�h5%h��m�/g�٤jZ�ֿD?S�Z�:��rt���4�>��=Գ�;���\ay��B�(�4�A��X�[�52Z<��!#2Ha(K�=}kn�l���eW���fN���QC�<|����"�Bbh�B�g��,'�%� US?�X�-��!'e&� ��eX��XDm�����x[9P�5+B5�W�?��f���w
M�7k xxPXlxVHYEB     400     1f0���q�}pC���ȵ�7�������x�w��AT�6��_�*�c>�,ݍ�00�5�H��p�]s�GRl�N�h��������8Ē���8���&-�EGw�����Uhb���U`���zo��r�-_��{ҙ��e�ͼpR��/_�G(�6�i�zlA.I4s�f�w{�e2��I} ^��:޳����i��q(3ݳa��FF�2[�]�5��:N�Hu����d�N�s�R@�����[B��ן���2��G9d�����������A ��j��	�͟^igvP����bm2�-�`���������b�I��+��r(�`+]&z-	�	D7�[���1��9a���S\��Y�����:�!���e���!Pjx�$�Y�;�8޳;ϻ�Z�jW�ٖ�C4���"�C&�W/�E
��xI/z`~�
,�{C�����1��u~g��Jŀ�~�ˉC��O�Y���EX���xM�#[��20��aXlxVHYEB     400     230�U\���8�G�Th�,����2���œ=M+<�=�Z��P�̻�4N�!�y���� X@]ۤ�z4�y<Փ��i���}��
W�r �N���a33�7H�@���>�>��E��Ū�Z�9��Qf)Fڂ0W��B��B ��&�Z�2�XY�6J�ɷ!�	����@�#8T�Zf���2^�k���[b��߱��\��+lqbX惛�"�Ě��k&��%$�p9������������'?;Ҍ���-��3҃�0��,�5��dTf��e��=S6 cym �-�`}i����^�)jb�n�ϷZ'� %�d�u}<���ֲچA���0�*�Ea���8oK�Jik~�����oh�?<W���DGj�	�}@���] �߇֥�����A��z���
f
˧�j`�!L�DH�ȹL��Ḿ���x�8C��s$haN�U�����iJ�]�H��ލF���ŏ�Ro-9cn���O1�ʙ���:f4j�ss� ���� ���ݡ�K1^��v����,�Tb�������Ş8ޣh�m�)� ����I�hXlxVHYEB     400     1a0^���2
DG��Ɉ���m٨�S�@���]�c:Hvё��mWڀ�!��2Ko��+JZ�Mr��: �.zG���_����?ƿk]^��N�J(���ݒ���G��M�z��si���?"�촊��c�_8tS�u&��ER�c�I�F�teb�1!�38ܖ)���!rQ�NAj]ʙ�U�T?UG掛�\�c�/}Z��ܱo�'��|�t�y+V^�×ճ�M�cϒ`�2���7:Q����k�ka <3��'�}iD�2�gt�2[v��"���,-�C��w�2��1�������exҸ�A�؃�c�R� θ�+X��}g���o�&���$h����BTo
\?����;�ps8���|=���iB�9���,�̉iV����jB{�	�b�	�Ӌ4���WVXlxVHYEB     400     1a0VH�^_� +р��z��Z�Ct, �x/޳dџ�8�t�B �Q�o�+\z�@#e+$��0��ɴ�"Ke��D� y�lf�(,�����r��u���&��){�rH��Q���sH��v_O?��יz�S�ɳ,)>Y��!�C����6��l��#*NK�H�2s'^�/"��#dϚ3jZ#�5vT۱��������'�_(Cw�ʘ�t(L�/��Ylk6�b�z���eg�2����:��ň&�s8��������&��v�-Ȟ=��;+
\�/�����q�I>�ٮ�h"�g\Ц�~�J�+&j��5pQ��͋��5�(q�F���q�TG3������U6~��s���/(��|)b5~�-i�h�.$�=k'Ҝ��6�N��%�k��miXlxVHYEB     400     1d0�nP�ߔ���.G����D�@E�Eq��7�l8�a_�����	�k5�a�ղ�B��A��=�Z#4Uޤ��4�!pՆq�
9_�R��(��{�}]\q��G���K����$���:���+NcϹ�w���!�*�r�T��)�ϡ�P�2����y�9� m�i���5�������������*���)�h�(lVc��+��e�ҟ�O��A^�{���-��ȸN���1��B҅#
�b��Ş�{d2GA�ʗ�Z�H�Y��_&#OTx~.?e �Z��ES�a�4���� `<������3%jt������Ԓ"Kqp�|p/��Z¬X��XYQi<�4C��?�k���ebl�>`<�\76e�F�<�#���"�ې�s�fu]Z�����rN����=�
�	w�����vR[��z��m�I<$���)��fػ��8XlxVHYEB     400     170^_������m����ry6�_�>t�V�W�Gج��M���8�$��.�mn�$��P�K.
�7��P%Y�ȉ�
�-MXa������d��H"8��v��O�u�D�_��"T�/t�*�,�0W؈yiN�G���쑟��1�T># \��/�ˉ�γ��#��E���i���$@��g��j�x�]�.5�Oc�#/?��?Z�����H��r�%c��Xќ��D\�5�̧)1d���G�����)N�w�2�BC�B�ɑ��s����7f����~1��!2]�5/{Z)�0<!�2UN<���c�kJg�c����=5�يa�n��>�y|�-��`ł�<�J XlxVHYEB     400     1c0�[��d��K���I�U�IXE`�my��l��M�����;��U���m�������dH$}o5oX�vˉ-#��X33����������.n>�'j�h%{�}�}	x��D:M�������˚�o���l�-'9"��R�뫴�
�_�q)턂ob�E�.]r4�b��*p�{l||����ՎƈrM2)&K6I�^��m�R�F���2�_F�a�y���V��?�i�(��@�*B�����S,�W. �pN��̖�o��`R��y8���^Q�<�qzJ��
30����X�ް�����l`�B��I"Mas�u��D�(ܷ���]��nC�ַ��V`��E�L\��4X��M�T��E�|G�K�J=+{XD�6,ۈ,�yF�S�le&�� Z�����2+3�r:�|H`�z��n�0 �g!�d�q��]L�dFTXlxVHYEB     400     1a0� f�4��U�� 9�Ňt]햧Lpb�}]�}����*����+�S&(s��H�]eN��M��B��iS��.��H+��QDP�;�Y�s��*�
RA�ɴ�Ҩ���`��fQ);Z�0YRuI�OZ�m��6�!��m�o��]Ґ�B;d�p~��^1����YW'�lC!��D%��w�2*��g��a�7���8�a��ޚ��'
�WN��ja2�/.3�y�R���4ʂ�]�f�t���I�H@�|�5��?�
�:����H�w!�r�����* ��)��؟�y�EW5��P�LF�����a#��)�Dm@WC"�~LѧJy�-�O���ČV��c;��Pù�����iy 쎙�x^�ƈ4���'%Α���n�!����Tz@�>�{dv���+��>� =k��XlxVHYEB     400     140kIIy�x��'^�� �����vb:�J��TD�s����<փ�jY�X1|�	PYG�j���$��"��Q�(u��э�975� -�U�u=�]0�N[k��2i@�0fS��NV��;�ܽ2=��̸e��쀻����b����\�pR�]�)�W6+4~ŉ�}\bX���5�U�N��ēk	�����cF*�N��{�B2�b��38�}�kĉ�j��q�=�W�(3@��y(�����?�I N�K�&��̹z����q���Z�n���Ҟ�R<a�H�e�6� P=a�i�
:=�5x����12�/���XlxVHYEB     38a     180�?,PM/
U�ոpԧ�=�h ��g�ܯ|@v�w��c4���'bW�X�U퀡�= �Dq�ɥ��x␉F��XC�fR��{ �!w�t'-�Y��ͼ���$��3P���St?p��l���b��8:��Z(�f�����4�*�pkq l�$+~���58�T����~AwY���)�S��iڿ^��K���B(�T����V����
��v�C���������EX��x���D�����+����l������	�3�*z�(�x��4���W��F�'\դ�u)�"j�Sp|� (�
Wkn^XY�jp�V�9X���z��/Իs`�����QW��dv���\�G�-�H�$B��JÀD�!��8��|�