`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3088)
`protect data_block
bbiyeRTZJXAqTRYlWJxIsFClZVVtULK0C4k3TIqKl4RkpZDfvwHIblvDtE15G/lO79hJIIGP0Ws0
tAKI3G5jDgqmENnVVhHRDAi4wDMGoEgOBQOklCFLNcrVUTPLiLT02/lO0ra89DPUtCkePDw1B4iq
u63TG2IppbF2asEH61yYTZeOQQS6T5hfKS2Eq1kUOUv9vGXrh3g49wd77A51iUQ6wkzjAVW771mv
ZyBQ74DOb5ELNjfjYvRXEONEkUpODcCn9BW12U87zmwIKwUvk5iBghDaJQQE0XuzpOTL3QifcK5x
8CYBlE7/bOXbNhrXoczKx4wjEg41Ouj7EMXRjj5JMx4YOFuK2qJmbRXSMhofiNEKqWT7MpPNbcdq
tGqS2yqRuPETKQGRyCgpHc1T0SNmw8oMuXYKyztn9N2f3afpgxpG2tfaSYbz6P8c3Ph4xwWNMjXb
ffv+IMRszI8DmCBxtUi1djuUoAAlGifkn/c9k8UVwTtd/Ma8NUjGa45LVDMOMVW5h5oHRp46/lRm
KWOpJqiUMNLrzEWL9bctwLM8b77MFw82fZERUr4o8/YcZOs/Wrz1B/H1cKkGWegI/E/Tsm6Varlw
MVnFATEtElx6DYeVrW/IaNLffUeiQvS1FGmBXJIefzoeBwHi01w2ImxUGjbvSPbmqsTdVcv+piFC
arBEBx3GuobjJKkRfd2yYvKKubZm4mbcaUa60tju2LY2hv2k9gvjMFOZg7n6cd4UCV+j0Zj4n5Ha
isL3oC4l25ZOYcQ/55aV2guz2xmBKk0sQ5AO9re+0nzezdE90bgz3ZI48CFxtCWiW8bJjAMTmgmE
LwBFlRjX6bhAvJlFtbEl0E5kLpBTGWsXlrC/T23AfSlMAe8J4Icyr/zFmTipGYoa2SkVuHSYDXEc
TFswmF8QbKUXUFwdO0XxVoTFx082NHZaif/vJhKNyMW9Ah7AuFeq05DgcY/j+g1fxZkBtrw1MbEj
omqmEUnQZQT+Ga2bLYd1KY+j+2Is5CChadfmZC27Wf29LTU7Px5OO3W9K5CTAp87nHnScQqep+Vc
yE7Dc+KheZsiZvm9f9X3x4DgDwokkTmIZWfTUIADMXKW8TeXFExHATL+XcCGkUUPiAqahXTqNaYD
+OPhCaXe4boAJkdUefEjSlkCBcQPIJ7Obz9BRisn3aYo1hjIAUaQT12uA7Hlg0kwowMVjqqVeD+w
wKnMaUmHIAJWjSrBnIbcGrjXLCNoWP1kWgtdFq+ldhhQxe1+66v47U9OFSJFWGDEmrBRr9GgtOMr
U+xZyKcOEZ9LFp0WqKj6Nn1UJx4eEcRHWdRbL7sue2HrNF1PipsBjAu/LaOMFxoHVicWm64MvTLm
l1XM+XGWQSSI33mUYlWkEVosdbz1X9SyXJB2oTGJ1rn8Siqa/VIx+aFYpcLPZYvw2iSJa0sCfksc
DPtWaTQZ0S5XjzPm9gqOCymALnTP9gxk8AACmkqnHAqZyH/OsznJ+dqgI2WIUMHcpc3rDqTs24FA
ZCmD/lsjqfIqXFKiNq4Gex7DEpr+vmu9k9ErE7RsSfjU+D/mU+QzpviV2EM/np9Le13om1yr5kbd
/9Vva+zrehYG4FN0pJlYaGnNk26jCqRJzTnvfoygg0kHL61OKjdurXzzHFV4plB7PmvzT9EVW/Tm
OGBcLCrU/zlxlhoGfG8ILJ8bG6Q8aOR8GpwLzbK5WsmiITL0NYQ1vYzQjDWHCnL6Sc/TB44J9IUM
XAmVCcW8xSo0wWXfi18F3F9/ku9JmBYcvf5NS08+XbYef8k303gX6pXtYVxhrtjzO9vydsjYZqhF
XPkn2vod+VLJKk8qahh/gSYsnp2imZIP0sG1Phsjt7Q1NvfS6oayED2VJ3fe/yUpcQ1/+L7SpVVT
23wPDqOjMralKDwPG47AFYNqqOxxdYfJ+t/4FHYx4Vvot7pW9s9OrhDYoFlvyKMNA6CuhLq1AtjI
uUT6eMVA4mbq1jUihNB4kG1XSSftFKv11p/Ojq/XNCHyg3wjerlzESETFlQmdJnYthgN6LG/vNl3
8/lgjbahnaqg7KQNTCMgNyiFbG8MFOJkozBhRcydtRmgrA1P/PMrFlH9j6HKO1sU1fKcz/HzWl4j
hdF+FMszjh3YZ/so75uViVLvPKUIpTZLW94IoZdRFO8hoCVCfuB9KH0PEnOMVBdi6CKKEJYHh/3Y
lTZeSekxsISJU6Y2g1TZ8xvhX60z214P1jw0Ttw8fhk5PHuM71fT4xxJiQ1YVUnUHfDG4wik9zIn
pNHmXMy2lrctNnXJgO/Cknhskqg9R0Qs4Yz6h7IqJ2CF8cg0pgM8wzApVPvsJrmfq8lb414hXH1F
Etr4aqzB8zBK5aN0ESil/yJc1/y9XtINOy5SxKg8vTXqcZYC6aZ6Q2MAcD2KWaznwwRzAtjdYLJc
BZPJ/Tb14SE32VRFvFcCj4OSpbL3mTKxVN2eGO9nj4d0f5PBTnNrp4NNI//aU/FFh4yMiRP7dt1M
EwxNa+mX5au6Pi1BDsQg0QP+wv9rvfXzpt3eUDeQ4kLqejmfJi9YIuoB4cBKnjY6JI9kF3wbfL/A
Ebi6iQly/Ne8/7rH0/yWvfvBCFsS3/+vGaJVxS35UZKX/ak+28AsdtYuZbcVKIvzCsvWsudW9wWu
7L1nID6Nb+zoQGsNK1g2Ie7ZiHeBC9T+PLmbiq3jxpBaAkHZ+PNVI/siu8NYDWGk5Fgn0JzMRd2U
gcBK7YqazhBWj/9bgz5hrGq4qI7EBvqfpBAoEC/0p3ai561+p4Cf51GY0N4GEeiElSZ093xs5zRi
Vjvq91hd7FkS4MQRURrTWN24Yon8D1/5PDr6mm6K0Ve8EIwzs7ALyq04cNgqhgqaf+AiYozNuztW
9y35J4X9uctGiar18kbtTJRvDZ6lC7EJMdEfr8+6hrH45zEdyWo8rkPpZiw9Yq6O/1Pyn1sPEwhr
sy/phTZAJN5LBfiZvaTdxF4TOsHOU3S6gzqb/QaN/MfseBxS4VmmBAmRaGnWzoPgiH4hZbEGif+f
QGmMstUbVpkYKLzP1KcaqrPc4K8xHqTMQSDt3sQqHUKB6HGYQRusuXTw58vURIkYaznBWWSnzPWC
IrUSplcZ9DsNIYGNbHdqJpzrpKGUpzR/J48lh9tsgemjGlhbt42Ft84q6uM/DRueNnvJplDcMpu2
V/BLyGgxG1qWN4JgONny/ZKKodQG8Pzh4CSFabfwNEeA8fPk/76qzmglQ7b81siw5lMMusTKM9ur
br8J4vSdSPgtqjywRtSt9XJ8Z2CwHbhX28NTloH7R3tB3DcAANno/f+VVMG7/dl/MyGxdNHmmtTh
Rg81+uJGGWxcf5UGfTEQu4g1RoaDJvppRITmps0i6aqDkUaScdhfXq04OzKNEjjx/yHyrharphao
Mja1dufwNu2JsbTGTP+TvIInAPsrDVRyv5fInlJ1wC12D3Bemx1kdp0al5CC2QlmQbcEaWQUjKrJ
fNGPen6sjF3u0aiFEaHFNMAmbg7WrHmY9USPodJG8UEdLacQrC0lXFbpNlV05OnQqKPfi2tzi1Mj
ecdNEY1jDevKACRzAIK0DzC9MobqqPR4nthQid4YRp5E0XdpSgy/4w4jj2k6uU5RSmKalIIwsuiF
fARLjwoZWuz55MbejCejHUhUUU8fQjvfv02tqT3H4NFHpNO5TRIr4i53jwtvozJbhcVfh87PHLu/
D//bN2OeihEWmPsJVElPdrSaXp9k6Ed4S4PHnTWOWEa2BR3oXmhVpCjcHZIvvKgwn4hfGDiZor/s
Si0DX1TFLm1FqqgrC03R7N6qIX5JkHP2tQLNLw6aWj0wvXZnEnAsgWH1wTNC1HXAIoD3fNR6/slp
i1WgL+MhSK7FfwNIFV+XsocS4Kn7oyIAp5jw3mOi94PHRhRosKcXSOrWqlFbRjJc+5gWn6RAMUxV
AfSD5LoiaeBoWHrXrIIXsN/6WciFe/HnW7gb+TOP3kKu52ynlO2ZLrQS0rPrtXwWp9IM9FJKNFft
KJdOncWt+Xx1Gfe19pxVoLYYt0pzlImCpZZy2SkUj4u4O/Llhia6gzkWWg5Fq96WKsbIwxiBv9Jp
BoSzrB8cz52pxA==
`protect end_protected
