`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`protect data_block
UtZQi8paiBUOE4GhqcKFxvAqY2JsdQaylA3UqRff5zdDHXbYaMSWWCY343vWN3bLqfar+62Futze
B5+2F6v6vaxpx1T2SgEWG1qULht42HvReP41NGkXJtrU1TvPPndBv2jlc/omM7UzxaIWsXt3Y1EJ
dem+0KVf6Ah4JMDQcV6rlrYrfexQqGPa/aIF79RVUVvg0vF3psZZ4vjt8Ryg2IHvwnr1qPSCDreh
WwQ8iSzHIr/t8aQgC87z3WTBfehQMJzjsEh+lh7ye6eLFOGDiuLFrZJn4ZEaERuR03/r5w9YT8nQ
xosKtY++oAb2+8vA8oexF3By2ZEiloA3UABZBMGF88/ZXFPFl5sD4nW/IsNXaaommOsej7ZCxkcw
QCF5Zm2NA1y0Mw2mOM5Ddv1hVgy+VkCIWKzCZrBwk16ty13H7aKlIl9+Wz1GS7Q3LHXNP8F+gV7U
CTs+iiIzQp5WQQ1ErdStgCfu60GhBYyOZ5HCkFU7088ixsmmhqYSJbLwdrJRPM5bZafX9CtJbZf/
4P1TTVQraa/jDnifdsy4pF3YtKAp68tQGsEu6vtkwcxl2I7/oZVPYzu/7VkWQAg4BAUZMmD45m5w
ZgDfxT0fG8biVI+2h3zfXuKTTjJZkYGfaE4X6IRK/fNh0285OScOFQIMU9Dzpymoy34PKNzmljCe
pH00mBOcdEFPnSUXrxNqDkBPEGGDr+069j8aJKfPMAekHCVTyKUY6PoaGvE6rQhNYIN8UYgrKtFB
3peER+Ejv4ptO6zF2U8Lw3UcX/NbyCjOTjj9ii4zHwKRQjwwBKJ1COyNWZn+3ldVDYfrYst6KqJs
hDRbeJyQ58b0aQjvfauNn/OMZLoIeC5Eb2mbdkuJ4bv25EHDQyK+caqm6kpEWOc5P0rFVLYrmMOk
glX3mPVwB6LFZNcIOngAzpAlCgEACv7NHJHI073heszEEg0sLiJbcwfJlRg4mf39sNiFtUthMbUY
0Ip7+WYNk1zr2WftgvmShE6/3JjsuSbOZaZxAAGR/Fas/ipygNXTe2dyMleIgFnc7sLGw4znAGqa
pSbKQFG9jm9nwXoTAVtc/YecY/8F457eXx3T0SQG3VfKDd8IWZIcajv7S+fwAkC4e54PzXmDjhVf
YHOgo65ZnQ0UmaR/8ov0IRqdhwi/Zl2fr/wwXeg2lMcTid49ZuF97S2tlu7Ay5fVJ3r66xIZYVbE
9U9slEgVHJedSSONJMovc2oxSleBL8a1d7/f3ec431Ev8cT2H7MMU9Epd6I9VK1DUGr+/PunZVOL
PySR9e6Wrlp9piNmtY08DMpS7Yy6wCu1g/Y5EUCZGz1s42a06r5kmMNwWsh5PTBdx+yg7kC9CiLV
Uq+Xk99lOdq9IZ7v+RLQRXfnCkmD6elhackt+EL/6uN4yxR2yixvSef05Ejb786d5Ch/10Fb+sY2
bbYBzfnKzmYA6TtgfK/rWCYZ4SXa5JnTKoSZMP/lJWRf4tJbgcwJsXczOXuXjqjpbFXedeUEkHa4
WV8LLnQKA5A0yrljS7lIT+L1nCf+XrnDoKaY9DnZfKSeSxGb+Nx0G8tnoLVrIoyIvCv7g9S0AhVb
SrqL4r5p19RSbpO7fiauLmwFYxj2vlubfBY9enZMiDKNyLpNWhk3rNfQVIMAGUTtagDCRY4kUM/p
FlOW+D5+71AFU5KQPmfDesXWoM0EGiOVnupv4BXNVCvw4jg0QFClEOH51sIg1Q8RGEubrB/xseJM
U2Yv+Ja0kXFMrOkcGkpjKOZLGS7WXzYoFVHS2gxIgXZIs1HtJ0Nw3s+exZKLMEt+L1/PTjD3sk8y
53ATpbZze8xw7JH0WXc0P7AMcXvNMBcVByNFoRZ1U4p8Cr+4h+r1MoPmjLx05DqvLbYVjSh/zcwH
1xkTkriYHu6eGAjUkwNdVZ7JPKLhyt3BDNskH20CDLiwEpmjwCFwNvk+aPcJks4hEMUdm+nPqj0M
eG72CC0oPVu5fbf4BpS2b4uYtRp2NZZCZKW7tIY53Er+qzVf35bDLSNaSml+C/PNczpNygqHm5iJ
honCDbpD9GcXy1XIP5fhFGLCR5Uyf2DqqpLVgrTvXcP4vhXIqw8TRY2EFhCU1G2ZzW0Duwp8WWqB
5Mmp5ShiEgfZ+wfxdYqb6Zo7wdeOq+OUTU8bHwiz1KqT/99h/k1zruFDSvFcS5Y7br1u5FCcM0SE
GcNJjzee6Ref1VBovtd+zG/cv5P+mhTfsr6ga8SpZ2Bl/DULqkyKkDgkocSFXAl+jYCR8VkSXRa6
CmMR8/J1ToA+4cRYmeXFD2LfBgANDDhr0VL96vARC8eL8jaUgnqp7NOkUD52kmZsqnPKcCqUJ6dA
ibP0I1xVri2HgEAOWq7j3qKAqfFP9D1vEmwA84xth/h+MD7GHLzorN7yRqcBwOtVpZQTWGvj/9d8
8C3efvdfeU94MqWZHhWFQQBxSHTmu18l2Aijlu7WUPtZE0h0UPGeYHN9kkqJVwKLJySuvKf294Pt
7f3fUVdlBuqLY13qZe2i7K8KdKzDF1AqFTocCc4NoSLChLj929QVaL8NEld1qDciE2Vegzx+o3Du
717mnrwD7UVj4v8Ep41okIpRfVThTHbEFX+RUiv53UIgc8aS8uFKptGlfSnVuMkwUCEcEmrkOOIW
WaI4nzN0TRGocLMwkVcEDf3R6Cpgpra+stYUNW1FxljmE6r4sb7aWu7KSSacZqVt5vNht/wVmXAu
rKm8Mm3kszEwYN3FsV0Jo+jrNmw0vx3LB8FXcPCmk0sa+23gbnYiSPRrFxfftsacm6uuf+bonoMG
pYWBU5G0ITXFy1NABC0zxV0I4s6ABbIf8ivnPENp0bsT+SZm0WtejBeYfjhv2Pe4MBvdGIw58XsY
u8x9YwXUS+xr3Q5RlQTFtuL+V8j6F/9N+Gy/t8cI2PD9PWrQFuRZwP0E4dKh7lKmnHYOSdREoVCk
LLKEpb5xjR5OmRryDWaocXR4esNhzf4ykNBDDD1lXCIfmPonkSQBcZMYAdUZlHpB6Bt5dAPzIOgH
fwEIJrrqXtB3JnLHm7Mw3qbwp9dXiPAC4ib4X7/K7UfWwEN9uGfc2SynzB4gPQ65dUHlAoLXuYfw
w0VgKEiO665GIaF0lYn4l42WzfAQoBBfBZZq8v4iFA==
`protect end_protected
