XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����m/�s�r�����4By���Nb���v����p�O\7<�$8�@d�j��EV�:%����>!-�i�M�;�����^	\F����?z��r@oE�@��1�[䂦�.�x� �J|�:�4�.�`8����ꏾ̔�t6�qQ�[�[�]u���<�M�kJ��pu�ve��4
�r�����ia@�������|ݰ@�^�!��8�H;�ܸ+vm��~G���o�N��>�����e�d�o����Ui���#�U��iV���������Utp�F1٭K1��N�/���+��8P�w�����>`Է9j#L�B��V>U,d��T�n�8J
�呣�Q�R�e������a[��`�1���禍]Odc�8Q.�3�"������qs$x߭��T�f��Z�A��4Dz#]�)�3_���X���&��Zx���n�����l�����E�hޚ	�0=l��߮�(���.��/��B�-��f�j�UF
�%N���^b4�ѓI<�����U���O�(k
5��pӅh���pt��W�l 3r���)i��+�P��?�0�=	����E��B�j���������>�B���'�y^��5�&K�W��C���Z��b�O��J%?���ֽ�d$��c{���q��^2x����g�ʈ]��־�e���|��4-*�Y:wއN<���+'�1Gs���a4>(p�*�ȋM��q����
�tDa,8�V~�F��_�U ���l���������tOӝ7ŚF	XlxVHYEB     400     1e0�p�'�p���Pw.W�0闚ᜑ��fmx��'�ms��9��;~���V�o��Xf��c����2�jbUe]�B�.��Z��>fm2�i�� ���r��Y'�U�$�Uܜ':,2`\�UTѽ���d4���=��J5C�t�q�j�����Hʇ���/���9!<VbM2��!C�Zɪx�dn�|*�W�$N���,��pl�k�q�H�ָ"�K�p^~T�}A��?���&UX�|�l&���\D�k�n�8vXo$�P�݄��\�4��#��7�'�Q���D�~���؂�$'���/�J�|ހ����g����G*�X��i���V<-=}�YhT���e��)�q%�Q�ʗc��T��d:@k&e�����H��$ DP��uW4N8���'�dF��q,k����^�X��c31��M���@�$5m�܄�U�A��uF�b����.92���䞁*�bzSXlxVHYEB     400     160�z��t��;>D���6䖢g@>l����m�ad�������M6۞�)��G���yx�&��B�1�
��Y�W�`����X�K���eNc�&:U�������z��iM��ҭ�
�yn^UD�����������R]y뒗�Pk>��{���Bi7��>O�^�&��V쮞�PO`�@��{E�/K�o8jc�8D�Z��k�
$ u@P���������oG՚Q�F[�b����Oa;�M	j��-ڈ�|!s�L)"
E �*BmɄ�ޙ8���pj�Q��p�B�S&~�M�mϊ��,�efoܘ��˧o��N6�#	���#�]�|1O���W�?��	b&F�XlxVHYEB      50      50�:*a��"S�&�˫R��c1S~�e)K��7�v�㪄���E}�vZ'��|�q#�&㌖��yk��>���$����-