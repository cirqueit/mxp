`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9152)
`protect data_block
97enig4e6/+P430MiOnZAuPHXKHBnbfWTspKRKIkQnTYq+145DHdNqHCsyaFaXdngWxjJP8nkWMw
cuiyvZh7L71yfoA+Of2sEsXbzE0xH0puxCBImO2hvk+pprdkLjKC1E2Z06ffh9JM03TRJfmylRGr
TKgCcM5bEwCyR83Xh3rb+0Zrjuzf1lODUoOKWx56nhESbY+9dZOod9peAHpBRCiuapfNih5fDUyl
6TwQY8+YxvNVxy9hHpbh1Ro7+cQE1O+C2VRTgLBE2FDouhsA8SwubxBKRSCMU2i+PyaLrj7xa4Gw
D/Ht5g1NX+dU3S6dEKMYzCycs7evRSPQYENmypaq8qAuJecdnInF89gS5RmoqnxOz/5PgrCvkIvc
+fVy6H7xk6p2neS1BZTsJkBrqRb8hjfWkCyvZdy/tDZ9g1EI2yE/HYH0GoAYCfWWKNWDjsSxhGVc
IwGV5jahXeiyCGlF2LDg3xDwrVe9SUv8KvdLyLK+Pjppvf2WxTYKPPtdGwy6+XHpbDGYfjB/UMVj
X4hRuY+AoS7XdNT/y/zfwKY/2QsA8UKJEjDUS7HbvUVrNfZKlDoLW1/AUAtqmBD/SE8EcafqY/fy
aVUwC069ZkUn7MUcd00BXM5p8WgFpGXmVaT5NFfFt6UagQOwsvnhzde7ijWYFhRrzMHvD+/8QGma
/DEwZ56D9wxsc418TQotdcO+HimBHzDRrbKfe7yzJDqHtSMRhg5jKE/Jo9GdpjyhSid3aez8VOUC
AzSHwCVqqcQ0ojWV2GP5rwPVmizF7FOqj4XngAjOzKR7e1tRSHGD9sU+R0RQ7Ugbde/EQ1KF5fUM
k9qgpV/O1Dkx60IrpEhQAnSB6hMVmyxeMmaTgqkqruiziSmn+Bs4sqSs1MfrgBfAt7Ewi/bGNDIi
v/iXQcOFux00x+MewKT/UuPtm0FxfDpgHAwnJ2Lp1Tx1jJ0D7yDfKgm03WGkrrZ5x6fXRm+l2N9c
RzI/eZYUVKYVR7PXFgesRO5Z9qJKGZM3a0pfxXcFz6N6v8xr3dlpoICFGjgtxNu7wlG2kkIihrMT
IH4JCQvSHxSyUiJU7Ls73e372FK0QgMiVo72Bqvo6tAsHnhrCrFNe4I6ejAmcd51Ll6Uy9NZdqNl
8PGJuGTYKknZiovUFXMnQ9Sopv7RXDkQQXWdJmpZ8n2yRgjF1OMXzuBpqPr91qyGEhEVFlO3HSHH
OTP+M/QKtj7p+F3/gj1bCLYU1QcYqSwdO0fL+pSancbwbsNTi9gKLgKSZahpbwES2hW6wOyIEAtO
p7DKZ5MeS5wnJgrvIaRWWJcCZ1J/UtLT3Q60mDSQ1DKrqMsLbUjnKsKkISq83Jvxp6Nu2/lL5SnL
Xmq+haTVOfXT9j7WRnHTmlcLoKYKBB3eAXkQRonmvPdz6LE1Yd/sbfZye24HJ9i0XMRNbGUURRBL
CYc90hPqTpApAt+QgMo69CBge6Nyemx7qomiI0v+vDVnG6PvJ6NH8YzEuaL5yinNgF17tMJeG3nm
eX/JLKVfT/yMBRF/BHMFtLjd5SEy7jX/vTYPu6HqMYAHgw5+vnMyjIqELnLo3UN5Tqvb0ESnImlA
GGMnY8IDCVYrwmD478OQ+EtgndbeYrZEw4i/ExGixrkIWOHpCNgQuqWg8tpSTOtcvvoks9+rtV07
6aNP0swEEkoZE4I1AvrSoPKpECEytooY8SVNBxMGZTlpGmyt56E4gTuKVaWp4pfuOvXI2Y+IbLrZ
W/ngKT+mW0OTCIuAHsMPIW5kdlEiGjjPtwbJLpj7/4fQVEgRBNcLQnr5RTW9KgUdIHb2GUgQy4DD
/Df8+RdUU/VsHb8tQF5dXVzZAWJN5nmp99FWIlnMzH3vvLUM2TcvBAJaOx0IwUV7QpJqKnsd/x3e
aT4iy6lgx57iIsZnBMd+rzR9Nd6odD2yYcg7pzCQVhPeRc2rqlYyZhn5yhgBTd+PF6Z1ZwOcYPxE
56Jj3pVUZlGsoj+3+ETDc8k121vyiDvYgyy0mkaZm2Stj3I0nrAkGgifS4ixbo7vf8MbTkpte+k4
GoOXuREZtlyNDqy2joTLmyZC8Q72VEU8Yvh7gG53atev+T0jEQopQ0Yx8GHnlS7na6nmWr6KQjL1
iHqsNpk8bNWaMoAdn3yW9HohpjdIXiSLFUzFadk86mRbc2zbkGl1NkOnuCtWgyiYrcrZ56+GE4xw
9qsUbtEY97ivQSe0kRfW6qSeTPAh1m5GHyLSeerb7QXaPx+r+Rtbn77CRnc8FvBx6ZLi1WxIN9a0
W4AwfdOqWRlwjOhN9SZJKtn0JFRZJu7TmuUv5LPGpaUanGC6yunGu/+mE8tpHLaIAAc9aSlDVV/6
NMrgeb+pa6/4Rr1HW9yLeXlhAPKe/uC3ONFX2kONba7l5r+eeb7Vx10kTKU+ZhlITu8qO7e/RAsY
B/DO3inT0J1Ea/VwGjLeRk7PPRfEsuNi3/YwpWGQ81qXSAltq+Q87e9dnmrGVw95E1Ao5IT9T4Cb
Sy4ATpT1Ua1pIQlslr9hOi4IKgKdxNUbahvaPXkqIvSbIqAy6hOj0NfMzTdWwddsLtJdFtY6JMGg
d2CaXsEirLXxH/PwYceUPDogjd2K1WJGK1uamzSUpp02P+idcgXra9D3pxKAZhfJP85pv8w70rZ/
xsdDBsQtyyITSsgOEdQDeQ+Cm0Dr2FQFgTqT0PrMDpNlju55KapzlhUpx/7NnjW5QK9xc9UZs24C
JTs/ZD/AV9w7X95R6Ra2K21yDMk3s82nS+00FHzkrbTv4oSsEPntTrStOErDXVgQAyj9zm7fUN0p
o0IMn28mkBUKRAXKZ47duSeDsboTMLYj9lDSPAh0PmUg3ssMADJzXOE/IjQCsWPquVWfEyWD5KYj
+OuVZ5yDiTTQHKu65kmeMHJA5MSGyArrIhgclUC84/oIYJjlAVX8LvLIudoYVc4TQnL+p+DIN5dZ
zOd6hvVMtBU9uoU4/cuMlEEg7Ort8ke7xA4qyQzvg9eNXxmk3Gb/flAhlzoYWpynhuN2ukWoLNmd
VNDSkOPgob2F0K0bJobAEGyxKam+nn3XykRGzDcoYe9FQQIvlfjiyL14O8DhKtvO5QBssZJt1gPU
gjN16G5n51H/U5xFyM6szE2k2Iy82Syj4GvyU85k2IueubmIAi7zVEj31tCLEwBdgbmth9Bg0fQ8
U8qIcGlZ6G08NRvRGCMaryafsU9Y7n8ksOYOqJmjOx9v+SiQfcvk/2cyD1V7FknIkwjs6HjU7b31
Gt/OxsQl9bMs6gnl8b8JR7dmP6g09yLYaFyB+3bHvWC+AK+x/emXbRI6sBkU3NQNFHhHEX8qRfsq
gXiGKQK6EYn4jtbzeiP1JrG1N1P5G3zMwKY8skhQb1h1kg3MAEtBHy0VkyuEH5D74UECWTScvFKC
dua9+FNjA+wbMbrLM+2mVMbXewdNCDO0hH6UuHN2eTxHPExeu7mZ7q+A1JESzhHp2cPLnJ4SNtoF
pTVHhob+1JrIEqdUREYSxKL0tMnNT5zdcXb/df+t1SOTNNL+OKcHdfPpBRq3wJ8BZYIPwK+mRdWy
xdbS/U0t0m4vomPSJZk9QFJK1CFutDc6WXlIGBATRlWBmtrIoIzXlVD3SfVF4jPbeAtNBpDZBIRJ
sQC4lGUrvbr4K5Y3KQbcDecD3U++JzpE0t1y38slCmliGYSCXsXbT3VzSdCR6eYsk4ztodkO+MKJ
Dc96bI5RjPGWDcpLo1GreylVA6WTFS1pygt49qImkX8+AjIqhoPgckOvnYT2AeTzPK9hFM9H1m/M
t86Dz68mzvBrDJItTqXAx8aNNyCnNQ55dSaXQ4aUDPVa1W/QVeGyern4y+6eMx61yDv/KeyxiiVT
2azAuiRBrwwhptuBLTDqt0pPLeoJr0HwUyUfTTE88m/d8NbuCXjljTVruRZiFyxlpo2wzkX5Cifb
UjfiS4D0u6gwIS6mBGwlfVebUb8ueOlJUt3b2uhLI4oEJt4/UEqDWUyB/mggQag8KlMTb/eJoAae
sP2nJeYqmnYXptiA2eI4Dog9zO3JcWWDC+QWfjJE4s6WNfZyp1LGDEQdx4WLe557wxEZ5Dtm9Q3W
ARkBWaEUIaQcaOPGHDGs/eM8aLbQ7jq0ienEXK3dLOABOKTzr7tDOgiv43wl5G7x5EYoFXq/yVgV
08m8D3Nqmv+4PSnAjWwqtuQlxKlkalOF9RlSs07FzdjRIasvbwu/rbyMcYX+bUXt6kY0io7nBPaE
YQVvaPmvIaKWTuB+BsP3irDaw6bwZFUAC8BKiQ3IICeZ0usSg9LP3/soqu51HHsFF37ugM0Xu7rl
cPRZfGOVk0zRfacR6HQ7oZJGuJooKsScjqI4H/3F1ntr5g3lg8ThW9ZEQ3zdxkFrdUvCjWAZlZka
L0t8wZWCs4pNtqnXrjp+H/c6l5wcZ5hiVWpWYp6Uocoz1EpuXVsRdZJoz1Q2oKcHRnX2qK08XgAg
0hX9ANnwCMKzH4+fpk48oZ+HhPfn7omEM00owa+zfVGX5QOuX2T+W1Lkot4TgjZuuw/GzbJXch4E
zqpqQDvXmnxQRYSGwBdJ5kqyZry+BGZb5QRiIkNCq/Oe8fIiCBp3mg1oYvSUt3S40BN8uir/iRtG
NIK/kMXyLZW27yWCemos7HFQzAodrxrq8njQLN8Ma4z7kjgg+XpXqm2/tlfMWWhzX1kPuwamY3LX
1cU5205WDs9Bd65wtfnDLG0a1kOhZY2buSwu6paBPhI55m5CECTNsoO3MSRBueqsoXA0rCOV19Ps
YweqyRGq/RS4hCVAZswlvlBod3I+bfreU4uf85HOYtNrzKRXV7i3whdlYWo+/jxxjFedMJdik+bg
weV1S6CJHjKaYamddtrnHqi/UXphMQHGE2/qzt/Ukrajw6FKTuQwq4i7kVLVv0eNhwHM0QcPNCQw
unzfx0frV5ZGquzBIMm/PGf8xgH8eXjxhfy+09DIa/suw6+c9XSLs8OOeeDYdrxCGnSEuGqzm5KV
stwDe2kQveUweloi8ZR4xkwnMwuwFRzblf7FNvWFMmYcMCMsKCQnss84PvHmUNnvtEbViA8bHKLi
7uTBS2WRkCAODNu5qEdz3wby4VtlGkQnApmOQezEJ1LViLo89wEcs2KxLtPSmAk4R9lunwqvynJ+
mzQNmGoYEm08zajMD7ZG5j1chBpvSOxa8eLx2lWXwDSrGyd7VJYvkwUG02DFpS/OAMnTU2PiBZNC
48UhVrlb7gXkGf0xyj/eRi0Otghxo4K8b2+Y9yioh8kgDSox5b3duT1fANut0X7EPMW42/reOgin
7aEunZolInTiU3m4qnsAtOrsp3iW8zQzkRrc9ka4b5fMxGk/32TZ8K3uKnjOulYX5dBadcwjKmMd
oJQUdlMrJ5czitgewpaNTOe8ZyuuTLQm5jTV7gIMHiMMK0ljxKEhZ3IPOzsS+9E9vXp2s4yVle33
e1YF3AkshqonKyEa+SCVoHFyAOuIl6KwiF1xr5gsSiiMmBRsEKMZGAfn93EElTgBF3T1lkf1yjg2
No77YZhCkcq1M3ykDf3QYhzb8K940nFCbDSTlY0C7KY+Zw+x9Af43bHAHtONdfe9B0s5yGwtMPlc
OdoizCZ5UPI8ulR1NJAGa2GjrucHGJlXsJzk3NWYjay0DBsMiXom7psuX7QoDOXI7TcDipy2TPpf
yKYnRxe7GtZc9IzNNSx9SHKE5BX17hURzExzaCDYD3E4jHfLinPUpmZz66/A7LP40O+pwjtg+xlI
XTCaRi9OfdqUlLi6k6UWAZgOo+UVaWWQLGgPowHmTo9eq4FOsvl3dMPFXfbU1xpNpNolItxVrfqX
eF/Uk9qsMfODMRQgz75HXx7NubgumVzHmd6GvTNqqQtTu2GCUcjM2vznsth2Bj6KMjXdj23NG+q6
t6vQKrIKpNWGFa+QRWo7lTpx1x4hK6dNu9fhkzadytKDw6yB4R3tC3X/U04omjEyprnYhga8tiSV
X5TTFHNPYlwAOSC+RiOy3uZeh1bNPz2usf6hlZ2E0h9eQpujyuEgQiPMOKXLV4jq/FElx0MYhKYz
jaBUzSlMu6cLaqnOa+gQa3uieTrjAak+IoYqcS+i68NcN3CtrHAcgWYTpAgpoGoOiOuNAVB4phML
NCRAXxP3LeEtVaiqcVLC9olXhSXgEcTzfVhrdM2T6w4zRnQyymXp0BKpU22NPosHV6+QeXKyeohi
sghkfXvXRcBGLPa6wfFPISbWYHGF5PvRS4oUm2hKi/5pyMDc8YcjG39cxiDQD/oHdLialhuFBBc2
ZEHx1ZE1GL9SlbV4MbnlTSv5s3K7+VVAxIICXHlvJU+TwN7Q9ljg66gTvjs63rkxJ2KEIRsPA9pj
2CrG9d/Z/MYtNHFx9Q/0ljztAQdea+ExKYr+uCSVZDKPh8veCl1eJSNspg99c7RnJMvQiIoVnrhn
xK2V5zRXupiYe0F9Wk7qtpYPUPRDPet8SMbjx2TPuxd3xTXjffZa5T/ytvONFRKfK2ArHcMByoMS
/vly5Q/ktlznKJIl5gSyKQz3FkN/w3uyN3w0grH7C0DysKmHiQMDcXqR4oVgUSsdx4Pr/LV15S2p
bfUnkfuybSrC9pmAO1sJqppGloTRxVYFufMp69qv9HhXguZMMK7ttycA5Hxn56YXCckjPLw+j9YH
QhTnhsMWj0yl4wpKuDQDhN15nC/gM2GrUBzMNs8dqG2Fp3HbE0TM/436B6WUJRdbwGeTMaLzFae4
EfjugLIjzR3yGKXi3CNnBo9IKWWWQ8bELHL5nrNY3ScSwPyTYHSgUbDSfvpit/+kxQoQiy1u3S4T
hFQh4dKXuE10rTzZEUkGkpmAXu6EbbirZPSpRiTtkz/tTwyVi/e6vfddTAyV1f5Et8Inndqq76Y+
aG6ZKAYqCdP9hMA20ihvcV0wuOBN5ZMQz3ggKui/NHyeVv6Nvb86QV5QrHem7RKQhwXvNi/Dgpbp
G26QndUrps/jHO7Uqz5rRblTN0PDOb9aBNhMMOM0GG8dDze9v6xNewM28KsxfEv1DG4ZGyQ7K3y9
hWZdNnItShF+AjukajtioJphfWxk0XVECzqcUxvg6IIVnRgOWBlrCJ9h/f1hiPdT+w5YRrVz4dRd
1VEEyEYz6qoIuh/VH8v9o+A14sxCgrcZY18ToysT5HUrT7QxbkLpNybSprxypmozkEoZX+yg2G2J
Bx/XH+0KSzqwo/kbqdk6nHGsPF69/uRGqkEGSRI0FF5MMO4uzIUdO3OJX7SGUr8zEf6RwXHriSbb
cgRf3Dzx/9ewrLOc+Z4RAGVvQCH68sURFt97fbnVAjpyrHc9ItjgOqXxMzNpHH99nHZUfHyOgAVo
h9G69FM32jnXpCJe1k0OmfSfpJtoo6E4fD86giUjzT+wbRTVDF6hpxzY3SP9eXjZjgske7npOFhz
RkyzCHeapMyK28NapVIh1e5jYoC+OdB7sKCQtAxj3oHuUdJ7FuvJZA6rZX97SAmd2Z9rKFUVlLOD
HNg0/gntS0F1basdP/fNo+tCYxyHyD/usX6nBwdvaW4j4yl77WjOGbDRQBnBADLYGam+X3FmQPpl
1NVd3gE1gMtIo7Wr16qdOigFmOTyZ6Jim7fkLj5M3M7U0pBT2P8c9JYW7r7JA9bER9TUYTAFvMwn
i8drGUepRJeju83NgUvCyt4DrFclflwfm6WIsuhW07reis6QXpwaSrlK9yG58k+IE+yTgx413/f7
BI7jefIrd7i27V0jkEZwH9zjLqABtq3Hp5tGpQlOFJb2jGqq9cqGIa73no7wlokaIQxv7gP2dmBL
emPFoSsikxdqJCoibEfZcwwIoyLYW/oeeu1aL+B6cxeQAFos3QFLrwBimiQ9cuJVTp8qRoQMdApi
bPCD3JfL8p1CQ29s2NZQbMTUE2SRE6gNbLjD+0xKSxJTc5ZQJmlaTrj/dDfgczJLAZHEVLXZJ0Rr
uvjlSR0V0P5kfbDH/4JaHYpj/qNFuQT9jbPovKAYNxKBA0IGuRHsZ0Wr0J4l4/mjr/Hdxmcxpd8j
030sc8H3TTAjzvvokP4NiuQMKVzsHFcHfEc2zlnMm8yxM9rBdTOqbz4dLQZ3mu4gVeLUdO39N3LY
+fZrn7hmLvvc2ChwHosYlYrBlrZ/vZVsvVDRTlBNEruw/JiOToBgR8H10j7HYSV4QrYNDJw8Ln/c
cw+VNXWweB2lp61ujl/+phuF7rWJhwDe2TwaQFpf3+2VC8D6ScsEERWdvAtBaqH15YTWI/Mw9nwu
P02pMzaj++BTQejCAo5DNLMOk94qIt34QmH8IUb0UsPtnqJnvIIbo5uh4YQennhpNslAKmdflfbs
OhHqtVIWDL/JJBG0qR6pYIoGaPTAK50sI/5MkYAHmPwCKGlcvYWaWVp3rIPVsaC60z8vUSjKtFQe
zWCMovYqSwQcIo/cok0+hZF8TKcqyC8Hf29XB6+h2gf9x/dg3iQ0RFWzae4o+AE1sjL/8qgei6aw
T92LYhPFPh2BhPfx+wLCV11crXvS/OT+2Zov/H2TSJv7vi+RLhyNN4a/G6oQq9429UJkD6RB/74g
SOpiy9a2W1Xph1+zv8foo+12Jmrs7D1D4rrCzds3unQgDd1NvHWdx0m0oumWFJWCZNbyZoM1JhIl
WWJA7vNpTELo16pSqPWB2BexZIogkMH/i7Lqh6UR5m+N/EdED58jt1etYfnWpTxIZkxepnNib5ZC
mZIypufijKNqj72dQ2IfT+ashGdvSDu/IoB04blAdNOtgTAUA+O74oci2AN4wLOYK894WTGbfK4/
eTsrH+WAHUA03TDcEKrywP/Siqh6UKzglzv0HGJom7m8ZGUUA6K2iuNJ6lRP5N7DAMSO22XFljUi
R5hsZnnUPbupaFrTuyXqim0Dcl8wUtfi+bPHcjHxPPs9nIV3EV77FOkkd4/eaQG9UH2gKpMNsVGd
7m7YLlkfgEuyWV1AdLPgwzWnIFiiUE9gDgpSkLHRRHVVw9EnB9PYTBVTtAEGxdsj3Fe4cvRaRfI3
UbcJfYUYa9DcgDIBqaHHxGzrs9a2/vZNhdUVaR9KQRNWHcdroWRqKLiAzn61cOcsyGAAyeBhaaF7
jLfQ36l2G+83jzwNBygPxifDURGIQFoowGs/y2kPofBgsm3W2o96OigmlEoCW4FAbQ/iR1oshduU
Ecf6PG5aWvAxMYbBy86mnhDYwCwVem+IbbPiQQGc3gUUS+kqwZK6j9R8HzOKYiV1B8cUiWx6N27i
UPYv+/CekGOIBSDE51S0r7Vjo85jvO6RDHsr5Yofx8DupUPXnuF1x3R1UNCRGLsKaQ8dwb8hZPTq
fyBZGW+4FEuZUosf3EODHuQxZIUpuCkYRCauhd/1vaxIHaTSJjUVMdhPeK8GRdZkmf0BSHa0l2Xj
te/TahGqIYmLdho+5hLY7zCCtHySdckmq0u89NC+FNh2ioAHD2SQeW8XG+sYnvPtpArj7GreM9om
MSZwuI6s9StHn8twFeeSggesGsmDOU5YBoloTqv8bOTFf9G7E+f3VyRdClBsOGg6hJkyu26pHoWq
A3IzJ+OsiIX1fs1bzqfBTrOX1bb40J6Remqs49MCZYKvLj5rYDVHTBbu0E+UOHvAKCoJez6ARN9l
8xBjO6HrFfZTzcEm6kN5P4nXnCRRFg4ByjgKcD4WAk0Ylr5+Z91Uv0z8ptxTOaosyc/qyfUl1tl+
Kv3DeUf9hHiGMI5173ULJct4lBCaFnRccIOEbJYXcoGWP5mUxPVo/QSD5B2AkInJqXQruWKXV+5A
NRDZkM+tsQKYRLbKQo3W11NuS1SoqqnZYUWzfReZmo/pyOqq6FPIlDVUG8w6SGD9EdWn27wjejUm
enWZpdiA/QVhfWVp1a+Q+XngGg6BIPxGQPgrUytWmmSdxO15cyQYXN5CxxG0s0WPQQD7uNeyvrpf
Zh577kH80kFIDIS83XPLTlnOMhGvxL5Ja86yY4UFlQQcDx+jIelJ3hgsm2BuXB43SlKDDCnEGiBS
O+yDd4WSEni/yRMJOqkVg5o/g3UseUp7VqNFA8qJHKKo6G/9bgHm7sKSjxrCV98nVtfj0Vhzdyrn
WzAoSF2K5uiEqklrYKD9I2p2k3uu9/ibji5GmPry+kQeQqQeHqMbA1Vc+3adD92IcqROZpFrepXn
Fop8pxIb0G5rviN1f6kZRj4EAJ9hQAdvjbR3CzoOoaI/8cdEBlXnSJHxytdNh/ijI42wOahfx225
tmhNSLsuIFETK91ZiayrKxnuIf34Q3CSX/Hsd/ohBi1kbipfOlOIyLC+5AJN8Vqvzc5coqUCuN7x
PoNcymBqMuuLmsT0M+Rvt+lGyT4a+0ynbVrcHZPMwToHZqU/66IKrJ0wvifnuWVIhVGuLC/PDqop
QSDl2hI5YbLQcYSTf9wdCXC4HX+zEW5DQBtIg+s8Sm86iUvt58h3uubMK7qnPijbeayu+gX7JAsn
JyMDopNu5vDb9c2/4me9wg7VmMkpEyInxXWjjKGG35ntZGzTD4Yx9X1/Nxqe3vMslugzeUP0kg8W
I4JQ4SmGo02sgxIsqcC8wnhWxtHAadltnWpwlYdao/dOBp91GTpAH+Gw0gV4Inkk0vh8pIntkjbh
bydl/+R2K6XmpryUp3+exL6wuHc9TkURYIbMwjvTENVraGeUzLaNmmMO8ycgkmgGRNo38VQLePe1
g8xdCNnn+XUXfDoBFrP55MLPIZ6/fJAvWA7Z/saawIA/CsaIq3rGcYWV/GQgmpZ79XnDQt3G/L4Z
XHZJBbfXeeQT6MZZstj260Fo1aBBPiYwjm51clSKGODUAcBZbvTK32jsy+EZl3GUxZ+vIThdeXsd
FPOUOZBPmBP3T37NMaqKsU0Llef88/3LYpJvr/Kuf8hHGOnR4pH1N6UTXuuSWfCyFXfouDDG0vi5
bB1Y3w28BX5i3GZD9+UGaXp6FxhikrWnjOJBlsDjlulUu2oQedNmTmmwtChswW086c/H/QV1vLHr
FPYdEYRXU5+4ua9MN0WPZISNru6njqUyHM+q+3pMrqDhRyn4/3WMc3nnFU0nBPx1uYTmPD13jy1L
lWm3ae9JjShCnSxdH1M79s4MLbUqM5qf1fFY8q824AbA5Oor8m4o5xFYKknKFS+87AVLR/hOpkKh
mqfSLTG+OUrJhoXRY/PbKhzCaeOu/4u8bYaeuZ+wBlWvWguMRJNWJZ4+SEFY4vBDWc6UjBBt9H2W
oBS6jVIEAbtOrHGRTnE2N/rLFKEETlj6ENu0JNuQth8FiPCcjqg1YrvEoJHYE1JZQx/CjudcG/6J
Fo5e7EEZ9/uTBCFWeqk9wf3yWC23/spCj5MNr4QRj/KMlPCRRWLr665+hbtoHJLm6CAVPflFxHIH
CJ872D3Z7eKrtmhAX+F1sPbl2DNOepoE3eJAtHlMMg7lQX44FHWGDvORRdj6xUHsKW3AdBZlHCww
Rw8Z7O9sACJUjPPdps73injxj7CiXuC3YKxMcp6AIvrvV+BObt+t12qCis1aZTgV5FRfDrUm0Bf+
Ix+l8J5jZLDf2NXjt0n+Q9Io8dUc0fB/QBh6Ao65b6DHZHKCOrcUZwGNXrx3cfXXHo4GwXiy4xsy
3WZHr37/TnMBBREGLVVoVEZ9O+SRGe5/apmsmy+S+ncKLGiQdObMidABNMYqSxEN45RUQEd3eRAz
qqbIAl7fnHf+6XwDzJOmqXeGO7Ig0bXUO/YPCJEV1zCQ3b3wvWpfm9kHRqFaTCdWhuikmF+YhRm/
Tgi+HRPE1H81p5LwnpaSLjUwmMiBrnK1YRTvLzPgvrzlaS1JgepFXKN0FbPN/ikLrgiepLpHt1in
KIcDUo3KzDEum7+xSJwNa1UnwsrRX8+a/Thzk7QhN4UjFEVnsXQtB1ERHy0kVtvJPN8LnqJjHJqG
d40E7raOybvgVvrcDkCtjwblEGgwn4u8rOhD7aU7DbQWdg5bv2DKSDteHX0vaPEYFWfUaKS4KRq/
ZmZowv3yq6IDRRL0+/WBaATu3mFznEZaJTCcQPp9baVJ5REle6xiEndjgvmnBuBWM5EFFIEEHKWp
2nvchFJwLszkET6YbfnN25mDYMlCKKKdRld72MyJqNGjBhe3mk2oA8DvxhQybxSpfU+kzBfocr1o
u0ZRhivBpeiw+GW2Lo/t83IUrbR5tq5dVxBLPS+Ha+8=
`protect end_protected
