��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���ၰ�~HV�%h�G^N!����X@���\�i	��3IA��B䔹ܖIK�=6�⩇܍�����8Y��Vg���Rt�9T��������ig���x^_w��eȣ�׹rkt ??6�2�J��lXO��f�P����A��s�#�:�Ԟzr#���<�8#�^V��XI�)��jr��AE-�U�H�3_D�45�Z#3�j���;�Y��J�'���H�'n���g�$ ]|V��(�-��gS�����糎�PB�C�%�����"� �fk
١����koqZ}�HT����=H��H�>�/zmӡ��O]D�K���ɚ\�F�_��1G}>�ˮ��h�ʮy�1㘩���ݜԏ!C���NZ�u3�?&�Hi�Pؔ�cR�cXo��g��$~Z�QeA?U�����Ch�!#v,��y`��3
}����V�r�l�+�����2e����/���"�NG<+�o5Y��;U�����I1Y20ڀ��(�L2
�$IG��Y��T�ԽB0�ݪ�a�m
�;�׎D�Y���?�䦖+A3s�݅���l~;� ,�t~�"�t�������	�H���>�ο�،����n�!��j�%�[;��/���_��1�Β�X�p���!^ ^Hu8F�.�0��XM<f�b
^<�{^�0�*����@�C��ޱ��?�x�v�ݵ��qV�Bk9���T���4Jf��sxV�ٞf.t쭽C���ȅX����#Uc�T��$��D~�� �Q�n��aS.A��J>�"2�n��(���CR��L�)ޏ���Xo׷�LQE{B�-w�����6������r�j�PY>wI��hju�Y�E��T�u!�N@- \Z)$&H�D��:��z��#�y/tNv�QG4��;�eQ�0s9�)u�x�(Z]FeuBDn 5�vr^�����+&Y[C�1���#0�g�HR�E��39���8������|��ҧ�c6���.9�"F��{������d8��j�TZ��K�.Q/��k\�D�b��+Ɔ~f�Q����й�KJ5�ۊ�ݗ4��`v׎�&��F(6�*�fAa�Rk��߱'����5�����]�܄$7.��ݩ����t9^��X�'hi��.����2��J�8+������ڂ	�A���bNM�|� ����߱+/�}�2�q�F'-s|aSc��Q_��'U�A>����ž�6� K����}���4���?�X�6@���L��S���_��(EҾ����ڡ�	��Q�C^��Z���>1 ���ӛN��͜r?�y�M��<]�(���~#�� ��h@�C�xɚ�}�J�%�N�)Eŗ�zHe���n�u#�ǝk��>�S�G�TO����U~���I�y���]��6���n=֦���  6��)邵X�<�"{Lu���YK���Я��Q$���u��B$�L�G����Xɮ̂c�F.���O�1q�Ǆ�Kʖ����!lڕ�[�����B�؞��Լ���;��ȑ�Ni�yrI^+c[ T�u;�.s���]+�vq@�ګ�"}�R�I��sՅ���+��A�1�\"��c���dڃ��Bt�݌QB�w:�)����cŧL�x���7C-l��
��&s� a�O?H9@ﾟrP��f����K���[?W���ݯ�����+d��'˺�
ߚw:f�6�V��	�W�;���Z��S��q�8�G�X���/�OR��ϟw�RS���<E��V���9�A�N
�tn��`-�0�}���+�?XSo���_�Y��V�	@YP��q�d	��n
�S�w�����Ƙt.���=mؓ[�Hk�Bƃ��+���E�^La0UAó���MX&��ke��[@�=�n0d�ۇn��[Sb��dUB��u?'�4=c!���6g�SMu]�#sV��F���w˦I���_-L��(�a��F$���sR�9X(HA���0 -�xH���{L��9���?�Q��Z]?��Y��o���mI���o˲7=�W�pUb�c򻽲4�*����� ���3^|)D�g�`޵������|x'��E�_U�m��P�[*��Ķ�� #9Z~�/�����e�����/C��BQ*G�YIpuLlxF,�=�f㯡9�;B"��&فex4x�kK�	�*[>A��%�>@�_�6K�1
W�v�P��d:°3�N���$���	e�� ��.bǐ;�0ڟ?5�^�����$$�rS3h��c'��|�:�^ua��z{Yu�X�߾/N�� ��g��_to�� aX�9AR��I��C-�e�ӻE�����x6J���G�˼�>!��y�27�h��������2.��� V2�ȡ����m͡x�+�J#/(#=)�W�m��@"�h^:�3h�Ʃ�G�O��n��ԑ�����b-�'�S�V�����"v�5X��<��k8xX��J7�l>�;��L�02�F�f4��jTAp��y����6sݙZ�f�]�۫$�F���-3�����ި�N�Ug�+(�P�̋]m�����u���3����G@X�z�� /������l>�F
`_���,�&�Ȫ�]��RSfQ�e���u��7;=u|N�}c.a�+Ϧ�g�W�¤O�G7�	�0G~1���T�HH
�yc�*ȃ�T�k���Q�2T��M��#�Dߟ4�4�oKw�C����F��Ws�\M6Øm����%��}g_����}��9XF
�	7ꗠ�jRk5��<�VW�G���n�e�B�E��G�����zl���nS�d\
�O���
m���Vr'�R �>B�qqr�յj��B�3h��f���<4�YC�%ɡn㧷��FdTm�p�\M�/�0	��Im��hPd"���P��V.�M��$e�Y=C���5����̠�Z��q���Wc�Z�t��1x�QH"�DM�6Uې���l\��k=E���kfJ��C�k��t���i#�^�Ct##2t}��-[�kak�n�2�	�AR{H�g$��2�����͢��T�4�H���K?�r���E�6Bɩ���P(C	Q�Y$�����=]�H�
{��}����T��\�@�� u0͖���a���!}�
�+�d�Wa�t3h;��gPF��L�W_�Q�%j:�:�����T՜ߕ+������S�U"FNA����Uv�/8�Ӳj���/��ؕp��e�.y;A��e�S��ύ�D	U�ሆ!h"F+�	��^6�8�i���N�Ξ���K�b�4�;��<&�_W�[��0�$�=w*F�%�6FbQP�d���f&m�t�H��n��h���7ĥ'R�X?,�ƶ�0�T����Gml���X��b���LD8��E�϶�W�)����m��l��H��Iֺ2T���_|.���s�1�S܃�4���o���DB�?�\�s�������Υ&�@TZH�,�����͐�G��{��ۨ_�����];�����r�Ɉ��Kן�r��U�Ge�&�u������ar�.��b�c�;~������\��%�;$��@��]�u��Q~�W�͌��F0�o�uQ��`��3'�)���2�n�>Dt驲z���M	?O��ވ�N7���G�	o��+Nm��vT��]� �E3yqm�Sg�l�^&�����ۢ�,܂���Hv7�ޞS�������ċ,���}�� d�]�!D�k.��r��jMM����˩��`�H>}��>k�j���jVT=��3�ӥg輫cmȁ��CK�gJ��C),���Påj�{wq�.wX�ٓhvU��3/tf�����x��%�iUU,�T�n�dr��	Q��AU8��gsA Q�@�#���P�e�kީ�)E�R�ı"B���6}�*()q���!�k0Z�\�R�������燬`�\%O\��>>su�Q�x��g޺�*�_D�T�s'l04�@5�y�|�A��Y<���ϗ�nh��}
���ƭ������!6�������v�{��4��vRXP0U�k�h���+�v1����H�t�*�.���	�Wv�Y ⓦ����Շ��jG~R��fz|�^
�kP��D��b�ж��ڗE���ȪV`XH��
]�}�F4//n�D���?l5"_�bl���dF�f6�Qy5/�1^��*g�X	"�)�xLV�#��R��χ
q+>T�O!�.�?𲺷^	���}V���=wMp�l�h}�	��f�,4���[k�<��:۹T^s\.	K�al���Տ�&`Vcm��1@�%}�m�����(!��m�,񡁾C���zp��(�w�ΡCꐝJ�\��Us�w +��n��5H~$�R�jޝWB�i����%�d}���- 8�r4�yb�F-�S s�(����Y�ts�����X�֍�n@>��o6#�eGiD=���տ��r�,9�:4N�v�����O?T�̔G9�HlJa-b���59�	�qdh/�Ja��A�MX�7�{Ȭ��T�BF���e"�c=�Ǐ6��8�D��a)-1n����eg)�":?�:6�����QuG��d�"�[0��w�&����`�-�P�Z,��!}����eq�WO�*1�*�fۭq�>�z��6C��=��WY'I����<���ф���01�F��%��'
wa�"��̬±���&-i�A���\k����c�	ve�Ƌ�'�Nd��L���d׋�j�ә������kPTV�p�j����� 0�c��b�=�O��#&�&s�h���p�+�����X:1�YwH ;0���Ou�={���V�/}@��?q�g�Ò_�/���\$UXS���!�+�Hzl�;�fZ"���5�p�^<ܥ��C�rM��o^b��:L��N"
K�a�̧�D�o zJ]q�KoI�����!��z� �R#鏦G���#Mc<�6w_ߎIƦբ|B��!ő��)�E^��W%��N�r�tjy+%]��ׇ�G3uK�v:܈�MI��B�F豹d��$�n�~�2� ƧW��:�/�*�+:���X�K��{��.ߦ����a_��M����0|����3Cj�<��	��jl�ɼu8*h�DL�[�s�<�dԘ,ډu��W�rޑ�=Ţ�|f���(<+�
�����à�E�L��k	�h���o�C 3�6-����q���f~4���7]�~� h�E��;�z>e����0�j�}#$��ϜAz��#5����AOU�47K���p"�j�= μ��O �[�:�����mzrGүv��j�Ǎ��=�U�}������4���'�
��u�cbܘBn���NZ����`0{����v�J�u�1�K����W�5�C��UJzP@ʾ|B�)�U���7�������1�,e	�9�؄$Ұ�/�q�����Õ�F�8�WF���v��uD=C��p�goz������.�T�t�ښA�IR��'~`�����Qc���(!����tTm�9;��MT��19�9��0�S��U���;�4��Ը���{����W�]Shե�R�h�a�u��g��^X��~~�/#�E_�Y���4�P[�*6��1ڞ�^�n�W���3nst@�^����)e|�p滟��&]D�%��WPw[��[y#wW���[\-�b	y�Q@�8&�Ӫ�{\�z#�E�=��r$,`Κ�{.5ѥX�lE" �C�\ޥ@�T=�_`U�h����q��l,t��j��3��R��.3H$��\۽T['p�[�ilV,���D,?�`o4�Ҋ3 \�&6�aU((�����?=U��Q	��9F+X�%K��j�u��r�!�-,*��oEM�����z�s,\��{'�*�D�&��Ψ� �%UQ���+f/�61�a��w�uǤ�.=G,�yj��}�p��WW�3����!8�lGTЪ(Р��ù�e�9���'V��t!���a_#����}[��2o��l&RC�#H#ﬤ�e�Vaۏ8k'�x�
�Fm�.���-��.���]��g��F�ů���;I(#�P"�ֲEh�vuĺ��<���u� �z�Z9.=m�zeב�6*}�"�h!�1|o0�âEZ�]*WU�Ԛc*���6�� �ܽǃ*m���C�r]l��E��{`�ʡ��vӛ����@� ��w��������{�==ӈ9�j��
�U����(PՄ�9�//C�)S�p��e��aW�H����Uz����/���0�������VcƷw��Ă��]����ڡ�M0c��r�2A�)�)��D`�
�/ ��F�ԁ�*�p?���u�SF��H���/��P���b��R�i+{��l���\�U-�}���U���Z�֗�Lq����+��v�~�՜���9T���^�ZX!�� lu�%0`<���l��v��`�G>�I����&���6PR���+�]�e>����{_�$8�Q)D�1��h�U,�,� h��!�f.�|$tq�q,���W�a|'I�i�}I�H���eZ��j�=��i�sTÓ"|�'M\< ���ݿ�[���X��X����,�	/1�S�# �/Vh���F�]I�����(���R�<�:�XӇ�q�?,�{=���+��K5���R�"�	�U�˒�L����Qs1x�obμ�,V����(�@VŮ���	���:��nM=�w��|����z�����	yY;�C��}X�="y�s��$�XMH4	K0nZ�lI@��Ť�9��|B�N�|��P�t3k2TGX/���Y��%Y�����by�H:�^��ſZR��Nq���0c�ve�qgi���f ~�+�Ut�󖥑�l]
�&Ҩ�z^��(j��+�o�p�����"�Z�m-�{�QO��Y���ճ7.�eR!�X� ��O�ȶ������?z��5�'��{0�Y�9�b�G��RM���#��|�t���HD��>�c4��uD��.�E��� &@~d;q?5�\��K�h��B�]�������]pu�ܤ��c�R0���Q��{�y8���B��Jfb�i���������仌ˋ�ǫ���~t��ġ�~_�:^�a>��F��34�S
��?(M����*�8�n����^^^��F�ݖ�����.�G�4WG����9NŁ=����}��aGt����O��6��ρ�YԪ	����u��Ol������%�VY����*��%0�2Q�}���Wg9����#Im
MaA��V�`�/��?�w������Zk\��׬2��w��c�|S�kei��ү.ƻV�5L���6�;�BַF<x��}���*n��;��ϫ�ܳ��&����ц&ݣ�'��3� �jޗ��-,�Y!c��!�����w�-.Q��o��+�A$�Ej>C�q�m	�?��MZ�0�e�9���n�G<�iԻ_zm���W;��&��w{r������`�+v���Tю&QZ� ����\s��fw�d�D=�΃�\g�(���t�=��r��I%�����r�\~�__��^�C�����Z-�Ľ�cN�S���$�;�	������G��Omλ��������2�;�@QR8$h^T�)�VQ���H�����y%�#P�Oy�r���!��}�*��7�1�4e����[���hΜ�D6��~� Tj��|�~�*�6#�8∘��?zz��	X6�x������vS|�}��Ǭ�<w.�$Fб�!x#��1VS�Z8hÊ3�����
������d_���{a�+Rl���������p���pQV�b���#P NEó?�#.8��-�rͶM������
���J?1��Ѐ)K���l�(%#L��TF�"<�Pq�&�*��Bd~:��ʝ����,+;�ؠ�J����Q���	Ӯ��J��/TG�P_�+3E=.��%�{pT0Խ�v�5���V��ɘ5E'3�g��Z�?y|Lɪ>�.ڄ���x�[q��֧=뱃��D�K���x J?�����)�QS���.B����i�� h���~��#Z�u�
�"��D�D+����A늢 �aj$:q�ă�P.��/�&+Hِ���V[�ؙ6�����wMȒu`#°�)�`ts��f��'hh������V�Un!�
?b�k����<͹�����?(�*�D�������K�c��P���#&{n����E���<-�)��*�XC���d&(O���g)�������O�	���\3����Bì�s�@�K�	�[�a ��<�xF^�Đ��"�#f���׫����J+t1.�!M�g����b�\�&��|D�&C��gU ���iQ��La�J"6���e�
���+��A�+�k5L�E��$�C;\Ə��^�e-K��:PAݹ���(�84�[�ci�-����n�B�v�D rZ���6�|T�Pc��{�H�&tAZ\޾cj�:�+�<K<H@2���(M!Q"�lųN��4�(�f���=��⃞w�.���
5��t�	E��� �������y�C�W�2~�P��T\���y)�]���qZ���ϫm;E��"_���Q@ُU�: t����%=w��8No�>CD~.)���r�*�|haRFIǙN���#X��D�D���5k3e��q�-lǊ�q3"Qv!�4Ѧ�=��K-.w���
�@�E�s�
_�h.@�6��K���&��Û�Xܫ����K
n��ʾ7��|P:���%oN�afE�B��F��*`I��ߜLԤW7q�6Maiy��-���o۞��Tx� D�q�8���{�*WE�O��L`���nܛ|�Z?�!(ު�\�%d��q���O�uM�l:����6�q
)��yr�??^6�[�?�y�lce����̴g:łv���x��VLM���3��e@?z�>��܆�^`�C���y��ao��̭Cz}%\��d@k� ��[�.Ї0���6���Yy�J��δ�����v�Ї�X�@�'��@-J�+�[�yZO8�!P5��v�ɉ��Ͻ���\k�e`�X���� D`��tW�N�qQ�s�L�y�Zt�l-<}�D����Þ��XA�D�G �Y}w���Lyx4�G/ԅ�����t/Â^��_"j5�����[��J/W��M�+=�$�3f|��hT����0��J�qG�q,a2�K/XV�~��J1"�T���<!��ɸ�᡻
5�����k5,��g`��ʞ���T���j�G0Er#�}��0����4Y�L9���;�{z�(}cn^	��5L�ٕ�2@���.��=�HB͐C�����\�ZɧP�{-��|�mfv����j�f��U �@ر����T+�,��Fh�v��z�.\\��Th*��<���C#�-����gי�맪����{�F�a�vz&�E|���$��m����J3�)̱۫q�lh��Ѯ���>q("�^$Ъ�uBLA�K��&�g����@�<�"�����<��S�@�I�&crt�f��9<g�'���N�>��r��X��EF�;��c��Ɋ��lV�\��k)%�|Ա)8?�;�R�V�\	*����
Y9	��t:���*�J��F��w8q�ΙX�Z��yJ�ر=���8��,���]p_��0�uC�w�e�p�.�0����,�
uxi�RP�����Eڒ��r������S|{��w~ŏ��zi龣Q��hv��*���>����u�H�z�)�v����Oo�b���l,Lx�6�
��'c�P�
/�����N��D��c���×���
��%do�s�!}���۩J����c���Q�ߦ �v|��4���A��wb��^t� ��fߙ�aĳTW�����~�,�ʥ��~���������A=���T�E�mQ�o챳������d�Z���m���YQ4���n�b<���%����1B�*��x{%Rܽ�:q �ˮK5���1gu
�}4��|-!���Tt$����̷���IܞG�!�r��wA�K��k��C{'6z�HG��eTz���4�M��S��1�f��ª���>jV�����fcr4��}��^��F�죘Zf6����\\��A���j=dA��&�g_20"��4��);ЋlJlmlL��ߛw�
�`�jʆ���֏E��s���=�bA�n�, �xE-��{��ɀ�^<�o��\�\��N\2m'��@��7�M�mȩGM�p�Y.9�_���^*u���Ϋ�h����3J�ae'�7(��Dr���}�|��`��>�G3.�y ������\������*�3�c��bu5bW��|�b�'Z�I+<ttp�$̕#΂�=1$~-/򀂐7����w�Ƣ.��-���ښ+	D��y��ڑ��d)2T�Ҵ�^^ ��|� ����u�Tה������V��D4�C��_r�_���AEr�!2�/��%h�����T9�,�\'>�������i���ټC���#c�����@���U'�cdnp��5������ꑁϗ1n|i�	�C�7 ��n���ɡ	Ţ,�*������zE���})�1���P_�l�V�����ˤ��쇈#!]n�n{���^�(σ�LJ
����&s@[��Y|��,�x��ʮ3�D>���ճ��G/0�	R���V�4��-t$#�?�C���i�3�	XOu��s%����-����2��`���"tzh���3HK�C °��9o�ȑL��yPI�r҇dL����?����^��*���@J����ؖ6}ɓ�S��|�� (�R���k�5K��Y�%�P,B�(9	L��z�=��җaB�1�}0}��5�^��U����_q$0�0��F�ho�N����m3V�^����ޚ�+�=�<%4dk�1�\�;��r���#�ˠ��G�/h����v9jY����N�]������F�@=�_;_�ܩ@����3�r�3����Z�1�Q!&	(ߴ3I=�K��Z�M(��S�1��$��B�T^�(H1D��ԝ�p�4����^��]`>b�wٕ�ğ����V��0߸��l���Mz	qc�T�u��X?]����������Jt�D	\;�"5o7��W]o�L�ך���V���<=��hd�b����uf�ۦO���Z���:f�Ɵ� ��;'�5��e�Td���R��c����{>2��ۜD�
���*��tA�H":S��1�� �k���z����ҁ��
^�ؑ]�0�z*9Z�qC9��~gld���1�29����Y�į�Y�HP���+���#)����h�DQ;�9�_/Yw Ec1sU��$�B|f���^"�J�n������F'����� ���w�[>ޱޛ�������ā�%[��p�R
,���[F��;�Å�E�v=�hu��J"k�����S]�u6�{s]�A�e�^{��φ�Zd��o����\/�]��qr�RN3�H#5'��t�Q��W;<��QNw�5�f��#ɏ0�.+���^������Fii�fgd�?�m;�b�α:�Jy�e'�]}�j|ŉ���yz�ܷ�a������@HVNݦ啑S�=	�ܾ�6�}d6�b�vГ:`I����P����k��b�e<Xg~kxӻ��al��}��ʃc"cba�^`��2�2*�O|7
����YQ�,A�Zꏾ��~�_���Aނ9Ky6�hS�.�������A�h1߸�H՞$ɛ;�����$
j�ht�@gQ�
B
|)L���>U�J��Ix�(�@қ�����.�E4+�X�T|%�g�כaI��S�g͕�Q=��������)���y��Es5��<~ �k��o�b5z����)+�N^���ri������,	!��-HH`�[� �:^,o��\��5�v�Rv��S8��6*��ŗλ�x��Ds�Y���-����vq�Ŷc
#���8�WqA&�p�é��N6�Ƀ�e���휄�	|rC��x�;�=�s�k�oa���O'�����MC�r��=,�;��0>T�܏�9���Pn�i�{}~qf�S:��2
Bǚ>8�@�"�J��0H�XP�x
>(	�eiLW�4Py̅y����aO�8���d=j����n��J�)�>o6-�ɝ�-^/�o�L������.�������W1Z���	���et����1�F:9�������c�@����EI�HЌ�0SJ�=&����� $��݌Qʺ��h�W[9��Gxp6��`'��+&_��?h����^�e�U��f��P�C��CH��� Pu���q�%Y\0%�g���#���V�.�^��q����Y�v�R�X��./��!W�a&����-��";Y�nR�H	ˑ�wk͑h���J�d1�����DSpqO�T�c1�*�h[ɧ�lW�>�Qt��*;�;����.���ϛ�$��Gt����G������Χ'�؅�w��)W���1���\�"��,�ޱ"|í���+�E�g�"n�/�v2��mX�-�V�M#j�j7�Btp�}δ'ʂ,ŒC-/0T��Ϩ�Ժ�]�Њ^�c�{_��NB�[���3�U�6�9��.�]�+�杩����#�������؄:�����;3-����/��W���<~�� yR�٥�N'�Ҟbl�[5.���j�P�Դ�3���~.�9Tp�}jL����2��c� ��!�i���0�� e��
ČV90�L�\�WJx�B����z���_Rk<`hmʤ��V&��� m�]x�A=�E���z���V�M�(y��;�9�a-�"��]�T�E�)�7��
:GW43.g�J�Ț��J]��(�������v="K�A[܂��S�vW=|Js�!*�-��74�m�ʪ'r��2�W4� ]*Ʉ��.^��&�Ѷw��x���q��UQb�~ϥ� ��[詯������g
? @m�V�8�n�
ZGV��RFj�0�s� ��r����Xv���o�&d/��T��V��Im�~[��4NM}�=��c�R� �<8IH�v�XD�o����X�a�$�C���`�ґ�O;�@uj3љ=�m�q)�dUz�˳d{О�y���H��;�RB&��`��J����K�~O~��M1��<��'n�IM�:��̕Hs5E^��TBFB)���вk?�w�t��p��5@6���l��}�������h��<
ӃJ�Uc����Ԉ���>��#�s=0����H�N4Vr��_�y��}��V�f����i��<��������V���0�!8�b�U`M���Ӓ��*C�`�[���[_�������&���1���`F��._A<g}3G��J����Km��rM�����^�����6�YT�R'�|�V���)��?e��C�K8��4��^t"۪���[aNS[O��hy7\7�e0;?m�'ͻ���Nr���́^�� ��9�|�|��m���\��HKD���P�����>�g�aM����m(�?�=�1��7�������V)��?�Z̥�ɿ鼖h௺���{�aJ�M����}*��5{��a:/F}��*}�3�&��Z �	4.03M�� w~�����fLwj<{ေ�1g�(rsfU�i���&d⯷���x�=�ޘf[Y��@$��X<b:��bnf��ܸ$�]�epTr�e $�x��`٨.S:�$�ΐ�	����!k'&��C%��U�s��;�ƑDj���O�`nR8����lқj3"2~p�Q����j�]eH���gZb	�S�"U�.��s_�r:�oF������a����`�,����P��C��O��M�������|Wd@�^Zã�3���"���[6�Uz<��3��w_ʟ�-l�ҡ
������MyK���d:���oh� Y��R7uʉF�C{p˼kc/��&�ϑ�� ��3����9Vpn���ԃǥ�B��ۓ*$�h�ځ�l5�d5�~
ey�ϟ����[AӤ˴�PǇ�a@�	;�}m����b��^ω0��En�uڋ6�9�(���63�/R��ϊ��G;3��Q"S�{�Џ������\)� _�Azi9�R�0�{�wuJ�h���8k,�W�bϪ�6)�+�ٵ�:������ϱ$s�����VD�?V��K�B��7t9�S�s*i3���w#{�:���X,�v�;�ۙ(A�m"�t/*�06�\>�ٲ���5���s���q6����eSH� �Bj���U28�m�K�09U͟@�צ��LD\�.d�x��9u�ӛ�K��.��X��)6���	x��xe�V��l~2��@��E��_�ڼ�x�r�����&3%y���d��%��d`�%Y��}��N9���;�PS�6A���;�@�#J ���g�W��Yi�dr͠o+8dn̻+8��5X)y&)iJC����d?t3a�3�b��䥢�s`���H��d����q�*d�G��6~v�5�/R�3nC��U��O"�.i�,��M�tB��՛���MYo��ȕ?�`!���N�mc��
g$��#�~���1n�(7e����L'�	�FSW����T����j�\&_k~;8:5�M��j�Զ���}�l��!���ף�{2F�{A(I!�D�v718G�n�d�/�A�ڦ0�%�Zי8��M�j�xqE�����`ڿ��^m�DU8dt�5��q�T։NA�7���t=m�`g�+=��]>��*BSJ�)7�7"���9	�g!��
ay|y��3�؛쮥���X<��qF#=c�4��`Y����t��nWp���#�>Fp��#���t��+ F��g"S�&�� ��uB�3xx:�=N.w�j8�sI^Ǭ���,�����q8�TcVdNptDq{���k�-��Q⪌��J��e����kn-fòs�֡�ߩL�罊�zD>�G��%HK��l$�:�
�u��v&�N�\���e|�ҏ	c�,����NLk[�DPO�f2I�LH�iu}!gfĲ;)�^�)�+Y�g�������vG70��>ۧ�eF��2�>f�s��T̺H�-ِ���^�Tr�py^}4 �~��j�.6�u!ݿ$hx�w&3��$�J'���E��BH𸪏Qlc�LE#4���a'�O�ӯ��C����3X]��&j`Nn�,�������E6:��=ύ!������p�H%�@�(Y��R	��\ڱ������M��[J^t�;�ɭ0�.	LR\��m5{�WV���n���v\��E��I������4�k�����HM/u�3y�����I��}x�"����Ȳ�D�0Z��N̈́ԢYJ!qפt�u�y��l�;��@�`Z�q�V��v�:�c;8������֭V!5��	��'��f�X��;�� �6�;�I�$�s@|��׊�����ZR�H����%�}��mӗ���9�<"-�i�ks�|SI �a}���$�#�����/�� �O����D����U>XL7"���:Tz͆��$!�o�0;��-�=�Neb״��<� �DID�H�-�6� �Z��:��z6�	���9�x�J�_+e��PA�������z���4r���û$�iJ)����:�V,�M���@�f���cK�� �V��R���?�%�Ӂ�K���ej����+�W ��}�:��r�OpFh�����J��4�3Ҽ����uȥ�=�Qݠj;�$�4���+���j:~���A��6���ɡ����ˋ���HU"�62���+^ɖH�"��)�ʎ����.1_�]ndh���,��m��]�<�Ò&9�v]�)zF\)��\��l1��y"�v���Wz-C��Ɩ[8Hn�V��RLb�h���uz'e��N��E�3�F'E�#G9�
�zb%䛓��JvD��j�~!����b2�,� �ŋ>�j��mĞ������2�Wv��5Y�{�S7U���*}�� ��B��\��؋͇np������'��}��TG5E&���1l�O������3���h��I���2S��lx����o���zI�'�����7�^�b8y6��Y�վ>^��$�Lo�	]���-�r������4Q�j�Nc�uh�����2S���R����B�'�h�*آ5l��-�B�]���C�"GXz����o<a����� p��˃��O����,M�ޯf���jA�``V�HJϘ����?� = o���g�q> ̨�LΙ����
���^)�B7�[��"#x+��i���ZlÛ��7V�ν�r54�;�=+��d^BV�wO*�VJ"��Y�*��V���ko��A}9�KP��-���u�n�Rˑ3�����0z�O�P�,v7�ʖ�Z髈˽���("�EqW�Z�T��|py�L< [ه�f��i6�wgI�m]���@4���Y�DRS.��`ȓ�~�(?�i1���X��'8#��7� "D(Y_�2H�&��##4_߾��|u�KW�1���T�!��z��|�G�bXr�,�	�
�����w�g ;=��>i�r�v���Ϛ˚�^X�j������eV���5�%�=r����*��2T�}^_�|f�bBz52��$�|9̪����R�"�Hڲ��ˤ��RϾ~ȥ>FI�JV���?����^���d���%F�4\�h8a�Cb�9�G,E %{F��l �bU��
F���2�LH��zO<K���(1|���Uj/x��;|�Hت\�{/�爣Lj�]��������[W��nơ:
.%���֒X12�q@-��Q՜�Y�+�F$ԋ`�2���^�GI�J�o'w�:+`���u6i�Teά�1�t��5����0�1�ݫ��k�aҥl	���Dp���O�H�'u@�s!+�(��lP�D#�����h]���q��~R�Ȅ�l�M����R�q/�4#s��k�^ٹ�j~��
e���To֑���6��=(bС^qV�~�߽����ow\�w���&��:��[xO���^�J	Z������ȳ��t�/G�ю���-�;�q.�@� Z�Ϲ ���n���J�� �����kR�cP�8���R�:;�]%\_߆� o���ä���Ep��
��4��c5^_MR��I�
6/���U��W�n�"�VA³X����b��[R���� g����P���(G0!��@w���޲/�^XO�bJ}B�y�͗�^��>
R���q��}�0���\��DD�8-��UwC3r�[��ZÃu��/��ƄSÓ�$B���ɗzw,U9]��ӑĦ���V�q]��[g�gnI�3�m��A��:]�FƱ^v1�uC��9� S��nI�}�s��m?���ɭ��� �b�4����}:L�����{���,D��Ժ����2(��K2,�슡LX0�ae)�T�R��GG0N�G�	U��K��3+��c!��_Gd��f��y��~���5����m���il��'�j?Ԥݩ�\��&n*����ȡY���*k��w��|�(�ш�f�4��m�AD��:����L:h�Z
18I�!Ͽ���AL}�P���co9Wݨ��+�&�ӫ%�H����?�k���ȠV�����K����q/lD!�TP|u�1��YeM�����%���D�W����+X;��#s�F��,9!�bݖd�hN�/�����~	��M�7�q�}᪀�nF�\�+}Q\��L0����N�^�Bf*���S�E7�s�5\�%(�
�Ƹ�$Lg7ͺr]��3�r�ﭷ�k�$��^��E�2��(��t��ϨS@i�r@O,�Y���hT���]�wx�H�_p�e
j�c�&'D'�Q�X��xLr}9�Ή+� �JW��:f*�{'�f{�x�FO��XM�q#��O��iUY��m�"*��7IyxM76&�rA����s�װs%,��@� ��s��7�K��9�7oU�a6T��UD?��O�"1���%�w�W�#�-b����&>��̷@FJ9��eӐ���8ۻc봟54k<G�pS�	�֊4����IЯ >�mۜ�,�ݽCU�:o6�F)�b����Ȱ�e��Y+4�^H�PM���g�d�to*�ݛ�(`U��0Å�!O"�B��bAW�:R7	Aaɧ?�d�{��y��~4;�lItEjNC�+b>�h�8�_5_"���U��x�o�ci�{��1Z��:�0��?�9�u��{�1Eɓ�lD;�PI��jU�{Z�-5��J�������mz�5�j��=��7�5(���`豙0Uw0�\r������%��(��)d5�@b�r���P��vi��	B�V���y���s�:2^{7�Y�^�Mb,����5	��eܰ��߇w�?�T�'�ZtH�D#��M Q��*��b'�-��=�_ZVGu�.�?+�R���;M��#����W�0uE��k�tOք5���٨�	s�V"'�F�w�IH~�ye����?5�f���Ϙ[�����,J�!��9�j����!_qn'�tR�J���P��}�eb��45��|��Kb?]��O�t@T�k��k�?��/��2�
�D=|KU���''R�U%�K�G�I��8��%!���%����w��/�H��F�����
���XL,x�MO�)��X���O��Vuא�5i�پ?4Iut��a�C�t���"ڹ�A�JyX�>dd��v�Ɩu��9��P3�ʑj0b7�3Yݽ�^����(��fNʫ%���b��>z�1�آ��hT=�W�� (�g�ԍ�I�����h��1�W���b�N�'a� C��u��b�k�C�J�"��'`i�I� !#�z��z!�2(��㪌R�:	�G�\j&ux�{�1"<���A�_�G,�Z�P$���J�&.��;��o��*63�$d�C�g��ɚ҇���Y�T�UM���&���}M��ߗ�趚��v�C�ϐ�^�j�U�c�%E7�S�ަ.s�hIlN��.iπ�`|K�Fd�����9���-��+Ժ3�>�,c�"� b���QV��o�5r�@TI���?͜\�?��Ē�<q`���(�n��Wo�mrN+$&S:��:�����\�������2�����:B,+%3�|��Ʋ��xWU WO�X�d�f}�VVJ��}^�v�Q���q���	��2���M��f}�5n9!�����<6�~X怙��ou�;/�;�ă-��)V-8R��<U��0���v��w]�,URM�F  ��	�T�7w���טʲV]JD����$�Za� ��8�h�U/�}|GNG��?�y5O�q���_�i��������O{�g�Gp\��NcՉ�h#�VUܼc�>�;9/�Hk�Jo�^��G��MAq$�|K�,���ߨA�|V�v^�0ٞ	0�x�8rY���D�/�f�`߽�}�������u.J�3��ءн�R�6�p6ԑ���!�����t�*E-"��id%�m��P̦K{��8�)�����^q�������ZH�kY+������pv	%v��T�b�=�]0�*X��{F���E��$%�(��ǋkš��������!\9=l��E:���SB��J�������'�s�)D�N����P��$g��P�qX��A9y�1���XZ��;�ajs�p���uo���i6�J��@��޾�?�3�K]�eۍC����+��H��R�48}�Ǝ�@�mHO�´ܽ���l��[�#��>��Ra�����+Ifj�����S��������T_�d�l�r�Rq�X{�AYO���e�Y�gλO[`l?�6l��I�z���m r�J��?�Ie��Tt?��M�	��ˢx��6���l�4��}٠��<���t�p#(3ScܳT�"��/��{�s@�����<TՊ\��m�[�-�G�X��ћP��tL�CĵJ����q��n��j3�H�'�}��>`a�5޲�۶[�i�}��+}�����Q��C�O��t��?ne���!ʔP�ӆ��t2��ј>�u�9�����!,�^�~�flYZI���2�T�sn�z1��p�J�xf Aʚq�F㑶��Py-�n�u�(��ĉu�;�t�ڥ�@}��Y�+o7uF[�dk��/�|�I��5�?)*n� |�ʍ`s�}�c�QHM��}ҿ��)h�+��7n���}cM���V}c ��	N�y?�<K|���3c��ԻK `mt�����-�vS�d���xwͪ섀�焾:�j5fp�e�@}����-�1j��������:�~vH]���S���K���l��n|h$2�<V�֍ŚZ]M����0kF�����M���A��g����ϧ�{��/�a'�l�/efu�l|P�p� �n�!��@o��}��Һ�f�BQc�uQ���I\�Sw�(�ve��%��V�
�Ah
���' �Óh����w��X@~$���9L�&�V�,�v���(MW�����+�J���_���]R%�oB|;�Ը6�Ͻ q&q`t*�D�x/!��o�~�'��L*U�ҹ��}����`��ÕOK�z�b�I����zL���.꺴|�8� �,q�ٜg>�G�[�ʨqX�)�z�I�I�� ��(\��%��t�7��S�G4���j�f�g<L�DI�\����2�_�!E;7bv�c��=�:ަW�c�j����t":z5m�!6�<�a8��ʽK/�6��ʫ�u�T-�m�\*���i��0�C7)8O8�܌7�9%�=����4��%D�v�P�(��IB�	3(+X�ƀ~���3�n[�A����?&*�� ؿje�h4P���"X�  ��k`�F?�g�&���7����7�4)Rъ�L	�Jk�7�;���`��GY<���g}]c�$u��.������T}��^fr8/��-�:ˊm�]>]h�x@�����﬎b{�TWg�Ų�'�Ӝ�7s�^/��$���Eu�������Ug�2JVlrQ�/���j��KׁPS, ?�x�뉛�,rI��)����(��>-�na���o˥��R�=L��?8|5���*��P�|C�p�~��ת쭫_�l=4�����TW�"�?In����d|�6��:𴇽�F�4��d��aߞt4��Fҹ�>�4s���"��o0�؞#������ˉHѧî�L��!�Ҥ��Ć��(A*fI3����v2��VevHȬ#�vo�tVaQ�[}f:�cW9�*�Y�ž~�hRg3�C��	��B��D48}�@�G"���eM���&@S���.WDȐ�zp�s�fJ���A���=MUr�M�Q>�˃�(�ȫԠ���Z�m?m�=���'~|����%��=  �\�}*7W�<v�l�������m�w��_R[aQ��,R?��M�X�F���T��[w�:���rm1���t�3︛ꞈq��o�0®١���[�Z�P(���
*�v�&�
��"��:�����u��@+�yc�Н�����H�Y,KB����5����-���{�t`�g�a�[��D<�Bvh�t�jѽ�%s-���;�ܞ��������c�0gCcM��koa��9��dQ�F�Z�`�����U��A`��!�K��8�6��Մ�\c�qARq+f�0�LE�ީz:��]��6q�� y�n����� �S����uŢ��Ǖ�A��Z����~o�)E�_�c?S�����7�:ͺ�s�vf��^auN1}��cj���@i����}?W6ɡ,�y���$��#,d��X)�0��f�*݌+�Li��q��e������%.��/�~d�OgBT�u�&��*���j33�3���t3��+W����;��Q��z$� �cG��Օ�7L-�x],E�3�!N2��U�M$�*�NF�%�v!X�U�D+E�oy�x��
Gbg�nH7�%�����M��TD�mn�R!�e/^p������=G�r�����Ó�����-@�6�Jg��lg�|^�y��|5�a�%fe�W�I�؞,V��E�����ߓ.���#���d�ǜvJ��D~L���()'<���"�e�����j7��qF�ĭw�i��D݊�E�ws���R[��5w�H�eI�w�o8������(w���$Kh�Pvr���CL�Q7:@��u/}i����h0o��<�Fn9�DF��Z��c�eRE�Z!u�Eo N�%<�� �ʂ@��oJ���/�&���NC��E1$Ē(�(�����[	���T�����`�)W�XȾ��)r�M+��Ԓ�fa�d:%o�eK��!o4`�yD���I�c4CH���eO{_��ۙ��n��|D�F�C:l4<2�9���Ɔw�-U�ı�k�/�yԇ��I)=�yGL������۰�^�D�����u��@��{���6��gN��Hʯ8fE�'���J�^b�Y������N�,x���o����U6�i�[��]�u�[�Y��s�6�sGO��P�ѪF<���#B$���C)�_-�G��Σw��Qc��m��0��@��%�L�:xq}݋?cC�*Ȋ�%���+��g�ˋ���o��X�dR�i&h2�/�
j�|�/Fx�.8��\�v�4T�+�|�?�J�?0���%YsV�o��`����y�:����)�����	Ayva�V_���m۞V���T����Z����.뿧�t�=e^��t�/��H�v%���F>H��p+ݲ���M\��-���q�F6��]�u#s<�%��s�^@���8՗�4�'��.���7!�eA�A뤣�:/msdD�������⪶��I���c�e�vA�<�<�(zS*��[.�ZXR~iwD�������ɶ����&C8�	�aG��i�d��ɝ�Zq�]]�r���z�;\��B��x�`Z���næ*�����e�S�=�����u{��/�9`XW������D��la�c���-���k�v��5�=������愲w>�>�j�Н�0H@����5���&&\�n	v��P]4!!��)�H���(EH��K����yM�ǉ��t"UH�
^V�PT;L��}����"d9�0/P	,WN|�FT$�n!��qA���Ƽ���>��1��&��)R�R��;픷�@R����)��Ϡim~E�������$nl�:-��4�%*�,^E�f!/6�6sC-w̧f:��xe���fC��T�x d���-!]kM|R��I�:tӠ	P�W�O�9�|�˧�ڒ{�]�/F�O�J�g� �����Jt=��������k5�ʳX�;!��4�C���l?h5��-3�X��&��i���R��w�u��!.�X���Um�ۚ�D��_��t�@Z*P���i�<���7�Vl��8�tmZ�:��<��`�J�s��4T�,>
���=���1.\A��c�Vha=f�@�3%��dyW�v`�Ir��8�80����)W.+J���y>�kyw��UD���f�v7��WmA,�߆C���і��k�wf��� ~��~J��t�be{�
�`��ؤ���3��C��W;/6�}�;Ng�^ft���^�g^)����mZ�������KF�W��=_�X��'��^�1�Z�C����Lۭ�������������������`�����iP3)'z ˤ�0:�6���u¡�-�n=��hG�6[�����ώ{]�ö�`O�B~P���1�Bܰ�.�Y	ov �sy;DB�3s�C�VbAԈRo��:�2��
�Y4�o�u�g�O�N%:�G)��[o����,
��g�#�������-�۾cB���*4�lt���ߌx�_��S��
18���;	�׵�m�b]�3f���J�Xqx�/!��;3\.g0��1��ãf�/�g�2����7M�)�TN�l����N-2�>g~�m�sn���H��k�.�9!���b�h��~�m���-�:f؟O�����^;��|f_�/Ȋ^�c�m;X�Em ~Fxi$���y����k���]0�锨�޹r����f�Ҝ6Kɮ0Ҧg
(TcR���z�g���3uc[�&��?��_�a�'��İ��>�� �wb�S?h�J<xwз�l��S	h�����O}Q�|�>�,L:0{�'��n��d�`6%�|?;F}��#^d{��O�k"|��RFBVr�9�v�,ӛ|�E5v�d8|�O��{8���c�YP��GW���;�<�/�Q�'�������-�V�A�ER��4�N� `�����S������S��5t��$�؅I�����`RE�ʸ�嫡������AR_[���sB�z�=!�`"~1D*��!F�Lm\��G��zF�5}�;�2|~�i{��^`r�Y�2m�l�������Ӡ�zȫ1'f���L��[�%�~��芄u�K�۲T��3[���@5�)oX]j��]��0t��JQKüQc���\�6z͖E=��!bÎYH��Ҿ�F��{u�ĉ(������]��*ߏ8c0I�"Z�"aP�]��e/WnqI�6}��C���ͨ �n��V��� �I)2�	��D+�ꒆ�ͳIN����8x�yd�3��<Ku ���!>����>�{؍#��[ƿ�JkUJ��P�hQS��z��"�z��s������N�����3��)e�Pk@'���8��:������hVc�ȘN�"天���C<)
ց�]ӄ̶���pG��e���A�Δ�W��<i]����(d;K ]���o�x��d:�i�����Y௣$�EĄ�*6[MWrG��$�
��b|~��]�]�>���5�N.��bt�i,3q�<�[D.���w�ݎ͸�� ��@W!�#?o�%��`
!�ӆ�N�*;��N̐&���~�c��ᥚIR�R/����Cȑ�_���ul�%\��=_�7�8.��5�y�::���}��n,��s7_�Jƴ��ۻ�In�d:���M�Z�.�@x�������R���,�=-�]���@}U9��sY�ֹS���)����3�]���Ř4%& 9���7w��A��"�85��b��S�����$�<ω�ڝ���pr���@�t}e�VEC�?BR���tiW �uI��fT�~C:Y���A���!#^U�V���D���/�Y�T��NOl�0(<q�U��nlW�c���̓QS /C��SC���= �K��b�Q��9��Wym�!�~c���a�L�o%�U����[٠�P�ä;�lF�]zG��Fp�<�@r�-2�"a,�)��5�=�ZhbL-�wH=�%�em7����y�[B�߶ �V��S�����qNz嘲dU��^�� 8U�a�������g��B5H��~�|m����1���JNK�K����,&aD��=+<�6��O|�tF��0�ށ�%@��ci����
?䇱	@L����K��{���IØ~�1,��A5�tо�L��Sr/d��RN�Pf��e�x�u4��μ��ڄi+��?��L|o�+$@	*J���e�~MX&��k$�P�[�I���1o�[z�*,��#%+Q�T�;-�H�����fhC��L�>L���\CL��}�kV��	y]�}!�o�xn'��es1y��;�+�تZ-nҀ-��̟��l��e�W92
.qr1��ђנ���`	����~��	MN��bB4e��p2l��R�P�+U��sb���?AyU�*A��Ma�5G;
=H���Om�2�����ҫ�W���j�|@��#
�h�O�v�͜�~ �tBظ�
���#2�����L���_F	vR��{q��;Q��"�[߷H�r2_�e��IX3�������͐�����Jjr��*J�E�hh��U1g(��g�Ă��֙M��,F�,hu�U��R���P	T����m���΍A?���W �4qRnȞ_;4��;V�bs�bF_#�&ڕ�J e�k�sD0ɏ,H�\̲�/J�]cZ��[{���%+�'DK�~]1l���I���~�{y�ʬ�pb�+��}~��̓G���b�|���%��Yn}
����n���%e��B��.�o�%��C֗�ƞQ�#:
@u6-�HB����U�2Wq��w_���aq�rH%������h����ⶪ���S�^�_�֟�V1�)�7$�u�����9A�T����X^���4(;M ،��2=��l��q�+D��=�����WI����\��ױZ0�l��Þ����?}��a?N�:���P��uzq�E�G���ӊ�����|�U�"7���ӣ2=Ϩ	���@�U��R�Ĩ_��-��N�m��/X0���S��.�R��%er�S��C�7>��p���M�\@ �<����/�p��@
�:x%����1c�g<Ϩ�5���[�s[x�נ�Quݟl|��o���0�fUɴ��f�$M���C��w�:��S#���1�u�����/��(�ӝ.{�i���s�V۹q���Kio̷�-n�O3��Q��m�BG[u@R�l�00�K$�_Ԏ�t�NO����/f.�T�fĤ��/鱊;B]�����e�H�>L�ߐ��b�u����>��=�Q�Q���z�t�C�k�!c�lNk���]z���� ���¯-�)�+9�	m������ĩ߳~:;#�5g#p=4R����}[�]�2��F��KX�,�ʠe<4�C��BC�|�{���`#h�as��'9hCY�.�.��g.��<�V�e3���'�51B�]j�N����vl��̍�/�:�}4�d$�ק���3ҿa�U]V�4���>�+�=W�!V��A�=f*�g��r�A��,/�¿b[�j6��)֙�@���9Q3T7���}��
�c�"�N�yW��͋���6O�?��+L���~�2G�r�ֵ�6�9A;'��X|��U�m%f����0z�t�]��Y���J�Аז�Q�<'L3�=9���Wǁ��%��Vf�ے�
Tl�'8���Vs�0T���"O�2E�~2!f�N;r{���CM�GK�0]7KPH���,<��(���0�f
�.�`��;ԉ|��#���852ب:f��'n��t�[��k$����|&�3�M4��R�8-�)�¹r�Z��ޣ~c�T��4u�OB�l�x�RW���Q�-&d\QaJݏ� �6���ad�0&���i2����"@��n�"����"�ȯJP��	1���NN,΀ay��J2H�ҏmfs����(h��HLس���L�sO��!)Bt�QF?m�(�K$O2�HWh�UUQ��πG��Y7.%4CN���(Tz�D�2�VE^���ۊ��)��a�j!lZ1=�oԃ0�j=e6�mnSIX�U�\	ME���$D�����?�V�&���M���MZ�KH
���r����X��*s����y��M�y�x�eg��o\���F:!��#�K|��'5#ߒߒ�ɑX�fK�_
��%!|]l�n�t�e���R7�gD"����}��"5���)�f0� |pKp�#�:h�-^
aD�[b�i�މ�l;^B���i1�Ko*zkI�/�n�ޣ�%|�pݥ�����x.
���X0�\����Q�r�F�����$��~���&�c���E��P���  ���0��+��FU�_�mGޡ0�>�����k��������Ѧu��ߣ���W�2*~c�o��?Ӿ�^k�>&��g��$/"=�]<n��-r����Y�vE�l�S,(;
h&�A����@&�����B�I���QB����(��@*7t+^��@�qU6P�����=E�'�@Ɗ�A��,���6�� [<��˓[J�o��`�#Ȑ��+ �����L����dDSөld����"��K�K�q�b�T�ͷ����u�$ET��M/�(��f��H���\���s��5����*��m�?�8r�{�
w8�e)����0��>�xf5�i����4��yD�V�D.�D>�x�>�+��F�CI�dN����s%�:�f�5fU�lj)90�,;�s?G�����s���`�S}?�Ʀ�M���+D��RI�sY��I�J��6F�H��=�k^�]�4�#t�T�ס���dC����%��ڂ	�8�&�O�7.�,�>�9pQZ�mיd8'rn�i��"�� Z���:u���F�j��YCD˼�S?/�h��\z)!fc\��Q.�H����5�/�� "��vt?6�n�A|$׫�w6@A�HZ 㺕tzX��/:�ϯlk@��\��^��&{��2Uxg:~��3M�T�}fo�<�{*�5۳"P�xx��~��T�g�wp0���b���$�?��̣18�[[�:��~���7�g���'�dw�>���mr�L/��|E��Ҝܺ� ~�@[W�x����������t:�DƄ��dB�1 `��.K����n���)ҩ\�
uS�(�|&�5A��a�V�b��h0C)���:�;.�ҶSD�%%S��*9��o����\(ǋ��9u�E��2)�򦽬z���	Px�� �>)���e:��S��W�I�4ձ�^�9�����k��ɣ�X{�$Q�����05��g�q�j��Dn��o���=�`d�ڴ/�4��4.��*�W��qX�W��s���a(�c_��e�~�HB�k@�z�8N�Z��b��4b4�KD�Pp:c�M�4i�j��#(Oٴ�,Ez��g������ݩ�LRڸѠ.�4�RW?8���GOޒ��g�{G���q1_a+�[���/������ �M��г0E�ӏ�hcm�E<�W�t�%mL�Z�n�o�릙�nW�����K� C4�/,
-A�	�ױ	w	N����J�dݘ�pz{N��� 9�8l��U�B�p�X�+�qA�m6j�^��_RC<n�Xֲ�1@7�3�����$󕚫c��A�J]{����P��dm��i�`��z�t�`����/�#5#�#޼��&���"��NL��ū<ڻW�dABH�D�#�a�6\@9a$�H&�@��z'ɕ|�ɪ��o��(�qp8��A!s�'�$inQ��^��<V<�7_F�X/�[�X������&�{����&�{s5�"�鱓�%dfV9r�
Y����D1��y��E��}]�	����x�c�F`f� ����V^�+���<�K�"N���{V��6��d��]�Y{�	����)�~[j[:����w���!-�z���_��6�kR������(�G�{$<ŧ����p���������E�}γ�273����r>*/[{[[���R�s
�mda�8��3ҡ�!�tAV�(r>�Y�폸� 86�0X�C��r�-���?����uג=t�8-e�&��\4cZ5� �R1U�M{��BA�s���Z�U�o�5ti��#rL��<���Y:�����C��CkS6�:�
��7)�;̟B�����E�D4�� ���+6��6F����,��m���34�f���S���^�F��M*O���%�jER a0�

�D7{�ƿ�#פ��%%l�1�ri���,߬�;0�Ks�ht��Iܽz�Y��z[���z 4|n� �֊�qq��Z,����x��:"B�U�A�c�c;+?$��x�R��_"f�ں �8��q�M��wMg J��@�8C���:�H��B�zN�֦xȈ�`R�%ˮC3˺+��P��'}� ^�9��B/K<N��|e�u:Vd����^�0M��k]��Śي����Źc��[�<�v�v��Հ6����s������xL�řL2��/g4gU�ϻî^p�H�9԰�n�m����!�9�w2���)h�(���߾����[�wl2/B���}��0��)���m�� ;� �Kd0�5�"v�dN��X�::K��8~�?�kt~RX�JɈ0�r���kf4��+/"g<�`��n�hz-c����� 0Dn�kQO�v��z�I��%�BG�;vʲ�Ix=�|W�Џ)�&P˔+@������2'	���Aa'nu��{�*�x|�3����k�f=�JD!��&}����F��ܶD�48��C� ���S�y�$6|S���X��M��F;U-�����u��	ӈ�nQ8��@�g�?���ږ�u�A0H�`s��-�-�$����s�KPHބK�Ǌ��^ �&�v	Hr����Y@�J���sZ�����]�ע���[2pp�֍:���F��L�k�Ŵ��j���|k�����x?ۇ~��:���^4m�����,�C;-�@�%1# �����IR%� EJME����-_�{��}r�����:���`�F�n������RP\2	�0���"�#_��9����Uf7�1�~�Tc"O	E����v
�tZ�Rk�>_/���b��<;�Q ����
�%ˆ��D-E�W\ཡ�Q�1��f�vJ�K�mV�?��bpӭ�K�>�u$Sv<�~�7���$��C㇄pP�ֶstlmD��:U?�N��
���k�����h������Q�N<yK��YymW���LY�ne����E;rM���Rz8K)����eS�jSrqKs\3�m����7�cM�w:Y�f���}+lǡB��.�3�:-��Q<?53�V����YUz�mY��L�?�
H��W��	�[���r[�����OW����/-,���&K	d�%˯���=?��?���xL1���i��01W6V2�\c�,x�^Q�'����C���f
����pwf�����WBI(��q̣���ʺ��D;�|>.m�
#l��5/:�fBp2���������I��*�HG)#���[	V��W+����F�_���͚,�\������(.�3]�I������l�u��������ōl[;��;e��.+A��D6�������*��Dg9�>�2���z&x�E0a��X�GE4�@���wl#k9�$ES�"�OE�k� ���udH/Hh���w�('K�3��Cj[��v��X%�)�W�ۦYj&TSWg�]�Wڦ��Mxh�}��[)�vI�\&�Φ�g�39%{�+���*�A��t��Zc�^,�ڥlS;��|3�'/��3��S�H�w�cVb�F�Ui��F1����HK�~M���\�?ο�<ո��N�c�ik���-�q����e��_l�ne���-��E�fUR'-�2���&v>�u�Ů��hȐ[���g�a�B7��bGǈ�#�S���w�vpp7(�W�;����B�.��%ۄ�}@��g}� ��U� ��$���i���M�Aۅ��E$�}��Y�׎$�X��[`����݁7�a���=J�S��I�-�$����k[bh�k�Wr��v�5'rXYE����BCv����#�/P%,��Q�ӏ�$�Lq�F�+�9�#�`A/��S+��XY���%�H��t�-Ŝz݈ev_!2S!/8���`���'�@���#�@�V8ÛR;�~j���V�N����Xv�'N�����U ��[����%�Y|�c ���y2�ք�k8�!f,�[[��2�7^� �a��4�B9��t�}J����[�����F���[��g�-�v^X� �ͮ�s��vP/���P F����}��dNp$�6�Z�N��P����W�/K���ύɔ{T��n_�M���cW~�~) +I�62�t�8y���=Wd����b���˛'�Xݯ8�͙�#
�34"�.Q�t�O'�j���JJcr�i6�P�u�gEo0A(���9ʞ�������g����}�f����q��F��*�UD~�����1rLȕ�;�Y�Н�v�oē��g2$6����+�,+ER��=^\5A?�m�*�}FZ�t�6�~d��H���9u��Q�[*9�a�5��
�q\e�6JԿ�����B�XM�����N��lRT"���e�VȤ3��F��o]�"RvO�e���UpD��2���p�C���TT�A��'،��kP�S��:Z��qT�4� �$�h)$�vv�`c���.mx�T���KL�/���A~�߆;G��Η}����o�/��w�߹���	dżqc𦃛h����Ȃ ɉ���͚\��+n�<֌����Jr�9��x��ڮ´L�3$3����nKe��8m�o8��Ѐ饲�:��GH��DR�]�O�J̳��fa}59�U|���8g!o�}������V.v?+L#�"5�����@��,M1�I]���%m�>=�V&�����q^ŕ����3[�X��>�R�ߍR����4������4	�(�����W� �>����5�(������")}��YGց�}$����>��@���t�R²�̦}Xv!�R)���#�l���B9�,�zr��)d�}
�\�kR�8О�u��>��t�6�ϳ�:��E�`��K��sW��оx;� �6d%��7�51
S,���r Ȫ��e���AS�.O�C.��d��M��>�����<�kź�1���+�Ls�j�ȣO�[���,������K�Q�fa�\����D<6�8uz���4לxe�g�9^�h�����Z'Ѽ3z
���o]��u4�6y��d�K��U�`�����׭�����9˿�_N|#�0�r_1�P��h!�s<��V�B~x�js�x��}7�M/��jK�r3��t�U*HH����[b� 1c*|�J��6��-g�����%mɥ�I�
��U.��COnHaۨ�zX��T��hrV�X��Ҏ����Av�bJ��qƱ�'>����#7���MM�Ry������s�f
B�Ø�F��p� T��;o��7�R6����9�B�����bY�cklp�de���5� "|�#�"�<d���B��89!��\�#�1�^"�֗[_9R��
{;E�S�|�?��W��ʧ�۞c�
O���4�o�m��Z J��Â�?�w��xnx���
���d�ۗ?��~�5�"��M�0��/�_�@��(�B���aM��ҩ�Ilᙁ�W�Tx;~^��J
�d��|=�m�����AL{����W�B�f��n0��~���UA�+���h�+X5�/r�.y���<7�cl�>�c��!C"��7577\KJ1Ћ�@���k���`6A�5#��i�#PA�E��)"�BqyA�h�(v1
ʗU�̈Rkb�1����#��Y,�bn���x����V{PX�bev�ʷ	!O�T	y^��,�ԇ�DS�DY�Y�0�Zĥ;!�����FW�q���:m��-7�y.��#KM��!ܦ�����â������Õ��0F}�M�%�L��Ĝ�aQ����E�7𼧺��{�eت*�ld�L�T�9�J��5�"��V\�Q� �+9���ڊs�98t�c?�Vl,�:.��|]C[�t�yMi�E����V"�Ȣ�K�N�U�0�S�#����HИ�v�t~d���Qͭ(v��a'�;O�?�=�D�z�V�w�DTU>�$r��]qmX��]}������*�\#s7�c��AQ\�wGR�%�Du���J���,�Oqs��%��VT"��wp��n�Y^���)����F�'z�+C�m[C�ج��j����I�4���sy��T�����e�*��l@%"�ݎ)���MWH>ug/�f&���Ψ��˕�,�����j��{I�lq�R�y8�?�|���������-T�hI�9j����.p~�~NND�4��=X��=�Bf��<�;�yۡ��[f��'�����|��a�9�[?9+?0V������Jbslg=O������AJ!A����<!R���IW�A�M<� ���m�ݚ�%c]�y;}��
j)��%|`گe'�h.��u�iQ�:��I�M��o=�?�02
%E}�M[1��l��"9]jo�N�����b�=ATw�W)\^,]r��˪���b+?X*=�;�����7&u�wwU�]���\�& �ⅾ#��3<l�~I	���ԥ��������Qw��o�4��t�&�����>�)~*�u��p����M��OK��� T���)[Ϥ���4�s 7ر:���ix�o�G+�r9���7�N�z�t��}���������I��c�g�N��C�#(K:���Z�L�#ֺ�SL�\Ɖ�� T�6����9�v-5'�#}	G�69O*����4*&����V�M@΅��6���kOi�5<�}�������Xo.@oކ*ˡ�����="�@c���4���"��YZ��h��Gw!�s��]�r�CO�Sۏ��v駶����<`��Z����<���ӹM@���Or�v"�.�!��?�Z-�ѿL��gUN��@���*3�"�N[��M���l��e'������sMF���#�`��S�AkKU��6�&��@�hw
#ey��b�E(P^���`$(�N,�wǀ�Nr��ܡ�����H�`]�8�6֔�j-���K@�c�*ph4;��g�Z�j��T����
G�]���������N؂B�����>!�$�t9�F���.�8���I��n��<#��>�v��/�݉Xd
��:��@��^z����1� ��Xa���bн����Ⱦ�K�9�q��e�$�k6���c�Z׏�Y�.Ұpٌb�== ���J̽i�H�^_ɭ2螻�r*D���D��흞>�0�Á�$y��ѧ�͜� ��7�;v!	%Rm[m]�ʮ߫w7U=��J�޶$�^��� �g��Rb�Kt52�R��1�j�Ķ����O��Bݙ�_�{%f�uN� Ψ\qFHx�mT�_S���,�b�	�z�]��ޯ���E���m�P0�e�?ۛ�:�ߒT�	|���-��. (�ZM�p,#�0�1i�,�yzӿ6`�J?J��yM�Fӗ�����Qv�t��OU��I	�&��4��CY��uB���%�Z�/�Ҙł�k�@�k�c*i�%[���ڵ=DX�'F���I�lҡ�!�=�Ԓ��x
`��~R:Œ���-�*+���Gox�����6�UC����(NC��eP�?��vܫ"����-�9H�Jux��.汘�!�a�'�#�n\:	5G�W�-@`Sh،V�2�X}�:�����A��Z�����Z|�}U��h(
�ȴu����7g�5S�B<`�@G��,u��g�OD\䒇!p#���K5��@F]�KM�=��W�J��V�9�b3'���"���ۣ���R�+��穳(޳p�j��9����-Iv���"G4ަj�d;U�|�$��/|�G�q�� R�#�����G>w�ܬ����B��*��zg��֝~k�I&P"`E�g�]����W��=�̓h�����g�m`���=Ad'��J��7�t!p@����&
u4�p�{ϑ<0T���f�Vo	\DB�i�7���.?���|��h�4���<=�d89��v٠'2����n�:��\D^v:������V��bK�Z��b�wD=�,�]�?	b�{꜠�)w��>�a�dn��F�'���(��rД!7d�-�Ƙ�'�k��'\�u!>�ħ[�:�q� �P�m������.�4����]�|�w�8�Ӳ&P�G�;�g_�?y�~��
I�S�WI���5��9�
�����F�sֱp5�<S�t�gŅbN:�S��n�C�<xG��t��;���s�5j��?�0�F�J!�r�iN,'Y1�7��J�&J44��}��o,	�)�f��:��
eC�sM{:?>xA��Q�����Ϟf��7{���d� ���`�B!���!Uz9$���<���P�>ڡ*��k��F��@x�C��k^�B�1ik '��K#�.�����m|�B�Q>�}>2s=������Nk!��� V{�ڮ�<0 �Ս��=)�-���E��aŭ��R�N�
�2s����&t`y�ҖQ" ��I�-���K�r �2�2M�ki����X,ާ%���!SDa1�2U�LV�M�������g�!A��*qo����ד��#X
c{|��j&b�V�RRI!�@�]I[7�ϥ�U
m>���%:�4�$n�.�c���ج�� C�?�p����a��YSϧ�2�{�	�Ё~�M�H����O{�[��]�b~Q��L�t��(��z9.�Z��5G�(n,�%@P$tt�'����7�LZ	��<����ʣo��-�1�����8M	���H)Sa�����{6@�O9�w�+�$��،��z����.��hHE}�w��x�9 ��2�;���e�j�rꃾ��|�}Q��A1i�m���_���HwE}qVO,4ZT�9
Cn���Lp��Q���g�>>d��񽧺����.�@O�XH�e�%M��V����?����[��!�U]�?�(d�q
���!C�MO[���B�7��H�9?X�xd�º�ո��a���p����U�* �?�!)�m5��D���'��6�[��!���L�k ��n�`l�u����c�t��Xυ� �%�]W�}nm��#�DH�D\�����Cu0�d��}zQ�T�˅~( Ը�����^��'��K"�~�7�(< ��� �R�Д�s	��A}D ��ca���y=�����G;�����zF��x�>,/�U�:�����yԃ�4c�Q��U��u?	g�Y�((u���#	�a��&	�ڭ�n� U���lu��Z����?��p�eqc�E�Qч��S� w���_td�K�u�oR�PQ�kwOSd��w,�k�ٻ���Θ#���B��� �61@�<�{"l?���XhZ;�m�@�7-�����fN~��;d1����:�/�\n���x⩑��v�Dͦ,s\@�?ɲ�ق���T�!���8ʉ;s�6R s�o�	��c��܏�0�ɻ�ϖ-dy���mJT�Rgu I��w�"��65~n^��9��զ����(=4�,��ő�U~vַ��wѵC`�Lb��7�)��Pc�'�@,_6�Ϲ*��5���c�i��5�.I�3��AWMe֝Z-�l��Ck��:N���q@>�β������#� �GNٶx$���4}��xw�A�M�&�'1E/��'Gnk ��+���J�ß�|��~�]zy�{�)��O'ixi+�����p��p�l>pA�_#�(�Q����s��X���#F��5j��u�B�f�]@Np:�/��B�:O[�lr�У��M���Y��c|m��2@���0y�!�=��<�UF�S܀���1h}�c�5gٮ1�cXL��BRШ��;ʧ�g�.UV�=z�x�Ћ��" �P@�NF��~7�&���V����W����4:.H��0I���G��ϓ`�P�rW����Ơi�_�o�
:	z+�0&����4`(H�8��vnݮ���4#��[����X4s�o�c��nV�p�e	�1a��v�QxP.܎�D!�.$?/GТa��;K���U(o�,�/�C��в��'m����J�?��$o� `�f{}0�ҫL�I�>��#��T�pċlM.rm�����C�zҒ���P���UiGX3H ������eo�3�vW]n�#̞<t{@�;��4�S(����N��s����PYC��D�,�T��M��8�E~?Î��R;rE��P�����$<� L�L���]E���٦5��y���yW~�y:�}$(�o���V��L#�<��:�o�U�Pʍ2Md�Hڪ�;?�"������?���#�[����I=!밽�Mů���V]Q3:"��~m@<~7�rI�z���g��'�� �%�f�Q�ZtÙ��఻� �K�][v�ҕ9U���5�xgq��ǻ���y��%3�m��u��j_A%����[$��R������ſ��SV<��9V��K�	�d�Q�Y����T��[�j���� �/C��; (�V�O�Bd��.AB����!&\]J�GՑ�̈́C����#b�OC	G�m%��?��ɧ�&B�x�#7����)x5.B��t�i�Ţ/,�y����B���t��E������o��T	���n�P[Z�Ń����3��M~ق��yj�6X+�~]N�@EQ�Q�CBT�3�宲e�9���s��t�鑓ϵ
\�v�����h2�`7�A�˧���b9���Qި?��8|n��Bn������%W3~D��9��RD6Z�H/�%g)�G��Bp�?W��u��1«�Ȓ���|�ֹ�-��`�y�N4�tz�!ߓc����=7�:	�,�m�H�U׆�l��FΰeQ�j��(�Q�%%�bz�ō�L#r��
�w�|J�<�Mpd����Yw�FTH����*E�q��_����>D%U����#4�J��d����b�"l���d7���w'F���b����mzd��?".Wr���C&�͔��Bt�n���N�T�pu!b���Zfw��VBu��╺�G^���!��/r�������J7��:V�M�?E�>ռ"�,�u_�wkZg/�-}K��C�7�3Ձ��
v��2_�
0���� �M�)M>��@7�%�>{*kp3N~�Ҫi�r���a����SZL����<�c���3��Aq(Ⱥd��<�\��3[7%�]����O�*���;A�����k�b�R@Wn�F�ߎ��A\*��[��;?s78�o�1oE�N�	$H�c�.��1�r�3O���,�x��f �<y��#_�4ի���3u���O����P�m��K|�No*��a���0��Ε4a�-����{�V�:��Q���q�nsSd��sg+�Ei�W�
r�";O"���پ;��-n��Q��#�7�;����X���
s�G� �,��S��0��z"�&qܔ����+��X�;����8��{�V$�@��������U��?yxh�E�m�Q�j��0�Էk&d��/���ϥb�,Q��P����"�d�g*a��E9��c�L�5�c���g>Q���>TwiL��HXJt� ��9����>ߥ�5������k o��� y8y��?s�F�5����E~�^��=�{�O��(xx��ន@�k�Oy��U��@�=�5S���9ܿ7ʹzQ*�pFO&���E ��貚��7��Tٌ?4���A��╒��5�`+R������=f����{�@f��d5�-R�Tv��Y3Ҧٍ�u�
2���=]��J}x��K�!G�tc����Z�����@�N�^FM��=V�L�!T"�H ��j���^�7�L0?瑔sf��4[SҲ|<���X]�:(�E��*Ϩ���l�8�KNU�3Y���5�b�3�T�0�n�T
�n�z/0�Q5��o�:_�:^"3u>�4�}�Xg�C�4���nK��&j�M[V�$E�'RD��P~��H� ��$ b���(�.��2 W�8#�Ma��C�|��g9�{�r�< P����0�@8j 2]J�:�|u�f� QA�`9�������pC�e�o�/O�XKW������jF�M��(�_>,���*dؘF�m$�S�j�^m��v�&ׯ��JG��8�	RD�S5�����|�^�_��f�W�ӱ�m�K��)�O�h�`���~�v��2���vJi��v$/�>��*ݭ`:���Q /z� �̣u���p�[���-�P����xdY���lX��)��0B����DJ�g���C�w+D��m��Ɵ�98Dt������aH}�8�	�N�?��˯Y��[?�Z�?-�w��x6_�˹)%
���TDI����h&������iNB�LX��5�Sf+��v�h�k�7��T/�^���c�tVd���Mqĉ�k���J���_y���}�X���Og��TDM#0��LްGK�"{�/(����a�{;9���6��~F��*�
Bұni�\��~�V6�������B��({��y�8�45
O<Ii�h'�E��b����W��p,�A�t��h�v�h�c�t1u�R�IN�!��]`��Z~n�pQ`�34V�Sm~0�����>BÆ���bլ�v��^i=��pgTK�G*yhA�����)�.��g��J2���ih�l��M��:�T��@���Ef��-�j2����$�:�!X���˸�)|��͸ڣ\�.H�I�g��n�JDÜ�5��C+���?�k1�R��e�~ӛ�/�?���R��6ѡ���<���ʴr���i�j���w��� ޤ�B���e+�Ҡ,@h��n�������m�KlN=I���R�5� v�� �0U#(� �|�,N^��������G�S�����PT�~	��m���K���U^=��N���/�с����KL���836=��˼���\Zg}��g������ܴY.(�7R*�mAk�.E
�XW���>�J�tu��GԤO�öhu��Pe��t�N�xS������E���ttse���C���b_�RKx�ce��~,^�`n7|y��+y���U�~uD\�O)��5|xhi<�p٥�[�8ckl�N�Rx����O]�:�kO�P��O!�i�/ս��߯�/(�ܠ��UV������X�t��bB)B����v�F�r�C���$F���+5����S��O�k��$:d��&?־�s9бuh�Ҩ���I����ɵ�����V�Yjj�]\`�L�Ǘ���֧#0S�AI|$+ہ��t�)�W�BT���F�5�yC8E �����b7/�e���DC�����{�Q�����i.n2IY�*q����$�W�j�\�������oI�ݧ)�g��G,�*D�b�vwy�H�����x�m�Qz�U�z	w�i��Ű�6i�Y�`��_F$�ѽ<6F�Y\��t��iؾf�qһ��{}9�+;֎[�t�v���ƾhy�2�lg�iV�����W<�z�7�	#�#���V\�T��W�~$���7� �α9���̞��W'#��j�YK��l��D�":$Ô��\�zX�pկ�zai���sDt��-B���U�J�1����B�SN7/�BX&}����[ճ��h�.z������Syg��,{G^}��f�����l?m��Ky�(�(�� �iElC,�$�zL��%SZ:((NW�E�~0�>����ŏT�Y7��9i��%��N���<�������v����U
�rJ{Ϭ�ǩ�AG�6�L��Zi6��H;�[���g0p�#��}J�a������D��q�.�ɉb���_�$I,Ǒ��A�����������w{�p�!n2�{z��F,c��^T�&�l�P�w��3g����=.�;]��Z(�WO��'��OW�B{?��ٝ۫�ո+���o����e��oZoh������΁ວ�SӬ��K�y_��a�����a�Ẑ +7�7P�?:frDS���%�7�pٹ#��ǁDt�]3L���v  �~�ߥ�����.�?��L@��a���K� hL�h#�y��
��5&���ܵ۞���t�*�j�hN�<w��,��}��i"����+�����+����E.����_��K��8{�gp����~1A����������I;������iB�N�{!�h5�M�(�֥{������7Ow�]���.4�������W�� ��3z;[2� 1m�e=h���w��J���T��v�<su�����
�eMP��zu�&9��mܩ4��/}�>��'�r}���cŴh	��ĩ���~h�ܑ쵸��@m����f]C�'1�@�pgb�9+,�9]�Diu)@�^���W�m�o1�t���]������4�6i e�#<L' ~���U*!yS��e�v��6AZ��\>��ݛ���`5-�9X3H�B�W^L��.�BO��y��}�]{�J6����J�:{#����\F�ޏ�}%� (���d.���H�z�y�ѽ����_�cU�$�h�yz�W>|��P����b�7�Dw��uHKU��,]����,w�%�q���Ojܠ����ư���ؾ�8�<�O�_���+v1r��VW�f�Tb.�7H:#xWu��ʣUa�� �ݨ����
���i*����|����}�Хwv����_��Yd@4�	o +F<��I�n��t|�On�������k��y�?^�2.�ui$LC`GZJ�W�XBT��z����<��m�G��/9P�y �&�����|��s������+#B��%.�(��= '�jL��Yʚ�]�g���k��%��ݛ�z�2-`u��0���w����XэD��X�W_�e�$o]��_(	{gk-�T��������0T��|�^y��`���zs)~�B+C
W�G[Wv�~�0Ug��(Aimucϖ���߮�1���`�	��1}�B�m9��J�7��'9�(lý�*@�%�U�>� g�0��+�m���	.3E��+6Y3�H�c��Bon���:P:��!9O����Cg7�P�@$`���U�o�4�?��D��8��vZld�N'^��O�`4	�+�(^�g7�٢�˺w��yӓ[����-}��L0��U�3Kx#&r��s9��.�7U�YG�a��I�-2����o۪(������
vK(X�F<]:�33[̭Μk�=�pj����*�4�E׌b)js�zIλ��ÂA�>ri�~	��>����ʙ��vߺ��'0�}�^�����r
`��p���%c���ml7�֊�V�l�������2P�R�R_��&���J��l*'.G[3]l�Q������%΅8RsCI��Uvo��&�C�6/�v-�G�=Z�}�rQ�[��-w!�M	���1�� �Im"c~2H�K�t��$m�=�3@����r%�v�]c`�c�}6���q��ZV?�T͡F6�m�f�W�Gr�������P��+n�+���}H��������pN-6�	ȑ�}�d�"uM���$?����5#�F2��ǒ(�1F�7a�B�(��jN��%��E���V��Ѽu֧��Κ뛯w�6\��#�R���I�¸x�¾ڗ}��F�!���㳼~�5��q�����*��h�_\zpQg��WD���gS�8wW��W�5UC�3��錙R':�p�w�T:n���������������jMb}�8yhڠ��j�ä��_��M𐝪2b�M��h���H�Yi��2G� �Tŕe�;��X�ֺ1ln�����c7��w��X��R�`� w/�L�SA��H-(3�0;��*u$ϳ\Mתߍ��x�\��v���DVXk�O|B�")6�]�Jv-�TsIt��AZ	xb$�'^��������)����v��*�x.Ch��K7�>dh��BF,:��Y���bʙ�q������9z�	����p�ܞ-��c��?���]n7u�!O��!�V��GM�D��,���ٽw&�Q!��g:���V>N2�X�#�P |�P��!��R\vʥ3G!��.5�]�@y̋f�;O�]��*�Yu�Gª`�Z��XnC���+B��E�nr>��2f��Zh>�� Q�0�5�'
��P���A��gu��%I^���aw�k���~%��s�f��H�y/�}Y-��G�g��"a�g��qI�u$6��r���W��	�t��M\J����\�HH)a�$*�vO*�D��='I&�1x7t�B�����(���_0/k#��x"�/H��L��}��#�s��GfT-aW��!��H���V�JU
$��-]��	�Ne"��xT���Yv��|����~yfu#���j41-�rʇ?������a�'�^�R����OE��3U
�[�(���������:Y�'��;.ˑ{��>����}��j❗��R(��]�>������*�b��Z����K_p�dm3�b!ܪ;�F�\^�ib�Jɋ,(	M�17[�3ҡ~�/�9�T=�98-đ���4_��Τo�#SX�Fh*�"���ϙoȳ�0���7��*�v
?,�����2lV�����f$�������<<y"gf���07 M�A-#z��3p��Σx<�9S@��|Ӫ���G㔇��u��e�
ғ��J�A��aPV?�;��`�|����,�vWf�~�����Ԡ~@ A�?5�/Ɛ��^V�7�E~�T{9�	MN��VQ��4Κ�Ǝm�uV.��M��D��u]�[WI�-H׶h\���P�LpJ#3�Hg���.�"Q})�Z����lHZ�ti�?�|#��@Q��|π���� I�l�?��+�����9K�0�%���X�W����������Nf������u�Q�� ���F9	�6u��܀Э����j_~��d�%QMr��h��,���� �K��xA�3��M�;�9�ӕX�^hr	U���H�Y�Y$���	���� �[�l��\J��d��Q+�3��CNW�4:������A��t�%�J�݂J 7���	0%�9� �.Ȇ�o�.�I������-L�*�~!eIϙk#A�j���=c)�a���$Hw�+%G�T�n��?GM~n���+�߾V���J�u�Ӟ�A��(X����bv�vT��u��Ia,93
��p/xX#~u��W��=�vc��Qׇ\��>b(ԟ/��fWF�L%���<����W�)���UN�_��;Z���mt���AB$[`�Z�:Fʪ�����Țxb���`V�����Dl@E�tk0:��Y;�'7�92F�H̠��6��W S�05ƃ�x��v<P海�F-���^Ór_�D+Ę=�p4�ۂ{����b�] �mv���j�dG�]��t����`9���1H0��A�"��$�o�1�B
Bi�V��u�J�����+�I�J��S��%j�b�B��ǘ�~��x�����>?�}�{�_�[������T
6#.��͌���k lP���P���d��?��6�([�C�"*�l	��dIP�~�X��5@�ɚ�"*z��5�T���S��.B9��B�'�C)رc_����L��whnxZ��@|�p/}��G@4P8�̞{��L%�"�*}׋�6۷ߴdht���YnJ>a�5�X1�=r��4pt}	I��=֕V��!w��*�?y��h$y5�ڽW���7�j�_l��<͘ԫ#m\��/F��|>���<}�0*^I,"E:5|�[n�3	��_E��1�D&1I�E�AR�Av�$)��k@�V����Y�|UdN͗.�Oi�(��������N��=�-����e;�<2���]��W5�K������X����]�g�q�4����*WEC�3���jv��2��.Rf.ZB���2�����jD�!{Ϯ�����(Bi�r@u��x�|$��n��_�[�:~����щ'J�a@���eX��vf-kig���ٱSan��QGQv�8���<1�L?T�A~������CX]��XW(��x�q�H�Ѝ��B�A� ]1,�y��l���:!/0<���r��)靏];�hP��#�Ȫ`�(͉oZ%Ă:$޽^��WA?]�0Ʃ���J�Y+ ��s\uwӣ�9��#�a	�2%^�{W0�������f2�>TP�y3�4�>	�K�h"���s�(�(��O���li��[`�[cd&Y��� ��e����C��ỷg�`ŚDy�T����z�~��L$	����iT��Tk'��b�� ��p��Q�	`���^3� �n�x
�[��䎰@f��#�� �W`+ք�8 ���<��o�a�%C�<�L�F@b�l��2Й�s}�E�/�5G�e��T��]w���wT�^e�T��xFA'혴�ۼS��A7��OC��]:#����py"
��>�y�'h��"�6 a��%����4�w�{���n�A�gj=v�4g}��9-i�����v���y�����1��*�P3j9� ������()=�?�#'_&��$UԦ�`��"��|��4���L/p����	f�d���Փ��Tr�8g�����w��h�4�=	yAȔHkR��1=%�|%z�3��!�P8�g�����ؿ�A`��p3uE�]�I�/w�]MqU�|6ӳ��к��K���>`��<�1�%�ƕ����)�. ��� �8����7G�^`ne��"�� �I�Lس���2~!�v0/ء�4�B�V�H� �#�zC-k�\�so�
�n����'mW",��4�҆d�)M��F�8�A�0и��?WB��+e8y��qBZ.�<���0�����!E�e�����}�?{Q�oG+IگN%��0��moĽ�L�*�9��Hy�W�,����Ư���m����6����^ufaU<��2*�ۚ�@q#Z�(i+�]�K��^��`��9�ak��!� ���^�5J�m|�N�*r-�t!oе{B�		IB��uu�D�`��5�U�e�/�^�Hv&)���weHs�X͔�7-��ׁMo%��t��)V7G+y�@�\4E���}��J�X��kc�%�T����l�F�k�g�<5|�CMbz�����DSt�ļ� ũ�?�3��[�)�~�GE	� g��"���
T��طI�P�:s����fv���~	ő?z[�}�o�A[p��i��Lp�قD%�8$0^U���#} ^�	�н���1��	�I��X�9Es�`���B�q�Kf`�u�1��o]��>M�w�F &{R/�L����ap����\��s$J�J���D���%�탟��2�s��Z�._6�����u�Z�u�S+u��-�<���**�qy8�:w�_�wx� m�3����O�����_}"I��eݱyz�����8&�?ڦp.{hU�מ^0g��
�u���uH�G[A�l�{/��q��0�;�����-`h ���!*�O2�}��D�&g
e�q[5+���CϷƎoX�=d^i4��i]���a=;*폑���*�3�zm�j��D`�k��`l�%g��ʡ�d��|B"�=��Տ��������ʻY�vS�O�h�yyh>��	�~�"D�z�rݠ/�	�ù��k���!�WX��W����K��$�+U��9CĿ�!eA��P.�|Vp������f��i逐���̨��'�ƅn޶�( ���G��TE�Q*�T����)���	����-��O�!��9�T�a���鍁����ے:�]{�sX�D�(8�:{�����u�wf��-4\���m����P�w3���?d�=�Pob�����ò淦8 �`F3O#�o
��ǳv,�g]��;٣W��c�0��p�Z&����M�m}z2�.c�K�==6��F�R��/��v���q X�#�~������
���h'��|�v+��LT�yO^���L��x�Z4�Yi������hdPL���be�|T��r��p���]T4]�9��~�Iv'6��RH�`���	�1,�d74"�s��j�R4��k�P�/�P�0L���ٲ4v��������q#Yr̘������J�b/�]�����<��f�:��*�~���0�Ր|�l|p'�l�</�p��+n|�s��Δw<}��C��� C�'�9T7G�w�.e>�8Ai�R�d:8}��~�-�����=�#H@G��{]�mfn���ۺ���I�������}�a�^�q��Fz�#QUD�F���II�.��\�{���d+D�~� y����Į��nIX"���8�ؗ�Њ| �����W�/�ǚ�D�X<gRL1{c�P�|}[0ك����(,�^�;~ϤZ�x����R�Rp#�F�
"����]�	�I�gf�|�x�I�Oo/_�̓�zuܨS8����o�廍SJv�;N#_ �小˗��v-�H0p���B�E�Z�`n�����`@�Z��+����b���ՠic��ӓG"ë�+,JWũ�pyF{�߁�p�Ӡ��4�b���K���̊���K~&0
Ͽ��:���%ŠMD���gm�x�t�*?��~�_؈�I�;��[�W�!����:84�)ۍޅ���m���*v�֞ٞ}9#��6x��Xn.�y� Ŭ�H�\�@�gU����YMoc%�M	�j��D�"��fzUr)��x�����Ɨ.E�J�U����,�eY�P�� �/MT� ��N��Y�:,4{+���'j}� c��j��ry��UbȾG	p}�`�(aCN7]�[�9���.�[.�'FUf��PXѕJR�(ӛ8��C���ilt{ Ge3���D �]�XߤН{Cw����>A"Wi����ߢƠ�wO[�������K ���,�j8]�5�oz�E�2spp1�T�'|�>͈����B'
��y���I%g�=�Ҝ��j�2D�H���F`������5�kk1}��%m@����j�����rd-��w��#�*�}���H��Wy��*RGNm���,2�)g`�kR0��c���c���]{S����6���΂5�!��5.g���g{�yX�燘��9Pf�Q,8v]�"�m����\W���ĵ�����,��ư�8��%���<����"�+�,��t�j��̈́6<6��]�JVѣ���LZ��2EH,��4>�,��Eł�eճU7_$.�H�6��}J�$���~U �t#� ��\:K�'�D�`�{v��+���b�����(�j��|��/��K@��%E��^^W��nX�r�uYlͷm��S!��Q}���O�JX��}��TW�|�P8�r�@�ȱq���Sbn~�*����:�n���\ønJq̮��K���P�ַ^���
��9p5*��݆�ԁh_Q&��F�O��`i(ѐ�A�QaBm6ם�)�s0sD5�AT��0M��I����k����a&*�W���s�W��6q���n;dd5�����0qa�;MH�~!Ϻ�����{�r��Z8�ܨ������$�ܝ��n��Or_)s+=�Ɯ�y{"��g������*�tb���je�U�3�js^PƉ����-�����PA��y�D�-����"�7\�إ���l:�F>U�DK����ٺ#�[��Z���a���u�Z�%��B���S�4�Ukk�'$�M� �+J�]�4�R}��*�<�:�O�6���c�L"��z����H�	�L/���l��������D�U�:T�� ��8�P���i�R5{�5B�H�ɤU��2��%��3�`o�k ��H��{Du�g
jeS��mO��.�-,���Uʾ�������:�2�/uݬ7�ȑ�����t�o��A����*�=m����/}�*֨�,J�D;��*l��/��T���$yڄ���g���p��+����)��L�OL�A�ψJ�y�j��x|���X�^<�*�>�	�DQVX/0� P� ���X��h2,�
��ޣ��hp������i4ozS\>��J���'��[[#d\]�G��@�Rl��2�5�@�i�UNS���H(�/$�{B����A|(��L3t���֩Kan.TuAh|_�P!;�GW��C���c|m�a;���I�m�xY$�
b��7�EBhi�QgE��e�A@!(j42��)MK�w�ޤ�ۤ���R���Q��B����k3뿿�Q[3�%�l��^ND�W�0t*��Z�*%�[}��]�m�ȆۧfO8ǁ� I���Mf�zz�8�N]���qr� �3�������1p&�Ű��Ij��u!���o[�K�L�L�N-�����inM�7;��lϧ��#0#������ ���_��zy�$ �ĉ���rU|�� ~���
��%�;�Q���~��}����kU��ۚ\4�*��P񳭲�^߷�m7� � "�ع+0G+��m�a�緉�5(8�(/ĉ@2��:8������r؈�`�����w�F��gl
�Q5�l'L�wތi�P���Y<�d�F	5{�lW5�5�üh�����͋8ZB�	��5]g� djz��B5��^"�*(
ⰴR\�lTw}xĚ⽲���Z�z~p���	.������Ow:Ұ���i�RQ*6>:s��x�zBT[�����)%$��{T���R��q��+�p�j�MF- �%mz�QZ_!��s���=��!FV�������h�p�K<("��?��F��T��[�]N)J3>v�Ӵ���L����mY��8�+�E�\g�mhet r�C�$��7�EI���4�m�Q�h���ڟ��f50����,Sq[0�E�����LG�Ch��JPH*�%���ݭ��{=�!�V#;;�]r�7����@֝H��BՅO��&����F;Z��8�܃X"�k�wAf&?<UH���O�J}+�����9N�5Ka"�m~�4�Y��M�@U�,�`M�1��T�8����i��b�S�.4s�OӁ��sx#��~��!��b�*��En�h�Ct]6�?v����B~���w˦=�����$��5م3��/�M�j��C�srpx�<(�uoVi�P}����X�˻��Qjg�V�Ԝ�$���Ul��ر���8�<I���a��]{���Iв
��miƐů���H��J&!�W��׺�h%Q�����^	Ѷs����_�����.�g"���'j�F�BUSDk�-�B�M��V\sg#���ST�qZF/�aW`*yT���pmhW��z�u돹�_�³5�N��"5d>|bԃ! ����~��}��Ra*m�����ū�����8Ǧ�Td�'��15��ƯL�`��7^����䒆�%}5r��&v-���O0�;KY��ׯ�(�!0q�@��ąFہZS���=�%�����C�8h<O+S��~AԱJa��r��l�{����s���8/K��P�!��A�ؓ�#�NfF�i��9��g7|�8�+W�z���P���:BȔG� �e�����,�nHf�W�:��X���܏��5��)0�����?���I�Ma|��j	�X��?'n�,��\�q�N�<w�O�SF�����e����p%x��+�:��N��kz~2�J��/B�&� �}�>F���"��^I+ZǍB��WϮ�����8�7^��X�b�&����	V�m�4���X�e �E1�(
�a7�r+�X5QB����@O��ە��T�:|��gh�ޔ��"5RV�E��'/�,�G��k�x�d�:8�qU�i|��C��j�S�OȺ^Iig$c$[�.�8�UغJ��Ml�QL�R��R&3��S�iՁ����CӢ�U����#�N�RҐ�ě�}�s�R71륳{���������	���f�*��q�[).� �6�A
����*Z?
����U�>I�\$�ɵI.�}z�
$��"�\t8���'���q�������T�NG����<�⍅Nn�9�2�L6����o���2K�d��=E�>:~7�K@)�f��KQ-E���P��Q���A���p�wh�]%s�[�����A��*�U�*b�$�\a�ݒ�[����9�1F�56����bSdЍ�X+
d��������(_R;�}˅->�"#4���V�Xs��?b�X�a���"w ���R4S��?j�lM�M����/�5Ce�>�#���f^X5� ��~'~�.^L�3f.�=��8s�` E����H?�B�}G&�9��q��@���J�bӢ?r��k38a����y�0]w�JCr��<��m�(V�'�6�>h/��,Gy�٥�"R�Dg*��'߼����^u�(	L����oX���Zis����O\�^�yy���RPۊ��V�Syb��3O���Ս�
N���C��T�a	�,?h��34n��=��-
�y	�
]�*�$n�]n7j�,ʾ�d�PO:��#Η��+u�� �*vx�DZ~��QAMD�Vm\*��>F�y=��
El׮��}��D�k�t�D"2"2���X��/V�]v�Ȁ�珩���MV���)_��͠j4�+�V��a��"���hkӯ$�?g8�Vsּ�Z�c+! ����Do���,4�_G�͈�4w�^r ���FhӚ �gw�|R��zܺlQ�z���M~�G�(*��Ν8���g�i�z�m@ \M�)�wǣpЛ0m�W�KM"����om���p�x��{2���z R�N;�Aم���Dr<k���C�2�h��.lOCD�^ˈ+u��9��Nn�^w������0zR�6b��_[r�T��	���s�o^!��^{l��6V�ty`H�AU�(�[n�����:I#�������c���-ȉ�/lk�d]�V��^�<�AL  ������uO������ʃ�;~�/���������m��*OV��C�����X�!�"+�Xk���z����̀�tu����
�9J��ͷt��g}&��0��������Yy-�C�Y�Z�H�Jo�cB�p��f@)���"�������Qu����L.��Je]���W]�Gs�2�?V	Z�viCJ2<!Ɉ��zތ�o�O�0_޶�m�t�W+����~BQO8�@e���Q-1g��^�ʹ��ۅ���Q�h+�����ii���%Xs%^7*��j6/CXR�ǁ׎2�V�i�v���/�VjU�٣#'
�{�?�P��fՋQj��Ud~�����h���8�C�(��#,t�ےgN$�b�w��$j�G�:nE���[l\��c�|p_3o��7��X��wu�\Y�?� U`�[.�X���W�@�'���O!��&�����k��D['��_}`1����Uy=HE��"=N(2��:�B�7��BZ���\]�E,�po��(SC&t;I1{��F��}�tԘn��RO�Aň�EiQ'"d4��M#�Cv�
�Y��um��`R�.Z�|�a�������i����r���T�D��h��LF�ą]�4��#|� ��#�|�>��C�k��,/����E��[&Wca�δ�α�|���K�d��`�}�+�N�`RAN��޿�0� *9� R�_��ŹH$5��1��S�y�b�ʝ(�3ZxDC6�����a����TxG�'��X,�h@�w��M�J]��)Y�pm�ѲK'�G��[�V�5|�5^�����Ŷ���X��T�?��x��#0cQ�kbX�2k��4��*6! }�O����R�}�K��]:��v�$X���y�MT�>]�a\����8g|wI��WK�~��E��}�7&]OV��/p�3��]�XB���v�D������n��\ن��T��gZ��8�C���Z"$4�8���4���)��~�=C�~�9�e���$��O�83T�m�k��
������|�?~P�G�f��\�0������.�[pU]j���MQ�C-�~����"&#1��)�՛����>7e�Qy�k�#:�Z&��'P �Mn�^��
�U�a��%��@uAN�e��j�!��.u�H7��q�B�W�{���"�c��7�vޖ4"sZ��k�h4ë%b�Yla�����m8���s'�9X���>�H�؄�=a@���.vnܤ�j��٤����~�e�Nh7���r-���q�={�M����2�;=�)����2W��!{�V�l�=���-#i��'��ڰ�<����A;�(@������:���	�¯�RL��գX810`���Z�s%�%�<�x�f6�s�ٲ���4X("\F�u����x�hm� ����e�ņ�����ѫ|'O��/�����|.�a���� �|%��P��'��<�2=(X�z8�#	���*~�^m��𤱈~��3��@>"���M�)�%��űp����;���`b����h ���,S�c�L/+�� ^\��7�!l}:���IP����Z>X��y2�u�Cu�a�v^*�%!��A+�*��A[U��Ç�eP�y7�?�Gߧ�*H� �13(��}�Ԭİ�����툸�Eqn=D���J'	%l�?ثf7��d�?�ư:y��Ig������K؝���Ǆt�UMj����5#�M�\��zb?OFrB�\�P'b�SQ��"��
�h
d�WM\u�ĔÕ�9���ǈs u��.��l,��sc����+��:���(�W�K�c�xǑ �J�_�b�h���2��]�A|�D�����0a(���Z
�Qa��^c�P�2��H�t��ȳ��6kz�0 ��rK����+ZS/�I�uf�.��^l7N�p�	-f��cŉ�F�$��B
�¡��(`����D�2�S�;����p�+��ZQ@�}Ey�2|�m�f��>,���t��Cn���(WP��K�a Ŕ��׊����R�.���o矽XX�r��*�'�~�#�A�����t�I<:��&�Өu�;�O�G�:���,��ƣ�j�8���)���thx*���M��i���9��p��5�`!��s�w�

���!�Ri��	�h*��k�*N\\ƅ���+G�<Z�Ѷ�5�XgK�/�~�1�ε �_s���h���9���dx2���v'����bi��`n&>��Q�>�o	�
s;%����)uc�*㺶@'< ��͹Ӷ/7N�?��?7E�W�u�u����D(u�2�/�&�g�[d�wĄ���M谈��~�;�h{�\Q|D�����iB���O���L�;�����Pu��gic���棖���p�GȔa�M�����H��m6�se�`����Vx o#��v�^�k�A��q�HhC}��W:���q8_X���,�'�x^�J��[�1:>Y-��mi恀�JV�2��i�?���k��e��z��^�%4�w��'dT�!\^؀��{�#�lѓCn�/���#��\)�GF$o�0{��V�z�-��1+��S��g�e9�F5%���E��ٛ��T�2���t�S�-C6��tF���	E���7���7=�"P�ɷ#��K�@�X�̠̀dg��}m�O�Mf�<�e��e|�� �,"?iP���@K� �Ꜷ�ҫ�!�s��:0�D+�nB�E��yl�L���Jb��rF~�+�X�+"�2���)b=  '��WF}%mE����'p<Ql�bח�j��B	Dۄ�`�>�IC���̯��]��v|@�I�UY��~����	m=�5�-�WBw���a�0�1��R��OT�S;a��t%����ׯF���g�d�J�̒�IR����S8V0�'Y��eq���@�F�vB�F$n]
�u�4ڊ`�dj,�nб׺����X �8��蘿Sx|��9Os��N����t@��/]���%H��IQ@�z�Pf��{��
P��K,�\����q��8|��j�O��k��,|S�6ۖ=V�R^].�S/����$J��������W�E�_0�\!��v�/#CRj�����j7��7)�`�m�FHF�T]��� 3t�ZE��-��z�Fr�6%jX�rR��1�{y�D@F�d�at$��DCl���d uMb�X8^��|Gr�'S�B�Ϟ<��L����TCc�OVTTX���:B{h2`��k��w�c�z�j��ZW�����A�1�C����%��yc4\+{a\¥K&��ZZꂊܥw����[�*��ڷ���6�⧎ QQ�m�;O����^�l�?�My�!D�I|�ԏ��M�����?��L��,������4۸�����V�M��W:�ȹ�T�\7qn3o�$����@��rF�U�,����5�Qz�Ӈ�⚕ɀ3�z���P=h���i��
Vyr�ɥ��d��KQ�*��l���,���!�A}r��-p�)(!�.J ��
�$i#��x��j8
�{Ҝ��L���L��JKr[����$0~�8� W�]m�	��g����9)N՜�K�K�*Iv1��"�Vr"��<��s�gA���`4$�jA�, 3�~G;e�8�f�&�!�`�����@��2`�x�i�<���RЪ���Ӊ�j��Ě��1�O_	�ѓ�Ά�#��c�]]Wn���4��p�X�Qq�J2���ۖ�?9���N�1ю�kE ��]�qV�l&�D&�w 3)~�[�uԅ''�|�?TU�a)����}Y��UdSE;�����������p-@�y^��Ղbk���O�ًL���������9�PΜ3v3O�C͂�_X�Z�ڧ��CĴL�H�������a&8�$�:�̮4A.�f�c��n��O+��v+1�wzG�e��B��A=��4yO����+ч��?�KfJ����yg���q���}&�nUH&�|�,L��]��o�G�C���<3���:�&�������!�A�9��0��2���_�K��Vb��ql���KӠ
�A��4�C�g�ݺ`!����;�H2A]�4�<���~#rlt���*��3jo��,.��Ӝ,�e"�j�띷E����e�sg�Nޮ6�\6��>����7���D1�
 o����L�^�N9&M�x;����M��n�[�If��M�}-`�P�O���!`Iyޣ�M��c6��Qs��]B\ڛ�V3�5���C�`��9��Y��}��I����'�sV>k�Wk��d��d4<�rC�堬�M�t��0I��oD���qUS��U{n[B�Wf�}���� ��:@��4+
��^�ŝq��ù%8J˗�!w8B�l��!C�B�G`�wp<_��,8�u@�I%|M�����KmFԽď�'T����P J/%=����N6�nd��t�-�~�����k���� 5�V�/dR0���Y�&N��Ĕ��ek��߹hV{�`�d#�}^NOe�}�h�ĳ��~I�2�����&PHe0��L�dI��q��/mbG��i�A4�m���b����jk/�b���^�o-��ۏ��{=��V8�����˟�r�ܳ4Z+����Yt�j��F��8C\ϙ��yX��iz�O[�i��@�>~�z��fv_��_[OM=�:Fb@uGP�#5�������*�	 �`1ٸ���ؾ���_x�5ZG�1T�H�a�e��ɳ&��[��]s$2f��2�!�L�>��B�v�z��g�`��[��]�����>~N�ɂv�RŸ���e����,/��L�����O��x��|/Ł�� �e0��@$B��^c~�E��Z�u����{o)�ڸب���ߑ�v�>t|J�!�	�C�_��J��x����"��;n�Y#~ZT ꯟ=��X��D� ��h�f��+Q0����vpMK��$\�Er\�P���t�n�tROJ&o+��y"˝GEh�K�eKG�t��wc~��^$.����/8C�y-�NX�+��zdTtg'���]��PȺ�`Bi$�;l�2��T��|�2o�
��f����1d*�(g�*`}*X+�	�N\(U,��Z�^�c
]�9x��x��& ��VF��c�x��NA��&�����랄���K����=�7��GH7X��}X#Y��~��+&i8uo0��͋����^��&v�p����+�ߣ���_<+�\^.Tlv����D��w����0������Q��a�tD�����ICG0�jt�Ԡ<q����,Ϸav,����	��rU�"9��O��c�$��m��Y�
Qtm���ߥ�C���� ��n�2�v��VX���˹$��f���[k���6s�g�q�b�Wnc�T@��Ѿ7,]'��#D��aƦKW�ʖ�jJh�<G�GPf3Fc��R�{��G�<*�{�k(�=�Y�v����e���W"�Eg�6T�l"����D��c?�����ۈ�h�#oڍ�N��&�TL`�{�u��Į�z[�"Þ�G��v�\�f�8���`b�H/�$�P�K��9�Q|`�:�nt��[�>[�I볒蕴��8T�����*�#���rr�9e���m�1����Z���0U��l����W���i�:ᨬ��I�I(R��|�fq�(�F��}��nL-�刵kE=p���]��&:b�yJ�,�1w��]-�1Z�l��(���T�&$6j��O�>P�DB'����[{p���Z�����P;P��Y��T���9�sV9 �/����옍�m:�d�p3�����ު��I[j0^��Axl�.�#,�&D
ǆM���R�+�@�j���+�����fSG>�m��1[��o����\�����M��㺱]�5�� �zc����Il�e�Q�U|������d,*K4-J���0ƶc,���9��\-���ٜԀ���%���i�$+&�Ѩ11X9�2{�a(~�d=�x�W��5�U���*���p_�������=�TOu�&@�CDͲ��y��f�H��cO�ҀKR�wA�Wm�D��F,��t\j!6_�'�Y�E��QH���SY�)�c:�=|��� �y�- �z��[f�lkt�"��}��lsf%2��)\���'1���`�\��J����1�d��{Ս��y9EeD6��3�a�\'	���$hfD��u4I��z];��lr�;�u���d����"�:��]�ɤY������{ܒv �y���V��&����'��o�__��A<,�#<g�tռػ.�r��%%��qѢx�� ��UU�i��+g<��z���G�]FZ���[��ؼ�<n�n�^�}:z����iB���x
���T3���Iq�Fj����O����l����te�s�����a[�W��p���̮<fy�3shP�κ�q�ʟI��(kj
埪�y (֞����)O.�U�q��K�E�_0�\����O�V'�v`�U�u(��3���gQ��$�L�i}=��Ŵ׷�L�0�8�(�q8�!�x��_�:xA������%���щ]��|;;��K�B*E�$;�H%ٓ���>�*eL����i��gS�mz����-���t%L�^�ȋ��Q:�Ax���ok]j�<M��f%��Y�� A�!��^H?���_���pA��<wS��<��|���Y���������3�Q�#��!dl��5"�k���=oRh��}2Sg�F�"7Q���J�__��\�Z� �Yf����78��i'ZVIe���B.���-�'�Hძ��o�������Z���C�DxL�X���<P�sST�w	�݈�9v��VH
�u�(Q�����p�&�@,��G�")[�3H���7����h�W����}R�%�2-��F\'9��ܰ��!���]H���p�����YT��Lۜ@un-�M��jE���!�/[��,[������h g-���(��-��B�_��A�g�g��]�}��
q�(��B��� 0u�� ����+3w$���Q�����**�.���dV��$Y��I��xq%��R�t0��gaΡ�*TRի!�_���C�jBގ=�)����'Sv-��Ǹ�(���Wqj�Ȩ��9���V�>�GǄ����O����2�(��z�
� !4o�s@�_�~V�,i�Z�K�J�8��21��=�j+=<���鐇~����Kri�1DdI�eQ��`(����� �Ǉd�]�4�'��<��ܹ7k*�CoG��Pc+G�F���mP,��ӱ�/nU6EwȪ���=���0���1����7�=���Pi�?�J�'���Of�G#9r���-�F���p5��&�E�1�|��o��0�s8s�J�ÿzjk�K�X2��Y�q���ױ��@�&�Z�J:�z���:���1��[�)ui�R�����k�\+$��_��D�T2��R7���H�[��Q+]�Ĝ�BPoBUׁ��G�� ��˒[�ܫ�;�9���U*%��5���*&S<���N.���u�ke��c4b�i&�r��P�A���\��ō%��qԴ�t�[�"��0��v�v��W�,������ҥ��SN
�u�f��5�ʾɥ2��Q2}#�d�f����]�҄��>����v���t����M��:)�����lչ�Z��]���CIQ���/mtZ��	����i;f��ẃ��gYG�l��1�p��F�#�E�}����!�����o�X��}-rC�`�����t����)��2�n�\�d���gR��.�C�,�2r�4���i��w�ō1a@-Y�\T��a����Qi�&��{����i����{`X����V{�l!��v \�JT 9���*�6��rp�~io�4��.���M�,Z���w��܆J�Zt�=B�,�k=����ٔQ��"����G|�a(���>8������[�������ff ��M#\���Q�b̭5ivKk����A�EO6$�a������R�T���n0�nFS��l��M�ZGF�!�A!L嗪�6_
�h�)ab��zfB�80�vt�ӻ�]�w8��G:�p�� j�UO���d��>�����)�[y������������ �dQ�!���?F�c�q7�x$���s!��s��Z�ٮԅ6��!�kָ\�-�� PjEj����g&b/�f�n�&�h�֕�� 7��T�"Aw�㪮X&s6W�����^~w)gi��2�����$�AT[{���2�����v^ũ�T��Iw�s�m?���KD�"�^������+�;�ct!��
�ȧ1���0y93������T!�����"�$ƚ\�\,�[��/�M� ~#�J������� ��IpJ�5o,v�¥W�-�\v2���;�nȘ�d��0k�uE�Cس����]�R�i�8,�!�v��Α����ͷU�T�7Q-L�sԇ\��؂:/̺��}G�����,��u-�
����X��D��}2�8���c
��i;A�0��y����Ag�
�:��|�6�C�J�@�3��z���ljw����_fs��or�q�"��Y$�i�ot���'O<��Hd��$�겑���($�33� �	�i�E���>�^�`�K煂o�j*�o�u�(ӽ����ClU�􃵌�G��:��1,�?|z3R��8���,@�m��ͻ�c�䯠p����2҃ ��m����͂�O�~��e. ^��E�E��~L����������"�tq�*�[l��/qk��L�N������Z7�my� �{ �t���eKm�X3��=���6hȮM�&������ݹ�G�w��m��?��'S�Q"��vʿkHa��s+}���r�z��&���n:�d0��>�����C��CL
��P�a�{vf;�'��>PV�B�.���̩�Pɝ��g:Z� d��mB�T���A�-8X�7��N��rg	s~�����5*	��z���#�&?�8eW�H2��y��S<ѵ�������#"�GYa!ss�E�L����GJ����b��ڎ�����.�#�~T�\�Ȑ'��z�`%�@�\'���CQs�J�}S/kY�sx�jq��UOUZ��|�A�@#�,Z-/���h>�� ���ɂx�KyH��筝[D��U|"���'+��߈��"HA`#ф߾Q���yU@�ĉ������Oz׼�G;��=g��i?��&�B!�1C�8�M��_���b�k�t�O�\���B��*-Q4LR������\Uv ��;	ҘJ��C��@��&�&/�m�������(��<Eٕ#˗�o��&�~���--�T~�.'ʮ�z��#���^m\��w�"M�c�y<��qO<*��{����,wH��$x��`tmx��¿�ùk�V̒�#�oa��I���a�|Ì� �I�.�e�(,S����&Z�|z��q�U5;h�Ѻ�)�`�N�_��ֶ�j�j?I�.�w�%�v���}2h��5:!
��:9�u���3���Ó}� a4�{M	ST �Q��2^IG@B�(x4IZ���K�Θ�^�\q���4/�"C�]��G��Q�C"v���E9�����2ȗ�0��3�fg~a�I�(7Z�۝�=;L��F
#A����*[�!h&
������'�f��c��jF~|]�3���"�wSsN��R��[}���@��
�������EJ	��v��b?0|���g6�wwVYC?~у��s�����Rqd������9V�ȍE�(+��x�����3��j.��^X)�O�j�@�t�����Tw����u����0�rCl�!	 �0Czo�f����`,R����c4�v,��Y�m��T�F��k��4S��<58�u��������z��/��/�v!j_����x]���
@<q�U��� �5��,Ai��#�z�ۡ������$&ێk�V&��i=����!����[�0��J��W;���B�p��M�`�\�=抐uDӃ8{�1�B8���0i2qmOu`�7����.�y���_�@c�6���x���Ł���US+o'���e�CNm�rv	MRW4�8�M�-�����h �:ڰ�½�qdz��:���Ϩ)��qJ�
���!fwB�ڵ:��ܑ��J᣾�����4���FN�ژm�+,�)��_<@5f��ix�C�6���n>�v�\l�I�]��t�Q�O@�"a��[ؤ��eԂw���	��jqM���)`�!7Ӡ%~jC���Rjonl��b"��L�{+���&�Z)&����G�Ӧg���9^e��a-uk��̒�i#P�a3���Y�i��s�K\���|'��%Qm���T���=Ӹ�o�"[4M�꫸Z��R�=ym��wx,}��Y�#�E��c���Z2Ŀ&A/�$��h��3O'�����q�.RO��Њ4�wz>s�3� ��|[9�}F����iv�����<oK*�p�����K�0�rO
������&~���wfhᶢ}@�6~[dN�yU�t����N�V�O��%��Ra+a�>�@��G�e�'vʴ�Җ_�ճ>7Z4�Ie$�g�}3�T�4U��Zb��ʥ)�wB(���/�f�*b��S�c.��{m��.*J�~0��Q��>��%P"�G�f�,����,�KpT@��Rݫ��(�rB������G��V�C����Q���7]�۳���2��?��b�M:�D����'AB%����nZ�8O�\�4��n**Nr�m����9�jy���ҔI���?����ˢug��i!d3FX.�-9%y,6�����}�ۚ�u2�Ĳ~6�+�Nr@O��Y�v�M%��?z8�r��� �'��XA&7�)��݀c���R&csW���S�<-��Dt�L�f�!�)4~�"��ӴC�(lA��N�Xq-���E�~�Z�o:�D�*�":Єȟ������W)_3:!3c�Q����]��@^��-`�V�t�	�t"yHT��J`���A,Y���O.%�/�G
=��`��l���f]�6>�������*�8+ة!�ڡ�_;w���-1��еY�d�������4;���@ÄA7�$���I��9�`B<PO`Kplr9[��+��#5	>bdKͬ��܎���T-�m��v�����EK�䅕�m;
y� ��A����PEUt�/?<��Tg�10��"tX�"��k6�<H�B:��[0��j|s�ُK�i�b��Ϫŷ!�O���ܓ�2�Xߥ-�J��>ny9;0���ɘ��f6��BM>A0)�au��\ Yw4V�|��*`p?Z�	��\� .T[ �cY���B`�@�>[�"��&P�%��So�N��Wd��ޙ�+��6���m�3��_�<-q'γ��3��Օ�E��6>���!R���6!�AN�(��L�)�V07�p(��ܞ<����C��[�eR*����"����>����S�p� �D�pv�>.�WG=��>`�P���3˻fӬF����<��d'�g?���'$m��)U�AM�{V��M�-c�w��aEVᨦ�h��Z����B�z&�����,J��l��:�]�8�j*1�'1r�qٸ���7zWSE]��Zwp�CDH(MVל����s��>�HՔ"��Sx�@�Ի�*j�a�*�n��>�YV#󗧣�
H5 �<��c��U�&��<������⍳\s��G�%�'�0Ȍ�I�BK��V�o�@C�3!
O�y=J���v��qF�e����J�kd����ᠭ�w��{�Ȝ#�[L�-�ω�Q|�:�j�wH����Y�ґ9�~0U��h'��������3lEn	L�u���`�VUZj°�}5eI��~hn�:��Q[m˶���K���L�/�-�/^����b��1&ߵ?1Q��C�����0~���M���WX��s�̍�@����j\�0,$�qta���j�8��9�
��B���!Z�q��-�dԙ�h����G��@���������u�L�y#\�
��{����$S�c�X"f�����JwMߴ�^��|h�إ.4e�7�+
� �w/��6�I�i=?t�x��,�/�`��k�єx��ӑ�$
�/TJ�~iZ������W،1Xsz�NZHN��y6���+xتQ��A�*;���ŸmZ'�ם�Y�a]&�X�?i9\q�#�R����.鑩d3	&-bF:x ��F},��KO�<�<3���ɁsH�o�P�6�D��mOF#Δg�6���7v?���c�^w�n�M�Q%�HSf�#5�����SZ�'�G�UF����P��:ݦlz����#��NL�g���F�#ⷋQ������;�@4o���T-(�uy�i����.P9l��H�$�QT��9	�F���5*2K��Ih�A-f�)%>��(:��/w"�G��X��A�ѵpd����|�2���b��;_tV�P����|@gZ;j�Fn���V�O0vs�}���[�D�\�����0p��Q�����9�{�E�1�R�� g	2$漁���x�^~��Z�;�YZ3�~�
��t�v�u\.`�{|N����8	K	�=����0x���Ρ*���}�D�`����ߡ�zS`g�]�1Ohnog0�=��iهZ� ]�sH$�X��tU[C�Y=mq�v0���Y;5G�r���fb�J8}�:!J����uD�.�U�0����#�VX�ɦ��EQ�/��L"��ɺ���]q��S��Gͳ
�F5&Xg�f�ˋ�$HT߷;tii�h��a^@ZDe�l�J���N�Ub� �X�.�K�j���rlye��VZ�
�	��@�\�/���V٤��QOH$��s=���_��=�<����{��d{K(�߯n����f
Ԧ�-�4�7n����_����j�'���DG䡗줺�jz$UEm���'%1�A��e�l��|)	�����N��h��,��s���i���0p���'�T��e2&��`�ش)�~p�r�Co�`�D�+�^�vKb��8uw.
~X��6��	<�F��6���#{r�9-/7\�CE�we������u�kÁ����3)��ndR�Ml���t�=�0$����F�t��t8jPm1��wUPE3�ْe�����|�f��\���������gL�I6qq��?��>m-%�gY�$(l���d恨�C�ּ$�o�d����^�+�tȉ�(�|h7����d.��Qq�rg��+��sۓi�B���A��b4�!�5Z�]@�ܕ�0��=R���g��,��^%0`�=��CX��]�Hu��_��m3`��*�<.G�6�[�^��4��Ñ��1�>�\�~��k��vW+�����57�Ğe]>`�u����J!��c��N��wԔLP�i*:��w��\�UG���� i�~ V>e��8�t(�Ӊbw��
)
ڰ,�:��?c����xLV��¹��Pb�9-;"�`b����{?D�$�PGZ���k�o��0��j���:LՅ�d�b��>����0n?�+���4dD�f�}1EE�+4w��֒���n���^�0L���|Ţb	)̥��4�� �x�Y���6C7���@�>Ц�~�]�|C{�Ww�_�HG�A��7������|I?�r�E=�0ic����ՇoCq�\H5};���Y����Jm�����(�O�1��D��')�6��C'�ԿV�?2<%E~S��)߿�����(t����@�mɋ����`K�Jee�yT�хd��)��ZT�ʡ�*y�c�T�����q�G�%�C��_벦�.e��o��ԗ,���zul��Y�m��r�9�2��m�q��~��;� �c��e�V�O�"2,U�G����!t��z_n'R~DXFx*(g�& qf<4���9̧�O��r*�v!x>��l��9���f�^Ԥ,�蟕f�v��V���ΔHq������4\��^˧E,��c�8��J��0o9/���p�Gf ۘ���8�q�x�x>�ex�dA�����[��)I@���E
0z�/�{���Na]���o`����Om5Qj7 ^�rӹ<k3�ۡj��=�eW�������|����_��uuV�S �֠o��7�W3�w��/�X�] 4�v�*7c�T;�W��x5���
�L`�Q��P^�����s��:5�Ղ	�Q�HYe'�p<XL��@D>��C+�	�t�Z�su3�T��I�iY���l�_���c���zA�õT
�#���T�+����6���6�W���/H��[�&�F�����:iV�b7n�äZS�	q0��7x����;�
T���m�1��'A��������C�ҧ��P���n�yg������6���Cj��1C��A�p���=���ጌ��nK`^�S�x�^�W�a6�7�Z6��u4�&��VwW/���z��ޮ�v��6�_�5էI�6w��K���EA.ԓc��������/8<s��W���-�G(��f��IZE�/l����ŜB����Q�a��J��GƵ�W��eX�֩U� | 6�?~8i-���r�))��mID�],W�?шt�p�+3�s�M�Y͞�捒�f�x�<�]�"�D��qrW��&n.�nc�J)��ۧ��C^�~4�[a�|w�	Y~��9zJ�oj�& M]�N�GX�\��RT�ݔ[��k�_]U�%�$bՉ�7.%�����BS��l�gWhGq���4�D���3Q�qȒ�b�����р��}J*��d�7>�rJ/8Pl�10���#cF:�nR�=W���iD��#F!�j
�Qk۰:7�H"xК���"+ŵ���c��V���L��9Щ��D��I���t�L���=S��0/�!�-�����~��wUb�����;�s�=k�Nӡ�X �}�4��O�
�� s�NR\:5����O޸G���Z��$�iNa5�/�'҉�$��b=�A������S�D�ͭXҐ�c� �+^]��Ѓ�bul:;ct��y<�@P�k�A�e��+�x�ȼe��\�c�|$q�ڲ�!7�_��Ѝ���5E� '*��Ƈ�	*[L&�c���d����Ӻ��hF�:��+��z�␏�:'4e�x�+	����@�CA�x��>�C�Y4�Kဵ�A �W'�2���?gR�i�|�ɛSck��[6zHW��tK[�U)
�:e�+~���&�(^�8�T2�=7�e�3�Fo�k����3�+~Dў��H�&����P����:[��:?�^�p��z���UC2��5/��n�2�����)�[N��.ɋOsU8�no�9�}�N*]{������`b$�'q���};n��q{Lҳt|�A1���F(N�����.���;�9a�65S�`���|?��s����ne�i*�(��R�b|�b�G\��;\�7o��-�����������5w�wY�5RG�<JWЦ�Qd��R���W����#�e u���9ne+-/����4�"	6I�@���t��6!w&���J����Bi�CkA��xx�)M����Q��Ą�|l3A����s#�������*��G�?�c��
�����q�Tg[9��� =�֕�1�&gdɯmݾg�f(9H�V�s�O��T@ ���T�9�?A
��"۹A��ĩ�i^���3�������$MZ�v��Y�.��FQRU;�^��s�C�sg�=S�{���R9AT~A6[�iA�D
����bV���,��kܼ�Je��xgB�۔K��4��)���� �L8Ѵ������- '�e�\=��|~�玵�+����k�}&���""�����7d-���9_��z��?�Q-e�l��t�AKA�V�A��@�U������Gm>����\���	A@`��,��&[#naF�bC���:�`�Y��y	Z����e�w���e��q�B���`�ݞ��D�?�Z�9�D��ul��Bє�c�H�EF�@lh����a�ApP�Yԡ;��Y�UE��\z���%ꧥ?Y<�����>�%�j#��.:%�D�CC�����x��Qo�;��S44%�rN<2ā������[�b��i�h�9�
��n�$�7�$��tfI���>]�M��Ґ W��"��������˥.N�ꑡ������4~N�Q�ߑ��[��ƖY���<1ݝHۙTߦ�jeKV[�Q�t�������5
���,���َ�`��,���[�6����Tٽ#��Z��.ߒgh���`_��B�&�|���AR�׃���[�N;[��m�^X���7�����j�-ݺ|LP/#8؋j̖�E��j �%[�+�-�K�OY��5�N}�������ێSt>U��k�~b"ʌxb�NAQ.'�����"*C�o�i����ѯ+�ǊD�s$�F�P��E\�PZ=ݰ�$�Q�1����YCYɕ3jx��,���j���m�ny�Õ�'���:���Ջ��7ڗgߩ�Cv�y��ђ3�ܒ7���TD︪��h�)ϡ)�"x�SC������g���o�L��_�»4����h���}٘��_H;U�l���K��������� R�7N�#ミ�$5��@b\􈣛�13�Ry�{�Xm�PQI��Pj��o���3 ���W��1ZB6Y?��x�p����M�QҲ5�#!8��C����s}r	���4p��Giv�r�4�5Y?,���`��Zf�۝����a�F�<Xg*�:-PU���*&3H�Mw���EjF�r"fW�ó�C,7'�اmP4i�*i�Ԥ	:��6���;��ГZ��@�vƑ`Α8��>hi��bVs!/��oK��^o+�@p�L�#��[׳���s�G����&�J� �Yz$�7W�15'���C���s�mý�8��Ӱ�����q;�9x��YĤ���k,����h��O`�M�X��Y+Uƙ��o��������u�;Y�exkAz���߂�v�E:5v3y�@.��|nnļ����(	�6}8��s�RqV۔�P���ҹ�r^�o���Pm�?�W&!���'��\4��u*�<�ng ���o�p�U��hjdDe�+%@j�L~�U�����zn�A�(|��z�j�2#JuFa���0��5���T��%���U�1�;�5������f�}��,&��r��O������$����	�����L��C4����}�)�d_�<��ʿ7���!"\En0Z/r.kI����")ZGh�ŧ����Oʑ����:����"h�Q"�Kx�'@�[Y��k��ګ6�E}��������+���&~��G�WƹD�l�l�4����Y�Z~ܴ���;s�$��LLK�q3
��ѝO�vZ汅��@��Y�%�[�CiIiYD��"���A��)j�2�<+9 ���� W�E�}�>���A��b����:R�����y�.WO|Ȭi`,j�=�\|� M�;/\o��f&%��B7B֛8�p���}P@S[�vE&��	�!��k���qv�í+3*?��Sn8S,�ﷂ�����g5�??�����&8�1�2@�s�9If�3Nr4Մ�`����>���Ox��l~'e�2��A�6gu��1a$�28�νjNyx$z�#1����N���߫1䷴�J"��c�L?�+{SN�9K���7'V�64��2���+Q5d�;|��Bګ�ƿUm�K�j���5��l���^cCU��d��P�����c�.�
^�n0.����q'ޭ�Ja�F� �a@����#�Щ�H�҄��=�1�e��*�,�?y��cE>xc�9����6����0斚[=�c�>M!m�hǕ���#����v]�d�i�D~�<��,z��������֊�@�S��D��=�x�����}C$일�v�x��#�ڸ����,�"6`	s�KB��qhLPƹ��1������:J.�t���o�i��8|R1�Y�f]���E%,U|c�Ђ������"�Vb���:�iWN��(mLMaA� {� ��"�4C���כ�T9���dU}��{�xo��`Αi���^�I��<Y!��C���2rUk��x��ȓ14��N_g'Ҵ��!-y��"�<�G�����A��5w���6GȲ�ZD��V��y�m�4��Zy�[��.��~߯��������ǿW�HF.8@Fη����0��
��i#����+���
�K�G]A�7�2�aq:�����u�os���a�<h۫�7��;�&�/��v��Y��j_�sY����/��'m�[�mI<s�iHWS��O�k0:��-ǘH�u}V��m��zđF�4��j.�E���5�%2fQ�/���#-��:2�n��S��>&��ؚ��N<����ٲ�K�Jc�3�̂���GBJ�};�6m���;%g���Uh%���ө�A�!~U�n�9D��F����_��d ��S 닜.����%�G�υ������\�o2�_I�	�R1~I�1���i��ڡ��O����75`�����UuT�c�,��R�׎{3��C]Q���pח�������u�R!'����N��fbBu�`�5��$�
c�&/��]�rs��+ici���t�m���O��K��ӶCF�[�C�q����&R\١�)��$y�@Ƹ6M��ڡ4��,vG�*T�w؃��͏�"����	M���� ǖx�o����x1�QTo���Z�(]��ꊼ@ J��h�i@/�V'J+��CA�w�2��^�[\�6Q��U�z���V�o���9T���5���r��EN�މ\ۈ���wF��9*g�=�¥�q�q�� ��0��D��`/b�^�;6�&�/������݊N)o��C=�~�NJڦ�����_����fi����*v#T��ۚ�]!�ck/	���A�4���o��	�y��'F}Ѹ%�R��ʆM��v��]zӇ?�gP�.����|䄄o��Z���MԷ�&�ڑm��ZY�`!�N��7��i��L�j/5!7�H�T���$�N���3���|����V4\�{Aҋ�ת^:��.�Om �k
�D�Q�/%M���E����Eւ�4�#_d��$D֩���������K"hs�s�+ǂ��J=� H�q�����0���;�{Agf�$ߵ�����ɦ���� *Z%�Iu��W�^�e-� ���<�|Q���k:�R��*�)�"�Cަ�b�)E�0b�9;�zf�M���I��S�cc`I��{����Й���vq�[s� Y�=���0��8kC���S+
�U�9dւ<G���G����6�$����3$�<�8K=��Ei�T�+j;"���_�"3���{����/w�P0}�z*��9ң��Qw��Mr�G�!���U�#���aw��$U�8-v�m�:Zc�������#�㍼�A��ˢcLŌ�_煴�N^���l�!+˚�\�i�E���4��q��OF��|vQ�l���ہ$<��(�>9��"�h&7B*���W��S�܄��mη*S3C�Mm᫷��X�ƙ|(b���j����-1��*Jq�H��A܆�ӮJ3�{}&�?^��ÝY)���%�I�<��`b��6�$�R��%7��"60G�E�����m�9m�(]�:�VcG�9�*x���	���B�1qS A-e7{�rp-m���N�Y����xP��A�;��ivg/MW�Bk,*IGи�e���N�fve�m���!b�FV�,��/�ʝ�&0��|r1����r�YY"R�&�`�|.�H34�}�6��ի�'��J�i�uKnP#dNw�_� y#z%PQ�5���O����M;����H��@�1>-����F)d�du.O��;����c��UH��oe�^������ͯ���7dURߙi���O-�0Zܿm�*%g2I[>w�� Ea�K��M�=�GZp��ۍ��6,ޟ�|d;=ki�u��7�X5�}��Y�~�$}/�*-ʙ��{�,��(~^�Э��EL'�Q*Ym9�š��B!�0ل�hh	{w��4-�_ʢS�-!�3O'�Yx�)v险ȣ9]��c���]k�$��w� �9�'(�(A����1AAlÆ!L������oY�b��ծ�o��B�l9vom(5~�mN�#^̤j�J�k�3��$��L��ɵ˕Sh͍������T`ؑv��cdN�/$��ћ�$R���޹��x�]��w���u�P�rq-�C����ǚ����5�_<7�ꨎ���;_���>z�Fװ���ϐ2i/�t��1W�%|PD§��}�%�?�<tk��D.Sb��,�������Vv_�?�h�Ak���>�q�#C��I�6c�����@ cGu�b���lb<8�P��|z��ɏϾ�/Cg7�w��ɯR�.�v':���]M�ϝ����W��g+�o�e���C�G�~muԵxdj�Az;(%V�l` e3�U4�L?2�Kvl>f�E�x	� ����&��B�)�J�$\� ���ۿi����KK�	B�T����<�0[�D	�>ԭ���w�?�S7x/�K��ag�R�C�&�p�T 䃃�T-|�1����0T�g�t���/i�3u��,ɚ�y"t(��Fbԑ�ͣ}��K��(��!��]'D�~�&02�g��!)i�&��M��'}c���c�B�L�Q�K��|&�ġ�-��xb,I�Cs� 9���*��VN_e=O��et��6�=o�]�'Ҵ�$�X?I\T ���A��xZ���������`��=S�?`-�4T�E��!9�c��Z8�U��������_�Ij�7���oQ�M/����ѡ2��Y""wQ>�]��&O#��s������̀<���dz,�j�;H�i�J�-��6��w�P�|�x�������P��f͑�X�'�3��p�ә�Te= ��E�1O�67�<�>���mV��E,ݠ������U?�J���!p;��UO�5~\�|���)�2��p��@���)諭�q��;�u�d���'���mha��K)f��)��K�k�4���m���������q������&�|i��$��XX6+K(ǅB���������6�;ۦ��eJ�a�F���_d#w�I�VB��qzW!��`o������)[���E{����g�F������X�8#�ڗ�����>��V�v��j�:%e[ �Ol��P�믷ʙ�����C�p\01�c��<�����7�'�o[���'cf{ C�뽔J��?�n\+���|����I��Jsr���P|���@��T�����FE:ˮNq���7�g>�����M�w�9Cr���u����|~m��+��@�Q�5D�ҡS9�eHfj�lp<���Ӡ��
�sW���z(SV&�R(_O+H,�lK���N�Gh��	��U����4����-g��naJ5��^��&��E����-"��������/�Gϼﹺsщ�����(�r�װ)� �J|:E�K0t�g��R��"�օ8uTU��z�=gh�e���8�8hRV���n�tz)�Cg�˞B�R���]�_����F�(^S�v$*a���^n�3��u��o�nmO$��MQ6tP��Z�@lp���oEI�=;����Y+���깥��S;��� ��ژ�����}6����'����ݏP�G�Ɇ~v&���ÒE40�}b��Upl��n+`�c�w��7�1��͆��C���	��~�P鬮��;X�wS�DV������^�A���wZ��HW��CvJ�B_�����U1k?Tu����"�i$u��t�'N\�<�����>!����p�ZB��:���3i�x�+E&J='�nz����t�,m��f�g}����XO����)�N���
�������t:cQ����jdtZ#���jQ����(i��~H���/������-�;�ɒ	|��nC;��>+���U��S�W�!�ަ%m��/t�+Bꚺ���J|�"��(��YZ�P��/Ρի��	��G�Ê?���Z�v?Wx�[΋~uʑX)ĎH; ����-C���Ing+ŃP-U=*�ع�Vc��u��T�͖�)�g�t��X���:f�&kN5V���/E~c׾ц�@+�yBzS���6~'Z%gРtf[v9�U��5��R����ȸ&+��~��T�|gֽ�:c*���ݪ��FA{�8KJ��g[[�Ĺ%�0�댋A�e�I��0�_��Maр%�<�R��^�m�X�f><l +�x����%@������i�8����G�M-,cEݫgȣY�
�)�G 7��g�s�^%@ǽ��������q��f����C[o#(��\�Zg�(M���Y��ѡO��qGg�j����kdj���5�oš�F]���G���_�m;HZw�J��Sc��j���ƻ;Jm	}���)�f�N�R�u�|�1����&-}��]�v�P�+�b{.l�%j&c�P��R����t�p}�(�^yـ��
t7d�I�m�]�#�=��\��0���*�T�L#,tv�,����6`<n�y��<'w�ԣ�^�z-#�x��S���t��MP��gr(H����΢^� ��:��B���$�͏�|~f���Kw����H�Z��@��!�j�KA��e�Uj��H�u�RӮ(S���̓��ի����%�|���ZE���u�i���+�j����^��Z?��]PV�I�,+����)O٭^�B�A�W�Hbޮf�uK$_
������da��hڧg�Y��ب D�A�.8g��$��#ѱ��|7���o�Ǝ�q�/
~�Y'.�^�I@R�*X{19 ���K��j|������r��LK�)�t��[��OO�����N��B ���b�`���:���@R���x�f�|Z��)�̫փ��=%sF�_��:�I� �sx��YӖ~3���F�	K̛���ɑS=�;-Z'�%
d ��/~n��b<4��j��c$k,j3�I�������@�(�0!��-�>�/9�Zq�	�Y�U�"\x?م�	U�'��̹���݊`a� ���3��gUFy��f,!���L�/Q��\&ђ�ӭ�<���#2��܇e*c���>@p#��a�){��!�\4����-�� *�U�Im̭^#_i�Fh��S��+'�\H��N�4`~+��"R� ��2��w�3/8K?���B�2����ףEw����@b�<�0&��+��])�ߝ�+�+Ⱥ$�?��W߯�A�t[��[`��������
>:�f��ֲ����J��6q��+�w�r-&[��fd��sΖ�m�E�}�.�Hb�����r�/̎��i��2�g�`q�w�u���Gq��C]%����E!�{��
鉭��s�C�ح�	�1��s�/�@��!���߹l��i���N[nQZw�q��M�Cc�c�O��޲M�2�Ða�A��5�2�Qa/�w����iѭ�_g�ϗf��3��4��AA`��v��s=V�]BPC-�����{4�ix�ާ�K�&x�;�6�Y�yOmb��%�K�y~?���}w��a�	��+��kMq�uVs���P�Vx�c?�]îD����.fC�2�,T�s"?�U�)m�[��Q�6V�OA��As�f�)�6����L�++��R����W\g�������6Y��^�
9Ej�#�ӝO	B�hr0r���yB"��$�x��q�8��JLjn��hT�_�UŖ�~��q%Z���l�b��
���[f{_���[v�Th�qD���_4t� �@E\2~<b+���U��1���	��]h#I���o/����L[?�3��U�<�ÍF���^�<�[�m��Jk-�e���]-KX�����<�f=KSw��`�H���nE�ü���T�,�dd��}�W[	R��v��`]�o��YI�Z�$�l"\a��ֹ�5 ���y+^�P�&9�82Ab#�zv(?8���0�lXE�I��r����F_Z���ے{Ř�<1�H�U>�p~<���@�����(5=6O&�!��2�υ��N?�΋E���X��iTʋ��½�R����n��R�%��	���H| $<q�_J�tHF·����ʕ> Z;~>�w#f^�t%f�� �yj��y���_D�m��j��l,L�ei����W��2t�G�C��AT2������\�I���G�N�D����u��_�� ;���n��,40���^4�<u���(H��*Njs#�����c������g��~0�=�E�1#b����Tݵb�a�W�d��F����8���:�T#f�`�1�h�٠�G���42b!�`�����i�I�Nc����P��|}y�4�����п��)Cg�������lyy��#E�%����q��OM�*,��_0�s/�.��;�H�Q䜑-e݋�N/ҵ̸5��0m�:�y+B&��f{דL���㮱�N=��b�J��h���ks�
YOo'��O�@�%#��[�t,1�������9T��~sU@�ͻ|G˯7Lt�*�y�P	f��wu�8UY��>����$�ʐ���9�8�ۙn�~m#b�J�N2�"v��e�<ͅ�_ͮ�@<�9����NɹT���c�_��::��SF8�����a���|ӝaO���Y@�v.�,�
�VR���M3��U?s��Y$k������k��R�ۜ� �_s���`q[��Ū�9��Dţ{�"�?"��E�|cD/�t4���Ӆ�,����\M���{R� ��Y����o����O�g���	Ƭ���th ��N��<����bc>�8HՃF�^큲��ݶp���F��i$b!�D���Q/����࿸�m�`���g������c�������k���s�7Пn(+0�$��e��!"Z|�ȴZ����Y�r�h�i4g�ԁZ}��X�Pbz{/E��<R	����Q��2!Q�� b���h��J������3_�d�!ĲR�J�]hH){	t�j����
���MiغөÝ�`�@���4ɸ_[����p�V���Ұ|�յ�ў���/S:�	ѷ}ÛH��:�}9Z�x�x=�\9�;���߽����;��[S���iseû��Q��%z�^kj���,XI�����g>Gi�?d]��o�.P^o���\H��,?��;�-�A�5?��/�H�^���1\�PC���Y���)�{�-l�8�[�g�d�u��Y�ĕ��'~�j͆���k��y\#3"uíoz^���T�y��)�f��s��D���NJ��-�tf��f�ދd�슽a/�U+�|*��/2�c�b�yƭ�%;U�U����f���S[w���ՏR�hd`٢�|���� �%��ۚUr�����ne6�Ɉ�l����!l���VC�=$�r<�ø8��4K�I� �࠸_^��Q�Cn�SBM�<�yr��_�O��s�"��pQ���
��Sk�ɒ��TS��h���p�gRf�/:@w�>���­!Ue���h&OC"Z��� q����O��_ChɎqa��>Ƞ]&���|�v��zU�@нl�Y�9:_�Iz����W�ׄ�&������5b�5ƿ��[�5q�y�����������S~���4��<ݥ��գ�͡'gG��m=p���o���x�j؉ɇƐ�m<qF_��-Ny��C����.���0T��7#�M���{�Y.c�:�:���"�heb3W'S}�Z�C�EkS���7�ؘ�J,�&�7��P��y�4?�Hh0P?HԵ�����c�4���r-�u�"�@��=�&>ړP�b]N��=� O���鰒��`y����ߏ�ڟZu��_�)�.�UY�&QU�:H�3���.
�B��������߲������Y��2�������5L�b�0���$�� �7�^!���~�L��5����8�.K>�A���TAg��U��,&��S�_����p 	�ܙ�W���N�k�vJ&�K�C�I��}T�d8u��̃�>+�9�M�����'4u�D~ۋ�9'���x?,3�*��/����"c���j1�/�T�U��%�i�X���ݭ[�za��'ZL���B�I��fM�0��b!;���S�k���T)
s�8J3���T:ݧK�4��߁��K��$�̈́�b��k��g��V���F��vR_0���D�I5[>�eMP������8��+ĺ��D7V$��O�MA�Lw�DP����t=��%�Tɵ�0 79n���������V�m���v�|���jf�_����iN�"�מ��9aQ��7��j�!�p���4�V#Uqa�ާ�j]ͩ ,X>鐼���*Y_ G����nE���:�R�(Ј�^Uk<7�q�?"6��-6��X��`��DE������}�C:�BMW!B� �99LIܢ\F�����M�!�[<v6�w�Z�Ұ��B�kVz�:bO��s�^g9{�g-Z�O%�w�.G�5��m���Z-�	��w�\$*�-���'�؆�zm��4����u��jب����/s��\�D��G��#Ht(�FX�i�`�i�Q�5̃�����VѮa�k?eƹ�@!�e�iڛ���L>��8Y���e��f's�1D�M����&������cJ%+ލ��	6���#OëN�o�W�D���t��zq���b��?�I�����^��f�%{?&Fh�eI]��������w2��H�V��(�����M�6�P�#[�퓪Nse���R]T�If|.FKM`��`�X޿��sJ���h3���&��U�f��;��(!ݘ>�	�a�bO�t
�X�0{��-F����I�zV?_� /��v�m<o��%4��&��@ޮ��4~��HNF�|/f'�����o�a'�0T\�f>��n��p}~�d�$�,Ŏ�NU[�u�Q\��,�i6t=���#~p،ng���w���y�܊n���rk(5��ɉ���$ni�^˻����l(�W#�N�y���ë9uc̺�/T��6ӟ��K(o%�u�I��ц���$8X>�<� ����	~o�c�iH�⚋xt�w<qS�A-U˨�� U�����`��#*�]ư�V�F�es�[u�r8��0����#��9�x�����e<�Z\��q�%�w�`x&��]tt��\��d�њZ�����JQ%H��o'Ф��?d��G`��/���J&�^�V}Q}��i\ "�g)`�
X�^�p�xh%F���'���5����^'�Ʒ�-�����6��y�By������l(1S�%	��:����.&�e��U5�XW�K�+�04J��xP%���� V @� )��,< �Y��2��	;�����[m��c?����J�K�M�'�)S��Ӽu�����}�˳�m4�b�V��^�^λ��	0ۼx9�)CA����R��P[���-t�-��1�+ƣ�/y�v����Tg�T�L$�(63'#�ɓx����
��Bb�Χ#h��E�?Ok$�J	ִ.��}F��7����[����@R ���t��q��h�a*�txD�4>o�BjwHW��	� Ch��4�6pb>6ܥ��I`��|�upN��ǜu̩.���w!7N�m��|���4-�V��^=J���.}��u=��B���\9�O�+Hĉ�#�N҅�N��u��oG�NF�<<�1�ۄ�u;�����tH>�M\l�6��\'2}c�T�m�N���s�v�ű��Q�aW��A�c!$t� ��Ų��]r/�����k��2f��T��)k��GL�m]�G+���r��qk#A�S�cP�d#�B	zV��'���=���=YN�N�r�,;��b�D���,p�B��
���dl���{�Zz��/�����eR�y�����GM8<�(�Vg)�N@���,��~��י|��k9��A%���x���������	t�"���wS�� Mi�����w@c�����vg�<��c>�"։��+Ȇۍ� 8�����LVL5%A��z�(��F����g���+e2�|��P��F�q�0%UMh��@#�g��v�(�@b��h@[&^R�h���f?%1O�>%EA���i��ҼN촶�T�,@�yKcV�\�� _�D,ѭ�rڵ�~���b�s4�����"]�y=~�\P��Q�tcT��a6�o�A|#�a��T�]�dǍ��/� ���{�BC�S���ɮ0*�!i�B>`YL�O�+�8�8�e���37�y~~�3��D+*i�s#�?��`���=$�Ka\⟽Ã1M�W���i�:**��&�E��ױ��?I��-z��z���#{���_"<i�k+�X�������v1�2po 6 �R��e�8�XcP�*lswޟ_�������S`�:�)�U�U|��k@��w����x�Yޘ��'�!p�۾��d��)l���N�܍��-�P�;����t���%)�lV����u��?�{�`6�F��<B�P
W*/(M�i���D��/|�[b�(���2T�A����7�ӄ� ��%Ӌ���h! k]��Bq/�k^�M��q�׊֠�ܯ�YY 6e��fSm$!�^K&4�.�x���i�!�Pm��=W��?�T%6a����o��hv�����5���hx���M�0��
����ݲ�皩���0�IY�o���t|��L|L��� ���5H�N���:@?�L�Ϣs
�T{B��B�ǭ�ck�$&����+�^��`�gʽ�!���f��'�
&��#�:H_��%sI6ݕ�D|[�b�<�΢�c�k��|dލ�0�&�Y X�:yK_kWN�� )ݚ0�<�� @�5����%���f~�6�7׾I�F�n�]g1��o;,T�qn�{���&^��h��b�%wz���e�q�sC�5�{���|M50�3
��I`pFH��|��Ђ/�9S?Z,b(�ձY��=LÉ|�
`��bm���1�^W#k��>7�x�٦�LT�~i��8� ���y�#W&��to��Y���������8����QucƜ��(�_1������U�y��[����va�t���Z�sm�v���
������Ӱ�%�XP�l��g�'Q�,ؾ��;�Kԑ� �@�#���^�%���D�
�|5�9
�������Y��1�I��w�)�緾�~���1��J����!�� ������Je8!d�x�d�B}m|�����E�O�����iuM�,��,��Cvdc�O�Mj�(�5����AN˱OuvG����Faږ�uiP23ã9��j�ۤ��� 7vPh��,j�������=����o���ޣ�� t$P?x�1��^6e��"��",�&G{ls}�E9W�F��u��Of@E�S�1�H��y�/ܽ�����Ϩ�������#PNZ�Ũ�C��e�<�I�vN��C�L�U�ݕZK8�Ĳ�� -�������B+�AW��k���zK����X���Q�0n�г�/�ML ���V>����v�C�(��B�F_A���X���ό��&C������� U��k�L%��⠧z��[M�6bGM����nR�RO?dg�p� W�b�	����u,�*����h��FcF���M;�Fd�r��U��᤽#���e��=��"�ڹ5)"F �Y�g���Ѹ�e����[ϩ�Į"v��g	e7���Y@�x ����k��F,	�Vs����㹭Hê���j��abB���\U�A��#v>G���q���j��U.��#����U�ICn���B7����48΁��Z��GXG�l����Ֆ��#�p�6�:�r�wL��4��tpf(1�+�яU6D���"@���Y�8��Ϻtw�8�o5,\G���^p�9Zv�s��gJ��;��{L����$Q̍'M��td XG�F�^1�O9��|�/�r�3�tN�4����hCO�ܿ	ʹև۔��߹��5Nh�)�"]���b��=]h�J �㫃e�^<���:y}ԩ~�,�t��۟A��Co�ͥ�6ɑ�`�,�KɌ^uzpѝK|�d�dSi�U�^�p^>A���y[U�b?zcS�S�^�6�_�&����Fc����
��/.��{�˘��Y!	�Y)��-����F��ׯ㪢�M�d�+hd���24pm����B@�;��fI<ET9DبUq8L)Z�}��zL�x��.����:��,tµ|���z.���\%  J��L@��ôS0aݭ@/���<Çl���L���p����ߎ�8�4���F�=�Z�����.�n�gJ@ص�E�h�,g�dV�[^��d�t-h�������0$A�ȭE��+�T5d{�4���VJ3Fq�x}��p�����}�ūI+������0�4�B�;u�pN8j��5����(稁���TK��۴�$k{0��Zp��w&���h���,ݨq��<3���5�v8�]�F��^�8����-��w���Ji�)���V�	��y��s�!�Ƕ c6�	�𬂦`��3���u�a��~��j}��EI���y]$��W��䃞�M�N_��+���؆�F�Z�̨��#�=|���9s)�jy�p;Q�6�2V�7���TZ6�)��j�O��v��3,�v��璩G�e(�ÿ9���$j��〄���nČ-rpp��D�"F,տ���4����{na���/6�-A���\�G�|y@"(O�~�w�	s���8F��`�؛!��J��q�y�׿����F�8��L��
��ߊu<i���T:�Գ�(5���8'�&�Ze��ܛ`��Q.�G���%�x��b����ⱒ�jd��Mo��t�2>xɱ�nAX�>.g��?2�!�ܟ���S��Jƕ�����9fC����O{۴�Ք�9폺k� �|O魷�y`בڊ&b���W�~��kw��1�U��e��bb�T�$l��^F���G$��`+���:@�Ğ"e�ջ��Ge%��!x�BR�Y�e�2��~�dw�Y^�Ur�k�1���g����a�Vo덉�9�7��)V���}�\n��u�MN��_��	)�F�P�C�A����ъ�7�>HV6c��zA��ڀ�'H�O�<h,�98�\�˪K�/'��X��{97n��GL15/X�>��
�p�8`a0��}Ȓ��f���lh�\Q��|���h��\��7'L� ��ӥy�D�鹨�Ői;Nѻp���ڕ-S2�>���Ӵg>t��"w��e��9c�o��'0��ۧ�S������11Ñ�_���XO k�%����t�]�~��C׀v���,g��<��D����t*ip{?�¾��*q�u:��o��%r|R�
R��(����+���H�_e�(�k���iuL��a~4�L����y�I%�L�����~�WN��������`���5���z�<��G�֨1f^��e|�.b�����":����j��G�?Pi*���𴫖S�HN�Ú�ֆr�oܝ�N@`ӿ�[>��f�Z��CX>�4�ظ��Wz�Ɠ�V��z}`���̇�rJ�}k�4I �Uh��[� ^m^���=[�N��ң��5�\�ۻ�賥E�,=��r��̘�'���<��yCƿ���bD#��^��ŋ.
a$��_����@@�f-%h���>�w�i\N���7%5��v]�!j����nY5�|��&]U�r��A�0���խ����G`���ʫ�l�����ibQm&��.{y�wZwT�J}����g���+S�����	nAf����u� l��\�.q��l[�[��J��PB�A����n�ՒJ�2^�Gۦ �:J��~�����n���|hs�f�}PG�C���i8�di��ȱ|���K�*Ep�-���`]:z9���ћ5��]V!r'�����V���d2�Sp��f�v4xTu�5���B���wd�?-�#����א�KCB��J�7-Y���,�s��t�o��urVY�B�w߅����@�+p�<+P,�>�z���W���B��+��v2���eyhH3%-_�{KJPְ�ȷ�����̋��2��Ac�q�#X]��}�����}8��=��Ks�3����B�]`[�Ӛо֧���0>\����XkY�M�9g��|$XJ�+6��]�`�&�>|nJ*���4�_��{F��.8���Ǝ#%,26H��j��tsd������-�#�����[�d�Φ��dd4p�'�	Rb�l2I߂�3J��#KR����Q��:�)+���%	���0,}^u*�T��G1Zk�v�lp�I��W�-ց��F�u/�!�L�s�,R���OM ����-NJ�h��O�!g}f�	�Q�(�_�l����hV[z��Ą:nkh��yK�1Љ����2����aZ<k��;U�N$�x��Hh9 L���Z�P�>���tup��" �^��؎l�`L���jWխ�X=�B��A�������2�} ��C�����-pn	!����̀��_s�B��3O�3���6M�r��]�Mf��y)��x4=ts������O�(ߙC�=]��Dd�d���GZ��!}D09G�0g&|�e����j�έ�R�����K	��)�P���m-�I�D�v�*��Kn��s�V�K& ʄoN�ϭbT����|a�;�-~��m�/uVW0��FݽBA�����9��ɥ$��=z����F�;�w�y��J|�%��;�9H*�9�ǩ�k�1N.��C���N�맜V�~=�լx��hZMc n`Xa��1����}�m;��¡�q/�z�]^���/��G&��fX#�g���<@��)����!�"��۟�m���\S�c����|��r���j<&�&C1�g��6V����p�k�\ru�lRh��:�<�`q��o�Ys��MӤo�:��O7ӭʵ�څeO;�p6[�XH-k�	s��wmν�i�D)b��4��(�zJ�,hX�H@���j�^���K�FH�da��D	z�T�[��M_��mXrV�ݑ�G���G&�"���N��"�����>q݇��0�ZiJ�t�������_n�~z�Op�y}x����8�;Ͱ߾����^���w�&.l��d�}�;�p1j�-jIY��0i^��sH�þ�Rr�!��5�R��)�J���B�񈺳e�B��e�b[w���I`�4N�"�W9�LIb�����=ՠ���l���ʉ��` 9K�e�� ��=0��^%)���D;oj��X�|��r<�1�H�
��՗B�&�<��$d�'�([�<���*�,V��a�#������k&E�Jp6������Z��]��u�A=���>g��H�����F�jw0A�Qe)�c�:K��?��b��sD���3�S����9��n#)����}Q(�c�1�Y$���N2p� i�}b��o��D����m�۹�a6�!�L�Ǣ�J�߷�Ғ�"�;pL�9�~�1J���2�w�L7�
.eߥ?��:�2
B��+�<�H�$�6��hE˄;�@h�O�sf��lg���d�"�Vm�f�;���y,���bhq��&����@
�x�ԯ���s,��G�i���z�EcL�xs!�7B1 'oޕ]I�6�|�'�������[cCR�kq�?]&@(��!WBQ������
jr���X`�k�5-����Bɻ/U���Z� (�S``c�U?�����@m��	�L�[�{_�n��Cf�x�� ̋��a��L����xU��+/RB[	��%�e^g�:\1�.��{sd�s�0��>�ܿV�Ϥ���_f�-~d�����kДĞ`�H_� \�rh�Ġ���^�d�{��N���0m(��k
!QWZ�N�:3��v�:ҭ�/�� {JwV^�*�f�K��7��'�񘬯��U:�ϑ%�et��2�O���n`�/�_&T*��I����8�*�����f�vw�B��WV|�B.vC�`B`�s��oX_���6��:-:��rƚ���譠8w;�Dr }��=g�dk�j��*��O��?�(]-��4]Gl��j��g}1��9I  OA�=�ZFYL�5�HJ�E6q��q�~♁�v������_2�4��g�kG؝���c�얃����"�B��yR5�,�4>��Nߡ���^ĩ`���}/TEO	�;�M	z`�G)�����̭uT�x�ay�36������,PS��]��i�n�?W�{�������~u�\�1�.8�E�AVя�+e;��moD �RX�$�*>��K��'�V��0`��+y`���p�+�`|��c�� ���D��3�{h�P6ed�^� ��Ə!��nЂo�c�.���"u�=/�0��`�E�-�h"<��L}��s�j4�_L�SG'���ծ.H���΄/ilq�}C�:��7���F�\+��]#������3��Mr������R���4S�@Ϭy~��tw|��˞�J(}��ު7��D&F7I;bH{���i�Xq��&�#��pV��sAJ�;to"[b>�gÔ7oc:�������7���k��B?��f=u�m~S95Ѷ +�x?S?j�?�~�#%�Xf]W�G#�)�vO���I��^?1[�o�G�=dim�K�n!����w/X*��ޯ�QZ!�LE���KWm{�c���Ԍ���7Vʁ�uL�/�b�����A���q���)�i�W�B�(��<R��6S*��<ÿ�_Q�����+����b�"�K��X�����/�����$�����P��r�	�Y�Q>]�=�f�ډ\,`=��g�K&�`�� �'�3��9�dm�T��=��Ri���-;f�39ՉX����U2�gG��"��RB��C+�Hu���۫���	����]��N=�b�H�x$��)�-� d|�Gp!9xͶߔfF�܏��i�a��A2�) �pl�n��KU�M	}<4eW T�y����e�X�p��HY-,N���K��3�ץ;�yJ�H�[�+I�?]ڱy7Œ	Y���*��)^pY�mt�su�T�3_웙���Of���]Ǡ��KO�ãJ)3$ �w1^+w�́A�sҨ/iv�l��+�3W��d�����q�Z�3'C�ΰ�U��߶?��b��87@T9�1�Z�C^.�s�3~B9�[h-���nP�X�h���+��|m���8N�#?��#+��� (�:6�菖�'��%��8�ˀ�Yk$I@&[�oX�}GᏴb����s+��RA؂.��Kr��	F��;JFj�N�3[��HTs�ܰ-k�,��X��5�ߢ�s�G��ʘ��٩2h��:G��<�i�������:���_z��#���j��8�(�/	����Ԛ��ХV�.+.ھ'��dDVƘ�SI������l���N:w��m�n�w�ȹ;�����8*"��͚�v�Աa�t�;�冑|�Y2����=�������M�;�ln�u����.�xg���!���"m<N/���v#~��<�kO	s�1�x)��n;��2��>Tv���<�𻏤G}�u>tɐ�}�s$�M���L�Z��!.��;��s�WqY���V��;��@�Z�q>!=�i.��zP�Q������%S	��c}K\�����T��M��v�C�\��� o�^Q掫t�����=����תL�̃�\Z�L E%��8>�8#�j����Z
�4�B� ��Y7&�xUaQ�dEj`[ޱ�H���BZ��%����ٚ�)8.`�)���*�tw�c&YZ���Lp�%p�l�nw�2skH 
��Yhy|�� �!���t_S"U�R&�54x�_�ͳ��'�v��^N�����B�b����A[�e����,8G�0%-�?(�t�%%�����y��S�.9�+�k������@u���΃a$C�J�E�O�Hi���{f��]tK���=f��^0I�7��D(ڣ���}��ϩZ�q��B�,|8����x�Ӊ��;�����Y��Z���C�Az�C�@Q�	s?/ ds������y��~����R��+4��+֢:}z���ةR:O�� M4*Y��Zq�4J��8$7qb{�nmV�*�@�ݜ)7��b�X�A�0��Is�+⸩��=��"�(��2(?r�{�c{��q��M.�أ� ~�ڷ���vn���/<.��a.�uv�Mcf�W��-��d�4<�N��-O9i�Ú��ҫ��:;�����E�/�P������j���K��斏�S��4��-������;�����ET���)�V����Z�*�]�2�2��EP�SU,�c��'SG����:v�ɝ��	��8 �gT��bj��0U}���n}�}|7��\)/�h楶(�6p �Iu*V���x��v־����X��:�+��Ȱq��!��2+��{6p���cxK-�����@V.�T֔rvV�O>����ף�[i�8�#!G���c�K�0۩���wI/$g����*�����
-b�	��PI6hQ�� <Mn٬�"Y�&��ʨ N�9��>rwcR��E`�d�3�'��AZ_�jN4f߷@�( I0]��aƵ��O��Ts|�(yj����k��tr��t��� ����|����>"��F9l�Պ����`������6O�i�����:֢!�%@{��c�n�L6L�O�v{��J��VgE��> �^��h(���<�c3�3���E�G���l���k��m�Dqn�}9��ꝋ?>�6�C �|��4�S{Vv	�"E'�,���������T�\9\��hΚ����SW�f���wy�I��׏z�(|�0�C�팡ԯE����N{(D����V1��	~L��䀣�%����˸Mǥb�q�IV��QCK@�Ԃ��{��`���Q,��'sD�YF��~� Q ��|�)*؞��� E06F]�6�5�.�ÎvBm��#l����.Z��3�E3x�Ӽ]��������-*��T��]��H�f�2i@�D.j�Vo�^�1[�J$���/R���5�8�݃lG��m%m>�����h�/)W.ŏzj)�"��VctdD)AA���в�3I;���e%���|�,}PQ�C�ʶ�
)�e�<>b�d��ҧ5��J��X�kkr�xU�C-���cM�?<�\�@�'�s��}��o��)����X�U��=������V�%�^9��x(��qʪ�[�ۨ�_��Kæ��+(Ȇw�zӼ)����q���\+�nD�$9[������Mq���	��w�3�V�olGd<�n�.�V��Vg|������{�"dVC� Ο��u_H	�� j�ӇJ��zD�~��P�ի.�����9�kYեdr~��J9dΨ����=f�XWf�9!��u·=0z7��z!���B�륿.��&B�+�(J��6&H�X�+�v荀H��#����6�DFie|�,��Fttq˽�Q�\��)�-���e���  =o������*�d��VYUTY���\B�	n��|��͗�k}��筕\%,:O|jgv\Pۆt�ZPJ�V�m!Aq�u���i��S��H�o8�oQUI3	ȧ,�~���ĶS����Z�u@noe���� �Rbe�='�D��6���Jǅ]*�+�^b��豶:�
V���-�����-����
���?���Q����m��z���%��}8���VS��0 z?.�_(��#��L�j�P�K��+��K=��`+ �1�-a�%&96�ҭ�錁�R����p�O�O��h�^����c��I�G�_�T=s�����C�P�Z��45א�#+�#<�y�|�zӪ���((Q�#�I~�uE.�t��/�첚��
 ß�x�ْ����o���&F���[2� y�g�k&�w�!�oR��$w�g���}��B��"Cĩ^��Ye�x�2�$��6dC�s��P	�fm���1h˘cu&>�Xw���;`{�' 8J���a�Bk�w��V0גdg ��I�6m��w�k_hm]<5��q�2f��`{{�XJ�XH�m.�;�;����=��@TE/5�:3�k��)�7}�݅k5��a�;Om�A�G'ak���'W=SJ�}<6��$?���7�� ����Q��P���o����c��j���I�)�G������� 8aw3J�.�x$����3�����/��PL!�^���j��WWA߽�S(-/6��&�ˇU�43Y�t������$����>t�cI;2O?O�^�����3�k�y�r��A#�v�8/��R��o�1�W��~x�RI�Y�}�;p U�o��3M`U��X��E%�Zb�h�x���ZL�A��f�������*a�UbE���AΠ��r�;�A�|�K��J�ۼ�My%�)��<��*_P\��+d�\un��7m�Y�p�x'D˧�,P�ےUso�,P��I�W�m0T��CC�[�`�#��&����R�d�$X��rt�Ivƃ��#��b��l�);�	@�$��;�"�:��G.�J8Xp����}S��o�S�D礓PKw�$�c����Bn���?�8&�C��:誽:/��'���=���� Ws���9��X�=�=�u�� ��f�i�]�E��&�]�MA�D��s�\�	s;���9~��%CCE�Hly/�V~���)~uAi�E�ʙz�I?��.����ަ���������sHTmq����?M_����	����g�9��1�^�Ê��Y0���!��c��(�:Ɓ}�����o΅�',��4O�����ϑW�s��$���6���Ͱ���6�E�+��6B���
�1�
?�>~��┷b�s'b+�S*k��<�<�e�.��z�0���4���A_=%�<#��e0/����qU���+�J�_�(�iy����@�0�� ���T#xY6K0i�^���+H�S9���L��6g�&�`�K.��Ә��@ �>�fE����Fq/���t`�n�<����:	GPܮ���6�Ej?� qW���gu��S�I��!�_L�-D33�d|������6R�f�nw��$�3�F�[����x>�	������.�ćW�io�8�,��9w���B�o/����!�͜'��{�j��`M����*������[R�Q���I�	��9S5z��^�$����� ��ڥ�͓֎�cv}"�G�2ïb��E��Li]q jT����Z�T��@p��[��W�	ޟZQs.@B '��� �S��.[�����ӑ��(�9��!< ��t���}8(!0�(oW$�����ɇ'Zr�7���N��k�v��-�9O3��TK�&�Wa�?ʨ�ҭ�����S���D�LD����3:C��<u"������rU�O' kT���;��2dS�<F�'+t	F����'��_6�ߥ:��؞��agZ��`G	�\#�]%������TM���W�H�����O}�O�(k"F�vҩ|(3ݒ��3�&�$�1�pO�o㡍�@�=�#U{
�u��!�DFRޏ�!��'Q�7�f��w*�U�!|��`�4ᝰ�뺡X3Ȅr�0fv��E�Ql�܍�
T�|��8E#_�������8S_�n}jnG<UP�۝����)���5|5�S��8��a�4�"t������j�Ѱǽ{'��E2-j�Ε�ǋ>�0�ںd��>@!}�X��Y"t�N�A�Lꔸr�.y%�Tx	��VKͬ����Z�+��g�'ڴ5�S���m�E�j^��©��nn�)Ò<��:N����_�BnT����rK s�yB�j< ����/O��z��y��b>��{12P�Ìf��g��_ݝ�Sq��W$ǁ���"���2psM�h�wWנې��t��МS������"�'
F%�?�Sb�s�<U�Uuz��g�d�O� ѳxk9��/5]���O^l�j�^8� ��1���æ�{l�j�j}+���5gWʤx{�P�H�1q�k`�1x�-������'	y�� �����K"yy����p�����}��,߉W��ƽ̼R��o�Z�s�x˖�ރ�:]��jΥUy�v���ÁI|F�z�(�P�%��R�>G�y��p��+�/crO� �v�Γ21�#�!�!�R`f��fZU��7�� 5�f��5�Y���#5֖�v�Lr>�.�{9�F�G+�����^��L���r�E6BFVW�R>��l�&�G$mJ+�}�gN�L�$ׂ�L�����n�ë�uw�$s��r�>ܲ�nf{��͹!F����H�`�'SH�ea��Uy��Q���M�j��]���4K%-F͙99��ϣ�/�&� ��T�)+�#��tv��`��[������֍0-�+�3R�f�ԗ2���a����Χ�\&�E�!&�}#۰�}�>�0.�ᴒ٧�T�?>7S�k#�+:pFnenk;������Һ�6�����f���P�yV�ʕ���vl�������G��`.�n(�O^OT�x���!$x�6�i"
T���3'̍�4U�(���Y�"ז�r�H�� 54�C|���Ab�:��M�)�_#���ĦOj�{���@���9$垛�����~]��E�f=;%.a�!���2���aj��֟,�i��-c�#�Q�p5c �W���������E]�e�!8��Pq�B�4�>,E�w�@Z��~�ҦN�%Z�Z�]�Ÿk/p�`�x�ǎ���V�N��]
$�k�z{�Um�5�E9Jl���u���SWh��f�UM��:����;�1}�	2/�	+5�
j�.@�gv�z�`�U7Ꮳ��J�+m���\�ť����C��������4�e�H��i�H�a��W]�¼�1]�5+H4*k~Q����J�/�ᡆ^��Ne�-�Y�U�����4��5x�}�p�/�ɷ�ͩ��5�Μ�Di�0y�	�Z��'(�XsF�(%���nzY��]��R��ߟ�&� ޱ�o5{Z|�$�m��	��喣���-b:�G;��E�v��k���:X���=�h�[�!|m��57���Ĵ�=�Jߘ�L�ӱx��i��a���J�k�����5�Qq�?������?�s���9�d��F#t�,��/����?zGO$�J�KP7B�
�*���=�"!ȜE�������"��[�GaoM��V˅�����(Rڸ��ԩҰ<^���&_Cr�ɣ9q��.�N��;,C��=`l���E�zq�7�:�v|3���(�g5��f)�J"��l��I2�?]�l\q�������Y�!�w6�P��u�H�!F�X�� i�}n俄���j_U]I�O�^�ΏbA���X
Y�8I�t�(Ӟخ�ۈr����E�Z|'�^���w��"�4�P7��j��Zbpt��gO�k9����Ӱxcw�hA��
 l:��� ?O��)��'�\"k�c�ak[�R�Q:]�?�V���A���=�/�}B9�S�Kn�jq�Wg�P�gVV��H�� ��}�~�ĊL�n��HW��?�WbJ�]�2t�XG�Q{�Q��"�Ʒ�U�����{��U*L����^�\o;o�s1n�H*$�������E6A�21ΐ��Z	I�_���L��d�nG>�������řr��#�.~'f��9,����Fj�r2j�Y�!�#*l�7�Н�w�'�#��W�{�t#Y�>aāl]o͹t��YbV�N��$Ś��+����c�])J�t̜�j��:��ܦ�<�8���٧�&ZZ�Z=�\�Z�V��EҬ����
�b��L�R�]�@z\��__o�M��0810��'7���o�I�r���(�����i�%�E?�j�n�m:���6�%��J�3���m��Cw���+k6�FS���ζ���ߦG��	��!�E~�sBA5 oF��oZl��Ɖ���q��=@i��UW�}�z��y�T�k�$KSټrAF��c��~�-��̭��<��>���t�.�.��\,C��@����-�_�
�@{4����H�P>�/���,4+�Oq�;C�c�����{|h]X��۳���&&���٘Q9R��vF�4���O��I��l��DZ��u.G=�H)� ���V E�TQ�M�?%B6��Wƻ���|����f����0�#��c�{d{���R�l�ѿ�mm=จ<��(Lq0���+c�ʴ�"+6+ϝ��v*�&�� dPBwe��d��̓�������Vr����b�$�莑���c&Fd�F�{�`2̬3�_�0����V�el�f�TY�f���"AP�����
y�Zw��Xt�]s�o�G�:d܏	\�ݛ�	+C�����E)[���x�=-.r��#©�������iuCnʞ�AŋE�Xӝ�����ߐ��6'�E����T�y�zA��
C�~5���%�vX{�=�ޚO��Gy�G%;��D-�a-d�8Ɛ"�d���.5��6�TI�\���7�����հ&�WB	� �Տn�*��(B��Z�e�����>�(|����]�s�s&�.)�ц��x�r�26�Y�8��.T�@�3h�@/C����Ŏ��I,�TI �#�s�c�B�Ɋ�P�zu�#��&ě�!2���=��b�V��$� ���h8'#L��;b��9�*(O�mH�q.vu��it�V@쉌M:-4́����<Oe�[�[u`��y!��$R~dk&�΂@�&� S��(��nY�$[d��,@�(���1my�}� �����7[4���x������#��ݷ-Ӟl��0�&,��HPV�}4e@�����	ܛ�Q���E_�7�s֍PC)�#r�\9�3���F�4`7�MZ�qr��>��(%*hI����N�:E:��.�� �~;���ꇉ|�9-m;/@���<�:�Ӗܱ���gRu�~&�1o�W�5��7������6���������8�@M�(��ʑ�f�Bi2��W�R����Ct�t`z&�9E��Ǐ����>���P����e2RTYx�3�_7C������X�]����������m�vY���eO�H�
���u `�����G:�-Ɵ�(|����,����(9+&�fF��3�Ɛ_ñָ��A{*w}j��22��|���z.:��F��RlD�Utd�'đN�fL�Hd�8f(B�5���B��s�HZ���Cs��	0�6#^ăl����Q��y�؇Z �X� �xī�e�M���
?n�����@������a���s��/�v����K�؀U�Yc���>�ֺD��Ƥ8�U<[�|+SF�#�(�ShF�?V��(���X��������$1W��k2����5��l�x�&���0��p@�E0C��d�:�h�]��8���'�/�=����/���_�+�hv��S�Vr���D1c���B[?��ξ_3���e�&�A�!xV��B[QR��4)R'$<��b'G�K?�����e��2�"���ܫ����ƃϏ!-xH�6���!El��Y���oM2����(�`�Pr��؅�P�����6��c�E�ڳ�{�L��(�=�X�s�j6��@U$��c��l\|	�i� �A��J��9
"yX�[��Z�~��;4��ܥ~s�0Kθ�J+�2��>c�SvK"Տ�#�Ǚ[�̦/\w��n��X���h\ʯK(�τ�G����AD+�������&ٵId;��:��a�hr�"Ӕ27�-�ˮ).$�t6����fx����U�&\�K)	3��s�>c��a[CW�0[7���[��K���7�n��E�sM����S{k+]hj����u��|���-꺰$���l._���T�[q6�T�����~�(oX�Mý�P��D������r#G��߆�'�9Vw?M��=�:��g�@2�$Aq^��m��eb�5z�
�����^ح5��Lu.'��V|��)m��yJ'x�Pl�T�����7����+޻�"�D�y��H�f�Z�	X2��QΥ��۳꽻6�6��S��`~04�Er�-�_��F�����|wO�?Jh��Y��
�~��P�����-��]�Q��H��%+��.t��l�B*���n&CdLG�|#�B�j��\c�?���S���pl�CM�o<�_G�=cN�?�= �������Ǯ _K2��M��-����$��L�5����2�q�_�}U3���Y3�s�3C�P��1��i�a�Z�ˍ�o��W���	�1dj�JA]��RyaAN�z�&�������m=:C �ɑ1�����j����x#Y+X����hC��*��0ٍ��[՚���)uL5������x�|��T�S����>\bxΧ$�b�i����]���m��Dn�!��N�f;��$�@KX�?%��˺�P����^�!������)J��{A��%4�K|�do�e��*�
��4;��w�L��a����{tD�-�x^ч(�@"2�1�,�p{Te��_'b��`mX���������RK�y�p��f���R5��mJ��Q%gg9'0C^m|���!�2�|�����*����d2�J%/�7]��[�#���S�~���m�3�5	y❦r���{s�o+��u�RFϰL(C��f�.�ގ�1q?��k-��	����ԝ	2h_�0x#ՕD˦���3<���M\�;Nbw�;�v���q�@�ʘ���7��S�m��k�+�7�=B~ÖP��u�V;3����Z<�ֻ [&��@{��Z�=i_.a�/2����h�{��p�Zb���k�^Y���p�lHD9����h�b���{([E��Y|d�s%W�%���#�W��7�r�� &�V�<t�]���~���j����34\\J+�:Uf*2 ɥۘ��z�� ���*-��5����#������3����i��Ҕb/D��O?�mYsǡY�nY�q�G�H���6�1y�"mI���J��Y![��Oǟ���f�@U:�3�*�r䥕���<X\�]?jە�2F}C��HC7�R���nu%F�ڞЪ8�.��y��b�~�e��	�P��^��e��;�
~��8�I��m5T��i�������͕�Gb�#+��ñ�����ū'����Ţ�}�X^��"�K꬈	�7���� ���6��x���;c��48Hv�ei�ե�pUoO�ll���W�c�p-|% �G��a;ݞh3��\z�)���γ�6��uի����w�{�:ӄ+v�ҝ`�Ӡ�[Ab���}Z�k�_��YhIn��L������w	@�/��%'ڠ��@�Ɠ��sos�,��N��$2C�\�;H�6�d˸Nw������y��:�[{M	ciߛ=��7�/a��k	�@���2t�+��E���w~d��M-���Sx/�(W��"
���VÏg�z�ei5ނ]��Rߑ�����5N4�f���DCg����g�@+�>^3z�]T�<�J_�ȡ� �橠)�a�B�fw;�h�|k�����s+vK�@��xB�����9;}���.Ƈ�u�C�}���HS�xV�hXβ�hn @�Z	Ѽ.�9�]���q콅Qk�'O� F��0��99��3�+K�/X�oK'Uk�;�F����1��sV7e	i�8�'�R0qJ��*R�8m�d�M 9QxN��d� �-?�[����c�*e��P�� ��˟�֋q��@̕	hh��2��)�tC�������:��'I��%`x�=���$��{?X]�+(�\�1Dv�	8��[Vqc��z���ej�q
�Hn�q�v>x�-�o��[�:�	��������I���Ə������v"}�1���>�,�ߡ!R�<WQ]^5��fKYtR��-�a����;��vZv%%P3�r�4T��W��cK�s�9scC��7��l.����� ���17ÿ� ?�����P��Qٌ�B�bJv
�
�%�Т�.�d.5�zr�����|s���|�z��;�3/���G��  �z�\�7J#s9�D=J����9�3I��D�Sm�5�K�5�+'�]Q���M@�I%ꔑ?|K;�ޛ�=4�k{�m@�9�;�z�.�h­kڷAQ�֨�������'
������(�_
2[#��>��>t1�$^v���0Uu.%�i����!�n`x��u��L�7^��Tv�]!�H�3���7U�f