XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"EPY��v��p1j�M!��j��i)8�3�?�O�mJ�VjX8d�����=fx�J���B�(œ<�f�F����X�y�X�~���e��{�r�vw�����r(��:L�,;W���[pol��}�X�u�z8�{!ċ���\�	��sa��d���P��0T��Ũ�ߘm��Y��B�dj�0a�{X�k�9A@u�(1��9|N%8�9�sg����`8ÝV���-���&���Ĥ+�kQsZ3�D�����刱E"�G�-u(�������Y�T�����i�m�\ڜ�П����"*�N���S ���1s��XԾ�A�!ܷ��4V�A�y���c`߈l-?�,7�Q�\$�e�]��W�8��^n͞��Io0T�s�3��km��h�-�kje+*XF��X��h�j�����Z��T�7���8J~��Uc�u1����9'{Xm� ��R#uWA�Ԭ7	�cfv��CN��k:���
S���<�W~�ax�5RR�?��j�0��ޒm�LEF���ub���eS ȶE����&�$@��as,����D��$�ZIa�`	����А�E3��,��(bG���'���W��`W��B�g�1ᤖ@����9}ד�����7��/��(YHg��e�=�+��Rw;��&_"/E�m~'	\��Z�x@Y���N^�����4��ј���` =a�4�Uè/�#"Wox�~�[@Re��K/z!X������W�J�$Q����D�j97�m2T5�T�XlxVHYEB     400     1e0w���.5ڦ�D��%���@�cq"O�Չ��8�/�m�]��'�=7��W�O8܎���Q�G �*��*b�C��QO� A�8'�4>(����M�6J≓+ǀ�ݙ!W��,��ܨc�s��s)3�������!���sP2~0X?d�C�g;���-��q���>��E��n�YZ�&� ��<�u��yMY�eM ��c�.js�H��fJ ��j�o�h��m�/�0�q�}Uof��}�^x� !�� ����7Bpe"���u�@t�
� ���z��r��j�U���'�{q��&bx�*���:�#���"O<R�Ǫ�ʁvɎ�Ը?�f�&o���nо,>~�t]Ϯ�p�p*g�c����0
ܜ�M]�7$eO�`Rv�&�� K��,�&�I����������u:[��Bt�-��K=,n���c�頿{·`_�k÷3P\�u��݄��o2�l��Z�jKXlxVHYEB     400     130�#�-U���\�S�zW�m۴��8��>C�c���Jf����+E�ɡ�Q����*FJ�
`����
�e�����`����t4������^�]V��̴��_�M��q2���T�.���>��x�O8!�{��[���,4
���:`�#�U�P�@5��	�I��	�k�rYQ�fSA�Ga��DO�B]�A$H��x��[%��j[�s�[�M����,Ľ� ���x@<�<Y�yz"�9d%�Ͳ����,SA�L��3��0	3[�dj�⭝T4T۾h͎� ��è�J�(�������}��Yc?XlxVHYEB     400      e0�*֤2M�E ���sɳ�J��}����=��L��-���Un���dc�p��294�KtbY���n�+�a"�pRb�vS�[�(����o1ե����;L��h.�X���BZdR�f7�a�D�����}|f]�!��V�>���'M�ΖL,{chð9���u�CA��r߾��_����^uIe*�Hm �VV ���B�$�>�V'��~&��q6E�2��XlxVHYEB     400      e0�oORڡ�
��<.�8�e��l���� ��3d���#�I0]Z��A4]�̌�ĸ�/�0�HCމ?z_�ʉ8CL�D�����vdUy2=��E��_8sv,��+� H��<��H���Pי�Uo��npq2�\����W��cQݰ��|���sG(Mo>��">����&"��lpj��>���{Y�,|���-a������O��ӱ���f�Z�����[XlxVHYEB     400      e0`S�T#��zN���,�V��%.{(@N΃�	ޗ<�䬦̘���om{��v��j�r^�Ԛc/v�ϝ����]N�����O1��i!\ �������b!d���ر�+�X�i��惞Ɣ���0�1"͌x�|,^w���ί�Բ�-"N�j	HoW�{&I����֤�-	z7ov��	���]���z�'�0�b�Od���/ԟ��"���-H�t�@�XlxVHYEB     400      e0�^�['�����脚	1���e�-�(�xp�_lrѡ���צ�cץ�2"�u&���Iڐ����G����%�ٓ�?vk�lc�_��[�/mKg���z��R7��]�I9 J��ߦ
������E��Q�T�^WDxk/Ȕ
�F9��<���c�w9�$��z4�8�͗�C����\��LO����kyj�(��t|�f��.f}U��XlxVHYEB     400      e0�3nnk=⑐�F}u3�q�Z���n`��V(@T&J�[����s)T�9�N�ò.��3���!��r��B:(�H���+u�^�~$��jw��rF���Q#��#�T8��w�7g�(��0��^��U�F��]�oV�:2��-��j��`��|�!s��z��)�ʽ�PVl`IP����c�2ԍū�_#��=Ra�i5�R�A�𩄱��(?��v��XlxVHYEB     400      e0��?��'���>�cu���\�^����IB>�l������Mԑ��	Y���N1��`k�����o]UT��-��_�'�&�6e�sp���c ��ne���AG6+G(;�	�mD���N��O�f�Po]&��K��w"y���1��С��J+?tҪ&�����Y�s�}:�Y��� �M���5��_�k��qct�Crp}2�{�~�WN���f�/��n���XlxVHYEB     400     1a0��i�<���+1Q�cɏ�($�Y�ް*�3�yG˧Ql�-�	�y�h�-�I􂉆U;N9U$�f���:2Q��mV�Y�j�2Ց�u�.���d�kD��dCZ�=h�
�^����R�嶆��U�����?ڏ���8|2��d���ȩ��2�F�C�����B^r4��������8�gu( ]�*
��*0Lw|�ԨL�����,vVwUg|b`�&��l�c@=�r�2� ��V�M�LW;6�o���P�p<�ƿ����F!�RK?�B{o��m�g���3��(pS��_�����CM������Jy���@���Xg��H�������-Wy � ������C(g5���!,-}Lk"�\�w�~��*�N�5������8�Հ #K��ײz��B2�M���wXlxVHYEB     400     110����+۪�*Zqa�kS I�0�d~`���������4
�����a�n���.�t�ͼE���@�G�ɭA�ssT�Y��Q�j�I��J����'�CY�A��_'>���ߧ�	�MS���D��LwGtj���/�p}p~����%��q�(�V ~I}�c']�%��
��%�'ӫ��-��\�x����d�N��Z5i,&�N����Z�h��j�־ؔ��y}�F�n�&Map�~�Ͻ��>f@�[�b�y�J�n-e�XlxVHYEB     400     180�TwD�e���I�E��M!�'�n�*�2����MC�|�{������쎨�0�r��ʟ	hW�oh��md�Ƈ�W}|Dӿ��d._Z���%���@{s���[iY������?���rr�F�Z;�c��� ;I�o�"J���ijZ�e�`;�H�0�j���� p%�HA�sws^=��� |��D�F���܌�bO��ȁx�	;�Nٹ���Z3�������)�P/[l�RMx���xNK��puD8����G�@����K~�4�H�^*�v�O�8;�nX���׌9=/;֑x��xN��i��D�>��E�}����Y2�^��6ж<ҚB���ie O2u�#���vxvR���_���W��^a�߬�{/#���XlxVHYEB     400     120���/�sJ�$�0��:�6V�"��ݛ�¾��
�b@�v:Y>��fj��>���h^+�|����g.��V`V'����T%��������O_��}R<��K�m3+l�/>�!���� h���]te�N��P���,�[��Kp�� F��Ъ�����e�o��IM̔��hX����ƌ}�=Ҵ����>h%0s����w��&Ӝ���1�98��uj@���KmY���lY���@G�Uԁ�����r�A���ȕ��.�����:\���@��7��CA1��dXlxVHYEB     400     130f��8$�r��H���k�_O� =���k��:�j���B�`����4u��D<�Hc<<�	����F����Ц�ϋ��7Z�G�]
'��F~�3$�M�6��w�{1X�] ;�w�	��mf��
t�y�9϶څ_��u?q��$��ބ��B�R��`�̬���bǡ�s���:��AƁs 8k��*t��Ax�����\3����g��n��f|���M�d���GM)VI2ի�Ow1{����܆����Ѕ�=��X2�]^�~����=J�_�ο|��}b3XlxVHYEB     400     120όa�,�~<0EQ��7nȯ��s�bd� /�����������֌{�(�In��$ڊ؀-�%�N5�
͵�g�ĝV1��G�4�)�e������cM�[,�po�L�?�鍲
f[���8I��4�*ݶkl�9nHR���"�S����b��Z1��.S�]�:��p\��2��t]�eb���_ŀ��f�+<kq=N����
�:	����m�D�,`�l���_Q����A���Xx��Y�H��{���Tbb���\H�ݬ��f�B'�iTm�d���1L�r��*XlxVHYEB     400     140������ԧ��,�O/�b@A��~tc ɒo�Dڠ1�����!�\נԸ��V��#���3��"6�W�3�L��@����e�d^���*�h�S�\�5�3�����պ4]��!0��zr��*j���,$@:�e3�9]����A\ ���ɉm��{4�@=fI/(�����`���rZ|9��އ�V1�g�������i���[7�5_3=s�qo��.P#�K߃�_�L*A�IIK�ͼ����0t�L]W��.ϻ��!G)�ʍQIL�_�۾�Pt�[�W�s�:j,�{?h��M�� BJ�q� �^����z&�jXlxVHYEB     400     140�"x>�ۇ�W1nC���x=�1���NC��	�} Z"�"=zÁ�S)���Φ鐽�&Ԃ�O��˦r��x�^uao�#7�b�*X_M'��ZY�,����Kl�O���@�C�_wz�y��K3���cL���p�m;4�GQ@@���i�%����z|]�X�Ͼ(�f�z�:?Z�$o]�03���>E���g�	�y�,9��!���iY� �.������*�|�5s ��i,h��ٍ6캜R&�Ύ8n�m-�ǋ�v«ḥ�׌����lep��]�t���� C���j�[���Nw[�?�E�����{O�e��~��ĕXlxVHYEB     400     120�-�w�oǛ��=��e`��)~�CJ��D:<jl�\W0a���@��+�k#)�.�4 "���f^c��Z��+z�@�0�CS�lh���0��6)��-�(�s����h�H�L��=/4h��Sb��pY>a#�鹣ӁjIșy{E���7�p2ķ��Y�l
^��j�d�q���B1!W�^L.	�oc�3�`�5e�T���#}��#��皽�����{C�q��.��x{�2�Mݞ��ѭ_�b���(Vu�v�)|k�� ��h�������48;$�����ZXlxVHYEB     400     140���@b�0�a�B�s��tt��%ԉ"��UF�?$�{g@Ž��)��o���
/$y���Y�A`w�vTп�;�t�Ϣ�#���m�������'��z�t�w*zd�n���O����n�9�?ob�\+����D�a*��)���_$�Rpɉ�MJ����pԩ�i�&������X���ʛ;J�_� '7��Dʠ�elgy�b}�̵�;g35���Gw���&��75������)Men�zv�.�q_h�B�y�$
��M�Ұ�k	Fz����Ms�����0��.��,q��9+�[oW�N=��XlxVHYEB     400     120�wE��f���o�;����f\��#�Hbe�"
*2�Z�h4���\�5G�"��+L��q��!Hxo@gj�[���O��+<L�ջ�Z5A,��?-w���t2�b
C"��B$�PeE�sխ�,V���`nz7Ns�o�֤m7.����j�����������`|\ٶ����r��lh�|gS�C֢:���f��F%��Wn"�B����� ��Z�.<�z�s+5=�$��_c���s��D��Mǝ� �^$rW�#��3e�#�w��<�l���L�ZXlxVHYEB     400     130~�ݕ��'�A��~7�q�:\h�-?BG�����`��f��j=�'��4��8�朓�x$ѕI͙����҈X�o��dv�ҏa�'�_z��ũZ[䬊�����|�[����f�b0����x��l��8Z� ����Xu�{Be����ƾ�-���X��6��j�:�����xĸWS�;���d���Xb�G�b�Z����ݪ�ȕ���P����΢�~ܬ~��fN��i&������}�BV7=f�JͰ-��~.��1���$}� ��<���h����W�u��XlxVHYEB     400     120���a����m{"��,w/o�7�^�Sv��0�S���X��z��:��ݪM�u�E+F�wZ�FH$_�n�O�|P��0�UG*��A�o��Kf��\����0%�	hO D�i��'xOi\fD8��'��TY�cl�<�+��w#�qri�圅י��;�R��;_x��E��q�����Xt�����'�S��ҋ��;�W�L>�h�-d@��y�X����TqҴ����Z�	́yr,�BO��6� =^��3� ��6��1=�5~I�j�[t�F����KXlxVHYEB     400     140ҩ6�������;+aЬ�(��n����:ۂPo���/��ɽ�e��g�`ma����L���Ǣ(h�<y3�ys��_D�1���ڈܺ��Z=�MN�>��)�"�u5{V��i�p�|r0z�FZwp�k�gV�W�m��X]� ���;H_X���E���>>uü#�����];ڶ
��{��K70
���\�l+�G��ؕ
�{���~={�(Ab
yY�� �2�����jx�+�c"��n--�����V���+���FzqW"ֈ��qIa�@��s�v*%���RuX�h��XlxVHYEB     400     140�"x>�ۇ�W1nC���O�� ��"�o8��K_�9�!�$���y�0�ᚳ}{��]�P߮����@s)lC.F����Z���U��|P��+�����В�����W�<�s�Ս��g�V �T ����|�C�=�%֛�j$�!����(h	`�n|�A���B�^��[��zhྥ�qrn�N���[H�r
*&@���,�|>��=%��;�=/&�͂��)g�;���&���*�Nfi0�S^�2}kP��VڔY���v��Yj���;H�> �! �"��H�`U8�~���,����s��HN���܄��XlxVHYEB     400     120	
�}�/��``�����w��o�is�Е ��F����n�L5ןY�P��7
��f��&<8/-��
�Oi�BjI�l��$�ۤϾ�)�b��$Gťp(������F|=��p��>�`jG�X�N|���;/����t�(��ؿ��M�>��_G��i��T��#�ɗ� !D�c��#	J&Ԟ��P*�"�}N���-sM�ΓJZUI�"���Af3�>}�4D 6 DU'����l��g�\��LX0�Pr������/M^�.sb�ĥ�7��.Ö��LXlxVHYEB     400     140����Uv��\ka��މ�i�6�2�2��-.8;b.dH�N���j�����_��=&��[�R��� �X_�,���� ʢ��͡b�k̍���,�p&g��.k�	������h���.����3���<k�e��>�gz�N�����@[�(��WW���i�����j��ߓ	��H��Ru�s+���[��OY��#���(�P���D�|ҹ�m&��2�$pZNMQ�ｏ�k'NORb�O1{��D��DaJҗ+�������؝��4����a���6G�Q�ЕJGi$i#�k��(5��Y;i2�c$��XlxVHYEB     400     120�wE��f���o<�kJ���ܼ=�iY
�y� x��d��'y�g�	"�)��2PS�$0[����*�u׌���2��Ӹ9݋wR1��?t��n$	����,��k���CK����s	��	ziJi�0�oU�-บ]�-�L�#�!��<�8_Q o���cA�&J����xI.�3C�����hZc%DO�V1��<Z�P�r[ް��~;D�-����7���L���/�Ի���c�Z���uP-Nl�rc抰̚:���D���jg�kA^pX�S�XlxVHYEB     400     130����y�.�.��)��pѵY��@?�ע��T���'�bϞX��^kY��W���褪�����\8�/fԵul�m�2���!�Y�����%�٫�#�� ���7=܈����&���b����6��vz��dK:S�LB~�	`*)؈��kA	E9[i��6o�5��n`�B�K��٣Ō���̪��˂�ñ��3�`���K��W��B{v�mvӥ ަ�����9U�A����Qŉ��r��?��T�����<}�W��H^Y�Ԟ�Ek�ҹ��� �(a��ϻ�K�K�kXlxVHYEB     400     130W4�N³��%L�a�l�.GN��-�l�g�Nr�ðj��2�����YY�	�&��u���ʣ��l!�n?y�A+t#�3Ѵ�c�? %��T@7�X`w�
2�2�r5�6���*��Q�3���:<J�(�4М��@"�ߧѣD�|��\���C2	�^��Ɛ��0��T���I��0G�1a��}�as^ɳ�ymk��D�e�\�g˵���X�;#�f§�1��Nӭ7Χ�B����G�lB?a������w��3�~_j�>����h�N���(��r�z]�^��1���1�RXlxVHYEB     400     140Z%\=���>9�<z�Ǆ��561�2�g#�̧��BF6���g2*}$�J���I�gy�T!�H5Rsv=M p� �s�p�N%}��Zl�������N!Zs��������Z9���)�^��K�n&f��2���g^���%��߷��b5Lv+�ѰA&�}�őT�G��A�t���µOX�_}"�����
�H�$8p�É>�h��<��ހ^j'0=��	� i5 �D>tj�f��� ۠m�h��`�v����7�u��V~�?Q����rnxU�~f�F��Y^�MKo�SB,�jBm����Ix#����Γ�aXlxVHYEB     400     150�"x>�ۇ�W1nC�����)no?����^Bݲy�N������ (���޹�͂yp�-����a��j�>}4��`�n\+�QHQ�g��i�"�.-{���Ϫ�Pv�� ��b��QӇ5�HC"���v?�d�Z2���8y�� �T��,���5�T}G�˫rxFҞ�XE"���Y#��o!���+���LW] z�	 j}��ST�e��X���O���C�;z]�Ћ��Q�H�<�=�Ce;���Ϸ�H���9�H9L�	�!eВBԚ�:{��yO�to�Qe��>��+|���'g��ɓ�p�0XlxVHYEB     400     120���1��+t!����f�/?+M,��w��'N���V]W�'߿#)  %Y��dga�@c�=}���M�������'%:0f8C]ԃ�x ��V���������݊/)bMj� ��0B�̴��ɑ��u�p��P�d�룞�\�[�(:��0��]% �٥U9v��|w�Q��*��7|r��C�H���L�������L�))�I�#����'Ek�T���������:�C�<�W�����aN�m�-�=</X��T9Z�J��IF�M+q�΢�xtpbjy���XlxVHYEB     400     140ܣ� � ���˲���^�a�Nf����|ƺ}D����f`�9��@�a{Ĉ����͡u�i@�g�nKSf����Ӈ����3B
�Hl��th$ܰ�mW3���%�O���`+�����W���O�:_4cڔE5�QVع�!u��%bs�MW[DҨ�'�|��{^�`tc�����w�<�a0$�Z,�A���,,=˟�P�K�u���r~��<3��c]���L�X�{ϑ�D�R|C�N�������Ztk(��O�'�?�`=|��<��.|���j��
��s���E���QId��ܧ��U�����_�#�?XlxVHYEB     400     120�ώq��lԽ�`�!4I1����r�Adi�F7���� �� ��a�#bn�H��t6(�E˓p%�s.e1���T !���${vY*��~�~������V�;���� �G�h �Xc��č#���Z9�~&����^b�A��WN��O%c
4ס/4���Eԟ�+�8��f���y���JD�v/P
'���f��w=�h�g��� f&��]"9�)��8O�	m] 9�����·/>�F^*�O	R�����b	�EX����[��l�V�?��-���Ɣ��w�9�	�TXlxVHYEB     400     130~�ݕ��'�A��~7��kG$����R�I����Kz|A}�CB�9����xv��\���ݎkF���JMk� ��o��#z-���W,���o3�#��D?��#�����m ]��6��g���٬��M����nh:>I�����Y�=k5����=����)y�Z��]���J�qBTG�w���Q��>'oC�����}�ʍ���56_����w+m�cm+̟��&�~�,����.�Ak�w��#(�s��� ������ǧR�e�cf�2>�uܣJQ��I�<i} z3�q���׸zq؅XlxVHYEB     400     130W4�N³��%L�a�c����(��Kw�w���)|X-q���۵l��9��YĬA�(��� ���O�%�Y�
�b^���-���M���9,������h�pz���h}O��Z��|y�_h��~Q�Q4~��U��/��L�%�*�:W�d��������/�M�#�VM�&	K���˸!���q���o�>s%�:̺�2�s�K"T�D-{���2�V0[=�}�c_�o���䥈��Ռ0�R��\tr^���kn/~G�Κ6���[bq K�d��і�7��ƽ��i���XlxVHYEB     400     140\��K����9�"��D���Fg34�����|�f��N5.!ѡU�E�D�?�񥽴W��	5��J�@���ES`LG97(�[�yFǥ�����Ip�l��{�`Ym�3y�34��a�~�v���_^![^V]�/L�����x��s��x�0n�)�����`��<�w�J��-�e����S��9�~HB��t��=g�c�U��������tZLF��?���}G�;i��]F�R��^2i�Qѐ{/n%^* �����4��3�u|X�T(�r�3(�2���m��&]H!�2rn�p�O�eMa�Ŋ��9O5?U2��XlxVHYEB     400     150�"x>�ۇ�W1nC�����T�>��7YpF�e�+�2$�� �z&͒��4T��WA�ńv��K�bݰ3]��Z|9��H����a���
<�}m���OO|���n�M0�Kh�����?<FB�@,8uk?����!m�=�ղv56��$���k��i�o�e�l�W�_V��/\k��Wä�����;>T���/
����
�Z0v�׎hB��3˲�s����
�jz;^^B�^�H�S��h�)�4�����z�9XS���r����6�����IR$������y�k����e �7�^���a#�����*0��¹�O�Q<��XlxVHYEB     400     110��t$qg�`�OV�����Ϩ�X;˨6WJ�����&�����03y��h�k���դg��\Xx�~�_��W���J��S�A�QSUHZfΚn��@hg��8�����h<8~d  ��]�9�w:w�ǧ"%L�?l?�>T���]�)U���E�L���L�+g�-4wy���������S��z��	(��\�*V���:�^�)����Q��ٸ���.�H1�q��z��nO��G�����U���(�o�>���x-�v�|+8��|0XlxVHYEB     400     140�&�_�3�8fO��	j�Q/�s�	�|S8�x7��ܡ���M���4������(�z���"�-mEA��w�B�U�CE��Ӭ1��d��o�Ž���j\Д��Ɓ���d>@8��.��^�4f��PR�Ι�����\��Ƽ<�{4�Q%�preh&�a�!Ů����oo%�=@*Y��T���ԍ�y��+~@z�s�9c�T}���+:��Gw����H���p�n���2m�g�$q����f�D�M��)x����W�i�[�H�9��:6�nȧPjw;/]3[��tC��?r�}6-�6�+`����_�%�%�(#�XlxVHYEB     400     120�wE��f���o���twm��qv=Vj�ʑ��!#:�c��ycZ����_߁�wEAt#C�M�Zÿ]Mc1�5fn�<�a�mT��x!t�:�f�OKTN|2���K?bO%��,����w}PHQc��:3��J���+N5ԛ�5(�<H:�B|�[!��P3�C�n������V��6+R��I�8%�ϊ��1�Gsm��f��lՠ]�N$�&���M����j=P*�-�7��}*@����>Bj"0�E0��P�3��h�>R�'c�?�u�D�o�Nd�ϑXlxVHYEB     400     130X���n�g�r�"d���H��y�Wy�D������h�^:���"��t���H�����V�H�G�x����`�y{:8��T?;g�
��"�;v�8���C�47^�4��8S��+�]���0���"�"C�? �$��ԏN#��k��@�X~��
d
�(��կQ�(y��d�a�* ��sP�7���?+Mm`��3wUB	c�6kd�����������l����Fe��<��6Y�r�Et�B���!쮽��Jgl��7�~��iye����V�̆�܊�YXlxVHYEB     400     130 �)h{���ɼ�>�Th\��S/i��yO�!��l�W��^M�+`b$x��F������0�n���Cn�YP�����X�\0�:Z1.��K@e�D"Ѐȥ�	�Fj�&M�E=8_�i�	I'���4����� ��&i��=^���2��_*Bʹ	��b�l���'ፚ[����ns������V�N�i)r��G�D¦J}~��}��><���C�#�~�0����d��K<���z��(����Qȉ?*^�=�ήZYH�˰?�I��4:�ɚn��i>3�\<��_�{2�XlxVHYEB     400     140��W6}��,�q�z��E�
|i�����tF'��5BSo�����I=���E�m<��p�� 6h���{�cð�5���ZY{���݀v"W^Pn.ҙ�3ۇZt_��*���a/�#��O&�ɢ�ܑ��~�޳��A���q9{���^0t�w�r�F0��	D+L1nU����C<�2��A�R���җxҤrك˺�L!!Ķ9��B�|��:(�O��ϕ�?��_�`-���������Y��D{���>ɠdY�:U]՘<� ���9��[�J[(�����~I��Z������ׄ�w�=q����Z��SF;�)�rgH>�XlxVHYEB     400     160fDP�R��o��f�+���o�ŋ����R�G����{
����)wu���c��0��a�l����kF�sv.B�8�pst�a�'�<�'=���d���&�y��ߡ�������Lg��Y�iw���ET��� �r�9K�b�\���_�26ٍ�.�S����p�<���HF�O�y��W,7��X	�Ȧ�9��������*�=,�^��,��97Dz츥�a��y7rV�O�<"Cy�#%��3�lX����H�1g���T�*�A��fg��w�}�_��X�Hq�'0~�=�+�o���U������qG�9SNF�`���޸��] �+�Ǘ
�f鞤XlxVHYEB     400     100�@/W��-0?�9��Vx��e-���s�Rz��f#�u��FL���g��[BN����]���^Q�\�#+������R�T�s���a����n�:��S��4@�l��s�å�.�ŀ���o��bF��2B�V-�R�+���?��u�e!<��k��V
B���NFM|�R wL���ų�w�Q��R��~�h���ZO��<w���>����{ewf�a*.��ܣ�D��lQ��O�;�{Pr��8mXlxVHYEB     400     150ap�]�!ȋ"�/�<]�5m��8n���$��1*�k���������i��:V�HgH�"�7�O���W���o���fW���oj� 5��%B=Ne�����^qƓ��C,�Cx�'���� �(vFY��J.ۍ����;��G l_��La���z���!t�w_/������������	f#<��r]t����Dfz0snW��If/�Fg
�+�NߣE�O��,����T��mi��'Ĺ���|����zsL
��]���Gߥ�ӣ�BH�~uo--��6�~|��k�yX���/��b��V2.�񆵒syAw��h���������%'Ɲ��XlxVHYEB     400     120:���"D�>�ę��O��t�UQک����;��u�>�p�"4+G��jI�j���� ]D��t�UUТny7���1s��9Ҡ|����W֠cq(��DPB����l�@�9��sb�@HTR3�����V���~wt %���f����ꊘW���ʹ4BM��Q֏%i.�*cV����(Hn-�Xܤl�}r+P@P�#B���ނt��TN*��,��$Q�{��¯|�=��ˁ~��@����.��P�n���ŅL��E�?����)�Sd�~�ҕ0�CXlxVHYEB     400     130���|��?�[�V��6�6�x�A�5-�^�pK��abW)�jp��Q�^���MOz0���]ʚC��!(�T���pK7�J��;���c��R�!C�ðQw9;{-��x��zKͬ����L�[��k����}Lf���;�'nkl��$�Ԁ:^�:�:J�S��~S!��Y���_����+J����״u��y�/ח�4@�c��D��Ǫ����d{']��mfcٰ$����P���Մ
��4i`���a/�u�b~^3q�$�$�v�㛢��5�E1$�k"��/M�z��\K���Ws�XlxVHYEB     400     120A�~у��p�_�����L�}M��8Sr�LGd�@uI�['���bp��Sa��sB��ލ�,H���0�a(��n9o�W�"��z��Mk ��-��{��/�6�S�\�Q���iw�2Ę�U='U?cJ�N��
�����`�!�H(%G�I�I�����c��c��KP����(=���*��\렼5�@��E��+��=�$ J��xEA9�b�u�[��'��eW���V	3����S��I��qTB�D:E4K�}[�Dk�ղ�1ú�FXlxVHYEB     400     140Ѐ�Z7o����hS��7@eY秲Y�T��fi�x�������b�?�=�L	�.:J����qddۉ���H$�d'��4��&Q"#��E���������5��	C�Hv�#��ܠ�>��Bm�j�hSn`�ْ|�2��F��=?3{��w�f���j�����L�TY��S64?���\@���˒�}U��I���g]�%�=H�Ih�ɼ�:�*\e;���!��b��3.�	��8���|�F>z�l;�#�|)ʿ����@���.�����(H-(2�yAK`��FdII�MbX������n��͡9!h'jn\ٙKXlxVHYEB     400     140ر+��~�s��_��k��t]i�/P>��N4q��8C���|e#�� ��l̨���(46�:��]:9JW999}�C{�2�ߒۄ2�'P��:�S$��7�d}��t��T�o��E�߷1c[N�NI�z/R��vM���b0��znCJ�'�H�e��~���=�8�]�'���@�O�����D9oGYR�
�\�V��%	QW�Tx�PF4�z��)@��K�|�帙$�4�btj����k�g���ڟގ�/@��c(�+F�?y7!�m�F w4��;<^�[�2E���GomX�#b)O�㴱h��$�6�XlxVHYEB     400     1201VK��uNx1�,��8CIw��GM��_���m0,��%a/hR_��T7���˱#3��r�HӳjwᎼH��z;��#��;�#It��r�Q���3�aL��z�Xz2?��׾M���] }BN�;���`Xy��5o�A����y�����y&>�ӆv뒙!g����{�b9�L��?�he'���o�F�<��း�zj���74��Հ�OR:���T�TN(�r�Y2��bj�cjh�8|`H�Ip�QG�u$��v�.�9��k�)ѴF���PgXlxVHYEB     400     140<y��c���[Ql���2�B.&��8�Vl���Dc�^�Q"JF������Ddr�y���?-ϰJT����ƓW	O�1}6huL�9��a߷@�ؙ��%V�D���1��J�yS�O�h��>A>���Ūǽ}Q��D9���̶��h��"Q�ů) )d�� ��J��$	�D"�# �Fe��=��u�JD�zg^��H��b�B�?��RÙ��������cW������m㉦�1����,�Vާ{,Gl�B?�"���`�)d�_LC�n�ӠgS��Ej�8$Hs ɻ�I�|,x�[ABt��XlxVHYEB     400     130�Դ��J�%�nA��A�,Ҳ-��o�-Aq���k�p��`��q�>�exfY�6I�˼W�T��#5w0�~`��_�2F��E�r�N��9���R_'zyR��uװR�#s�r��F.R@�6��z�d�vq~��*�Z��n���}͒��}	��u=o|blX2/��̺�S(|����Ip�xu��'�Z9i�'�,U��� ����jY��ր��j|���F�/�B�`�w�B��2�+<	�eQ�V0��-����)�[���/��z��9_-��PƝ���؂M���XlxVHYEB     400     160HE� 0Y2�t��8�1��)pT�����}{��S�YH3򤸆�S��d1�'�/q�R�w�!���F�
Y�'��«� ���������/��PQդ\@ӬQ���d,$z5��g���s��BG*��	��N�E9�Tg(Q�Ҿq���lO���o��(�:���A%#uߤ�Dm �Ib���3*�_���6��"5�XB>SL�|B��q��$ȗ��C� H�^h����r,2�D�q���l��Q5�<ЈP\PD�;�1�ӱ�I%�S�LlC����;*��JԵǪ�oJ(YɢNJ���a�gh̕|�������}H�6[Kݭ�3�����g������"�7XlxVHYEB     400      e0��sᓃ�S�k1.�۪C;������+��C^������ѯM^)�4!���ؖ{���$}=wy��������ڋ�o�����nĤ��G�Fc��$,yq`��Xkn{�d�N;@�'?G��mz�|9R:�J᫤��E���+�z|���I�ԥfW���ۺR��L"��Q���G*�8ϗ8G
����8]�?��P��*~����ĻY;�XlxVHYEB     400     150h/H���_K&o� /ug�����g�\��+"��9p����*%����^�Дp�!m�N��h�9��F��W�)��w6
 1Q�2@:o�>.zYr@HC���4z_*����v1CG0.�_�20>�P^7�'D�-�Gi�!ͽي�3��`x���*�ع1��R����C���K>��������7,�����2�|ĝ+�o����˖/{��͒�
�}˾W�����Y����~?�����P�߈BA�T���OS�Iéo�k����%_�=��øp��%@%��%�m�K�\����6���`�yz=�9׬V["�b �/u��XlxVHYEB     400     160�b��.2�y}PF�.w��,�O�uz��D�u��n�/��y�4������g<�P[��<��e����q��G�0IfԄ��R̆6�������2��� I���M�1�2oy�V�3J����z0N7��\��U��������ɵsA(ږ��
X��~4���B�ֻ�{Y��;�C1=��B�Ѡt=����"�!�!E����_��� }�u��ơ�+���/��eԊ�|��:�K]O�)���Ǧ����A}k~�+4/�;��ݝ?Tg	�ɽ�b{J��+ o�t��6�O�`�B(�� ��A���8��_I�@����-���f�zq��|��t����ZXlxVHYEB     400     1201VK��uNx1�,��a���F.����Uf�*�,U*��vQrBD)�k�!ٍ�d����zz�R�Ց�6���spg�a^�7rA�|��g��J�c�ӗI�f���Bھ���`����z<�J�J�hG|2=�(`�2
� �k}<]>:�hҡG�)%6�8r��4S�XY��^���{7��j��~=S�y��s���gP*�������n���_�;:�m�7�'U�.��	m��a�Ab`gz��K9"Xa)pw�Al*-��-��D@ '��l1]XlxVHYEB     400     130u��Fd��1�9�L���h9
0������v*�� ����ô;�|���o���b78H�U�4181V�	��N��-*��Bm���j�s�#o���V`�v~.P�v����ʼ{亁�YN�(��v�vR�Z�t�&��T/h,g��`d_\�d�dy�[����3��8�_+VTn!��|�e����_���'�G��^ˡ�j���:E���آ�^�hK�c}q>F�s@���#lޗי�0B���I*$���W?k<��o�/�,��IN�� �w7�*<X��*?�(�)���;�R����XlxVHYEB     400     140uVR=�8"9����%�m�v~ni��ߞ@GN@��@޴<T~��ǖ�4���Ʉ�۟$oJX�ʇ2ZN�i��\O{A�},>��s�=�T����z��*��~�L�ض�;nmWbUە�v�!��gf���g�^��G��]���t����d�@O} ڦ�շ�'�}>r�<�(��~��&6���U���ɨ",'��8Ȗ<恸=�*��SG�c]���'hb!���K�[x�c�w*�D����(������J��V��C"���1E�H5���l8����A��8�|ߣ���^^_#����qsUw�S_{�9��XlxVHYEB     400     160�8=�!�4u���	������(���.��1#cp��c��3��=�$��K
�9mFٲ�E	��}���I�
[3�dDk� �+�2�"y`�Wh�E�{'��@r��O2Fà�Y���&�q:v,������߲���"_�_�� ��A���Cin��Yb�zy{�9SB�8=��t��������md~�w�]G�=��Em����,Br�P�+��'�.��eqBo'��Χ���g����}�y�������бCL]2>/H�Pq�|��p����4�@n�K�<4<�[H�S̛ ���a�^�,�	1��|N������(�)���P�M���F�8��l�[�XlxVHYEB     400      e0%��p�Q����1��.wv?�-=n [�SU��C�*�ۣI5<\�2�����]eY��Ϲ��}���
�ض!l�O�%*?���Q���i�Խن�niߌ��6]B���{{m���wNh�krJ�� ![3�>J��(*B�z/ܯ�O��G����f����A;��UMl�S�4�M䵟Q	�F�����a�e2��o-T#�z4Z~��]���my���XlxVHYEB     400     170`C��DB�Ҩ�q؃.�g�s�$�����21��ބ���-��C�}'�'�oP��B#m�1����)k>3H�V6S(bE������"�	��{��/�=u��T2[��� �i���6�>�˦�6��/�K"�X��!^,��"��͔�O->L�Aꓡ/�5�#WF���5��)���%
���ڶl!^����ܺʴ�%���0]J�1���`��q��FGu0TKi���3�#UA�p!<�ȸ/3z�rdr �HD���.�<_oޙ�p�	��S�A��\?ͧ�!�u�1Os�g2A^(�˸JV�\j~i�����/��´3&e���i[]�ďs�S�+R�󋛷ݯ�Y����N^l7�2�XlxVHYEB     400     150�_F�P<�K�x�Q�=a%Ũ�
މ� WG��A˺�Dd�d�+vJ&4rc
�c*��/-�}����V��&1����S���`��(tgS��a.
&�$y�����կ��8?�@Ȁ��e*��''5���W��>�;�g�n�K��Ri��={��t���F��p�mƛ�E���ODƽ�/6�Ӳ��h8�H�������J��bK���U�8}����^��2kԦ��9�z�e��D�D�{5�n<��&h~+�u��/׫�J��l�AW��>2w�:v��͌�f;>y��`z(�p�nS!ad/՛��}�Ǜ�{B;7�]KJN�Z�XY���XlxVHYEB     400     130pE½�y~�L���0y��r��X��@P���zi̊��ó�2��%ڐ>ԛx�
�W�P�U��gN��?Bۋ�r�K�g�K8�����2��%%�(�e�ɛ����Z�N9��o$�F��m/ގ8A��jJ7�A�em���N7�%"U����u����va>�S$s�Nc1��4M=��A³� ��C�;\�����x��]ވ-��vItW�rZ��p ��s��# >���Z���\7�4���;�W�7�"��Z�"��.-�%�|�i{��<��э�+�(����s��'�XlxVHYEB     400     130b���c&w�����g�ɰo�����A:�S��g]�LM�wnC�̀?iឞ��[s�b�d
�4{M� �Տ!��g<�� ��N�xTI������h������@����
)H��!��>+�v�k�
�1=j]����܋Lf/P�y����~��c�RZq��(�^D������� ����h�3����4�\�:@T��ۃ�0%��E���~��4��@�w憩?����r��$rW��ΐ��H��x�ǈ;����]ϐ��v}5	1���5�k���(���@!�0�p�2?�\jˍ]XlxVHYEB     1b3      e0ͦ���!�W]��$>˓x+�<eK��8��W*f���;��$"G	���;���]�($�WNy@䢕�FE�#��n�BV���s+�ZOxН��W�<7ϝ&�y����$p+�����mѯ0�6"4��q���.�i���Ocn��gѰd��I�ZC�m��ae�C <��Ib����)��6���GɆŬ�U�X���1��(��0�u%�عʡg���