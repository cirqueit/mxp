XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���3ښ���CjF�XTx�r�8`�n{@��c	\�q�i�)�Jad�G���1�-	��~ص�]w��Y��{п����>��ӓ]�"��K�0�>�?ypa�hT�;��t��h-����+���Q�c�)0,R��ԐaسO2T���?�P��yI�	v�*�@�;�6���K�t ��+��)�_ʿ8^���P��/��r�?�q�F�	��Kb���@"�2UJ���Q������hh����w����*�"�d��l����z��ΫS4D8d�=WQ�Q78���
Z�s>qĊ�şD ��
�k]���9'��!��9������!RY���~1.�~6�Ν\��	��0��A	Aj#�ci�����N�����[����&z��K������q�
B�3��<�B@�oh�r�z���&.ѵf��ێ̵du}0�p��h:�ʄv<)�:������/.����y�(���-H)
G�F,�q_�H�U�C�5��5l� OTĵl
yC��M�p6)�F����H��W������nP���]Ϻ���1n��K�^�j��^D����+N���f��uy���{?$��0X`0���dm��|���F�":15=��w��#�l�Ы��/Y���ֈ�,��,_�����ap�\m�(p;Ӵ�g=j��=�q����k�iq���H�EW�~��+9qݨ���)mYr���'� و�a
��s+�����eƃ����g?HP��XlxVHYEB     400     1e0�B���aE������J��s��}� ��+�C�.Id��N6�c��Yu`q��)�"���I�&�ő%�5.�m�5����ʺ���#O"8��&�>�9W���[�OZn0���c���kZ��٧�%%�C�<[���+Gj�n)v�U�����z ��=�E����A{It+�A��ԙ�t�(	�j(��S����s����ׄu ^�g�9���]����H>�V>�ؾg|�&���Ǳ�h�plË|��?�ڊ�ǜ���(G�Xc2��`s$�E��'����}�2Qi_��P�M���g��z{�K���6v�/<��Ǝ�RM	g|�P�����v'ۉW�,w�Hd��fQSC�Y���W3��U����`�Ħ"����t���XSo|s
n�%D���,{)�F��bvZt�d���g]0�.��8▄�ׯ�#���Q��崝0�铭8�P���O��z
r~��MkS�9�X��XlxVHYEB     213      b0)H��b��scl���\��a��J?`ZÖ���x�3�]���q�N�����g�G��z���}y۾�.
��b���h�/��n\��<⠍�Y��g^V�8phO����6� ��ښ�D��\~͠k�tuV����䡛����_��J�.��I��X�����M<xY��xs)