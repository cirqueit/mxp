��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��л���,������SE;��QNt����8����K�|aZ#�%��I��$��A�t�|Q_�8{��c�٭(���Y���,��Q��>�]
�Q�FH�t��-�GM�C\�f�M�1�/��楮���ܾ
i�505�^K̛�����P�G8����sUm��}�[�>\�E�����&/�&;���>����{8g���|������&}8!����ĞFJ1"}�uiP!*�uj�z4?T�K���
����gr-o7�9�� ڏޕ����$<%�+�Fɼ��Iù�[�~��9�SeG�{!t��O[��@"Ϫ�jZg ��;�?\݌��!߱�~'h$BC��8ݳ����:�{?����W͔
�iئ������/�\1����[��`�B��z�7�kd�Mӝ��p&��H����_cv�o�V����Y��cr]�8����+�k��=s�	�l�b:3R	&V��e�.D���I0��F_+�t���N�b1KU��Wn�Hބ�֙`Ov)�М2�{s�E�'^Nq$�I�<*+}��cF�1�~�p��+����m����a�qZ���j�/l�t�a�&D�p{\����nG	�63���u�|�2���Vg�,�Z�A���44���R��ݹf���q��@R����뱛����pQ
p{�id��bz������5��O<����.�Ei��R$�9HF�6��m����578������e֝>e�مA4ȋ�5�<t��ǡ����Xⅷ��'��bq��kS[m��dô;�bC;���<G�ϩx,'�[��ǐ�mgz�S�|�7�+1�5#���h|���𾾬R.��9`�nu���	]C�A�2��}�+��'/�v���+%y�Y��	�8
�04Ġ���W��-�;���ǐ�|	� �qZDYf-c�ɳ���7��H!�����D��C����	�W)�eF��.-/�u�;���N|�����i�0���fjw��&�{�����bZ߾F���֝�����q�!r/����6����L��(�`�h�2�LzW?��ǅ����0A	
4��v{��AY�מ��jr�ɶ����QD��D��q��l��&�Q�
��)��hFYb����[8��K׶���mK�+����\>$	G�x�*�y���%ʦ`�Z�q�-:�,ց�����Y�;ԩ"7���.x��mŹ�5TE:?��p�GyNg7�òm��G�\��<���ܰ��-�8��HV�v¡2q�R��&`p��mk�Y�C���	�_�t@���ƪ�)'�
�r��t�u �	�\�i��=�M�B�1�ٖ�*7�2}�U��n�g�Qū�P�%� K���*�-_\�[��x�˥x#���o��0B���%��r2�s�V0��R�]�Lq�-D-<�{�����^K�i2�
[D��[O�RF$�3��比�5�����ʾ�����J�K3��B ����5Cm���	�B ���%�q����E;�Jl�V���7tV���a-�v�<�yb�Z2�rN��VJ��:FU���c�� �D�x�i!W�p���63�~%%K$WHlļ�!x<s��o�%پ�9���)𺨈�i��Nb��!�Y�׬�Vyy�B#�-
���r�,N��~}z����4��������]�X�M��Ig�R���i�	�Xq��b�~��79:�I#M�<�F��k�&���P�3����Cmôr�}�g�T
X�x#|�
-i��n� �x�M�HP7�
X�x�qjA�H��8�0�Z37S ��K��^[vеG> ٫���׋	N�:�wp���5����jI&p-���� 	#ȅ2�0@�Є�����KKr��7�8�uS^z	�'h���y?E�*[��?1J�<#.]2�l�l1%D+�ސ^��f���JA�.�v�!�ٓR0B�m ڣ�i�>��[���ɭ�Z!�iM��Lm�_