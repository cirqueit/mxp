`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25184)
`protect data_block
htKPebm3a1XHEw+hSdSp8qBpXd8JKisu0HrE7Ng3BIgL3OcD1fMu0xFiVgWrA6FVror7VgQ8YR+A
muU8hCuX9t4OKyRQBA87wHJzOn4kgcHNmf1p0O9LjpZGUHPDhglPnvS3GC8pHHBs8PJBKbkjBVY4
mOeX4YJ7sdkzFdHdbfWgGxgZmufMoos6MuLdX8DnjSM2KNoR/dWHOndybNMlaCjqvgSDs0E0Mue0
M/FavHLm5aAoK5ZPBsE6Z4N5Lre1WX3Hno08+XULTT7ivIDLrKgEwc4iUqjalkoFqi6uGCAnRNl2
yjkCVaRw0hxE0n4bdKDAGVmUQp5bQSyFUijPjH2knoF/t0xa7gq8H0vyCUCyKWrchadftOv5/em2
Q55hgQ4NkxXyA69Gq2BuJUvgfjaZwyepNwKsroOznZxJw/rgOX9qkC16qpJWSpDZeSewaZrXv7MU
B1MYLtYyMYbD1yZ7LY2pM0zQ8S6mTfQLkzRfMQcojVbciLrJJ3jxOg5Q6bHyUV6G9q1BlnuMhDqJ
9JQ5jVB3y478FpG928ypIdlj+ltCaro3AHUaQFOYMSpvttGugNpbj1lsf+EeWYpjLe4rve3Qo08E
CBjMEyMQk3gprkfz3CuJVT+5i/TaUhJ+xFLe+f/RUH4esH6qSt3fEykZJ3SBZ4UYgQXinVKEUAKW
e2WcWHhFTne58osiBIc4BdMcF2WMWJjSx/dCKZKJWzujc4o99TOLm3tsgdXjq3I+HxFSGk9trNbx
ufEXIWvYXC7TcB0vjUAkaftiBSwEU7yNmumE8GaVfjyXoC/COCYxAm9y4xSJVJkTEi7WU1sWr52r
5avAyG2lzhw1dezXDR1fFhm8HGv3/fjOnYy9QHEOIM7bUMNURv2glDQfqIelaocmKDqxdaObvHnz
qukOdEWo3DhtzLSto/LEDJXNFjEaxS0DasFsZ4D9DYjDlRrcxttBSS69aE8hH8CLUJQV20aDIOb7
F4dQW2ww/h3nFH0qQEfFg4EorZ8ev7ykVTEkoiUh/tL3iGXqZ/IlXSLWtp7/6czVvKPWUGGzmewf
6mJgM+N6ufz9Fs1A5g4gGn618LyNVhwLnafyAzzndGxp51XYWwLw7cjNCH0zJHQhzqF+vZcoqmgn
Rvd1SNHWEXkaOusgnnDvF/XaiZKgxRk8+tmuFc5ZaFJw2uOtfqaMENLgpwtuMk6KPMbos6Ss/Mgp
iHK4gFw9Gbl/8q0ocBI23OIIAQzSnTtBVF68o1Qjk+vzhgCZAYVt6PaBVHpvFUik2LxOGLmwyoC0
8nRVI7wnt5u3JMDbZ7f0OfTJEyDr+y4uZ9yerMQbF+Sr46PaGIBD+TeRMcsIgFLe3xRUWF7CgpAn
kkID7Xhpl4axOoV+KMmT0/zIYcJPCpQWllOXVXS8k3HyTJUTdpABKFKTthE1dI+dxRr+WdGjzP/U
xSBjjGxsnS9D/VdRhn/ArhgNGtijWHprg0S/xT1DjvtsN3LCt9UZTaormUU5bD/d9vy/nyCkMJX4
s6orFzQNb2j/9J9z45IB1iVBIm8XqI03OTt50kq2d3dx6mEPm29vnmo+xqjb643uxEBgPuElDUv/
hsWBK/QHy3CtsLHi2WiviOz0leMeLtJz0nHLDuuQqgI7oxxgdOPAF+3y9Kp37T9w4ZyDNVzClfND
L3JgxBuSF+RQ9aRg+UoWb/uekPmCFCuHgQRRtERE+gm0KoOWJQxOPnIm++ZdLZ7VskD9668CMeOu
weJk1rvfZaV1XfyZQ1dQz3ousADoi02H5oIwr+X1BjDNK/ySF74wP4u1HVqticEe3il13DY2+u2i
nAfxsG8g9HF4+sTZtYb0grJL2wzx4zrJPmMvaIt/s6jv1nauj7WonPTBM17MQGwKcB/DvcKfyK90
W1aHfNDHnEkq7KfzorGwOJAYW55zUSULsKR2ARtLosq4tn+REeKtYbpho4qLIYuAXE5k4Qt3KfRl
WfG+JKI2FqGJ+WQHtREgAVjL0R+1VAvKE2KSDwGnotvrznA/ZAjtlfYTjJBb8SfDLfh3LldVJ4zR
SWFWjy87vJOUYaWgAyGzXT0HQP9rlGU/w6zwgyVcLPvXC1f1B6bIyxDzvXHBSaz4U8dTbR+SHwWa
b367fPWwZCe0HP/1aEkGQ3+Wy+vTWP4+aVMNZsrZ1H5GAkZChkgasq9mcwe/OdMo7Lw1RXRnV1bE
d34gQr49oo590fOgiS1Az2NpsniAIgDSC5l6f+Vl4eX2tmJSD4RIVOwqUseSu5dYvS2O3Xc2whqp
rTWr0nDTudtZeS2o2/enQp7aj2UW0QoIDVOyN/UJhuP8nwSCmuLuaMna1VyT62lZ/bkr/7MfTbfm
olV48P1cdc+tRttYQoRtE69NDcqoZT5Nce0Rmi1tMS2/08qvS7sb6sJn4lqjJG3wCrFpffQCs7QP
YT9EMQzMx96Ugn6mHeDytBNaBqcEZ3ZyEvO74eS/Zk+0tQFU3oTwr8twyTN5nlmZMkbB6Xpozw2U
iSvjWaRWODuJ0TBmB8gxHyrOBRhb/M552AZOEYRGIbGRCKa6HBun1igjAlf8l/nNTD6D2LdBCsP9
SQIpUgmhoeCb9vnE+HBFrQg3njEErXtQDYr7YnDU6uHaqco7oFgaaGEaUAqOKZsosHBAa4lNgEal
aXNTd8Eimeznjzmk8YrJDpDlF6d89RJXsM9XLRX4YFjV5YRb4d9SurWredswI0Kx1SXPmIqb7QHK
1kxOqAXXx3it55AsXWxCHx+mRxU4xO2ggugFge/vSyBzm5ufspeR2/gELbDxTD2EecaR8Df05HQk
7bJc8LBjAXsXVDNPDiajfcwnbGV/1M+InL00w5ne15p9duJhlSp7u7DY+TsOzOeOLnPck7/SjnEv
CgPy2fWAoc7cQGb1MO6NjVVojECZIPUuflrRjF00gdViYOleyR1T4PBOXs7ZqNDY0xRmg47D6EwE
3I3/UlbnqF/gSCrQk7OzP9oRMj2sR+CqqFFvEbh11lugkhJbG6hxSLIFSQG2JD2I2k6Z9TCHcYyh
5K0pCHL4ACpr4IT8sjhlux87EJSTebdtKpkdI0paIlN14lKPFIwmf34A6cGKM2rbxHAmGNJWcgYI
KoGmzXsn4JufR65TeVBdkCRXuvKCDYQ6HcDMerS64pJaupCVlP9MfJM02uTJvc+IUiIFPa/K2TyS
eAmud/wZg6rQykT2yoykQ1pPfmcoH0bXb7SDd1imHMmMteWh0Y+rpeAn4LAF7b5Zoi7fqk00HLOo
IM6Rwog83m4ySVJAuXBXX6GxA0vLI9AAwH56+zJtE1uML1OaDrYrTkEuWxqcblWsZvQBFFi82n6k
K7GEzSjpYrokzZpmZpWQwzNNQVQc0sz+hhofPKXKeDBdiRRQyTN6/UhSq3qhnQHH9eszTPAiSS2a
Mv6pQFdne25D2l+YikK8SUR/LH9B8SjpwYpERmtswnuP31ytWI2eGh30q62wRqGaumTFr6OUdwfD
MEY6lEx5dYazLH5yW7dHL9jMuZDVWs7pyjXJitS6dMJzH3hnb+RSTHkSDESsZs+T5kx5bff6gTM3
CKMsD9MYPqWFgNJzHpw6usLTTVVtM8uoDf6bucEYLbYmo7iqJDeu+eAEYV3BHRNTnsC39jI8bigB
xxOGT2WXJkxzf9SULEkWCqUcCbk5jeUCkwLwXTbx2DjicntUYTLEsqcOFN1xbtUi2c2LgpXF3Oko
ANBYD0VTiwpr1rl/VFHLWXw6MIiTXdnU82o3gTnU/rRIyjhKJ6nyu3O31YY2m0oM/ODqhy3busXH
fBg2U8u+7dfYeTxdCEbhQ6kScVMmGZK6spp7Yt4W1S4lDpj6CdnVRP5VqeM8pa5f01yyNsb31QrD
jEwzopMEuhTFaDIGYqnVcp1V3Okn/aK113fv55ICg71sMR2QS4ofvVnLY1YtnIZa0u3YoMEOMw5/
WHGwdxRLxmFLbs72MDYQS9ciRwSgrgVoZX+uX9TPcAIzxwlzIscFAeUjylTqowWWcoXI3iSYVH3k
hWhTQHf53RAVi5GYK/twPxFQzyshE7rtH2azBLBkZJhSh7d0OtxncjdJmLi3xY9bOqLOnYGqo8F2
hmx3uU08TbLsh8BryE/j0pbUvw+vVOCZ/Xazivj1ToCRPHhuo5o207rgkzhbRjj+VAgCGsKHMcoS
KZAict9YgKsbnW/sZgVjuh1aTdKEWmUIEGXbRUSuTpx/AhVe74nS0w5Ij1ceQJb8YLtweIYcwVJp
HCsDILeVd7hyb8W3w196v27BpGZo68in+CMkeci5WsB5DLx7eIGlW15hba9ps8medXe6DCTKJwOR
mGViBWii8tvLbwjr7a8mm7Gz4B5KeREg7Oi0UcJyUxgZczsM85NIrY8D/JPm5APMInKpYekI8P/t
z0bC8YhpFEWA5Y/reJYemLvIb1Zk3mXmHU1XGExcYRlU0J+T07y3GXfc780Szm28YGUNFKzJBGFJ
+jG49am9/chmNnrJKkQGj/eMPsbagRfyXBpCdeq1ZAn/XkPKFL9BWLO3Ccr8u1f3I7ffVGcKIsIt
Vj0S0Koaz3i8uLPcWAdTJLsbk5t9VIjd/0RJKNUP2aTmVjizksEiiSYLC2pJ8u9G2knSBOvEG0dr
cskXIs+6rqfnSMDXkG4og9ADD/s5mNbYwFsgGneXsYA/YGEyb/HpqxugWfkDmfM9ecF+bSQJRRbr
gMKejD+ciyokiX7jECvwniIVoSnYS5nyaDVM5k12wS4ZNjU8mmaI0F4tpyP3VfbOpJH7vAkcWjzY
FXG+MNKY4l84/CtU79bfO472t/JtmTKsHKDyrVFcoUrWYTMCsShg0l1F5Wb6H6/NISGlldSNL9PB
XVNoNp+KUALXIL/BaTgNrxrOKU/Fi5z5FdR/ZKHMSUsbQAQIymibvSnzbXzm49NtpaLQNDg9qHRX
nUE1SrombcYGJgL1xyPr7WDJShjDfYAD4RIXGftt88Ktpfa8jxXxW6Sfg4Q3zVgDgdBwoQhrwGFw
czbLzhKNQgkHO4hIcGAt43d+m1/8Fyt4Ozl2UPksbqrt7CWFYhLHXoR84VXdWat1ZyZ+uejwcbJ2
Unhh6dCO3QOkDgS2YDDCn4O7YNsrmjoVuLQ8Fo1R8qOXloqzOe3rM7LjvojXCUtVgaO30E6rrqTL
2GJ8mgeDKLKEWyCHfE1S+DPQ2VdZ+yK0CVhj20IbCUTcz/xKlkj7Yakr/zIB9+V2xq6oGvwfBDbT
XRgpDIaAmYqMGHXI5C+Wk4iPpuSvfx3bbsWzyzgt2TTd0P6zkeaqWImpSvQB6ouZLaFzZLvd+fzC
y91ZEdIeDiri9NsHx11hVeylxUlP79t3s9BessFQp1SAild+tXaF05HmbtEDWfdQS5PhrZ8dowgG
SsQ30GRYIFgapxloTdnb5r2wYbfdyRW4+uuw1mx/sVxEL6fpH4LplRsesud4QOOUS00au45j2697
RkNhtfIRCgMIDspUA6Wfv7t8s2YuctM1bIUAtyHRgrxaVOyYCTdwmjGJOftmIcHuNnGy2jqgcV9C
vsm640Q2cs7lKj1p6m8lkZN/RUEzKImcENGGyh4vemCEJVsl2encsldiz3pAhuwqzXGVMwQn65tX
4OJ1JWWCc2oLfSvK6Jl50negNDzv0NCdZv0rDGqvdtZiuzHP7qJ1gBY1sCjbfCf0AP/O+P4HGi6y
59qWx3lSOcGF3WI8YcAQlS+WhbB0RDCBVRnUIyHwa4EQCrQoJqQfXuZmYu9Gagc3V83meplUxDzm
YQRafG50qDVZ8Q/B4nIEUZNeSAb9H7zscU7bxSTilc8gVSCG0LykeHCiVkqP2vATFdvW5BD+ez03
O83boxctM85wfvAdk+Owozss6oljChKCO6bKG6dKZYQkUTveEExZAGw+Ark7eV4Sw1+HYi9HGadR
V76xEJOn7TjGszuJrNPVze7c1vEdkYLOgQOittjfSeG97kRoLt8Y+A9HGZVU8yOAnCopjBnMAXLw
iCoa7Pm7IkIU3jfPU1aJXOTxZe1jxpqPoHiEU8j7x5/JP/KHyLqWL2j5PIT0mQmA4REPEZhXyTp/
+JbQB9h/GJbBb54JmelGxQdWgUb2sEIAjfV+Bc9MjLQVL1gUG89lbPqiZGPLZJPvCiEnODt8oBBU
EuEGJBvLQ/l5Vk3EWmyUnMUOEe9UQzMzYpztLoq0GNBTtXuKb6Qi52JN5FyBONk678w6CWYu6GT6
DOiGxCbn+AgBvdlJJINYI3HTgTeq5thT9C57Edo1ipXacuY8eJTwTCF2ho0d9ulfHKEGuWEVkmIj
BBX9ApOrKXs56BNGncNtpL3ofVVjTLEBC8rRGW2bwkDRUSzKVUt8pG7KCkxrueF51CvfxnvD4YlM
oQLHKmTm/L6X/iAX5a7xBrESojSDGocpmhYeEF3wxaRj5iHDR3XpBUKQ2z1L1HgsltF8yLHI2Q4e
OI82KROuMJt1j9Ns16YGHgnHO08TdfsP1KFjkM0zol21izhMKyiCJk5V69HGwXGCNUenPt5Tc5KP
M06i0/IOmes6xNbCUayKZn/SsZ6bu2Qb4MbKEug9rGS+4+/9OaH1vNrZ1XBbGZzfv2/AmAlxknzZ
NHtxS+nMsk5CJzlETE8NfgcOAivuLBA1qiVsLE+HX+ICwm7HFvhchQ6fn719d0AEdo+Z0UIuQK3I
4eI+DBfwWaOL8LsFWoj4YiBo1hVlWIxZHJODLC1kcfDP88E6H0+un+EJgRLikojJC6A5+G6ALmcZ
ncBcF9rGiSD4HJZ6X5EB3lFdV760oDW6HFz+aNpTGdqSbeIN5COfrtDVmDBwLAVmDPsgUW1+VM/D
3tCRbpAVfcM1K9nVc93xsqpuFurWYqsouHDLFousFwkOCbOPRqttpvus73PfKXC0HGe0q0W71Myd
8s0T8M1g1Znqmki8Arz/ybEYhs3TsqA6pgWY0qUODs6lect7z45uKMhHYCJzZDw2+Hwli94cloDJ
neNz68r/HspvGtUzfOmdoQ2BirVmklQ62rhuhoEW4YcL6TsTpILQDHySmh9Vb2axOcHs2JGkOY6K
P33c10YkqT/aUMUbW7QlPNC+pJM4kjPOEQ9IWmQt1dnlO4M2zKXJ+ufFkXl05sXrDPt1ALo1iw9e
d0jTF6epmga5ru97yni64+bHEuSPBxVHh7GhpRR443V7gT4fwP7lb2vSChIAmy0CIRGIQRyZA/wD
5ijHHD6KKJgmxA/nkVx2WUvodnfWtMscO1FIbFT192bRJA9g7qT1gkS+iuI7tTM0OJWvISaUykdy
ake4j8laltLKaOxAAAuCpwjCPmSeGoukfCcuiMiFAiq40xa+f3Q9dqph+s3g2VLQe57rQNSQwO4z
BaRZqTL1Fpqo/kuoZAuZyV9xQ4tqhE5fmnnlnOob6uFfoyqyb2X/F+WhLGqMp3a9rk0UyFkaLhcE
mXGWipH3V2lm+AYKmWZvCp4aaEnHe0tfG5g9nFg+s0OX4sefTaL7jrurJUa3LFt2z2H56e/iYZxW
CRHW8OJ0YfB5ejFyH+x3G7bjJpySCguHYvdq1zgjcIvXdFI0UxFWeqP5dDq0hZ68mXLN1lwWr4hh
l8o5Rfm7xUGrL+4z7IiNvr9iTGJSrjgLCjTm+93ZIbKkf3c4RfoIPVBfZ7xfaSU/P2K0fh0jlU21
GS+FhvYnBL01doP6dmW/HlhBoRV3v5yGURD0e3zI72ifmUcXpi0ilzam3MhsM7SRsXq1tdS4BDGy
4FBMW5ELCZvn/XyLFeAXLrGkKy6ROm5tAvsqvgAgur+T9SSoByxLkaPwSqaztHpJj4S1zTBb63kq
DsB4ZDWylgYVZzBNmH4/YEM+nzwafwgGCiOti469STSG6Gr7Dl/+e2TPjYoEEz4XvLRxzAh5KOVm
48RJpvFncNHl2Ajd4GM4CSEzd7WqoGA5+up1TSL8KJV9t1l9e95y8sIHv+uDGyE3mqLLfLm1V72t
RMStKVKEzFAgZGdZIduatDtGKJfbGRR+VaKeArZU/nlBjflvM7Orxn4BuGbfVjlIKdl2g795AxvP
EExU0M5Z3UkPsfJglP7Qg1qHr9RnXQs8Xgj7fzI9GXrH/7MvKjKS4wTFBTnv8b9pfN5Rzp1yV5W9
rOK0Lc4BoXHfhZDJGMZNbS+25vZ+IsaJ8R9YxMjq6ETLCIC9XdbqtoIpqZxghfKWgKGBtqmZK3X1
HdG1UDrtAuG70qlR9bORfKmzej3HX8yNw6ufX33Gj5heFrerRqecLj1gwGFYuZshGr38jjR3Zlq/
zRaxo9eVnRLAX53lu7a/L9Nhviwm9wh/qVDIhw92mkwmoohsycPo2TSZYRfWSCG9qrjGWm4fV5Nm
KRohV0xOjGjrxKHNdI56pOCedI5fshMeFoFZjPh/Ko3oOzmy5I+9l4dQblNMUxg8wxm0F1PnrRxE
g3Lw+FD5MCXTKJs+ZO7wTSRnjfTjojcGB0dBA/pjLfmmG52bybuTFddwM87Cifea+nOd4D2oN6Gr
Eb+LpYTShf4Lxad236dRLEcKYMEUR2bEApbuBiuAOLByn5Rx0c5oBdmjVGqweo/SsJGiZm7y17Pm
D2lU16mx4e87lJFwcCoC1bIymKqt6b/ra/hrY9xf/jj8csb1T6DAaqK/s9Ez2zyiWrytLMgPWIHt
HMQzKQTTG96b7/QYSMbouoWgsIPwgUa9bcDxRwIExOPgNwF8dVJ14pBsvcvVudb2HYj1qtgTcrF0
VF/CnAMWBmb2RSDVr8e44wI3m9tVCd7SX2YR8kBxHnRPdZdsyUoDYuNMOKaXZSPPkRbKtPCtjlVE
KGnlRwFzuVUUDIM8uLFA3NtaYbg0TshM7kDipB2Mtgw3xlAKwWsFsArhbRtm8o2ECVfotwpt9hho
OOk9AjxkR7SU2cjMNLCFtDx/qoOw6lLQGbOpqHLHPmPP8P6HM+T9NjrZWns9OWlUgnnfMJK/HcUe
f5CqTuKcwoMNI+KG5M3auoQCk/rHyl/hbN/Q/IjsxpBoJI+XczuzKb66qRugN78tg5WN6F/Kkmx2
nDkwZU6zwWFGCORR1TBPk2yNA3+eecPPsyNh6xda2qL0U2gTNanV1lOgxCYFbNrt3iAMBB/QUooC
jQTXg1LA0DsC/NRz8DV1PfVRGjTAkJd4IxLS8HrD/abaVHJlFz4jA0ZYZJ94OwbO/rmXfQN3r47Y
/Ydt2A2DWsBlnme7mRn68x+5h1n7Fc1upURte4161NR+JJsNvW0RBHdRRLmibuKcYtA2W6/Fa0U1
NP2w+5Cc+vjVKocqHf2vdOVUe6wExLTxKMfDetFjCbV9cx08CgnQLb1dSdkoiWJenuuHYtLO3TmO
eMg2Xvnu4rzPp/dUiOtGvi7BQ1ndkzgsCvabtFggEpQdK1ytrjWqLf8c8du0X/COgHBUbPqIpVct
SP2UXGaH4ARdq67fsFP6YdwtjuDTI2Wo7ydV3SCh46quzURjPJwSwoczKBimwZdfq6IKjQ9w1SID
PSTwZmPKJRBVpIR3NB/PBHLmvrlG8PXsS9jUt85+m7oTv9TvBPtq8CYATC+xFM3uaF3knsu7Lzjt
0A0XRTL9EkJGscpwVN2Qlwywn/r7+nOpg1cLnVdZFQTKAVIHIB6o7TNN0qibrNqVLOWA7vosX8nK
4ObXuyX+3Tv0mup5+twi0xl7wKfVl8o8KHyaSolroMtEaHfqXdRA9EEdH2TLN/0U+ynhjee+xmEt
AhByZzuc+NoCJ8ma+MmEkAbMMlhEYwoL+qtWHIatZQsdoQmuljxShwLxw4A0CkMsLnk3Wzfnnbti
2oLOv9UNrcEJjdbPlIJmyaTmVBrdE8KpG2yYpPP5/ScuIt4rH8QFVN/zFQqu70bIhVYjLogsOOqT
wKYaHMb+Gpgrw/stT3EzvOjTorznDaFubFFv5a5iYp8S61ReSSAWcDytHDoaJAgjGN+xDn8JT9e5
fmNUiYzZtGDVnjfRSUQ44WGuPx3qivEcgZEFcYSvPnuTjrG1oCoy+dKiUqjuRY5giZPFnLpajLXx
mnPwEL1QEFl/520xRBwdr1iM+cO+R61r2fRkb3I/4Ah82PlKZBs72tLuIO6vpX4bvPeuB8GSwOam
zXDyToC8TXFE3o6yfHKQnYDfX7VVKj2aJqhSjUltAhilQD8+zcRkT95pzn7oN1Ei9jse2/bBIe5W
4gtCwh3ggJcMtKJidQuW1An2DLtV8/Bmg6W5fKe0IwydgDorWPVnX15ltNURI2nfRlBUMMV4JCC4
pplvbiaLdhyyLg5furUbLhLEzbalmCB0zzjGePLKsj0vxM3bZrDFx6XOFZDgv3ztxmtqZrDmu3oT
vJvRz4/PaaUwhzjiBdZnPbn1smoQTIM/inYNIIP4zwT6953XL9rgV+XmJ+VunZ/cLqPAbK2I/eOb
tFh5U7AJ9sye3hx7zzKkos8N3X9z1Uo+sdNM8kuuQ0mlGP+DWrirBM3Z7y7TK/B7BMKJVq/uYsPq
czX9f2YDvMmIoqmqsUztUTcbG4CkLHip/ERTmFbcqAKkKULsslSQZ81HdUZRfTZ4WtDROCv6l805
DslyBnP59K1mTqdXse9BX3X/RNEMG8Y6s/mFk6e+yJNtvq3szbjd7oVEhCRgthDeglfJlSFm3BsE
dD4wrOt6KDS17AysqVSqAcRtyDLz4A6oZVHRd9qdEeSqMKZrOy7dalJCD80oPGKVqP5qJ1P0y1Wl
NGaMaJ/nWnlrOKfXKAFhIHv9s7n7kzPnZWEdoiaTNX7Eyqr3tJE37N1k43YxvL3kU/3r6wDEDhbm
laqL6oYlsCXuVTndHYYusJHqU8Oh4PETRhDGVAZAPZTZ4V+BuOLr3cHSKprpw98nFsQ5Qa64tDFy
gDhNvGGeHNxT2ZULd6CCWKo+TQRqMS8IZ1qFPOrL4EP7cKmVtVSNbeTKQyfMIKG+LdPgAW+XOv5Q
vmigkSWx0CBmgRZ177p/jSQ6B9CIyxjwczVibKw6+DOBYV4L6ebjctyZQO5P2fLFegFuLLrsHk7b
pI2SbXHzbfhzr+oC4L02XBVoR8omGZIMQOF5XWyKff8WbNlyWQ4oNhSBcTlkxtQcE/yNIJvt4Hei
eoPOi1idyPtGHVfy8v1JVoNqN9H9KxeQ+erdYyfjDP65BCC0fONbhAu837YgzacKd8LG8rMbPvho
ghMjUTT78H8409FejZYMD6lQsn+rryx1db3y2Hx8vZ74AFmZnoNLK1o1FO+apKniue9knHUM+e8p
7FPL3s5SQtvB4x7l6kHvSGsE3LZPuLahwufDEG5N+n+xLy/LZAY0skLAiqazY0UkTT9N7WFruRZ5
JDB0g010LjCBeT/Xpn9S386A8n06J0XmlIHb6E1b/Xe0s3NPIDq83MH+Vhc/HDqFkZKwEUybwxtz
lTL34hihmQR/oTU7V8ARaN/bqRgel808w0wsjihLeUICQ8wqNsE5j35Ic6i5eDt7QoX5btvnOi67
En1mWQwsAEY6dIn0xO+iVvilEck1VHfhvsEVe/2Li8LY9YZgfbhSaE+KEFphCIlM1p12H96Glydx
BwcU8s3BtFHRLeZors0lvmzF4bRisv7iyyz3HVOdTAw7tQVV6q0EVEERlTZa7NfMx5QPx5wnTrBM
Ra/SV7HOLExD7piP++9akrJCBBhhikq17IadXOM4Xgy98vpxNfFGrFag7EB8fpNTx8J7aLU3eZlD
8CTMY6c5K9oeAJ0unRf9HlZO8x8LL4NbGxMM+yYRCJR5/bfnN7rLWAFd1kG4Od211SZIPwzcwdwc
AJt9d2hsvRz1W2SbPFp01+xCUx0IB1yVEHqD1HYCqMr0iO6Sl/9hWtqb7nffSQyMZNwaUywIgEcF
WQxVzJQrzZKTP3qK534Ho2IxtTILWwLZTLF8NspDCMxbPIBM50OVjis2pFKCyS6v+4ROIIJLPxlo
uN1M05V1q40oGl3it0gNa8mtWDwqcRpd7jQlmltiQUbGA4RMYF/REhwDQD5g8up5qDmOBwByFOWN
XPDDp0zENxn/AMfyNY53gHFzvzsMF3YNlRP5BpJwDtcID0WqcnHC6s6niEmD7hKqBZjpkyCNss7X
GqeL6BXpvnc2fW+S2Y/yUivkJiCWIU1WkKSuSHH/8yRRwZdjkz7j57RkneuGBSrp29/j/hHYx/QA
JzrLrp8p4kB1JdI6khxyVvigunOpJzcY9cTSIRJj6rfycmv245zHAoa1/oQjZB4W7AHgqFFvJ3q1
Lzla4Dab4f/AiBWPoG5z+8DfO9d30rEHlX7b1ZJvoj1r7/BWdSkQuV+SRpHSevi6o5m8g3AvEPUC
XQdbYSfwMfQ0TmAlf1wCJnpYkYSc+fmzmVEw65MbIBn7zuFvb8ABqmh2yJ3R5vgnDvVEdNZfRXY1
t9EXHJaRNvPMmnSBMaS+fkkNPUsEDImiWHg4s8nrgz7Toj6VfCBgc9LDAL/X9ZtCnphG6vSvX4//
hvtogIkVpw+I0n7svh/bePgzH061ARTfbf7tbaGqZb3qu4Apa8URrOTVycV8dQa4qkg0VWioWO1q
roSeH2q4qV2hCRSlDPKPnV3BvrRcSaYo8xh0IKNOl9Wej+w0Mn3qJrR+ZkuPg0+sUb1U6svy4Bsk
P+do1A/T2MiK6qR0BRhj1c2GKGM3e2TgcgVYvK5sSWm4b/+eIThVRx+2MfrPjM3x63EypQlxMp+x
cL+J7Yps5+pjmHNOKktXK+K3e2aOBLtK7AybbUj4GPL77oqsvCjPACj+xXVHnBebTdOXWA1SCGa0
PEykFm7AeGIH2757vtiBoX5v/plc/QPt1YBtYypuL6upIS7n+ZdJ3cRhVepzD6bUzI5vUTKt9WUV
RAKf40mhWK2k46E8bus/5oHAAUCMHIYfMORtb1WdkgEPgHVjmr2Z42C8dYl8X+YZ19s9PN0e8Bas
otXhmb+1+Y0FANPT1ht9DXSjTe5raLQoniBk/HkOoHgysZBskXrkZ4KjJMNwuQiLmaxel10hmU0y
DnYJe26vXYPuGU3riSYvJat5j/1bpaOpFrl8PqLTNn3Kt+20aab+CgUuNm2KqWqm2dDOSjF7Blpf
H6Gd59Ln00iei+8UWKGe0S7fGVaxW1LJdjodrSkuL24PyDpVL8ZtJTL93oobRb+4PkIgUQr/g+XR
m2wKs/XL4an8FahNe49PZnLefpJHkttQ+35X8LwYVq+VxsM7s6O803QGQCnnRY6+who8W3wlNfQy
HqofKagxUCVwqJbwjNvmo/aAVj448+cHy3hojhoQgif6Nln0nxX8gR0iwZnK5C2YYYmB9f+vg5dY
dEEUrNhXh/8eF06Em3IZLTH+fOIlAQni6c3ahOIvPwHdV5x35vkuvVJD71qG6TwebQI3tJBA7oXA
XuRYkC+UgQY/3483/vkIgBZ5gPVrYByZuaP3cwoHvob0D+T5ylp2+obtcoS9X0ogcdvwV5QdgnS1
TqxsBEaTnwxw8otL1q8fQPIp+6Z2uNoadgs9UsZysByG9JvyGq8jGalhjbEi5E8r5+XUXs+Esg39
AKsJrFIS+r6VWifo6m9dv5XsgFK1ERQaYTwFBylLryJIviuslAg2iaJ5PX/i9ZPh9idKEbKaVKJU
nFR/qjOCu0M8q0KlKgx73QtaelPZAv20gdLQNmd+9P7cTzajefLbbi+2RtXihH2wCo7kXMtA3OYf
hgDflbS2bnOR2zkN7CVGLEGsTL0jt80nhoLAkviYrHW6nlxAusGpBq9gRbU2kXqiAsd2PD9JgtZY
Pd/XnqO19JDvGduD07Q5ayp12VPNBQfWkh8BMvOsWoKNoxmSGRP+a1atJcBOEaPIcG9Tj/QTUiVe
i1wadFjaMRXkmznN3oH9V6hYhx7smg4mjLbinugBwSaymRBN9Y8CCnUQc/xtmY0hLnkIYuYoRdjC
Uuqono6UWTFi+y4sgcbuQheL6AVFXUB1C89J8afUWPwg+3JIZ8UJu5KEP6cAlz7ZBVpLTxr5oZaf
ivb4iGupmNtqseJhqHH4LAjWvTU3tWbiUE66e7bhQn2w2wNN9c1osnt5K+CvC9pHgis/QyuKZkD3
qOrs1gF2j2emXkUsS/AkBcdkKzw6TxFLnXcm8g7gEwZNpFux1cu9xuT2qKrv3eC+SV/v10Z9X8e0
VfIqoETuS/wXlEBFHksla4Ti2Mm6CRB1by02Nsp6tz0Z66GdNw4GNmdaF4mHkdTU4skF1FAOMg5V
XLmswu3KUHBvWkWdJgYskYLl3O3kRpVXM06lRO+jUbIsNr618OyMqmY3/qOEjMkCWYnVaH7yddhZ
tOl6v0Q5lypiyVybkwy7GeD6fdd0aqzu+KraIafn5aBQFmON8c+6k50eOjp+PSmI/BgzZId/A4OW
VwrS198zPgLLeNWEw49C7iDEH21KWG9xAilrQRuf6Jv2/BZwsEdoHu3SNg7i7rMhhKhVMrlS0/VM
BtEh7lH3VxAzom2ChBn5qFZzM4vdfxyQbGfmgbEGPSoUZ//7CpRoHosaaktj1hvsju+B0RTh1/zF
WAcAVTdHX4F+ooKaNijgxxmTZawtvVyzbDuDyls+5FVSIGa3l5VuNMwetCR6ptfndfg+hVc17J6M
P5GU1Yux6D9b87aFZVW2FfRlymvqEK5yef4pnOV7KyEDxtxfAmilyjKLjk/1fcGerN7XV24hoBk+
A/R0jXFfBII4sw8pygHXKbD8VV3oaK0GoEs1GswK6yRstzrZy/ZtDX2n/bnOMxYVgx35X39OWFgF
NTRgM5P/VRbty55ingNg/qp4KLE2lBqQ5gO2YXS+SYPs+0SlePM1neh4R1BtQCMcVY79CzHM6hnq
SuWivCSO8eUhmLP8cQ8uA2KnFkO6B2zZroCJuYXd2i9Z2egSXD/UNgG+kpwTt9GPWDbXUgSImJGV
ZmUp5ReN65Hu+oLCXgScjYkT5rI8Y5g5aLpdTOO3+r3G/UJ1d4SSJZ0Q19qp1EG1slIuqQhCn4jz
l6r3QrUp9nezgftn4hUcpE5PTrqYPmkWzJQtYvyS/uQa6+6sgpHjSzE58cw7DwhujXFErxFCC4pk
gWWjjJ+w40RkEFr9W8+ZCxRNWIJTrTV2KQ1qVFf7OK4EczgfgxPC/v799GftowEanuyHaVb6eKrx
1keiVnhu/H89jXRhwqm84VIPzECjxyeDcXTeyP0EMfY72EuE7MoJJdLW5leA4+Kh2HeVJNLOQeV1
PZmh1cjfgVoXtg+yA1BLUgkUbdhbDutgZk/OazrW/yzy8j6sqPGZ2pWsO2C48jnPizwbOZmBMTK0
rKQThb2VRnPCrS0pu841NurNDjTT+mFCA54P1pvIgVK43+stvsDGymKSGdlGRDTDEO/4VuXDOw26
TU3PH0TT6N71TcHaVZbxgX9Cy2mqaRjAshbY4BDS8CvgABBkKiwsnYXMRwjPQcmJk8RhRySN51/V
9/ErfFKS+JY11QfgjiIRWRDxXCU4gkzqYJA5gLK+KgDi37mjCu1k9Ye9c50JinIAWUlKyaTlx7+0
tYsCwdthX5FnJcEgWOj6jkUG0R4FniMUkFVdAYqvoJzhS5sQdTpCefXOmYWh8hlBdsiGFikO/SFI
QGmxj7lc7Q+vNJbvtjUBrR+i3EbbBARtNxP2ymgjO8aJI3p21m+7SRe7osnHJYsr4xv5Jw5bgzKf
aNdFSf6Km5mpg7Spx3CEV7A8MFCvm/wDdGtSucuxve+ppTvZ/B6xgI+HTv57YAQW0Ji64/n/c5nR
6B/MBskLYIY8B9Uo16Oi4VXvhku6brTKFb2fvLvwufgRHTg5A+iX2NA07knqGaTQN3n0tTOCdIcq
6m7G23rTJbggnwjbvLtDJXpeQFEf50EJrTMCJdBIDcX5Cb6m2qBb7Ghsk2+8NMlrrruFd8/Vw0Hd
colP5VL3rF+Tjdp+RRkJveAhyhmPrXZwu68C43xf+mY12JR3SohjCv2cEWIJ8KzhUL+FfgE+QdnO
PmimeguABcOIxXb/xlhp1kko7XUOvYR7TKMwJdXtr8EzcwDMla/Bj4BsQzkT7nAcY5unWKqAM2X9
bfCV+B31y2N1YNUFScVtAhgq0XLvuHPUno0V1M4NYzbyh3uIZ00CNmNhADx/geW5xWSmIRDpy1ta
dMstf+gObN1jPa2ewszXuai+H3aW7C4aHqaY/0t1zVSe0wF9Y+Mu8+GH0aIn8JABb19ta7i17C/8
PFDa0+ISEaQeQUO/FogFymEM39usV8GYrJX2Bhspy9UkTUc6q89hXigBPEy102pt3IhJhYHNGJup
sMUl8/t/9WFhRxUMt1fHH+A9b3xqJvgKPBOHQ5ja9QiwhEnX27E7yfF5QbUuiRIHwPB99iRAXu3N
RplbTaRrCwlNHY/Rs5qgCilwHLm1GqFTpzMNFrgHfTFiNVMGtR1DPJJeiCFKtL7IVXB5UgH2eM99
oREXJrzdTdygdKsNYPMC8J5YkT/xD8O7AUITQJLCyjyIPcwuZOVkfO3rn1PvtviJNpKKtt1Y58b2
SGhHViywX6cz3Mf4Qgym6H0HqvldLJYWDPYJiskQzWEuslO6Z3hjhjF74CjySjPOnIiFYqnSNwZv
ZrNUdr0XX4eeaW0dAcihO89VWRCnExVJx5FQdRkLi0ZHr9NWho4YjByRFEH4jhK0qn2VQe6KGqwG
WFZpS2fHfoMks2V6JfNn1GWgCYB+EZrywLrrmHK5/tqrbvFa7qNIyKMJnSxpSFlwx1bsAh73sA1x
hIlKdBtesFgmCNq1lpYQTtAcqJyI6dCDusmZGcxl9y4MCo+NcSn0jS2b/OSjkCa//ZyjT20Ijsg5
5q74tYyrK9PV17ot2sPsc1Qzwz7ZADgrkzuTWtBRFEDWIAp+k1Ijmh3bnxeFC/PSSafmISqWf1m/
Z9AaqToNjAgf719owJmM5ZLUeiKkF27F9Jr0PRMV/Fla7Ktr+H14DTRqYpH/t6Yg+t7fbG2tCT5t
tBeyHUhnmFnEGi3W9eaky/N3M28bZA23PBAk/klp+qjHoNsSiUyvwr+DeqBUH1gNxgckPQgX4+Lf
iSgZeIDJMHh0fCC8c6wNOAATUBuCe92iXbbw4gr5D+gi694Z8HmgZFW7zfeDUfSZkcwlwTvnAupH
LClTQeH1QrCDDf2Kb/TQQT1aB92k1DddvBeEQo74HeRgIU5Q3obGSSEwJgNHRF9BD5fYXvgkbPvF
ivSz7qmi8d61DiJQFqBMMUA4qZohZCt23aDKgFK1hihZy9H5ZKYm71TCjDeAblXZ3+Kf9O/sA8AY
2YiwIUtMXRwGZgUdWGlVHKARV5BUtZ9dYwf/akbYQSgrbPUnikOHZ4qnBEBfVzSz29gtVIgGSXFP
c/mZ1nSVxkHyoyZGxS59yp0t0t7ttPeeCg58x5pEt2sqIhhq48Wc2tdQYoR1P5KJdmWExMr/H79M
LPCQLy1xvl6ZUQQXrVNEE314CRxM5Sg5xLg+jIP/2HhzquO1wQ9WyQG+nCJzMZ7dKJqQyhADlUA2
F5lbqT4mTxWcyGUsSH561XbpbXZzgK/FiebMZcB2GXaZL6D5kEnReEofHkCiNz6svLFgV5chy14y
VyRtpXcwBoAk8YQfvqmVoWyQiSVzDXOJLJYW6ww/an1nzfS3t0FuXY0N+EiKllw6XJgUix0II4ea
1CUlQmBkMDQYjym35g3REhJqTJSmTRj2FpydM5rUwNXKr73Chh5iqnv+mR759ToBUatSkMXHL3rK
BNjYbcef1R2Wy4OaaqonD0iE58pvS/2Q9P0dnbFpcDjw/APJmm5NySPhO4YKsBOMHAtMrESbwxfy
jNAS7f6gWqmARoqPutw8g6Bo8ZDfnJ/kQQuZtYfkDSPl25MOEVjpdLBwndNP2beF6Cd9s0mgGhT+
7Q6v775Lq403xaeu85HtMHOBC6UuZG0my1SuAonckpBByVOYFZx5tSCqVIPAzDErkPhsen87AFad
fUjnlCEXurfdRxpy0H5Xgke2ju0J/9itGd69aNJWdo0f9KyfJvhtbrP5F20+/wIsjL3oa68gQAnV
lUa8rH1TEGyCkvGyTJqMhHEhzvuImtX7nWwe3EZNkwEAXQ+6jz18snLNzSkLrnmfJYCKaK/QdKSA
8RBb7AfPLV+zDVG7oviJ5CS4FHdaBcwItNKow/TOKG06r3Yv/Ch9J7rcKsrJMj7stLVo9SsXkdtE
wMuMOaL//QHktRsNo5t6lE62IW0Q6B3qyZjY6gTqiQk3Gfx8n2TnGlYbpgM6xJFBk5MoaZrkvGAZ
OPNObKfEiRbYyRZOcmTaf/jUVorkVD9Ux3LCpvEi1yo8MUEmOB6LtqSjXd0U9wo1grsWupiJGMcu
+eSxxM0DYDqTrEBVV+1y1Uu/kZYwgJNxj4Hz7VInX2+iVCKtVtao2druIsOyzuptjFcUSAdEKgFd
P5WULVEORHlmWbNObUprU5+REC6EaQbDbwm9aLGjbyszqDiNQUST7XKcz90OOxWcmMVYCtBdkOYg
kP/aHot5nieJTnOyeDPiwXdIVFZ45MswRuICUqWP9zVo3JTLMGokuEBjskR21PFI+PqeYuLL3IjU
v2lsw3UCDhbp6oMU0cPYLI681ceNWcdpOWLDATHmZQNhSBrjfITzVMwdDFfEUiKMmiurjFyDWpVR
SDpAsbPLk37aeaIv2OJFhhUkxbpyYeqlD+UFRINNoq6HkX7rxJ+xomLUmXHF2NJsMo6PbBtiFYEP
nTN4ul08S1iU4RKQNUFpOgeYFvcp4uYHmDjEpSGjA5Q1Av7Lo29K7mAsD2jrW4ziJ0dsbCkR0Bhx
UHFlFKca5bhEFgNTy5FSY4ip3SjrvUZ3DBCtpgMxDUc0FRxZEksy1grAwvcayNpCdWbnyqG7/Sax
naR4ZVscOw3nw8PMUqwAOst2IWphhQBYc1oCYUWuippsB6oM/8v/32URJ26PjAjrTmbaBs+NNAUS
4oCF+IhIrQ4wQcY56F8AtuWxWjedrs8oZMCddugH1g0KiZaRtbXHdsKgIeD6iP896QFGa8kSDZdp
CUXWcQV78Cr/u+BDjcmxJyDSCVd+etBRFnXkG/Y1xkeDTNTERm2xr61JAWYCk4ySITuEQ+NvzOoP
kriIDaklwtZUI5+ZW0CsQxy9KHlLHOH1qkDtJ1IOLab0awYIbuzEVzywRwGcjQvKcG8GglNAdtyu
Z9SX1mwvW1+AACHk7/I2u4FGbgYIPidOc16Ev7wZ+YbGWKziUaYP0evzIHmuybsiG5KzxjiXV9i5
ktahYvWxtuHqmuqgFkoNteff3b392JiMt880Y0lK7pvzRqC7uzDWWRbMQ1wgQDeo9Uo0KjnssxFh
feSHEA6E16vuzRwDb5Nw8qd1n+ZZ5srmjT0+nyZbzJVVrksnMXg9nzn8EP6W8jEStU1zQ+wodMTi
K+8TAuLNAl2RBUbS5wn4VFE1Qzg5RBjLItOqxWdQrR5u3zr3Nlj7wNpIwwv1FlNpaK10hvDwXtrb
+nTFfe4T/7LTCYg26cTJ5GSN0KF343j2HcNJ4eHZYb5kxOJ6APtsUp/oFjv0Pf6HK9ld2j4Z2zXo
W9wDiyGJ/BDuUTBbNRvoY0O3GlRui7B348IPmnyC3b8dih4dyWwkplGPIrwk6dRxWhGetLS2BLo1
G0njiwUclYDOudJnAyQqJMxLtYHeNqPZ5BNRsoW/jWnal6F9im5ASq9JkRipJNvGoDR7z5fKL4u9
j/hSH2nkpA21brpOuff6mp/V0l7ZYFpoJLpJWKW2powHJeVUXVL61PheqXJ8l0wVGiRylvTvouaD
FS/lzA/vLB0XlOaSceqBSsFX12kxPLT7wVZxjHLLpNJQ2GmaQnjt+Bzd0Iv43q13liF6vWRHR4bc
ZK8W1mbCR2kUQmumu6NpsCDfQL3CU17Z9++bS05vkew1W3lWtKco4VX0608hKH+mTI0fMssZu8Hp
x2xjRDkoSZxP3mnFOoVAP+ocKrvxkDu9pIB1cT5iRl/cUxu7QTNhhyJr7s/OPEOoHHbC+68FaxRe
SR1YLlFx7ULK5TOCpybC5XnPz/JmJ5ub2hDcuGJDSE2NWmxuu3tUfFYNpv55M0W6JaCeG/LtgPsM
HTChVeTbMaQVTrueY6PaCVneCgkMXf3PYcu3MrxYvnpvrs2AwPJPNLP64d06KxVNwgVABhoV45gP
g44uXP1EHzOk+T8mbfJ3HhcjIYR/Mzo/pM4I0UvIx+60RzUHuEyE9gyzkUhaROWtzskXOiV6yMuH
ztxYffwSThJ5wVZKrg2xj4+MKigqUf0NstvGurpQXuTc8BG1e2aC2CY7awC6leOAI+VKlQ3SF8lu
nbxfSVIl4V5uEXRNX51RDQo1ydId9lbQg7rbB2UxyX3dxewsKqj8CqlfEWU0sidfdpQSoj93gY7f
W7KxgnpbXSc50YvwA4BXH8sDYsJFTDGR1tRmpQb8U3THzj3y1b2G2+HXNVXT8SCi37zGx+x3s5dm
jHdjfiBfajgDR7YXO6XMfs7o8+UlbPPbHMYKF9S26rW71xeHqLygjNuBQdMUdRmoP/p7umotCRB2
D5GjRWmchjoHyXkLB5Kz9hF01t5FUfmD+rOKuEbOKzItnyXZtBAeqdiwkwQmpDUHpHUQWhxfj08o
wrKB1TjQSIywVUW+/emVICzCsH66jdMjmm58rwmmMO0rgzKKMcMxslULiMtIaJWMouTvRe064pxw
FN66bw3Wm/fdR8szBdH8ajoQsWWoZwnw2UDS5RoF+tI+vCbBfRxLT/rF/aQpnyhc1etARNwhDN10
K2T7/m558+DZinA82TrZUGpcNLE1Y9T/Z8C8zwP8uOJPEpsy+wpwSQWaOL5yvFLBZkjjr4ZAMBL1
vfbPyU1dgCQQMnjqmzG+daA9/dv7LD/osTfDs1ayY9er5/aQulA8aA3ht4R6/ESH5hIcPxfZw4eA
fWqf0igL5Y7uh9OXEzuVeG83APT7OWHCf2S82TmfSlN7Tvn6mznMLKBL50HKggASSiMR+ZuiqLz3
ttCixCEwNTHICKxVx8uZHtc/+NTA5BRrzJUUY1LNPiVVeK0pTIgdoLxMxDLUDYT77w5D62HrsY36
lCu+Xo8Vjjr+/clLOPUmojBRnjmT5zf6TP2DkLbQtU1Tles2uBN9MlE5lAME8Ky2tvuVIQJc2UD5
j8vADVY2X6J8dWHBMw7sHWpoWxkPhFpTk74ekMT2k8rtLiSGVfqG2X+W0jS1QX/gZftrEqTzH4Tc
XDRHe8qQ1sABRgrmFVj3K2j4+pk0Ul6IoS/5Y13I2Hjr3y9wxMp8BquMgJnSS44MjGjqHIOxBJyR
IXl4CDL+cz8ZmqsYrNk4GQwqBmbiS+4Wb1vYkKCdaLXPeDUDhz88aZGIWJ30gI8UJur1dv8eRyyV
qz98uaGHMW8GfmTsPmU9r2JAmxo3MbxtLBRszE99c4IRHQOIHan3nZXLn+3e1OQWD358aBgLMFMj
EA2Mx340eegHT7F59d2V3dx1LFK6oVh2qn2Qsnzmn5eidee1LfYNKXcmuZFOg8zGR9PPv34vLl++
aGRJDkcVGljtgaLXLtyREpwip+wEqGEgKbZhJn9a6OwgW04aPhc7iPAswsQ37nZbt6clmPRReSWb
LteX8H+mo/S7Sit7G1gu1wo4NFT404ccXzHlfgnRXzojv0nDo1Y2xVrYxGFvbwUSmXRpJZo2B+NH
sSwscEsUvr2aD/s/RRqfcNgQh1z3Qu8k2oThF9KGQLaZNkV7icuL80B4Di8u0NZRL0vbL4EIJzMO
+WAbgPa6+pvrLcOA/gXLNhYImb9eEGDWftgvwWUpBqgFizt32zP/7xdAMGMji+so6lr8U8Nu6DGb
exQ2ST3xYdAtwEWfNMikidkOGfOVz4JHtY8KYk5lIFDQAKmoeCd5TFLIh3zBpUYKgWahF4AP/UF+
Yxf3hDIp7dUi961Id0IXdWrq/lY9DuCBEcJWNPmQXllrlo9Tl6RpwfMNDQczE7ZU+FerB/f3QkfU
AEvtOoPi8HJDeHckOys8NHiMfy3afVX+9v1ItxB3DhVal4Ocvz5y/h0vfx/w1UYMyahxWbg+O6Mj
QNuaNknlmqG/H4tJDqV3vUtfpb5YkIJIaCG5l0BSy0Kp7shsGtbzB6TQxZJ4VcJQlEp3xxMO3+s3
+2PzebH6VePwJuRisfi2Q9OLaairIY3LSFN0G7JtT0GCtd0XcVpB4ADywBsw+rSfb/UaNCqC3/qS
H2PqoEO+KOs8bDuCpoa6DNp22eXWkvPruDMzq+6AOgN6/8JXeMaof4Ab6fe93/EYdeyiAkpgeG4x
RqVJq+fjJnC/2T7iKL7LYmsoBR47gJSD3Gaog31HWC7PxRZ3gZsds/EywQI6n7jbVT7gclJSYJSr
wc+2fW8s3uNmchL/ZI87qxIUIywNXwrAOWMRSrK3+EHpiGs6MlhfLSPWIiCpp9F1+7w4CklRXOCY
x+yYRpWDiuA+c5nTP3QE0UY4yrWXsE2UR/1O+GfK2nceYk7TlCGl1qfxdw60S6k/8c4nq88a01Ok
p+ZD4zEfmR8zQk1mgQH1qySubAbVgvawOJP6BsGV+/SkTEpWInPnXk7+oluZv7FQ6kx48OzrbpLn
sF5e0r7A6XiI2/SSbAxp3b8JhjTwZ1S0AQXnhwLSvdneCOTtsy6Gz42ROUkHzeVq2KPXRjiPimWw
2xnEdOTrQO/ntzVvCzji7aQVAKebqnSmYytPufBViWkfBeS9EX+Eq0Lqz/15HjRlwXFxRYlTpoW2
t0gNYUsZCo+lbduRBL6Ezqrt4hME3KMmNhs5qYC/pUGDDHDBUmqH5kLcieKbWP0/370VvCraKLDx
SPE/cfuO2ZtZTWMwPJUhk5vbT0RD9VDCfisVbuIJkVt7p5LBBGVWugK0bQG1ZC58gkjh83PPoY1B
Uikcjp7DCuzupETUg1fRSuBMQX+VxE1Z4jv9hDbUJacfkjy2o3a+xZLnntJKktWfUchMbnjGrowG
YssdD7vNkWOFYkT8Xkdpqmr/E/5z4YNvpXIgBbEYDzUy10IQ1HSpsbUoKYVQc+Z4/l+uthgCcAW1
YPLIgwTNa99eNgh6P1QTHqx8u69eRzd9GRZp+lOou1lssZJKzZl1zugibjKxQNHYVl/WsAyZNTBq
zK3ilYYxn7Ydqz3Jnbgt/Etekj1m45u3rJ113msKIT8BgY+sNS9eicz6Qtn3tzsI7dpdZ32HLmfu
neUOeW7NXlRl5Qkn2AcrScV7FW86SVQzdOe7VXUPWxd0I/SqGrePuROy3OP5MiE0FY1jnaYlgQ+Z
xwkfCrtjHMpjyyy2v4SyHl+ZqJ8+tc0Q9Ju7g0aIZ9LN9GbM50+KQhodcnVOjqgxbuTkHPP5X/1w
4OcLysWBKn3bOKfK5DOfAiMvJ9APoNCnTnneTNhbU9nfJu0tOcH/TOVBSn9Jqr7RL+IhhEYvaSFo
8XhZ44ACKJmpBlnjomrg5mS84dclBWbIn7DZgz/CAZDwLt478dcLFBYWiX2HPalzt680nv6CoCgV
iVM5oh39EtCpzFlgryjSd7oM4uO9p6/mJY6D86jvQPYLrFShfszIlhHrzNH1Qhz85AEXrIcoOmlR
D6PpyCji3HIacfO3AjEAnhf17jM1sALR5fPtucQyeVRq6URIvZNZFSBec/4NUHwNBSUxBDooes56
C2Fqy2dD8QqqRoY16gwp1gUXQ5/LLNUAPQe2qLBU/CQZcIDt+B0VsUX6a//xSdwQ0l+uTsSx+JD0
twPnXJdZEeq2e0AWDcLtO2CALMyazAXvz0gc7Etcwr40nPYeA0bndT8AZ5tp00oA+zVg2wUHjKXH
Dwk0Q4YjYygpPJE6+/EAhkD3ikuFBuIfyxo4iKnQzuF9uuZulC9tMKcd6ie8j1rnkXgRQiq+cfJT
cdCpzYGSRnpIxNnnuAymGZ7GedwnR1pWp1Y8iqgMq91KoSSKS3dXfHmClF2x28u7aH+MIYGYtRhn
v2nc3nVrfl5l1X/iwVtNIutK7NBrPL6BGQEVVSiFsOoA1Eo5xyIzTQFtepUtDQl9ZWKAexCqSZQk
ROrPJMUOM9bLPNfPVfwFT0rJ2H8T0Qp1UvL/dQsw7e7EJomkY7Qn5NIaC5V2csT7Ggwb+Sx+j2Z9
dcunEQrpSV5Yj4KVPwNcMBJ4mWDfBihzxBLRoN8m1mNdN8sCVc74vEdOP5fuTQLaut4OTOl3531f
Njq+4LoeRJ9H/oWTmPtzlNN6RF2Wkvj7VsfbqLTIdFQuCq/Mz3La9Y9RymqBI7UGULlyrUOqrOzf
aBphwajEA44URW9w+xC8mqkFblJk1soyPQAr3D0QRnryGnlO+MrihCfR++s1rlwv2z0v8vb5D41F
ixJYB2rV3dxACqjxg67kIpl4j0pyqA052viL8i/4+5APaYL4mWipPJMH3wZCAMhZmeB2dHv7bGJ7
TScaw0+Z4W3c2VS22M/S907xeL2M5qyxo4+TyQU/cKs2gfz57CmN8nOSEj4n9IpyLFyEFF/RkSWz
GCY9mQ6OCCVrlBIS5/2ML7R+DtpRqHutsdavKzMBScVSBnkW0D3laD5txvwJwNShq9Cc+oH/1c6E
TAlp8wYoYtZj6fAWjAcIFPoAEH0yA6pMVm4qitFl7KB662+9nVOJDcKMgDgO9kwopFPFXcBJIBnz
pjatA1nI+6Ae0mAEc2HfVsvG2CjgEbPLgL5h9h3dylPUEc0Iy5SLuHWnyAuMyMk5GVnd88HRx0sH
jbVFMCqKQUwXcOEjm3cH770vOD3FyJ+gfQQEfx7VIZt+CxIGcq7t5Ulqd/NvZEvDwruw0sRuS4H8
HzopuX74XzBJ4O4yPFSLR7wfxU/INDvVLtsVnZiJhLA4objJmGm4u0TFzYUVHKoYYh57abggjx+d
XcHn3kuMnLYYqVPX3EsDcDzslJVTvGCCRp/nszkx9EJjwqeKo6QSJngZT+zNSp8g8PQ37QeUmsq9
JFOqlb4UvSXt1F3cGGB4H+pFPFGsOvbEmbTWO1rdK04oK42Lcp5+ibXEYZxL4kVsMtEAqOQI7wQk
IOFBi/u/wOWTZCppKgI3z3V3zP3a4MspqO12JKBBMdh9kwiXNU/YC1EAkfkNZMAvZLa4WI/G82+N
F4OASXQt0/hQ6BWwtUCrJ5S9P8/oVkB0x/D3edbPICVgRCX+FG9TP8Lh85McS8TTTagtfkzSEBiL
yjlOe1/au0BF8oIiXhochNKJoB3ciKdDa4coFnMGiLHR+wPpBzO2CjB3+VOAPc9R0Ob8UntXwcw/
kfQTez3tpa7AayR1pYvznPYfE7lSotCJ1bcnesbOBEgjWvGHWkCx/VmYHbj2bSqcZn6Sk504Uox6
9vfZlTa8nw1UBn9trnEiOXbbsLLBfOjoaxbPpVmgzKdLZ9E+Ct/IUGCNpOBy/c6Yq20Qc6aOYeLJ
bafwSRIFkrGeD4iE7poHZihVc/tUwKIyjQC1Anr40rf4fNYt3rVt4MyM2DQBdNmWAyHZdJpuAiBJ
fOXlkYtrRX50xHBvxYpp3sF05R5jqlP3XKN7yXMPDw4RyJYIlFfaaaR4vebTD8oIvhoEqEu+qWCl
PGvhSYWQVg/db+BOi6Zm5ajSS+atEbqiH1fLWr6iekMuJWaHr8pfdawRHnwKZjj487ae2tbVk/et
ojUaQeAlH+BUNyRsesJMqHZQLtxuOEHvCWN+Kz7/9Q6j67p6wyVQzTttzmYGnQEfxDBo7yEElwso
HRFnHFPn5BiqG3pFegjcPvWUd4ERgdQ2yCUYM6PhCSZ/Df+kaUtdrvm9CIKpgX5tLQ166StkMUJ2
Qod6igTYp1xCmjtnHxSl3r/julawJIky9hiialWtwTWXlnLjGTag4rP0lkiZaJagqhw7ire3He0J
TW/oKtC4bYD3mDrfe+x3Flp3crUfbSBswEa6veBtfGzDpGAGX46/aaA9tv93bpo2CvMwjux6w+q9
hpyt8tYPE+ttnnUkS9p4UGe1vJaOEH/GeFQ2/XdxMqrTvwzMPnvhDZx9IBEyBr2YSzXzmjgPBMFi
KrA77nFfZW8w6H5kNbjp8wPwDeixLL7f509rCjjd/EylhHxVzbjYWvG5SQ5ZziKKY6URuT0rCH08
bMdKjaoRFbowP8TpCFHMbwcCOj1SZfF7/ydLTFzOa3EV+9+bm6UXnBJqNSHewLqr4pa9vEdcGqH2
o5d/GTLgyK8JdXnSEGsYO1qgovVQeVFYKndA/oTIt0KO47guID1ZLRZBNxEyR7zq8Tvgm4OHNLrZ
fjsq4tPO9H+6PlzXyyD86on/pryU7L/54kODP4mbRhJXGQOsFe/v7R+SLaTWJtgrUYh0dUOSH+tW
6qw/ZemP2JZzoCBrOcaTUH3Ds2Ivo6efdA+sIQox0zIQaR6tXqwQ9iMf8cYsLKDsOvIRubL/1r6c
60gadnF9///jwJhzEuTqJUTYqVYgybIHm8/5EH9V451Gi+vXvvVCwXDgytYTDENdOVFr4uiTtOfL
g+pZGxZINaHxb90qKtbiO7ovHJosHN1qCVlXBpJKHxAE7JhThWTfUDY6mkEDdD/qJxdxl9AN5+TP
rAmNmZU/rH+grbX0fYpXxW8wopOkRPAOtyyffunWWrlz0873ou2gETESYRttalDh8LQd6Teb9a4N
kq1AS2BX0sKnkGlSwuuM03XFtEiYgAmYjXDPrjkTHeSRyBV9cHnwJotY4NeWrl5/Des8YibrOUmk
Z1b9Jn41ExJS0kBiu3IH7Jr+4Gyxh4+K+vNdB5lNEwv8vO8ZLKyny+1vBPp4oZRn1p8r06UbJnm6
kMSwR5tVpb4gQsVn1IOZOrj/CbZuzSCJ/0BuvP8ujxmnkpIZGdzkcqtzgHIAdHU7dsj4ZxcWh2x7
Xg3pCHt4C5R2fFnLBy71Na+UDi24Y5JwgVnrTBcMQSDyda7qNcOQ3vK7Q1VTT6AMn8Od2pucvTGO
M0QtFQGg2OO0NRRVVTZJn9i5OgcHSxAYOI1bOTa9S6LdjEgEihBd48SCh+2LYH3q+fNGpx1HAayX
BeBYotItHoCn99YGBmSHBWggnmvzpRYqwarCwQafgXnqNTuE70uv/7N2Q8tSBivY2G86zsyDAfMP
AlgY7Sdt+SAgJPovzLRRahI+ACOCZf+l1gVTEK285HNxHlYyqgEPQUC+ZgUR9VY54MURpW6BQVyH
Syce/SPuu+fhN6VweUTE4MrLGqposs7GKK1PnGKbVGjc2R6pjaGe2dbxSAS1ouVEtb37p2P8/fkx
B3Ak8RjqDH3AdWR8SBwSU+3v5qBik55yTqC0K46ISZv3y3YAnehu7+QTE8a84q3K4SQcWZyboZfl
3y756F6weP5l+Hmamxi6o8TzBIabub1oe6XSqFXGatk1q5ianzp2xS/oMwBYO/KK79zBoR+N/zyN
YGytcWolfx8GtRUHkPHWB2xlJOP0or3XDUVqZzqZhw3SIOT3jquPUavFoW2FC6KvRmJ6WTojIdI/
kPiteIgBZnizsquvOJ37FKTNKwABFqQxaMnENJo+yrz1FiEhOqOMzo87iKWvGgO6ZVUwBbkbh22U
or1Yg0AZcS4beEZczzE595z3ZyhDz9vUqMyTlt0eREHxC/juQ0MibKbu1V9p6I7rMKudw7lCw6Gn
uBF6lFmGLhPanLLkSKTsnjf09HMxPHWhxzzzbWnqwP+4b7bKMoebCqNujsoS6hAWMWj+cG5jUIjN
/xJnmo9TQxGLnQAF1GMFFpktlr4QEkjYkvPaiULDTvOZbeai/rz1ob4WrfPXP90m8I7JvafwkFxu
beAsfSbyY5F3wYk8FI6KQUVtILgtULGv02RysADxA/mE5Gc4VIkjzwyIU41aa+qU3nSlfv+FPtAP
T9+SFtECkYk4nukzIJNMJ0uC4uZKI/qkHymb7/JeSTZ2CNe8+YW916oXktiaRiuARqaPzMSyVM4l
J0gtgkOLAUeA2NjFIrV5teQVXezV1Lv35rMSf5mdmqx4oyOmoTweL8x0kPVjAneXGPVEICsp4o34
BYQpFqfrFkQHEjcsmbHXruErC65vLxhiyQF6zQhCJxEKvA26iCSMcx5J4kjrGmgjs6LVHbwmslm7
rVOIXyL9845JXxPAyWkVD0qqQ8fHACsBotDkibNfnkcNgVSxlMC7xE122WDjQTkiO4wcDnIp7BDS
N6BDJMdNkeQUbbvbSevAEgxIulw3+MNRXuKeETx+LAa5WwIUZlwHXbWkofOXAJ6gn5PddT70psXJ
+PYYMe8GPO+AcuOZ0TeZMeVvx8RWoxrYbd687d/hhpwlFAgx10u1y5hhpbvipWksiBguqbEU5lEI
PIwdeOVjKaN48NEXTz1mqX+X1PqxjQP4Iv8ivJMn5eI8uaDfzC/cUoM3tWE79UCxd1/F4uVJhGEL
vttvqibaKkvnN2/KCKYkRbok7WTxYn9BvHspZg1Q5R5wXFmIVwsJzQrw0sB9DyYnATiNr20Og1lu
el7AbSu0TRMZ7UwhH3HAeeM0p7uleY4jxdIyEMU+jKa3BCOf/rACwe1iSciKgLDvMouktGQnBIJD
VynDtevekIdOE9C6ysoZaApQGdO1uIjuVNTuQsBmLtGqhVZn4MBeR9VoJB7LfL/mJFFGPVjx/yvF
sql2I1HN/FU9zkWvT8Qtu3i+0yM1ljtZoHJZiobET20XzDvAb05FVL4hnMYz3mtZ1sYpCvysFT22
2lrI2t9iop6GtYlHYulaGf2ny0xAZNOgt+xTA7NES6T8cJGWPKh3Avuzc2c0mFMM34r4SAxZPGKs
CmJ8ECi2ApfNW96yYAKuKBI3yDjf5RG3C1y9m0r3cUOpkwn5kS6sRnhvM/Jc1QwMXXa6CVLerIpm
db1RLm0QaYRV4X/TPaz99VzA27OME70gjAsF5+Lwz8JB0tIzfovOu5zD2DYKm5NyDGL8oB0LAi9c
iP41aZZ/ik5GRXTWe79pulZSKP87WIrgHfPfdtyYM4W0IAv7UVLcnZ2YPZPzctf6CW3IZyJJfytR
WoLxaBj7qj2tsJm1P2tdN61mZKAGSyZyKKVsog6c3x+GfEKi2IsWRowVuORWaGZdf0k5/pTIgeo4
S6vfTQ9b1/GQGIOIeuYIlWG5pAEc9RbgvrRClfGtJx/Bso2EFJees+LPW8C3KH2iTreXu8UeySgc
A5Ul4IlnQU2o574MIARWfpB6EFrYcMAbQWTCLaHb7dzCVAiGomjmBkal1JdmihEXeaCNN/hUf6Vh
2bhM44SyjLcQmgEGXaJVgs5LLizDAAbdquLo+Q+ZBMoH/oRL5ee5X2ZzGNaAo3ochvOyC9TbLaEc
tHUdNbhB0YwzVj2WqaUSa7IfZIlO9N0+HUwlrGykqZ+rPsIpdunscHWI+J+KjwA8Rv2HSXyI9vJ+
kUQOcRuYPdj32y8KLFQXFBbuOHgk8Y9sj0UUpD3QGbvhWlulcgR5XLvcmSu0/+44tT4fUuCxd+Xa
0mvLf556MI29laF2xKZSWKc/QAt61abVxNRgk9KwsFaFe9mCzu0ypwrF8zToeSt0WlmzVOYNsnBt
+iXanAZ818r8cksMj7zGVqHMLEi+MfM3t0hREdGyCLY9W2vHkjXKnC/QWNCX+naFYzFdZTcBvkhg
BrVtVMnFjHMPb370UVhJJJre78KdXKMJbdC4CY0XDv871gI30fWbhs4esuUDVM09pBKYEfKgLsyo
yPBfeJ6y1Yc80+FCAdcWnfUgc2bGlcqBxvRLwkvEIyt0Lh2LRQhDtk79+7szRPGQIkyKjjXsNv8m
3n8oMo98k8LPVL5MKkzzBa79xcPBmMfQ4HIP4VxBWWuWLge5CmDQxnJbb2OQPYLUGh//QpzYvdjX
W68gQMqvHxOZ7ZnvDN7GNYZFXHrzDsN+JtXPG0L4GuYYGwn9yXmk1PPDPITLjeLd9GobiK9EXzOL
ZWa3Idg+0qcEzndm3J293chwf7ZwE3MUu1z0zRYCcnb2ASz06PiYMPXvhBXv1Ojjd8722qNXeJgA
eTR6CI+E7qpUz0OsCzm9ysSQUiIbR0XjTmQpYE3366t/fyijoPFcP2R6FBu2qCvRJyO4cPC+Qjd3
qmB5zhjV6xmf1AcUOt1hjrWhzfXf93o0W53H28vTDBbn/b/OKPwN4oy9eD/YwfsQfwPVXEATEAhI
+6NAdSfIzBNF2BkQERrC16YKP9AF0573WmYahkEto7uTEZst1V98OtT912kPPc8oJDpxqzIhqPRR
7Pt36UyVnf6cRJyoz1tVbOuTaqZlbjoa7dC15bM8i97E0NH1QhN0V3qw+8p03lxlZIwHEtb4mN0F
g4QZtOppxgmoIvASH+VXqRHfkQoljBMW3G1xegjij3qo6bI3BGHASmdCroLdzDgXe2yo43iKGT01
1pYgHRGDc8HlSllGbGVB3jdfp4nw5IXl/aU07rlWkD+cHN4FOBNRq3mxJlN6Dc4jCJZWtyIApU9Y
ysWpVjXnYDcb7LeezrNtSMgfK7FwYgSq8rWQMxFP1+v5+/KY6MBVBcIAzbkMztG7d6vcj6JUNVDF
XRhYMy+hI8C4S/g63ic7Vgp5xWV5DY5mJ1KyVWoOKRLka6b/EVXEIQxnL4jOaZo5fjNUS/SqpSQa
1bhkN06z82Ew6POtlmRfbQqt5YelRfYmUDwN0aGu4GMR1AEfNf4ncq2P1X7KE/zxGqNzb+G1hqYO
+XNpvMO3/KSM0A3j7yXQCxuDyJLnv6Ikp6oxgCA6fx6lDqvBFBecz+LevjYjSEFARfZkWSUMKNy6
XYPxXl2+MmiPNbbdPLZ4b8KvZABLSLA21g2puS898miS7oVNoNUJC9g/COzY6WslD2kC4PID2LSi
k8TNqhoWdoANb+zWwXsAA+kUDii+g+YTsNlP7+QHvaxHQMBOGnd/g/H629HA9lDlUddhIaBjmL3F
AeaxPvV8n+8Am1ISxhmiEmFjuaAbdAD1Bbk7ON9LBplCIm10dQz6ModEwHVfNiZEf9uzeFVUuC3B
TsU7Ag6RFS1ySGkeel8sKjvF1TQepHwmgZCbV8pSDo3+K/IAb5jef4uO+EbAosjUgeFtAX10Yxn0
YMfaFlToQ2vPsuzCe8NqHUWGTG9Y4nj8xqzeHxHcWZG1Rc/SY5ssLHASAo50pzKRbZwczVVCfXIO
kRjSzW6af06jKMzdXLLEJ2Hcr4nJ+tLOfilUN6DZ49vsPbwr5RP2X2hJ6UrnSCR+f1RwHTwLt8v6
oMv20RrUxePtXyb5P/tUr7+zgIPQwHl53fHlz+W5wOiZ/mDRnvyL3hNyf9Jb5wXvgD0dpAj745oh
19BHGByyULMLp1G6O96f4f0tI6My69/ZN5yCUEir+OPU7lIG9zPtjH0bA3Zzo1mob4yzh/+WNiWN
eIR/YGrGFdRfz1ZgJGqCCeAIscYGsMzawC8XgW/DJxpEiLhTuTC9alcL0m1rpqAfcn9BCd/jIH2q
bd0MQpyr3j9gOadCkXBmdfu1c2N4tNET3MH6rSp7XwSHeOSmO6UtchrAX6gkeXaQjDFzhq/W9V5o
34rYsT1V4/g79IPERlwGIt7Y0ls5Ct4YiMLFOOAuZ3rUqS3l6dEsUcdD38lhmt8UF71kVtks6roI
6bbUJ7cC5PjFPX0EJW0NFTXqdirWv97boHDmYdyEBaFFu5rNUUJDZGHM8Knh3JuXfiIMHo0aLz8q
N5PbhOSm3CcEcJo+pzROkibcWXn5IemGbAQGRkBLpWCutWOsSjsiy/A9D12VDpOVPig6Rb6rLfms
UUV/y8u9mOQscA/Ol2SJwZ+ifRzlkmo17KlldzoZbH8MKLo5PT8iq6EES6GKPDMBviJXrxTgsJpS
CMWPTrLoV9jNKP0wx/32Yx4KFLAMLUTEEz95O/o3Ir6nnIvVFpbuL57XcrwJWDC0+ppMarHHlhN0
t1QvzH5EdKVZX755sSSQPCBJF0te4mYfDMcxb6E+QMk4nJWXe41Pu1ndA9Ud1OaFik4lXMLJyfrC
muoNvsIBjhmlLtY4tzYb58cDxc5ohe5mKjysec8U1ym+4WWKvB8Mr10afloGNWvQOwgq5JFeMSB3
GvvxqJHpHihut+ltcv7xj4jh3ybjyGD9LLgJuIvrZOPPTvlkE6qRbR3BMVQXSh6t+41GxzCz45x1
7xgdy7SJdvrKidFscEY5UMPV7ICQJQesnjfJ9e3yNDRlR5Ulwgmugglz5/UXzZuV7IHbF+0z6MUS
AlZyROg7eOyRIcrQLQ1/nvikSqc8SWVBcxiuxWv1RKBnBCqQ6wvVDmKHAniV4FdDDYSxFh8Mt2v1
ghT5kbMH6xA7z3k+JM6G+eEV3IOwlfPreMQ9jMn6c2f0JV/yJBiyGnuV1uWCHNBhgsFqqamqeZsW
dg60sgKDmWJoxsLpY+PH2F5Tj2g32U5yxKJiylsJw85dFKA66Ph3v/1GnJnwk7Jh4yG89QCIhhQL
X1jfF9cCNFlREts0d64YSzXdkR5vX+U7MQpSmWb39cLnbNa2HfuGhfGgJ1HYsiCWXA489omqBfMV
sB8lxiGkCxAW12mu4SPvbL/DPXWJtcR/YDHbYk1UE6SK27K+FmdhqLK3rUwF72XhQIj88BsRb1vf
MYSJFA8LLI/OfqY5U2g96ouhRbb4HPiubuMqZ48j6jsU00N5W/zvaR1T5chwZBLEmq+2N8H1xMC1
9NhfaLWjyBGQ2U3hiSjzWAQcNs9yHyuqkE+ZhcrsBXMuDvMltzD870y7vXbcSdRz+4+ds0usH70u
v3AA4LZi7Q/3342RNvssMFmL7MWAkfuXQD6srH6GcdZMfGiCN4Jf6Ir95SHFmSt8dGr8FwqR2jk3
pszQMosA7XOmiKKDtHkteEWvlRIPx2C1OUzfxRyBDs3Sf4xY/KZgyFmOmKuubMg3uGWu7KZjFC2t
YAi53+Qt7tt1uv/ZLxKSuoHG+XwVcy6UiZfcVj69HK/R/LRvGrEpcsXVKDhoC8co8Am350aj/ZAl
mBVmyihibyGaOhMrBngkXyP3sMSHJc3Da/h7kwppJYBoHE1pC/63OkhVkUiqLlphrM6lU5gqbdvh
YzSh8vF3Yr48Cvz8j6UyvLZLefih8WZC8+/WY+FoUISgS+ezr49L66ddSpmdsS6q9VV0lGZiQV06
k+dhflxNa3WOsUrLAeMYghXyJKUYz8u7/tL1WU9Qy4TIF7dmP0gl2oL+LDCK+uThjfnDCigvYxH8
TQL4rBJhpAMhPN1y3nklTWjEbgtOl9IZIVhzgz4RXpMnnsC50SoKm95hQ4Po1MW6fCEvkNfGkNNR
/V5uiBr0FtUGHNE1KhpbkdfnJPiye8O0oRL8Au9NXScnsvyWM6KwKfKxXUyFKdqNWmt2YTu2TTro
gqsWvCQmR61WPsIdgimZdalJyIrCbQ+TPaafJsIcdaxYERD7gyba1I1DYx2cC+efpFttGmlILX3b
RKJ1XhEDVYJN4yBSh0mtLfc1InzIjdKj1ugCfPHUbHqSSgddi6/ILom6q2KBE4WvRK0YBcJY8lBi
bBRLIY5z763XeFiZLtVaQAR7B2TZ840v9tiCoRqyeI4JWJBUC9GukE+e0R49ld872XLGTYfmZ/lB
/zNjht7Lvp/nldwFhoxtFZ7gO/k2i8gbaCAsk4NvmO8SHDY2bpEo8IPzmVYsgjc=
`protect end_protected
