`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
5hA8a2BB3Ekbqz+YL9K5f9eR6f4tR/OhfdGQOZuJSllvqD3KbCs/4bicROPeU9763kxcSoAxztHe
Rr4K7KyIjoGcjzXr1uIudbprDNNFdL+Ot9OVmcrA2e7dQ7461/rrUt/kicmGhDoOcZIF3giUkMKn
9e2Jbh4sVJh17FBc/oO++UdQxVYiycspcjlCOooRrFm+f3YsiD5KJf1HiI3a0EkRwSzHDC9xJf4p
o72CBUwO/HRCSHL5Uo76u/fHNJQUvmOJm7B4B1mQmsSdrUd1IfR6sAKvtSG//66eJ7tSM31DDCwR
7qD+SDmEAD7w2vYyTTJqb6ND/kuYtmgKg3qEGvCm2VhZOixv9OQyPOevmZfev7ktL1MKy5NQvcGY
xmKPKUD9I98gKcTpXqy6pxw24bRzllYHNRGWFKRu1v6fUVYo5ka5DR4cqtXtoYRu6OFe5o76oCp1
7o/bffGSaL/fG1F3nCoG7OZ9cTvIyDu87ZAn0YRBelQ9YbwvWjjMPK51VXcmZI03W9agOBGpigTX
3L3UwY7129K1cAW2FgSnUKFRdjc/iRbQW7wJ3A1BhhH3hWtIYrWZ459LySofVjNgKgxhxI3Xe1Vv
ffBFvIDEXMJQMHVo4679Nqc7WyE83IaXoKG67JYqRixMaU8+XLSGl5gWjsGvMyHSCYxal4ZiCm/n
+GgYDViAtUGCBtD2EzDKKQRoCBwMdRD1ijBUh9OFsHGw+mO7yNTrnzbuRtEI3qdsp4Ae91f06g4e
VI5AhY01DEALiNtDHT0BBZJPIUg2+wOV9WomChASgcf2DqFefXPQsqEbGPwK09W9Mk13XG+WTpsx
ZoUPkKNYerrGkU7ZlGFRKMctCZBEgzN6YjAcrPWJkr//cDlfdcMvMUKFnZaTtpLli6jbepmBWF4e
O+0p5/Psb0Yg6Qv1FDnVupCKWaKHMIodRlzR0Pr37hZU9FgoHSNmTdrEOIxxOdjFv5ViFIm2Hrpf
t0egYRu+uGN4ZyUhajIlKdFb+kyxY2B6TPHwOs/4f30xsxY+xUMrl7GeHh2gQnEZ/OPB1Q/23tnO
CkRcSXDGbx6DVuLAKIEa6Q3ThrGH9YZFWb+vDhhScwGk6K6smGt07Whhxqz4AunnWtHYt+WdzWut
RSu6XiajmR16SKEkf66rS/nUWuEgAG3n+CCfkWSbAALbs64s2kcxbpT0U76cX3ZlhG/MVsABsMKX
zvZnqHajvRl/LnOLoiMczLU3GY95+xcwuuzexgy9A02beMQTr9oZ0lVgNfHgxnLU8Jpxi3pr15Iy
KhafGaadgQIl4SY8nf9rSCmzm+a6foVRky+GAGSDzdQdBAljoc+pR7u5MeI3mY2UiZAdgtQFX78b
4u0ZTd2thYXX2ZuEAFv8ChtJWefpdngNi9i+5bVItNknH2VbE+isem9nVGygzwp4SLb4LJY09ZCJ
/XFLKdwFyekf3EcXwyRvqMVwzBT26a2R59AW5+2WqrY0s0i6wkqDoijMlOylCI6GIO8MWr9G41y/
YW0jFmKjYCA9stIqBlK1c1UUcp/RGG2FGx4v1pTyLsQDqw/qGELDCyJbruzRqde8dZEa0mM5ONj0
onetnhQk6R9f742xEzbplSs8arhpNBayb1+jLRm8K83XiStG5TBdWynmbKsDaqS4Zr44sxnDiKvR
J9O+j2HBXV5Q72hrqvPOVXgzMys/S+hkEkPvFqhPEUTSeG8Na8EjQQHFxuKg4ApXzZqg+pILA0ur
OlOD7JLpTu7R47INhcauhcAbv91uBqxpNiM1lXwiEbQ73eiQupTM+hR8v4yGB8FA8PB1FSSU0JlA
xFppqKPoklxnQlEEhc/bsitpnPs7bOZTpHmk1ekbLVRCBqDUmGGgrm+RPOyvqlPrHnYuk0aeGinN
XIiMNV9ZLxGJljUlVILe0GnfBc+z0E42nASZlBaVQNJhO2nZEtvZ9oySDZgqi+IICVduYNHNGk1n
s/JuTCY38d0y+Y9CnO6GVs++F5N7oc+N4lfymJ7u3YeO28DAMs3trmYneFWPDZsWqXAzrM1FXA5b
PhrrrP1S6buizJkTl3Xgeig5KF7K7eFvGUuCK2Zhn/W13KJbFnNRWHoq+6Rdv8GcoKKPRet8AGtv
y18OoCInHeTHEP1vJ3JzL0hay7iaKsqhGrxITN4i0hYcSSw5JMrJnA0EOEPvx+My8FHXbthzNXjV
RDNOMA6kVW4H4wbpRWvxjjI5bVHv+jcqSl7aM/Wg1ykpbZ+9jGMYje3t52KVVAFAboeIFoRsET90
V51jwgecXz76i99WvxFrHoCWfMkm5iSjVPiHHkz9/h4befd7LR1T48icVyd7ZyCYgE96pT77kpZA
URS6hmpYEc5cwb6QkKS3akGoQFdL73EHJCpnXxT/AfI/EjadIx1JakR0kt+dvKfEyPW4Qs2VNCDm
cHiE3x1nugpioSVwq44H7Adz0Vgj/5Ey9dBLFdNID3lDWfnUPVZKbypaliw+r0e0hVqE1jXFPkdu
AgyewI7OJX5g/P/5YSPFXGZPP84hgtMhd7ktyxn4xWnwv5pDxJRrF11IMrI4VkqUxXSpJQK4d4Wk
pa385eKkpesS6xqbp9Ux+ECCXhkhE1dyjdPDtP9kuIGAkvEc41dBiAXoVqTaYtUmGZCC9ssJ352c
mF7NVPoGYMLrskoKgx8ekMvKGmWxBIC37NfPLJWrdUZvjx4mqrZBtku1RXAdEtoKBVW1javHo9h5
pK7derskbCl2N24BQ7oNbe+3oQ8zPNVxu9IEtB60R3ZKJUzpdE91slpo84VJ+SMTVBQVu/2/bLFd
6R5W62IYDpzYa7KeQbbcYF1YFFos5cLb69m4BqhN8GJjQdhreEDRGW+NQTg8KOu5Z3ZO3FXkSnKL
iEZhF0/hHO1AvWxj84Dpp1kPdmk5zRKJbOdYm7+lRUzLkH4BEhx09UeDXGEz+IjXmJqfMIgPcGNr
TIEBBis5Q3ZVDDGAkbeNFNJC401+awfLu38rmOqwQbyWwWVIHGv+4tifFx+JQ7k+cJk8gegOt3GT
4oFe3j8/G7u1dnpg1lXFqDUCc3K1bg6nUDWky+3jlnLRnT5P5LpH7QwlaeMadXDEYOnL/0ohH0jy
BP2kNsvlVGoM298Jnq35YI+YPJcLGajTAIH75Rs6Cna44NsQ1S1KX4W16J/kUi1nNtSCUtM14inO
CJTe2s6tSSdjaOTJx2bYAfsoSJbENfPmBiJZCee0bnzYx6GVPtlLzU54FMWaabvDtS5onW/pRBDa
Dgjeu/jVhOIviQ2RiEyfxoByS6RKuz5uAzvNHO0tP5m6H2G4u0Nrk4ycQLKn0lN5NeW0pAF1LK1M
UWAEgJb4pzp1MjE2AsPwEd1KamIXWXCKuzSGq1akehNQ6pHHBhReB5CBtZflZH5j/nv7qewQyE7S
rG3aj1Q30JYrNMB7S/209JnbetZkJVMOCmpvl/O1t71HGVJBLcQk5K3HC3a2/dOtqiYHvk7AT8kO
3ltpNrDUQG6PDlN3rCk4gtAK29cCmaYMi0vqZLfW4DV6SjGyDwXJTllBArwJngGU5AwyDMBhPYYv
GnPnN/rhoERI4V2nj5mDXbX47AsPx5Uj18c0GqFTvY2XHczr67JGQQYegRoB+6daqVsOvTd5YEBv
xE31RwkQB6ogOB9cM9/MywY1dY0E51Jip+6xCYPrTsR330C+SieWF50cMOkFjVrD7N5gdU8CzKa3
dGK/j+fafsmkgWdDvsEXjdCA4PBgL4r0jpOH5m5tlr/YBhhJtS9lPu1ANewjKn/JeCJ3RihoOjFN
1HTKtAQiYsUuIRhDTMFxVEOorX4+LMV9atBOeLRB/GWQS4DWPwUjl2TmNrLjeVnc1GKzHTcj57y8
KqnqyjhmsTVHKA5SWGslcUP5fsvIRQ4NMfWegaKcVXNIiP2tsXhzKb787w/8sDwrkLCxPciSaLQH
rGNpo0UmxSBsIO1AMYXtQIObIiz1PNbYy1Zdd5gpFFziXITRZVCXXNTKBMSwzMQ+iJmny0IDsmAO
nskZXIJwc419QBoAj3/8oL01+IKQ8KUklERyJxGEstbNi7usWt+y0hs1yM6eoVfjHhqqPObvALfs
UmL8ykVORFHQxf5lR49vKUVEcLBsuIHNRhjoPL2rwJ21+DmUYG9CyLNQnW2ujt0xgvJ5EYLp9bHW
t9LFVAF/zFcKPDWVMCH2bpVGC5hKPObYMbRqeGt0Neb+
`protect end_protected
