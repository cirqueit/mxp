XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j�,��ǝ�e����:x���P��#���j� �V�.��GP��M�-aX"h|0�%z�S�ְ�_W
W�nvz�7p�%ݐcy�����&9�dQ��N�����>���+��|bE:��3����LgIo�)���K���FD�o1��s�0I��|9B�����ↆ�r	�bo#�Fm�<d���K��Y_r�u�r9o��1��啵��|
�9�/�O�1�����n:s-.)jnA�		��io��t���O(26�u�q�Ƒ&"+_K 8]�� T-�b�x��~sԼ��wU3@�(�N��p*	�E�� 6��IU\�%��ԔX�\<���4����wu3������Ϣ>�t�Z�Џ�,��A�|��;�HRT1�����ldG���d��$u6�V�ٷ���jq?��k�x&p��}��\��]D���Gp&�C��E�W)��EɳC�:%fӬ�	@�OhNV5#g��(/pG�1������o�=W��g�W���8r�ur�-�0���z��-����鳳��]�9��F�ܐV�v�m�q����j�Ӫ�2���ue�eY�yxVIzp8����\��o&v�a��Qx�Qu�qǆk���*u6�Cڔ��f����S�V�2�����Wr��!�%��H�X/]��yKD�e.B�g[!�qDE�OqQHC�p�w�^A[~ߒ�v�t�c���bS���J�A�a#��F�I���g���HCֱ7���;Hɋ����ni��W���j`n��:XlxVHYEB     400     1b0ȣw-����ʹ͠;w���ɢ~"Y놚�|9�,�� �i�>�ϗiS���<�W�K�D�W��<be&���{���ȉ���mN�ʜ�:��
zn�O���e[��uo~%������fcT�T�*y?��#sc�?
����:,��p��$
X*֤�`�U�?ArO^Ŝ��o����~1*�� �Z�u�`�2�� �p�BL	1�l���,��(�����}xV�����o[�!�h�m�eG��Z���D��Kn�)ԹQ��}#� �6��6��:����:	DOP��rA]T孺�@ӑ|�~`�i��4	�]�H!�2�l��h#���g�4�|����EɻK���^��-&�F���M�;����0��A�?���R�x�G�I�5LcB���t���P未r�Ak|w����V�f�����sxXlxVHYEB     400     160��ܤe�#����c��Љ s\��x�ב�\_MŹ)�k�7�E��>���a� i���bx�"Z�'6p+2�:�� �CNo�B��E0_͈�30t��ę��a2����Z:{�P4`��o2���0�qF1m?�G����~L��|��΄�M���%�S�u��4 m�>3m.���/hZ�i��Rar�f���B8�k	�c���k���g��==��?p�g��N;��y�&�1w�6����1���+y��R�J�$�.e��K9q{(4��A7�o�.��H�T�}XGwRSb��
�nd$E����t!L�1ZX�< W?��7j7����wׂ*D�Q�Q=`wXlxVHYEB     400     110&�+K$��x*U���2�*���RMԊ�0��R[k�'�Q�&R�R�(o:P�B�~�G;F� !C	�:{��uC��q��Z�5\>�$�-�	}W>j�;`L���X���&CE��%���<'pY՝����6~|�����,Ο�[OĠ���Q1Z��U[%�9=�q	�0�n��Bb ��~=���i}Ԧ`��ƞVZGi�1�ٌ����K"o@8�:!���h$3��`�˥�ç�b���e������.����2�J��XlxVHYEB      42      50��X��5�:V�g/����ۜn�Ύ�u�2�K}��]���H�R����kq.B-�sOXVG	@�Zu%8�m<4��q