`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
ORbdU6CF47soCBpnnm6C7GFQwMdD2NoNxFxYvJ/t/k6IIqMBzF69Yxd/ocn8kzi1IKA8IzCi6+fM
tFwqW5tyrsLWW6ja5DVu8Zo4oPEhlC3r/BBPnzjvDYFqnUN/9593GP73jEF1XdyRVpChToYFJ5Q7
A4mueFZYyZHYiFnQ3+YnZ9IIcgLlmOuXDfc+CVG5IV9i9w/dr59Yk5u6HuQRRFT1RwgrOuixjSix
54MwPVA3nqtdZuyi8YpnYOS4ZIBFPkunsm0rjTr9yOFfXoI6Wj6K3AEPRQGdVkAdMDkyFeb7ju8w
GPJjquPtCDCW6r7+8CHpv3Z/iIZieej7i23oAuKy4o8SQfPI/i9lsqDP65aMCeKH1kSpkw5WdZSn
Y55F3qzddMcvef+ZXz/a6Anvg1t8IhCegHwloK5Odm9+ah2Banqp1d6VRlbtNVteS+T1Hi47cOiH
bP6HgJZQvQ4KRqF56oVL+LBwXQyOrvfG0xPlAK3mqZNBiTsWx9/sBSh8N1leoMdh/fq2S9Jy+97E
f7NXVAd21E7vCMjtKtEXAFbiXdnktv/klHrVlVDFOEfNixlXGU9NQ1u9G4gmodG6hgnclP0ocK+J
K1y8oAZ0A1ymYfPNIXdU/wAPwn700flUJt9eZJu+jj0eoPRlG1YdIiSRFy80xhOKV42zKw86aGOF
zq3pRSjvRMRFRCzBtlcIursZYvXnjN6M6Wa2SpSguARzPAb1iOO0XrEEwPZvZv5mDOZn9j/YVnDl
0d2IyCgh7HMpvk3OsVhg0RUdxbl31E7swXBIkUaF6IOsOnsQz9Oht3XzhRJIQPtxnszoaASOTKbl
oZVutF9m87r0LoJ2bd5tFIi/5zj/EJXP7eMoc45/OpHPBQ6Mj2zrv8wApC3gjPdb8ToPs2EYYgT1
6Dz268uOdqTS0TuO8D4u6lTap6G9YzgX83ZoQh9eEZVUcnvaRvoeX3a2qIbHapB1dx0X01DLI02o
THqbzllasA5unP16wra2LifGJhsNAeNArRUNixbwaHn/ObKariWjJrhdAU1hGctZX4hyFy9UNnhP
cqWuSSfQzsAg5aBXhcrbInaq9akdM5IbxF5LfVWd1KukNZBDSaxROhqat50J4ePCbVYpJJjAlJCs
LmT0uUabgBF/wPHUiTl+4RGvhuGlzlvBQaUdp3amhbCY129swX5fmtIva5IOzhOCF8oo0SNJY+yO
vzDJhjb4xLzYP3tvT4QSL/213NBXqOEB4wLNpI3tE1dQEQtDdCOj0FwQRnj1icSaqwwCCfzpFIwf
QfJt2QiqpWksS6qKZ/DukX8P3aDW6hDG1Ys/xYgXevJ/IVjp+NrByw9zK/Y0Go3P6Xh3fzNiAxCj
foBGvDPoXMcoThIYVHWZho5rKNAVOYBzaclo4QCOt9IRi5PxSQjf0gUYkLTcH+N87sBQioGxwk8y
KGxK9L0XwvRfC9Eq81fwsF2sZIXn+t1m9WlcK9LH9EmXpVkkIXhMDpoHtTE+U6HjQlQBv3BKvxgE
CfRP94LHc9W5rZf5zuRAPAX53t4H0Ha/JNJbsdsIsNvFjRXyp8XnBbJBS+A13QdjTvG/frL7C3el
/46t/GY+tDTLxvUfRAjLBgPJqrMGIpi/Bed2iNiGNCBpG9L6AB9ggrA6i6pwxsWPL8uni2XUZvoz
qGuMyICLeyKGEtl0PwtqYDXo6i1+Y1DasKXW0jr0EUYothLolCIPWvSp5EwIAPFG262XIvKzeV+9
CzPpmjV8K5Sjr3exvJONHotzEwFAUXOs7wkkT5cInCaczCRvXxbNWl3Vw9jaXgfxeNGYqMsSno1j
OluuJ1BxvETTIrA3Sp8yFpXoykL9ImVUOpak4CbGvJGeRTnjWcd1j66Z9csfCrdOBzLdKV85thMz
VDb5lR4XHTkO21p/xWrPHODxf7yUsBBeo+T6MQ9XK+Bwzvfv3+PScO5kJeeGpVrhIVNg7ZbZj5Mr
7+3j1wK9hrsnlncuhKlGuIICzxJ27rXsLwRGehJsAR4Da+2y2BNOS+ENfBKO7JmNDUnhiDbHhjHO
1BlJ+z5xqoG21S13bJxkjHxxJtVJ6M3QUZqxGfgyFjiBL9fFK2nQSCaCJaeTRK+hlTc3T2WudAIX
39pvv+lIIK8fE2Jp5QLNCp8tGJoqdOhZIV4CU+5EVily+oSs40hMmSgvDCWlMyQ8c9G37VuPjxvj
6Nq1t+0+ds8NvE3gpl8wxpqyG+7AzvvjLBJEUnDAcOyPzlLr7kko2i+jXcCi5QqHAdG1gIRbPLif
SNtXJhyX126zzONAZO2MIESZ/bxLSnT8jbCb91EU98KpQaGomEynJ0iTRFows7Cne+4bdpYsXm6A
wplnCjGC6dnIYKG5kyZdqixB3kP1Y9+d/Ju+NAkOYloflNi09Y2zzK3Vo+opQImXmLaArf5mG4SU
sKpapdyf0RCJitGie03hJ000gfO/HLYNncASC41fxR8GHTZzrSz6hRy9o9tACxKPeHbq7RI8Nod3
xf6xoOv6mO1csJeJjKCpGd19/Xmh6PCfNAovCst2WAfcJEB+yLOmhg1HnMbIR8GDC/sGwZTggHBx
JcroZi5Z5Hf5vWB2LIfNGGIzznDBzC6Jwa9WJjLLZOk5eKTs9t1u/ZxufCLuNFV8umktPseJgsSM
G/oNpTWcIkCh9/0pzYy4qrPXf82OXt+q42f+qqyOgzFIXQEf6V5lWjW+1mGrEnsq+S/r+SQHpAvo
FVfz71w6IpEpJWsfpdWeIkdiY/JezQkZvMewO3Hm1lAC1XbRROQKQbCZL3DEMwLrIDv282AZt0J/
MFSa+cWyLVR6U4Ck5A6bx+GMDAy5X87UU6ui2f+gQxP5PJsYPNI82D1LLNh5isuoXeC/dPJ1l1Ln
/E1Xu5rrp07bIuieDmkHKP+WZo2vghjLIGYnkhnfsfUf8i8oicFvMtg8WbZW7POvXT9R+ExUQNr9
WJaZRva5u0iGZewbuz7B2FUukpf3L/IhkvOOhMIGVtdfE7SDQdj1Mxn8tT6GzUE5RyfNNukV1HBR
R+WJqO8y4eW37gvoB7mWT/Qhu9d+JkbnFyXNUABuQVOuxamtX85P7MIrBJsD11pQxRB5JMpxANCL
wzzoIn0nepVGXKhtMuJbTgXmZp+IEAzFALXATPnBwA4dwLQPBUGd4erPAUBUKFO9vg2xd5jXwtj8
n5XiNlGQbTAUkEVsPZp+HEGDnqSebdHKPVj65EcYvdjPJGwZJGnYEMk1+EaRThdmhyNU3wEAoPNN
/3NcL737FQt+gwlJSJYp9zAU/IYv+UeABOJ7YuX1Aa0q254/a7d0aT+MUN3SqqGAJCT4/ZUwtEd+
UXjEEBPo17yJWmF/jnQ2Rks34GjI53tHDfi2AZjDpkq5ye3CT13nKgpPstPbPjT4l1GBjJaBW/LU
sChv76QO+WUYnPmtRNda2NA1dix/g9rwgrJunjIFL0hmrISACsLJKc4QQM5wWo3D/2EsdsJ+6Pso
vW99B60nMY1xqFtWDH9VlaL/svhhZcPlZTre+5AQVrmjNZfq0SMTOuaxmfYiZPy6eOrpzChJldM6
d/z1+2l/GNkw1LKsfNdeJnUClJGEXdIhFxl2aqOv0Zl4Kf1eKetlDfSumcK6dpmF54x7MIletZGu
CNRo+7K+RFj3zptfDgdE9/bY/DytnbT+Vum/VowKU3gg8z8t7IBNXZPR+0qP3IFTuOhgqYz2xh/a
JlPnCyiFT74sEuDGxzDYu/JYgMM3oGeM+10wz6lYBfY+OJDDw8wNmHn9U6hcXDQEIVX79h0UKLAt
obckIpL8pl+0jHddK02rB2Fi2MizmgUkwnUtxcvgezGYDsiKvvnnPXqecr+Pc3lkZfuDabphpL1Q
CKx997Cvd+htSklmGc3l/SdzZmS/H3m7cQePle2l9AaTG7O2huEYbt2XJdjpuOMNzhgLsqAINMzq
aQEhKiscnY7vKCAieQIIq7sHUEIQgCmyHy4P6HLLaKoQgnwnjptirJKAgafhGoXe5k5SyO9eiRUn
GLcAse+3Yu5bkBrFH+FMFm6DOOtw3l08U7K4O8oN372PBRQtHbTgK98Kt0w/u68KDqGd6vUtj40F
1NE53Iop2VryzKq92hUPV9UAgZhEaesn3AJgwnAAid/Ch8X0onPqsk2a2WA9uogXDBy3HAU8qtP1
7+kU2lj9RHo6tWBVxW8l+26ImDCGLFf6u1m1Jeo9lGvgOMLVwzN0t98ueWgjzF4ZEjuSOEX1T874
phHRiW1+zpbBeEdgTGH62mZypE+amg+8XTeYK+4hVAtt1rOzwJ7sC1aXHx/Mzkxsdght18omF4HK
EO0uc8qDDT6si8VeFO5d27PcmTn1d9AMU9oFuRfpndnA+ekFg3FAadHLkQFnnviDn1wRUayciMDz
1O+IGdgSX8B78ovTS2V6vwOVRaOKyUOuuCQGNWIINtIarudIHHge3uDhyamZwhlif+tB0IBoTO7m
TaZY6jrLUTlWgN9oAjn1q2y9At/fC+TnwdPpiM3RM5sHCxwHZDJxmFH0WNm4k7FpLkhm99ZlN9h1
Os7GzvArrhbKDVRhdbGxpvwtmVT6F8RXKNlhBTPeLU5njZZM0hEHvpjadLxaQKKHaZKNph3uS4Da
KlxFlTwdPBEN+0Q2O5XjNfVaJbC6Ah2461BohdjNZwRozrMf6X/C8CyyaEMeioeo7817jEvHZxQm
D+z3itMjY5pOm3XpVKts84jdm65FKcpEdoNd4oCy73w6WV4v2EHKdbTj5rS9WtJRpz1nAJray2yV
HQa66DO2AqBCZdBslMljJx/ohpCDLHg+N5+jK4aLjVflwW8khJL0fx1Ea7uuBE5RJHWtBxFO53b6
podvwd6B55EobxhrqsUXNkzl0/O+AEBNnVO9wEGD9sAofmAH/Wiozb01Hez4LMPVXQslemUC20Dy
pF0bWooH1XZToFpyhrblGSwpXf6gevCxkDysC4bsj9PqwZi44ccEdsUZorM7abIieoLfU9PPrgP2
UqNz8EM2u6R4etEZxYdhLPF8Cth03SkrCDfLqhb1ZxyG7uecxY1CU8MC2+2KLqvVRQzuCxB9t3cj
Csf9zizWFM16U8UrxDRb4a1Ry/vmpJumQ5DzmiQ18a59LM6/kNcRYwylFVLOQftiStnmKz65ATy3
X6jv758bihnsG3lUUkc0dBHaKi9VUNphBBN8TEOH/qKvVK8wjQWsrWUSmf6Gc9xT/qjRT/LlpMp9
BtCvpWMNn0yjiAHidTl0WjDx14UKo7RrgvbzoJkCYtp6m6Gj9m5ydp77XURpA8C0x/N6zdWda1jE
UlZLKQDvdT9VLE01dXI0kIhW6CbIuqomCV/YihCwTDCXpDNNsyDj7s4XBTCd4F4giR80mgTn5zow
5tSGXlnRX4bbz2fF/nM9Pflpl0M4FmCCy/OBPa2YuyUqq9RsCQepIpxcb0LR7zUmgxtfUGGKD2nW
45ybsBw1z3cSFy86Y4S1ivwL7PAaMof+HZ7x+VCHD2k06Ezn8lU3FHxYAk/1dBxauoxu0asT1s5c
B94ASsJ+fZTtNv63j7H+sHkJr1aXDC7qd5+hoSUC7vKlzc7+l41+IFcB7+399BszB27x+h79IhyX
upykjNuVmpdqIXpFF6hUErMaD0H8UXqjSmU1g7DO6T/7FVboDm5nsQlcnA8nuOnsGiBr/lBtRYg9
fG9ybKfCmv/9AEWbjRQRmQUXWYpmvDi8pLGAT4WcjyB9zeOHPGFS1OGZIlltn4UTKsrer85kAy+S
9EY6/pX9/9pDpDyAp73rYLWAIt1CdjgDUE6O7PGJq+njhJrmfeLwk7SwpOpeQEYtyP3nxjyheXyA
1JnEJ2cchpdo/OWO1QwBYzOF9yOeA4EwepOq1bMi385KyChoZodD1hpU69lsoce9ckOJBzF3HJc7
NMz/fhrKOF9AIrU3OpCCQW+CwT5a+Gp9LCLLv2pxLt/RhrOrXpDF1Ze9OEgG9HF59zxkOH6B+TeF
LWMlraomCXwRja88Gl+6DLEU4ktArCpvp2YWwiVUDPL0f/ubQao6xtBXg/iG9LYVC5Zdks7QEfsH
+uIwfc4mpOvKSaiL3gJkdUVIkrgA1P2kHzafGbGPwdudC5mobTjgaznOqsEmuPI5TNRJT1hdgszq
O/JNh12hyn7UBKOsmY6jKGOpNRCI/I8AMF4ewHdss8ldsy8W7ZViJ608ERXGyA8UYlllNyxZiLyQ
loxKyZRsrWeIzAbKXevcDH94ylSmOXnpaCdC7yroFoMfO8eOHtYuxJxzv12W01xoFf4fFou+JEIy
VLkgEa9WhGAOBZzvGuNqC24SN6Gmi0SmPh4I92mocTUkoIAy7hqqRF1Z7hB5vmtHVIwLajINNck8
KDer29WxKSbjPPGlMqDHOtiahlAnB5bCdlPaOorRnB/hTQjwnWLDQ9HrkTig1m/f9+a7sUS38KSz
LvBki6SHrNJDmWZsMuTs4x41d23aCEYmEP6rEeZkexvkoKksO271YV9LiQjNZ0tSFD3WX+mW8kvU
n0gaCQf3Kw70+vV9OJ/goCxSpZOtsoAfa0kK05aA5mgI2wTaHtxN8XMRhhp7LYMd/CMnQzXzw1v2
UTnxD3ar92PmXDeYbdfnkV2tUDF6am6+RBbK2dpCL5zJAloqt6GQkPLVeEyrCASCT9rBbOaTRTyX
BJCy7V7QVXrlERJdkvZfNA1AuJM4eo60v70+IMOlsXieuEy0I89E9K5/XgR2Kpomo5vP9opEwNGK
4KBwx2ptfIfcEO6C8FYvAETQtaSpAH5OA0lkkeq9LponV/mgME7jHi/+vOPCKc9j/1w95lQ3FDaN
WXYBVqqlgbdvkX9c+WXwpW6KN6sABaPrD6BAx2k2XaksYRsGbX4SilIRPotCZdn0EYd0H9yaNqp0
ksnEhEC/yryryV0C2KllI8M/0TxZFOTRF3AbsB2UcZi4w9+RiyjRuuBKNBov7q6VAQsxRDgruXxs
HZ1TV6QxhMfT5/O/UH5tQW+Umysok+vwTk4noaKcxxVulIB/iTDlDisuvLcILOGk9/9ebfaTE5on
/02LnN10sZiQOo7phcVtibH1HKidKTPbV7t0Lktq4poJ4xtTfZ7fojMTHTleSQOTOk9xAiIKeSxh
nn3ck7YtHXCkgGZO6TrrBdVXLe9isDxPmLv00hX5gwvFVfRLbf0c/1uxxy3fugZ6UzJQWDMcZbyW
EDhk64gXScn5dQVwd6pWBz2uxfZjJHIKDuJ67Wqh1lmPKLsoXF/RXRdzJqfypUnIo6K+5XkWbRiX
sSxl4aa5b1iZXPE5Oo8SFHFRXQcypCiRr7qIOsWguVDD4nniSGhTKjp/RFvxwBV5Rddo0fLfDB1U
WxMj+uSYrZxkU+pnaWc2s2/nIw7eis+61ABU0LTVpZ53u9ZO0KaL2LAXo1RDw/GINz+2UX3LuiZi
FtOMhCZv11WcCCDRV3bCgLVMASMOaTKjyFcLor6zPY2md7OLNpuUq5Vq4PNrXPBwzqB+aA9E9Dst
7iXb+nPVflQjwzq0TQ+G+0j8J9jadV4fXJH7HzINBoQV88EM2BYNJfrt/lnnG3fM7W0xUfUlKJeU
6fGlKZRQAO+2HV0175xazNpLe6VKOxfibhlrxcNiMlVKop0Bumogj9evJz55QM+tRn7EmUBuWDCZ
z7K5nZ324sST3vLJ4pK/wq9Py3ZTatkP+KGncPyEVUfyoOWbj9Nxqq2fAs2w9p6aGoAcHqNnSg7C
AITXAnpoXRKtGaZxuOcDrP1prsg0SOh3K6AZqAZZW6wG5CTco2wPbPMz8db4pRlnBT48rALuNEb1
mn/jsABsUDSCMGNtFvkhT/jndUy/jAw2TqPK8UJ19eAmI4+7ge0YGUg7MHFjl92UFlFKub+BPO9z
+L/SkXSPuG3goMIpuWQOZauDBzx/8sG2KUN6jye/ebdO9zWdph1iy/C0U3/EEmIBC1ts/GDRwD5o
WXn+x/C+XsczgSd+kRMT6euVai6wQHK5tm8xPuAoJwUbWGjM0waZ0u29wNBYkO0vPg/oItGpGJ4N
6ts856km6/FMXMbDWpKyXf8XXZybKOsTiAZx6PC70A+gnbN2y07LxUy5D3hbAhjISdqKvOnk7nr9
zPX4Ds7waxnGQigDhhZiCuU3CLczMenAn9KSTMiGcf9geH/7O4NdyP37d6r7veaFVdW7x8uG1K4P
D5vZ0yI4Nl/zBb9VZCdpQZHSiDMvu5mgCcUQYTzOBoKH0WIdwUPH4Dw5c+sStpXrrr00/x6jeNEI
s/chFahJZcyZfkDl+yu/Gcq9tkVCesanlYL0F81X+V4lWVfqFaVZ8XeFgw==
`protect end_protected
