`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74304)
`protect data_block
OoJzMukU1CD9Y4zNcXTMF059TVTM95nX7WtoVEVo7vjj8z1/3bFl9s8LRr3eUVy87yHnrq7JbaYT
UQT6F4Syp4OyvaZ3DVLmNr2qykFscUFNg4bNyvOuIKK30oVcNgQDjEGzICyl4xGfsRzY1KlPKPJo
Yv7UwW8WzSMOcc/tC/Yt/nq73mDlfSiEjnUXUGqxtUL45Oy/L0am1981ttBLISrMYZxRHTOVH70C
wLEBvukRVe7xIU8IPKh4pEdMDpEddHAnNaScLUSY5Iq5mAuT0SlAYt4oXj3pL3yTbJB0uRdgz7PJ
njPDWw2S3Ul7cJnWbtC4tBlqFMdgjg4+RcdgjgulTqMYhEejZxxNwTDmlH5gQm4IdstUQdFjAF7m
pnEjZfV/avMF6BTer7QitSFs+8uihtyhEdp97dBQpxJslMXXlRzr5NyZ7ePJ3ErZFIj6ZpIdyLPp
BjM007r2VsGLp6LSOgwyFB+fLQawB0gH7H14MLAm7rzt29qv1Lgy8K4/gEK/5wivFNikQbiE8MP8
eSWyUbj0QJLxgjrKHc1PAA79paFENVtF73xo62/TLazobIMQXUXv7KxwBRvs9ZDBmw2hxFoABrV8
ijeJJd1RJqq4jCmTkHWZy9+tDV/dQfZ/08jNlvFsOso3436TUQ/UwETPj7P5VBPimzR49ffOxTpq
tbO7EMM8YHkJTAPlD35rJTlggpbAWQqYBQLMyi4K3cvR7ZZdtSSQHCb3PHA9pKv33P6t5UcK3YTh
Il0/hI6agdSj2KH0udwYfNeGos2AW+Xe72+WMJix6UH6AE9ZT9yrr84Wl0HmIDcrNnSeWhsSBgpH
ex0Xtt+/ekSDvaoKwY/wG4SzcOaKPdYVc7F3ORRxEBI2dpBb+mvMMFb/E2R693m7ccIw0eUV34/q
H5K6A3RGuwNBbc6MsrUyvaB5YvkxHtKYFdDu2iwT8mi3sHqRg+H6semD0YG56aRaU9QNECeBGMat
DBe1Y2C/cra17E2EQPB3ZN0m7LBmXf+T/kO5xAx0/ig3kKW6AjHzJS2P5trncoNHHLZYTcvF3UWK
J5wEGlKpNeSxyQOe1fsWUs7MzzWNsHNJs123ceAAQEcx0tbV525JQfvIo4XApPy/tIXu/gWi/9iY
egnlKQchd/wtw5G4rVzCu0f4f7zlG5Y+71BAAZHx4Hk2a3U/rK4wqStpXgAHXsWzO8AYNe/wZnkm
3gdJgyti/LiODpbsKWsBSsIHGRikTlx5Lxg/wd837ClBXIa06Y3foiR04oPBsCFDRMNylNIbt0hs
9jsuKhN3oHLVq2y/pE8w/WBYn3NyNTaVAEGuNgU/f28IN4uyB6aY/TJkxVXwiNtf8MJPMGQby5JC
1byhioRfIWwJQx+aPpmZYnt/oUTU6cZy/Kr4y2VGqumi+bhmzLvAmxRzdcKQlIhvSE/y13isueut
yhZKGZ7wPZE0SOHlDIsOBnLBMIytB6fZqhdxOfNMX4GeM2ImYGfN5bz1et8N/wEvfpbRR/UlnvrO
5HeiZicFWzeTpOFOmJEvQ/cbFEG0aDjYor9TFPlwnlojhezUag/NNGD51JLB/qyT4igEtIYIoUlz
vVMoA2+RjBSR1zy2CsctP8eCMIhSaabEiMqFauEmKo8KwUc7V6rf8QjjQrz+TQEpqF+tHzQwJu9j
eBuH1Gc87n0AtF5zv1mM6Bib5iaBHMuNeWNA5jBb489z5jvrmyHv2EQigstO8azRSodmlexH6zdT
ElEOTTgRaU5XUFIHbxiVSALbW831cC7PEA/fOP55xkHRv99dwKojbI8X11EHMwjL7X5P+Idpq2S3
HxkKBOVkKqTFTswBKg/mrNkLSzdJxkY70CFxCx/Bldl1JeQMJmgXDpFaoa9u07nhOExNIZmatZCb
tzHBciAjbeFLCSdmhX+h2SICyu6EiBTZuWrfe8fqfjbyoDGTVlaOfxMs9sCJHJ3dPld0T57oj81C
LrZl6Ketwk626JuwEUnUskNIrH165h5S1FZRqeftDOQ+GEBOzNHQWpcRJ631ujXwo2OPQavM1k/w
Mv34w34XWqqIfP/JEve0rdX+i2l7uUexZ+XacF2e9ikn6xtC44jfMF5z97idyDDkgwxVBdRRs/oM
KLX4tf1sNHQlzRH0F424qTC/ggaPbr41AugcSEe8B8buTCUTaKZz/NZ+dDN93TIvylXDTFCQVsI/
Y3V1nU9ycG8yjm3C1sLHF/ukyp48DpLQDQ64qCtN0lR3NZLHjD4KxpBkJ6yl9vvFtykFFxGcgUQX
8MWTQ8P+3b640wK7A6nuf5Sf1q8Id/GK0QX0caKA6kpgA1+IG57ScjWRP/pB3BtIfI9N0PqEx2VP
fE+RLxz4htsd/IN510WjIke//n42dHPSBN89S2sxn6l3cvHkb5w7qlOQ7cCUkVYnRwxhw0hbuGMb
HBxvg82re4DuLevsHr5HyXMEAmBjsgn0bjRuIE+sOyG0eQipRbOLWOZThJxax+4tskAndc3ccUhG
d6z3U3FQEPWouvvm3CZxr8LK72ChU1xE0zCYeIFYcB3cJMyWRSC7eCQAgo8HEf2/YfH6VzUoiYAZ
uJ6pcVOElcnUOe0w/4bz1FQ9yB2rHj70piu612Kuj/V8TeORJCyFFBO59mv+q4IteVAeU01FIzha
lU43EZsS4QoFXaHlC1nXM/KoEVIPwEXk9LqZRdol3nD7tX2pNpUzcav//Qf0hxrhP5lnHd0uwQMQ
GT0qzbDihOsSxRTM8LVie5xDrjqRj17dwgPMvOu6I/Ms/rHuS638owHcY6spXv0bPB9O+uSuWH7x
By7BiAJZCxKVAiRKJPcWnQwNk/v7OLR+ex6roweUFrZiWUmtBsW+9gk+jOdEwTJkazQWVOeXC5vj
LbX3wB4eqfocLjM3I3gA8nlcgvM7tNZo90vB9vtzkYL+U6XMfjwi4L/k1yUvw/LyO99DhFAL+JGL
KIKjR6790SM76U0iqTLaQkAMniFm65VcOHiqsPr5syp9KLGGddEn2+Tav4k1BqJBURZd4Bd8/T88
NheaXpaBVTBITYaYfl5m9A8X/CXLLJ3jjKBFzL1xF4jaSAxaAYb6ZUNJOwj9ocKiPlFUbSXQVgUI
gw+XSa/CFrPA+Y7LeV4heuQZRgtwJ7tEuRq4dyG5aBfNBT/pWKFr3pwVDtXXdJq1f6kfnEvOhK7L
b9m06S2jixJmHGV7rj5U11ELrneLrCJDib7sAf+5p1QuR1RuZt4cfJxvdUCZImUe2nTw6s4Knl/Y
K0sdgAGa35cSkGEoEjCLbRYtq1EIFgWTRcimVYnjNGTB6YBZQXTgVYl45z4zmegvx7NWz0sywJf1
O74ejULmoqwRXaiYj2a9MM/AuBmbHoSyYgBvu8C/zjqUQpELQuMhgz1zNLC8Gdi9GHFse1NIxTbA
X7pDXA0N1MUp4dJ49nM8wYKzwFG963wSYEHlyZYMY8VWcwNoTtOfTDDSgfrUoZi3TO4sOrXLI+/h
98U8BMydTxXuAaZJtHni6UX95xVZOCq4iyggu3XaH1cdTk2PHWRG7Oh6CsafueHJDFojWU8L6opd
nswK14KhGYgo3x0FNyHM8cp7yZgFkVo6YT6cvv3cOUSHWAN9kkjWnnars5E8ligSBVlJyelA7iP1
9qty5vXEem0VsDsQLyeuhzkC3Shp+GJ5YH08HQuYrs8HzNPmmU2ibFXWee2jCSjteZBmmZLfC47x
kbvNlfEnTxDYSOBqjbxNjIOBKPhAPCh+c6Bemz/VS2PQS7EFVdTj10Ig5cdRVm3/Ce+0iTIY5ynB
3n5bSMSa7lrFPeVjf8b5jg3R/QjIiGJiJOoSyU8RLtY/W9JPlakFiTajJ+B/cjZ9DZ9CCECh8jwx
1pe826OgQTUxmunaX3hX08RwbFSNcd42+CuAt1sqOvXbHemtoAhYD+cmIFH0P+2/aqmWG88EjuLA
hsbgyJ6jC8SueI75nwNkt/CsgVlv4i8aoYbjRayLVcDAj0xj+32sZeyRvviKTHep/G4v4OlAEaka
tp/hVhU5yhlZfsU8JIf0JbgAWeYBwl0tIMcBfNRJdpiyAr6kid572STvP1OMyLcqnMeN2rbe26vG
vGxIQCZXPkfc+A9TzdRRGrSHx/6QuiVez0qPRyEOhk1tPKcSYQ3HVisz53Awh+d0prcUjLRvD2Ta
bMFXz6wH/rKveLgJfFRV2geOculHjO3nFSQcIuL3kxVEV5D08wYl1mSZcIIxPQWhOH8sdHufPgwk
VudUfRBsmdKqOipbujr3BwM1jHQG8FEBCkrnTg0wBy8mHruIbr5iTAHCwlhBQN31vFUHY7AH+Ejr
VzyseZrNBVHBh792N4tbLlSM3DYVrHI27tcDq4qggZc2fq3IG2HaBsF0A5JRsndhqgIOLBgGOeGz
AsZmK2REVLwpWL6sHsIfexH2fFoNEa0K1fCoZwUKJSi+QMAuzBoAsXXpTSyWyEcMpI1VGeDIDnmb
Si/AGBljUhX2TpKUwdDgZkFn5qdYt7bpnxNb8L15tm9MSq3AeURpMGyy9x/ZTBbA6Ulquxrh5pCw
MEggJFoRLsflBlD7PmVrOj4NMWj9+LTEhmokevrO6qeTDfOwejAJgXHNIyXcIEO9h3wNI7DkZ8QF
5yBovvZP3/R+o+U4I6CQAWsbngTTu8eEi4uixygmTyKYVvfFEDZRtVEkqTmhyorlaoMcMmgJhoKE
9sPqQCAqvm6Wiiy+7WnZVVd7kmLpotoUP5vfvF8yjAfof2UfiHMgQrn/6ZAVinmgDyCx/VpY7I+K
sh/qqgSIn+ot4h2SZC0X/B2OipSF7VVFJhj0maoA5kzZOheaAuzbpb0oaNSuT1ynV/gUrQIKRoH9
09RxV9wsfDHXuVmNlMYQfv7FsOkr30jNrWwY34ZOi30nRDwDTZGA+4mUs7u6CdMI1GvObxpyTVkG
qqP4ZOcX7zXExygJO0S9y+Pb5cfl+erxI9zGac5nSzJbNYk29UDf+Ew2MmUf+s/3CdV/neyodf+y
Cg0nDQjkmuLuJZM6PHstJExrx+2/mehV20YVUF4IVVkK8BB2IPY30BF/Uy6T8t44tKDDfKsNDQXZ
Pkyp+yPzGf4neSmAcXJc/qhlSunv0jHE5XhIde7cBAxen0M7f4wNyAQHv4DNE+yf4+7GQzlXIwsC
iEg2V+64DzYOjkKLKqP3s1k/C8fx610y9QqiKXDKO8K++Jht1TmXLQe72E366kRZGIAa7Ixuo72S
aoArNTXJb5f4JJOdWSJtAnE+cyiZtN8w4Jv5al2SQGrQeP699x2ErED2pR/17zCacu2+rABUZb4k
ohzFU6p2mY/flfzWvhXtd+uB0Cmqy2L03FmQ2yNWIp2Eu0ILxgqMLjq+7u+aw+o12LLacFzpjM7e
Bm7pho1Tljjlh0Qyu4mfhw/FJr2hduN9HB8TzLS1WpLb1AB1pU7E4Dx/mRM4eQDQ6FNarnJjpe2s
MVkeUlGJqI6PnmK+R+3kyZXSrXIaF2An5FQdSIkIRozIg9ngrA37eF8+l0m0q3D3HAKP4hAl1xJC
awDaFxKJ9wrPLmSiJL5eW93H+oC+/n9T3ViHQS9NURPttQ63cEIa3NoV8LtKFaDngyytJexDPCO6
UW6fhOeCuwANt6cx5R8JiIJBe7xOF1+9YeQ+htbxPPUsj1ahq4X4yao2wqwtgYpdPJAGF7nGc0Wz
H/o2n478eNunlpJ5X5rO/2CO6VxRUmOlXoobhbZS604/Bnl0sr+WbOZwcJjxQeayxOjdBVg+/g7X
zkkzTPE8exPDJYA5Z32S7bzDMO5u2WKzRS/oVlZB0bJYJi5kueyr1EtKdVk/5hUCdfJKH9Vujua8
jrmwglC4PcKKbyqtKhoT/8DxdiCtIXUDyZxqAt6Oh12a/6zvGrKQpTQvdF8PxOSSV5sZ0soW4tNJ
FVxnhq+IQbC238+zN/ZLdokjq1sQMnam1mOp03qFC5+zsd5Vz69ZpOWE8jSNyQuTat+kaAsKZo0t
oMl3ZJ/CyoQTKsnMruz75vjqdAwVFuuozmzEGpTmptTPAlOyoCnXcK33r+2uGPoa86blEbWzCbX+
SCuIX3rnJeRP3fLQXWboVNtCqeUxwukZ64VrMghuPUOGKfQMT1o1O8eKUpUNaCMD5uIFWrx8FWi6
hgpqCGghb8l3/CLhXdIr8JJ1kVDSYACvTNk7HF7WXej6KhLVMbWFY9KMXQ8Oh9/PNmOsycuzHYrT
4hDXpBUBSycMylC/MYAmQGoPPrZk/tfFk9IeUA0gvfE0RypzZhlkpw5grpZW7eiPRSAcCQI+DczT
aZD0hW5iYIXkGoJoxYMlNPVKKJjfv99JCs45eGJE0i73GMaCBTptWO1o+zJJyHvtNu2Jde0OvR1X
ql5TZHyRxafM5dVKvIfjvBVJiGBZ2qCMRrQDJNx4RTEe4f8D6OgKZV5lRJ/iaIZmGYiL/1YCZHid
5JDFVmtVcSj6PqJd9kGdPfo3FDJsiSXL+CbVFw9QFeYs8/gQLXtfsL+ZHfsjyA7JejZHjJZo37dY
cURXxspJDCvKaESs9xZwkBRpZBYKxkeChuBquiBf5ystAU7OCMNqDj8wiTZdzg/hLxpm6PY0AhyZ
V8bo4BGKz5JZATifokokC+wTHtr4mlcXLZOrRIkH7kOZqbsQGvS3eLQV3+g9Dkh57V10YdiQjlRO
XUea4DxA+AwS/zrnXdltVXY9TdciJVdcYkMSxICmUB812jN4pCxEQpWZfJSzmudT/iWeXLDlWYHz
/B30MAeuV64GTt0CQgNB26+EXX/5YDc1SwjcB113zzFWu2KCxAXrhATytQNE6s2Hoo1a+rBhBVQq
RmG47k3mf0Bquir94UKqAXUHSGCFmv0ej2us+38dG8XlNrbKTLDLqJijGP6qyVerOqhiP1zqY7UI
rzYpB9Du1E/g+UJcyas8Jr+7O0iRqxdS2XOqZjCwDu9w1BpaJm+3tuN+encgRqovv0m+X8tpN0SN
0hcDVArc4KOr16l6bxF92sQbBShMvHD1+iI0kxo+u5u15bUlLbPHRUUVlSGUP6eAt4aiPx+yPxq1
r3Hy56oiK8h8mwa1L9VpNNPVymDSW0TZMthteBLuXs9So+AUZTn6m1av/VoIsFVdr1XLl1g7LVWS
QoAMKpH0tojVAj3QY1vErf23DMC6odvihAR8XeZxwtXsVD/P/pxX0GgrQml82gS4QHwUlMG5ISFV
rBwkidwBARD5QaTjIDfq3hW4PWbmUln733yOXYt6MbBcfPqDvlHWdl3u0p+1+WNMAisDrST60Mci
41F0k+81+WvP5l86RSEu0Gdg9d5gKj/vat3HG1poIg1kH2Rl45ijwKkCqkg2+7hbIHWKS/quIaPf
tqea5alazlUAH9TdSTtTxMijxBePr2bi8FUGvEKvKRswgK+zgjuAiQraSgwx1CBGVwYfDE8AAjT/
E91tZe3PQcNWNZtXXIU9ZjS+5fm9X7V9b9LZxFYvmzzHECapNNBzP61TISFQjOzNuFEmKKtQPg1+
zcHRTZv1P9+E76XctOgor/c+cqEa1KRTOKVaHMzDv/tYGvIhCoW9g48O/2wpMtGqes/sxZDJRHG2
f/WJsc/FiaaA5plqkaoezEfD2f9MXLBbvCVLAdqVnP4+dx0Pl9thsB59ehxwzfA4DVkn4QOjTzms
drcMi4ANMsr1YzKbMCubisty/R13TKRfXAGkHeqqliXnqI/BtTWfZ43tfZY5NQv4KLtAgnnaVami
R3LbXusJ9RUnx8NRIZcqWWdTfbVU73wkYcQdW2ySZLWcUxIHBOrI5Kg5Xn5sJV2AjVFaoaAf27pB
K13+k3v4l/R3rGT0y0VgTl02FLkyd7NH/2O9Se5uKlMSOUBy2jyy3EN/k7AIFXcmiIZ80yIGF2pJ
Nk+CTuw8qcBlqLQWV6yIsp+rjAlGGMZv5OC+0c1HRGCNPbcOoQnpER7qyinh+sJQuP9yQ6M4eA+m
juWz2E3SJzL1x1CWo7WEe0nYYI65z63EWn9H0uW3l/QuAHs9xyIwDssrFpDQ8sfUHeXP/ijZ1PHR
kNruoQwUBFrEw6dVmj2tJgv1/1YpFmMh8QmkUbsCw7cZSHa9dbEAl1U0uaodjtru44lDuYe+ZcmO
aRUkUNRWKJpiX4lmnvC7YrTgxZjPfRFCD5hklGappry6Ve79K1PUUw3T9/Q7RFFFr8xjbM0mwg2I
PLCk7VpYzpmVvlDFPdlHZngQMTTgrGqieWGimfNoUwn46bEu/lbpN+3C0ptyUC3Mf5trF0Xq+g3H
2tuY1JkpQvV8gCHNHuRRSZQPqlVPgh8rkeBYN4PaCTVD3oKA1vn/JvAgJtVE2HOcxLgiKdtI5X2r
qRRXbMLJ43otVhjY78aeJUzbi0dJvNDHcOlGK4A/HuS62Ge11fmonFXu4w0aWzVfzLA8QJF1Vd18
ihBI0yyN5lKpQvLz3/3B+ji0NiHDrfy19fYeOpBCQEHN5NoawkVQ9LnN3xxGCyN3t1PEP0dy5mBS
2rkhF/jcoTDtyA9Ja+5EeU8n27jaUXBWlofGS1DUrWIJ/09HAlXT7pGkLqv2o3AhtNJLOQ2jbQzp
wLgVUn2ZmefyrRr+lx2gNN8OOsVksj6HtS7go2MkczgbTQgn8i/EparO6hA10iCs600vttBNu0Sg
10gC1qQS97FVEhyoF87aqrCQBNUNy4H7fFGEWQaW7jp94gPDfKcwBwasSMjTYoQ6XTq5J7swo8RS
UG9cgpko0Bmw2mg/Zt0eBHRNzd/wCod1IVmkWiONB3XWhTp/80xvxP7TYZTdf3JBZFKVh1P0ycoI
i6YjbwkTVkrNU43cayLWO6uUgxWMndGEteu/hOUH/YbCFlowtFQBmSN6FUXNLXkLSSJ8lamhUzdu
r4EOezf/nhZO3RwxtTIPNtYIGrlwNB6EpoejcsWA5c5KRVlkyeMLcMo0+VrLJY7v9xuVv+pA3Fw9
OgY9BEFghn8sk5rXcdGACky46FYl++6aG1o2exIJsplWefAgODK2cV2BAF3lKaQOSnspoQ3MnHTp
OhOa5CFZe3Oz29sTnjYg1cdliUWYZEHhB4Z7ggQ+h7j4oP2Y2+NJV3mYu9Hqafo08XLc7SZCBhQH
C+eX/4CqpIGWy885QWpAOt0odzimmXfWNWRnG9P3wLeVn7dzCQMn016tcTpOh1Do6l8tpxLnAPx5
puH2XejLlzawSOR3OAR/Xj+YNHXY2iJhQry14d4XZXOZuYHkkmQDkib/Z3Knwtstoly0ji6RChCR
Drq0y62YfPK53QYJbLuFaFtFaYaJX/kbIEAtVP7cnpqV6/WXgphgICcGh5si+y4HGONPPnu/UZUK
NY8NtAjLcaaiJ0ng8/mr8bYistxeBtPejjQjQb678YbMaaVe+a3ZtNxkjWRTUEgVdjpS7XcG6UTb
qcUa6CZF+ZV4r5VvU0q1rTXAbGr+c8mZvjru3JS3/JjuntafsK/HBrEDjvvEOwPfieUB1e+l4MFa
Da8SWcfOBX7B7u8fjM8WGRr1bdqePM2rBCgDKFiHn0ayHeii10cN6zYcZM8kEJa2fYprR/8XQza4
4Ty5vueuN5WM0pWlFjyTOP4QrN3y9ryWUd+t8cfnE9VrHd+aQ9y4PLh2yvQ+Pqm1S9CjW8BgxjNJ
i/jfts6HPcgDKQoHkXLV+6JJCSkgbGPBK+rKD9byaNe3DnrbLSHhiXHAcOF8Ospp12PYO6vvO0fM
hfKL2tNtw/dioua97YOIKxz88IW5s/dseibie9LozAKiw2vmxcfwCIY6/o5cYnwQwBZEKV/gaHqm
q/8t6tgBDxvVYYDZK1fRiviHbu024/iZf/WmazvqecPOn23s9LnHxzXQN5OJEtAkjFR/FJTd0bf/
xgtFGI/ostrQjT88dqjUCrLReAbieCdXGzBhyNO0PIHAIN5gYCy37Ey9sYfDVVMaBvDsln9W3Vi6
BOfx97ks0/2GHnmrGQGL1vFf4bAUD1iju+XrqELC/ANpKk7TfHRRfJNduOlyfgdvX2gk0owz4/uQ
IuMonzh6Xb3m1PqIZbTKpM9quhGUplXGZBXsk8VL6i6h/FIfvrCLbhBRdqhI172junIt/dZ+9Y9a
x+ELUhewwVM84SP0O2s881pMkWXMQ2d27ZYGMjP5Qoi9gM6k7Cm/X/8NVIwxj0Vyyh+ru+bjcedk
m3lsXD0QPezuRJbVJWGg4IE2JIBBWvUXmaKVjJG3Dqw5NifLaIfR56wIpbWCgCWLwS4C4/GvXLVR
2ENfe/cN7WdK2JSYu5+IMIqSqYONhWTXsip6kwhCzJpUSD9KnPPfJuj7P2Ih2n4gHskVJRUKBtuq
a3kTvG8NDVFEJkGpoNPejT/2M4OnEQ4503rK+RpZZmqnrU/zKM3uEXSWUD/OwWJdSQn6Rtx3D8y/
JdkS5IDUB9l/EQaVBFVmGIKNdEshpXfIWVvLmCX2up1IahbskhPg01KMVhmB703bJlt0ZMuWYiDl
T/gvcp6DnduQ360Nq6G94MIEaWeFQ8WdYa6rxm/nWF00l45Kd4AImVeandIKd3sbXT1HGnym1OnO
bbSwMa0fHBtkofwEySutZ8c0fJDa0+m5lNaRW1V3aGcJChgthKao8pjYNKshJkynoaSa1Wt3C1o+
9Eh8ZfWYxm730L0f+Q7/EqK3O4xp4+NzqRPEku09EHGqZjhvqHc6Wj20v5NCDuixZ5zgctqkmmPa
pVTBuJ6JiawbrsZIibZn9lRNssJCAiZQozPaNkB8R5Fny3PjkgE3JuiErsRWG7vztMuOVUHbQ3Bt
aWwUutz5g7yOvsiRGTvAKNMkIpJwDYL1dEexqEE/TEdox4mMJL7noE0+hCWWefV/lbd80lN0f5le
MNMtQnkSPBy/SimEZ2TcPwjSYMqq/FxqQgH7LK8aEjqOXvAKvPuP99fObXRw5eZcV8LcZAJtOEEI
i/4Tw6Pc4bhQOHP5DHyNdHytbHyZJkOcTyR1tD1k8r/6IQXrmfnIyNT0sXd/Vn2w6npM4Vt/oeLz
wyrTqWY8zJ4WhrrjfmkbCpUJerrgQmGjajLjJJo/z2ArT+Kkmx31VaiXiRlUDpPnv7j2OE8jZjzo
YtDbjeWmvbCI62PAG3AO5JXPx0K0nNvx/l20PokMlaC4fPpZoVtSzUuFwnT2T/uj54efsVLMKVV3
2XQHp97HKQC+T1LhtVuMZgJVqQP/ckyqabKHDbIWjVSZfnydIz4HSdy0/K65/IXBtrmbzA0fxI1N
/oQPZlvgIs1qnUkVmxK/Msyr7K/uhMeLVBaX16zB9ur6qBzsjWu/yPgjDAE5m9tZa8zMCB65fXiM
iNSdmd6iTlpIHIosS9uWhhJy8MYyGfplmDP0v18EUzJ3d96KHmPFWNfk02V7Md1yFa/eiy6GeHdS
BVo/sKtlNyx86fg3FqQz5qXHiBTBp9AOnJIhEautvznRJ5m8jDhEVvEG8lKQdtnpDzVsouBrhxw7
d/+g3WyDtoqoxrPTvZ2GyxB5gtTpABqVL3G4H1g6dyEOKVBKCPnvKoJ/EVtIhWe871KeaPbVEpCM
kx72tEi+oCkG7EwPuywHSpvgNf1L5ieVdS8ET467LI8LLEPkaZTy+4mBNmwPwMHV1rFjWt0EX5MC
idUrSKGZ7BSADKgKsWv7/gMnFiJE7Rcs4EAZGG6+IPOzuFVgHG0rWr/LJYsXjC28Wf8OeiIo7V4w
IRZKh9zUOrjqopRGYVBraQyar3uT+pCnQe8O37v1ASASI8Hslr3R81Ity2ObdW0EH8v2hTO79k3r
N51layZ/18IMNH8eiMLUocQdQG0BzhV3yzjm5zrLT6Z/J9opgw3bYKexG4BYGNxJliry488HK+lU
nG/NcMDypBK4RjwENcplgWBtorGCFQL9N5W8qYZDQmbKt4CpsQ4ntMaQPHjn1hy9I5lomA73N0Ld
0QAMS8wfIv6mcfjnf2+Ke7o+6q788acrnv7Gwg2W/PP0vJO60wQSrcEkvbLoSFUS1yh2pX643woq
5RoTnlfVFLk1qBujA3A6yrr9n3GtQjHoio5kfjKQhMuVtwWuVfZRgquGC2DDwnoJNTJa8WVqnfMg
4Oz2pnOQZiaGPjI4RoZqF1cek+jdVxTBu5OjrE+OS+ByL9njRyex6GigtMWSTKit/YzVJ4DK1PzM
PhYQHyEUGDPXuorFqtaEPya5T53LUWljLTF/cFyog2zawcvB4pvx3m4FWHyJu8LhaOW/ZF+lqj0J
m/0/G42ePZ1OEwMAlia3AlMdf216eUgz6Y/SRD3X75DaDIHULkjUSKcaRYIczq861wYFA0wlBLQZ
zFM041v+IEgzDeMnvq3Qk3FAlJj4c8TJzg3BqPJzClvScoL0tx26UHi8OR1AXy2uY8ZoiY4klNmk
v98e8ke2Ponopsp97fggqXmkFgPa6i16mcqwm2VmZDWUbHGiewJrskbE7zDl36EjUFE2w68ZconB
18592jcPVPqnf7ppBaTouURtYYTXQqtzIcZW7mM4b5nSjE0wP6VckZhzrwPpAjiQQrn2D7/gvehX
ewldk70hj0osY4w7OMzPh66o2AmgqdHkgNvfa1jWx35i0r45qFsmv0mQVSGJePz3bYAuPrwlUwVZ
owmBEXR+tqQJQPK9iUwlXgQZO0AP4wVPI7D9iE3D0yjsonvq8WRlZM8D84SksAVH+HMpwSbrMs6q
wYBnfXVb8hQqxK22RETMY34YSVxvbspm2l/o8E6qhxEzalx6P5M1pIdik1cas+gvAow2oZHAcwIg
Awb3aPDI8a8veHNo07xWepiVJzHp+ZpVvJXOX7kDKhhNXqZ/eOZqcEM03d04fT1H1Fo4OrIUGBO2
rZzKTzgMmHMQ80VraEvv9Drf5ZaZKj+sNf2gCV37dwURRkoGdqVUXFitY3GiA3CZrSv75VDOrjjQ
glkun1W3g134+czYZJLoJfyLdHuB+ee5aNZI/+NlfOZVPO3QQoOy+DY2lD5+LQFdb29JYdTSyp5I
92atdmc26RaDuecTGtn1Z69cUKOu/0EtHgsdo0uA+P86drc0azK27iz/bFAKYkww3OXeJGgjyAdG
xgFClv9xUA7n9slsLNwKbLyxUHEsqpEjsqdDoHkjoGs3Dn8GuWRQ2hMTSa6aoGmCqnO/yZBtC4iu
TSqLtoMciFxx6HdUmg/GpvklQYPrvYYmJCMNEnhazox89noJD0vtkCFDBJJqeWHxPJZrk1SGBO2e
jAOH1oV07700qFxCdaMqTKnQb/lSiRE1P8UJSr/PJjMqE3xm1cmokcWGU7KXLBeXh+U2P+Yn3/Tg
hAWpS5mGm3p7XoYyX0kph20miDdYFatd+6Ei5pRHqclrutp7k8xbnipv5ohCQYkxlfFCK4HBuF0d
9guWFSPvvFfiHzy5o7LPP85wwo3IhSG/JciR9HhgZHxbw5V3s97NiIl7jHHGedKDs3B4Ld9XtpUk
QdmBTdzHvqcO/MDhAsnTgYXHsKA+52Eaw8IRMWSCPpkEj0OZ0/PBrL2vAjg+72YT/UDEyMKC3Hf1
ULqpk5lPOH8z+21GqTqPESwqmRNhM2PswcKRwO86UPMEITYRmFftbEkATv0Q846/tb3efLEq8ZtX
V63D1zzDbmpduz6Bn+GWRGi6grNnKhBJ0PIg0ir9LkpX49715s4v9sp5Nnlbmt/Avqc+h9P9/oxo
Kt6/zy80KJIwl8ihbIGdSE7qPXWBf3M8ivDlS/91b+KYQCEptFMFfVC8r05Bj69q4FinqpXzbk10
4/HFcnrMXQj5sbgqdg0Fd4YC5hk8lMt5Fe1f21zxfoJEzWQnVLQtfiMWpG/k2Ecu5yMBK38MIfrT
h5CeKUBbEd870zzqXR1i4FjtdfvZGS0qAFI1ig79RLTah+0r32A/kphC1vngOrdpTz74NwzPiss8
IHrkYAPoADByd8dKOuIv3R8niTbe4u4d76C0ElOSb6q9qqzowOCDpckv7JCKQ6KX/8OuD+gr9JCm
pZ0RrO0JKNW9BY5An81rNwhMJIpv5iiZI3VXyp49NuZpYgEaYu8NNZZXd71rZy9bBBkpe8Leadek
j+oArv8Nkw4aa+fZWLUQ2RKofZP7hEnIuXcRRQa8T7Mop9X47Gq4fsZ+S2Jv/941cCs9uhsJfKGt
Og/PPPpQW3upjVi0YmHQp7hW+1rMh49klCTrRCe9zL4N5kQ0h8/SLvz3/9vCYMPQhVFaVxvzIkmD
rtuFHTJfGS/XNGl3sseB/rRijT7RPbj2XhpVzGQbQz9W/ZEhi8aWM+L03OJu/FcWD+BJotirLeuI
5ohDAN3z24NiGfvCyTNoKxazUX0CPGbp7rI7YAPA/Eph6PLynpiQyKlX1qRD5kjv7zpBfMlXmOZc
JOi9AsU0HZQnfvBQLLYMJbpdfUdbXaorqlA8DTlahC9i43Qj9UPWCIhvr/FZnEpOvfPijp4U31WG
56tmeGHwmq/llYwvOSMACnuBACYm11ckrZ4Z02fkeEx0ctcGD1VkNp+6AzhsEcW8tAKpu5BldXwk
wnk5w992H/IRqZbgGaqYOIJQFdNyAxGwf3lpMx81BCv8IU2QoZx+ACXqOxPPw37OCIOdITyBs8xs
LGlUZv9Ho9iAHPACIdtx+/Xc4Rpt3g5wRA8mOXcZpx9MTA1L4kNau/1TtKoB+g+s45qy2HTsvnaW
meIaCImmFyNlDpS+3q2+/Y5HDxGGRivHzxh7JYzvbC+qTEEYbYztTHcEtvahoULc6umclt/xsYzJ
G/tNxFIDijmDUo2It68BMkWJT+QNrZk74PQSPCJUdW7i0DnltPXMQd+wbmTgKbrlKnQ0k2NQAVVa
ru9W4n8VWNhWC6szmUutJitMZKM5hrCntXQIcb31nvMg0/vXgnUfJJjqG3K2VJ1G9PA/8LEtpQPd
/fxws5RUtWpw0U4kgvspWaJnyHJIVB18KvGY2ibiw6WGMRlUlYW9lzmd+WBwPwi/xvA9ufyKjLhC
mJ/Y0Ce2X3d1CDF6Dc4L3+ZwYC0p8c5Zx+kYI/f11ix2oPz00zhjyrj0MDs3oxa/pwZ4ZCf8elvY
PL4yUdSapxIxyzHOR0X6mrAMC6kGHp/6HrGephJef/2JCPRBXQq0UgXfvfMWda4kWldyh41B0CfR
U4QFpLv6aM58hSg7/nkArGIe3gr8mQ8YuJQfDOCFAU+4l9BqXLbN5GzfGYK3S41RdlgASfmp+fJX
hWonQDQ9U+pjju+1Tr5KMPAzRa4NAJSJEkJGY8U00285A8M+hJKuDWxhvQmKxmgIURM586mqS2TR
JpjLBlGsHipOx5CAa/8AP93XkroDoWKNOkGO4F5vvwRlOXDDXWK1NpdoZ1l68TNrrUIB0QlaqKUX
k3wFwUwqHH29RDiWxSI89tEt9Xudsv48gePxnT+3qbWFA/zKXKBw/clgWx+5ihLC5qE+tSd5CFd6
dbZsdmbeRjIdgpbbMYWGHKlYpxsRe7NJy3BkA0ZfyyzGpP3LRPG1uT1dwJEMmdN50qLoAg09TQE2
v5Ku3/usocJsIZpEpSxrdWwj8zPHTABZUbc0Q44WZAdnSvni06D4yzMpUQXil6zJS0Ti2zje9xM9
Ah1AI+x0yZlljHHzUscMDjECHmQM2S8cU6LyxLbgH7R6BxtXHfkFiND1nqYVipk5a2NwZEI6RNXP
z8CBx23hetZUIvXhGDMn+36zTMno1wqO4NikUc/neN6skCHVDJSTzkJAlUVviAcygtWcK/wbVa17
6FZSQRGKAb1Ob+LusqmzTSoMpAmZkX9IpAQmDQda2Rvlw70nvJ6VxvCexQFO/pJUMasaUzUyN+tA
8lo3a870Vj3FtvPsUCfPSm0XWFgb/by7HPpHemrKHWtAKHScygjpMs2N/YeFWZ3NhwB1d3l+K2TM
xxFIt1bx1YDMBIu4y7jeWzmtjHn068OmADRen4sqhdMfQsWUvNL3RphK64XrWhhsdlKccr22hWb0
Sc5OEjcq5hucjFm8VSWfQuXeMjjP+seOXic5dGR8eAacZOZfDapV6ZMkZ444S9WnzTlmhZBJuLX9
e/kUCeAGT03pqLRlnT3t3pbcMcZ8m/VN8fEDXDOirVsuSVSH3QGwOdxorDXUGXcmxIiFYyxuvHCj
OpE5+xFwFz6qv+UmFeypNxHVU0O/fNCwSofRfMBq8NXs34FyHZsw91xxkbPxcDfhp1muXWHX9T4t
gbju0/5taAFBv8IRPZ9bByfoP6LXu4zSrVrNWNZ2Czs2S1dnBAXsahl6TLkByVvRkWRURsneyORA
1DVc9fCRbNi6hSFftpOHxEdqGLgF4N0cQisRNSa5WKPVNLb+90LLnJ04uac/govZpNdxyv1Cy9Hp
22RjlNjD0gbG2naux4YVW3K0KIrYHH8apZ0Usy06CS0F4mDjxR3NtdAkR3o0ZcJnDBEUuvqQhhzA
Tn38FkcWWEgNu1d28w4ICv//F13kdLjzLlgA+D74+X6T+b4NcgtRgqFobYASTinpaSeXv6p8CUGp
hXLoKct/wecBy3OaKgtiT4ZD5QMtejkjHqtvCnu7ptSO5PgEOm6CZNwIT4+pd0AX+SkQOoSAJr04
pmOliZ3arAZAuZR0yn/37+H9ZEAutukdqBXP5QmzOZgcCwEQ9hOKQd0NsImiDV8AKiQDoc69G1HL
XaO2Ysmm+jqVqEZbuwONEXQACDo/2MDHLKtSUZv1Aj/LoJmdWv8QLCrUVIBt6aQVIOWN0Uw0ZcEV
biJHisG+Ij7/3DU2QiHe2yxQjfV5E+VlGrch9xDPFfjKKb7NjA8TUL/1KyId2VS37DiE+b4bwYEg
Jr+h9nFI5J3Gpp7FYTW4D1xA3KodM2yQMHYZxzWTLtjjbDYJgmBqM5wc2TNUwLuKn1icVrsUnNmh
q/bCi7sNP5ejbQ0+khds3i5OYsJ4wtutLst7gEvPDdSTf0o/8E8CK+nfN0ncknqmUU/naQiqCKVU
7x7j12fWKaoI5ompvuW8f3q3yeeVAz3C06iyCKkvcimgqq66ZKe1sUEG2Kp60v8qn5XTVxw0G/T2
8oCw1liJCgISM4v8kJey0P+achbyt5NShWOT3GtSnuuiIzLPTAjruMfJKYqkA3CCc5T+bw+ep/BG
DtgKuvN+c1Q0ZXYG9a/53146EVLt8OEOtcKGNIdRgNK+dJy9cZ2a29WS0T8YQfAlnAB91M3sR6U+
SmqIq0BnyBtE1GLJ7HKXphW1W5KpGHcvU4F94KfuXi99m/S0A2bvUZeM/kIdx9tcEeXbjJXvDyBC
NnLdgdG7qw0mJtGP1UXo35A5VG6HrAS5Px5HLiuVPfoMjestnBHaPzo7o8aIO3gTrkCwpvNWmLMe
lyQfCedaUL426lARbKEtO7JVWzunSR3IlCrc2OWBzD8wVaEyalDoZgsNjYW9Kgyj9+xCWGVIncbR
e804M7uWJGLQSWmwo3EXg7z8/3tIrd5cWiE6OZb+XZ1wYyJ0TfzL0b1eijjeRkMYE+UPR+y4xIhe
pGPQhAQy0UwlKMfMRn2vLXQkOjfxenRFFx4WDK1gliHywg2qoY7xO3bYdb4b+Wil6D1/KvYxiOED
0fiQPs08z7P9TBqjUTHKH/c8V8KUB2am1dIVKCce2idR657fzFfl57kRDm4SJyXkMO0wuLH80950
UJyoumHKnA9kEypDbGtCyE2X1fS900aRApDWX302vzyWxLKAskCsWIjG+GxmW5mkt7kgbw6jJo5p
wr5iLvrJEwSCQNb4Uyu+OqW1M8x11FzHqMyhi/v+QQVNcZpk2jkvhnmeLGNeV6RgknnMDi12ltZA
3NEBR7ZSohFCRA+FiQmngaDgbyWOu38Bc5Xm507rQxN9Z6KipYm5CyuKekIJUPFoK0N/M+2JvKK5
WhZ1dYmDhht3Fqk3pz7yfEc8uVwze6VlO+UKKK5KFPuHl8MmsjHDSZm/OhfKppVVPREy+qLwWkkF
oZqBlV+0/vai7puUfvKtUxiVwap8RHv6picwK4yzuEPYe5hyLqhBA4eQuhVHlnXpF3vTdEBhoTRj
8ausxlNLMGSheawNO+j/vVQaP4a5V9r6k5a3k15UyIdsoYEwKpXknpiGQnPKCMe4oGi2SJhoDhXu
okD7M6ZHVzTkMZNba4p8jZCrXzjKIvHgSu2OLO0qqfaPC5KGjw3jkrK2GTx4wZyc1KEjGGxzER2I
d/A2SC4gRN5AwoGVJ81DRxHOadrgLeJmFQ2ZC6ibpaPb3Nga/SPNHTBwaVkrjYmTQcOHyesvRCCc
stb6SN55uolOBADUpaBFZmSQFVioRbiWruLGTwNOM2Sqo4VkaKVXHnJmV3V6gqrf89X4PJdkhl41
+Haalf022ukKlzhS1QGBIIFEeN360JnUStZQwSu2n/6orgL1nqFvwu7arQm+bD2TiONOBcxX2bUU
kg9QyQoNSRFDf02WNhiXJugLn2EIx8g6/bUOxdktLnPfoJ2v1QF4E4vNKLfApecxchs9a7cN8KRB
9Gxs3XlhoZFVjCHKUasSfn1bVsrgiyBQsPeZ5kkd3WNxjjaR4jHzpVfr80kP0kep6rOs+lV3zW2z
l4muuP9t0yTZLpRgD7SB2146FpTFSrMVjSl7gphN9BHnsDlO7qL7LMW3yYFfhoZ9jRvaAZ0XRbhl
hbFncXjy34NbIXEclVkH7OxJpeFU8fSP7b5EkjZjgTCDx9KBLjlqDACEQY9uMj2bTViyO6sev9Kl
L0H8Fpg9Wy5ihwso9FKnrmKjFj8UszpSTao7UoUMqUFrZWWs9zh5KPWeyGO8waDXY8bV0BI1ndhX
UB+E37KPznf/NsJZIc9MNXJ0mAGxFbI0Uf3a7qx0IldIXTqxgEDh+7LvwLTxDrmNKBtyjH997Qpr
ReozL2cnXwZG7GU7ydsTfEiFMHfiE72w1Nk6RKpDZVI+Sgk/yHwdl8mh903n/9pvP0Zv+uY8JGje
o/c0ddWDpWuLqZbxuraxCezVzo7fNfFWa+chDVpEa9y6uDgwhIKdawlNZWVKK2LnNbfx/KyRKfe5
AvMpa5n3PwJwWEHTk+g4vzRJf6Jy9b0E94UfTVXt7Ia8Ky3vJakTXweJoA2xzA0NJzI6yosHO6JI
GCDd0YdAuSni0O1evEBkVNsnGX/rdOlqfX7j0DksbNApqHH+/zEGba/C92D3/s0Tpd43gjeCIMky
HsTzma9J/8Mz6txvwTVa1RbwlwV2LP451BneCwe41MPJa6VrctgPLUz8AtydQR03P6IbquU5n2DC
iKwRYqCAYBUrdq2N7Zn+t/iaAS6/8QR+esXUfCXd5uNvIIGBZSIhD7xW/oAJCGjAi62h25fr/xJt
lcVvyvSeciYFrjEnRVm4K65c5Qmmv+2eurMincQPMEmo9eewe5LVvrjaV0Hpg/UpsIL+3P0mQ4bE
XlCHFtGeHXT/yxUC+/R9ccGN8466bBzx91Tu2goijRG4mVMXkYnv/JrfKBnobBQVafb53ezc9D9u
3HxSKEGJJBRVItM22+tU+kwq5MMUCsBt03HIk5pOraRPqU3/bn34TmnMDG911sEcCr6eFp+O/oBi
wwOf/NQlrZ9xckjFosgAGz+F2yizXH7P+/zOuTdcWhy/MVe26QA9A34mDh5yzrhXVzkvBT1pI2TB
6aDQ54suQCiprclUwMmWwWEEpf+oxKNgtKtVau293JRXTUt85luoD47oq2WqvXGgK3Qx7d4hGov7
Yv/o4xvBguWewYQG6WNto6oCXDdG19AS/BQzLm+4aHxd24x4S08DZy+plWioW+5OrHARCsmJvTU9
eKaaz3V/vAnj+ECvDZgJpvzNIn65G8yecfj8ZIddPlzvoV/QZJUajz/8++JM89shxxdiI81dY6ic
0LCZrV4aIeOrHcpaQWQmR39ylNCJrKH6C6mbc5+qRrdbIwfPipw7V+HgwruJK1O/eS3yn5/bBppH
Eca/m0ub9vt/mumCktDVfQjnr5lERqg5m/Np66YiLkNngeFq0aGvVko5D0fsYzPMTL/mM2SjPZ2W
dAB9GYbsUtrK7gDQRf1AO8NSFpaP0R0IdhTLWScNQKmrdBIYv4DIxwi8Tz1/ceeL4e417uBHMiKL
xI9fR80+/BZRvh478eWD0Ay9Bo/dPv/8ezsbbjynMtpuGoV2JX20C37mOtmGYWGh8zLDvCRqekko
z0SaElUNsSqFxTP+km4jpVeyVKLoO7MNyGPmSaLoF34UXatBD7FmtA+zATh1wlPpnVNgrzC+jYYa
PwNSTKugXI/dIGpNDgrGYQ4lU/LFWiJAqHC/IIWOTZnMsLOrbJf3w5fNnXwO4cTLrep9ecL0Wjqt
vaPPyPxSzVdkLDiEqipkVJWeX1phYqDNFH8PA6ZC27abmIBkXHkms7SkuOnndpiA7GaAgWcR25uL
DnOmJFdFA6bZo5fV5MMcsaLMxy8rx/hP8mzBQ2U53j2+2jkeRbsXR+2EAJcO4+XGFKlzDTHf3jlz
lgJxjc+lRdpzxYO7Ta97Z9Yfrly5kg9uePQo/aPrq46EC15RPZFctx94Yuk4fGy0A7TjyYb6oukb
DX0s0bQryfBKXGgRXCYDeuUdM7kOd6+Q8dooUFUETD4o5oqwiqS+XcK4lXm+M4/qFnp4i0Py6iK8
Ke9hJh2csIF1mhsmHlSsgLxwLTdV8TlEFf0EY42Q28U8xkT87dLrYHzRuPVCweJRqg8X45J4NNrs
wbZkRgEO969es8hSMqYfrxIgad7Sp1CZnBCU4U22DhPvHV4pF3DpIXLy3DxnRAG+H94IQHwtJVCB
Srgi4UNwulogNVTLQ6ZZs7/YDGTkAulTZV+bYens5+w/C1cwzxAL7UR9wMmkruiROEzMZxvLIl4i
e2I9hcGZBJ2m9ikhb8CqfNQ4HI67JAv0J1O2OztFshUFHbWcSnCYGc+dCWA7S3UPJiQ6iRJxvlD8
A/O/A0RNlPp13hBYApR7Vt3BM3FOJFSXeOpVlTSuofV+WhLdkIGO9KLOxqG4ZAKiv4J9bmAPRlyV
NOVnEJFrbhKo0XaYlliOVVg8v/1DgUX9NHtLsvajEwCm1mt2Tq3MLrMMsmqdSHlo+CAt9O8r+qJ6
M+ZJ3dMygTvUwA5/uumM3pEVPeDs8Y7U5aX2IZ+Cx4D78e99KuNGblKiCGqn1d5JAe2TXPdqm7sJ
vKgYKdUL7d7kse8DSeW3Q48fpm7fY+/E+BdrSnhnibqP0Bwa2G7DKbcXOn6gy6DtdwMK5nXQK6Fb
gm//e2FYtnRDpKswH/jnoER1ZhFXUPM+SO+wRYcl4R6uSveRem3seSNTYFuN0eOrmDDoHfWTGsEj
Xu0r263xkjpmclH2cIhmWrIVIVkd96jZ/hW7nzdkD54m6hD30Ew5aoAvt4dWh67EL4e2dTUdLSbc
3B/bwqcZiz7Xwj+qyNqmFZbXYDt0DLZW4/dXfqTp2mmm+zHDk42cHFccz2d2pMpW+vX37a2hLd6a
BTNu/wkJRRwrqKKC+lEy7W8RTaRMAsOf0MW3uotqZ5+DA85eHB3GzNHoHxiFf6b3CiMr02prqKNo
pBBIk48aUP7ufR6xV+uvCBuUE/9oqB3jHMLzku4pHg84RbOT1jtHZPtm4N/BX51/G8OExyUY5R9w
oY+wFubnacS5qCB37/pflqLPNU7NkxzhTU+MAVNYA9UmCRSQ+z2s5cKj0JI0X+w+Bgo+0LC/1TdF
Vt6Jvx8HI9JxxorSzc7VDaCbUVltQNQMOwFh9BtyMWMh7mvjB/EpNuXOCzGgxyERcgujMPLqpNRJ
J55aqZrveZrO/nb9sjbHqq/0Bi7U9062CByVSuPmze3YWgBTYKeJTQUu52iejwLUlB/7dm6nl4cQ
6reQLijc4IB6sbxBCw8NRdV0rQDKL+9lnbAJjy32d816NLi0MN2k19SIBMlqwSaoHeH5iFVAygG1
39t9cYQNWyXLt66l+6r2dOQlRKOw6Dya3E8FgfVGyq91hMzeW9buXZs3WOK1AbXGLr5g49btqzgT
qte2+2+2JvhMpECqQyOd/PyPydrugTfE2MIBE0idsYMnmbX88E75rcaSzsaBqlh6YxwjwbWkWAGx
le6dmeHnIX7MZODsL43+KhBrGnvHj3YTvZvmHxhGwRTTemhRZaSizlDceotSy9fNph9wq29YGRC4
b9vMX1LDBHhFXOIj8wCcBo7ohDv9eeKDCn4pzKq92W8UnPzej23h5DS1jd8RmRHgcKTtyjBTbKiz
joE+seImbsb/YuujdoCxBUs+oEgA9wQdpnkKm43cA/0lMinyTeJfb9e15OGtCMbG77f1Yy4dApri
cdKkxY9Hyr68CiiGrn/0/aqtS0mrIewdFT8TTNYJnaOyF876vLi0bjx0Xu5o6PGIuuMrr5ahIZSO
k6rYrYwQTGeiEMlAQFirCA0Jl2Bi9FBUKiv5osRpmBgvB9kpvZhTqYy7WBiy0HSzyOeEtyTAR8Kn
4JMqbA//1OQRcklszTOH2sdvAt+i1erL0qzyW0AFdokZnybisVLRNaALAiX7kIcwb+CpZnWPxtgI
Euqgm7Ml9JfNe6tKkIzb8XdbhsigP+F9MEvgCzx9y9ZHTlVwuqVV5CgMX9U5oLNNHP69tfTSVkMv
0QzimlObEru9E3/HTU3MH8sdFJplmDb2Jarooov9ltv8KdYNy9/auyfNG/fG4CyI0G3RaHDz5cls
Kq0M1MaW9/iGJy/NTHv8e+wgQd+ahvuHC41HFMjaYDsevX+ohzHTcr+xARwXqmO+HzUb9ITp0zkY
at+pz2l+89yKU+NoOF1y33K98PoCMbKws98oYgl3y/n0n18F98gWJhz8g67Cm72F/+EwEfzLh7w8
V0QD4+agVYxWQqwJllx0KWS21XAL3H0ZLP7K+M6TMsPjqBtfsLsG0JsehNrgQlxwQeH/gAF08MOJ
n944xMBRLJuZrmDmFRVPL2h9ri1gaZn8rHEIneovUCCb1+cPJgeSOKF3g2APenCICjXPV6cen3Jm
7zDgyTk0b0cJLXKonebRZZv1xnCblnqtTxzcqMzaQM0ZL6tCgLazG4PUxrLzZHza4XQVFCQxfQs0
5QrA2rUb5AiiYXLhrKfzt07mOwrw+t1vh/qhaaYXXeBWnayq8sP8kI4dMaMsmx1j49edmQo5LDac
nHevMHvsYhdbtXFCVot4Up/rFmCNuLekeJ1pXqZ3mpc2NPYNU/Sx6hSVg+3m9Y1c45HbCjcsxrNG
b2cIYgIpbGB11jrQQUOe2TT08yhXtcdi9evY2q5gCvsGhjFG9extUEms3mNBCxk+zk1z5VxALD87
X9031XJhzR7ELW5PM3/S2a8dwecxu2+AIBtV7G+pCxKXx7KGPzSZXApCL1mIc9e8yfQHRbAiBge6
dklRr9iTnqh7W4JeQ+HSPixbDK2OmfKVK4Oc8ZeVofuwSeZshOCug8G+IyEuPKz/SPDDWTlwCtXP
QRJuKWDFDo0YCYqYRqhyBGfq7PgNzfFGtbMnGUJA2IrUJezCq3X7NARN7ZMPLfzB60AeluHgX42d
iDyrovRuD4nRqvyas5MMTMvR8evG+Wb9GFQjbZVBubTHdGenBG84uw+NEykS6l1WOYwzaCbq5bqK
HG3dEOzrYuSc6l+JOtZ075uKAWHFnDgPp79IGsPlYKb9U+ma45c/T0DbtEUT6g+HPXnR/RemoKb3
ROsb9L7a9aGHVy8twoqsem+liDa6Pf0MY32/vb8hPzU9EsyL3E9vpfJ/LU2A9yQBzsRehgwlRc8X
LyaWbFqVXzh7a/BsnZ321FR+oHC2WVEMcFqr7HDaRADCOuvdz7/7IQfsmo+z1ig57So43Eo/3uwa
DrmQzk+h8fgoyJ/6SpLzMpw7u8ZXFMNkBrQmi+A7n6wEZK6WBMQpq2sbMbNoCYt7E6fAQaXblKty
H8dTGMRR8cM7ZsOxV+JFEU7NG+zdLW8Ypg6uxvmvHr7p+94OI3p2bhn4tcCqhCep12U5RALbnI3j
CzvuhUtugS//iz1DruRsc0HEap2Ql7YxhFyEZ4JdmyDgxVfefaT8Y1vjNRzmhXUcxXMWezDN2tVt
o1jJZEjgcVfigSplLdkzEMfCL9nVYKCVqv9I4Fcfn+0cPjNmM0YArORPxNvQtQbUhfF/jOozbPqi
Z8fLuh0WitaZJkXqKfggZ6nBe4kBmSQETTb2Crf9uHQ/gE/+n0sLjnfwGMLXqgbsTCXMXmD06Zbz
ltlvDpJzbnzujfDRS0s1gf6Aw5zGWkgXC1Z5FmRf7f+1OOP+7vLZAuRpbsCSlbcw3BZAziEBFiBz
ac1yGxqxsR9zL0LFwRb8SHxB4YnM43xE+WJjvH8kQw0CbkD2+GLjBMb3aLMEGU4uHrf4bRkmwFab
nPvV2u8/jQUsE63gE4I7DVVSo57Vshf5VDDeMFrYS0El7nAHZQ+X51PivGx/i6drsu7/JbEpHXi2
DwLshUdFf0BG33s0cpnDsHLZJS8LWJh5rG4A8tXDN7IWlyL4yXhy/eEYdePKt2YeBcacJRWkMUOX
cu/OjsvmDFIgzWeIeV9rRGPqvwYvFn/LIMq/Yz1p9a3psD/wVm+HAGgPmgzaPrHzis2LwMPyIS0Y
t6n4UlJqvZYguZoVNWZRf5FutCe5ocoDQDidHvYuUsVnkEe+v9eVJvgIneycg2BhlLEW6JsiKxAC
waGHmOoIL77ebsZG3L5zTaOfv1E6e0z0v0/WmRJwunBN+8AE5WX1E5jGj8FOFaMN+cpMRqzpP2bn
mDQabz5+XV/5a9i8hVq6DZO9AgPidXnVGtCIPi1pDFXCBYCEMmiI4P2LNoXmUFdUM9+hJs5fVbtP
Ksifs+OJbkJVr5ANnmOKEK20azJvKI703FS6gzUuJ+qt/jA3DjxhiuNk9Hs01afEh/wnpMVzhPRH
zcsH1kWb8D6b+8oBDH4h2VsQl1i+ySH5UBTm4UkfeMho7kY5VyyFbLqkhdHe9QrPx/twYo67XMH+
xr0enUbxf0qUZJuXxUr1BK6Y7vPRhuL+5x4T0iLH7KgjHI1V3bXSg+WW8CEUG+SN4zB4TPeNm4rB
DL0l4tJAD58va82mSoEsUDg00vW82SbwgJ0aAT6pIdK0kd/CV344ZOvQslSDAVNglDEM9jQgVc50
CCdMDxZeiaCtV8ZHTawzgIr3bq/2+YG5ERwbiIKflRO/j43iZUH6zWvj1IENoA3+2gl0cNQBpf+b
JAi4seL/upmBdM2nejkNp4lfp6dn1dSEKqZozd+Stg2hIjcc89k+zLcu7AfYlbdoqlTFgXwdatU5
LKV/ABgS8VUoq0D63g/bymwE7TqPxktaHvh1JFFRE9qmCMOw9zbSfU8pbNH594dkMjXkqlnhOyUp
Vi37s7WV4O+byPrBa5P/B1/S+106O119hODKMxLRgTQxs/zu06gbSa3uI1j+Mo1ANoULJ1MAScmc
ls5md+PVSo7hYU4GHFJ126t7zEkyRRTUssBXfOfqlAYih7nJAMdEab6uRUbRoVUNLEsBp9BpH9pD
rMJOU7ijQ0ic7YjBsCbmdcqT68KQQx+Ro5RVYI5OZUXsA/3SWsd105UAEM/Fcqhoa6EaEVLAfht6
Ii7uTnYUXK9glvMInAmRsBT22e9d4a05d6VY/FBiWo7VQb+IE0Sr/CBjvc9im6muuXLetnNQ4ahG
ymeGLQZYOOjTOey8NyX1wTi9o2vWanWaTSTfpxTneFVbdyNT06aDKr3kYSyF1/Uwhs7fX6iwPC5s
hAAt6k7MJ3Xr+t8zEeGGQ/6Cqr3Yf8E6ki6BkEODd40oiq+k8hkKbbjZIRB6g1cRcpnc0TOGYQbe
kHmIO8ABY9nqbBRyvyNvwMyfZUVTvdX3JLgSBcYLt682Gv5EK5q+XqeTvHlttKHcaqG+hprnuNTt
DWPkLN1zIXj80ExZXl225uxh+vMi5/H3S93cs9Ekul+sRNsPJrkf1z98e1Hp8Omau0ixzXWr3Whk
1Ulhll6RpAcE+bh5DfTSZab8IfS/DDBnm9g467GA83eBpXjlcsbhzd86npBI1KivjOGL/eCJqq1r
qbaerVaI0+zsy9OKsgPPUcYv9IrWXVh9HNIRcsBlfOQk1gDXbxxsvPXaqdq4RL8O7bQwuRlULFlG
KhjrpyKiJFi3nL5jRYCvOCcZ0Ynr8hnRXSw+ZKsYQBWcQBzv7p6W3siF3llyQ/iKZpUUmu5LmsGN
f71JSmNVM1UAmI212DddELITR53m2yZc3uuXknI0zikzHyKCbWkf/7tn8d1DjWgHsr01hUcybCNl
XgDJPO/s/nnjnRFXTQAdp1SM9VakVa3JS2bMxRY+2KfNiW8nFSDANa+dj9c78qxuY/0sWuS/ev23
1PI033lScriM4Ux9iunLxoWxLBdgL0/eL4wgbvGpIfNcDs/oqPIY/bhl+vgNiAf1iaQGttFG8LUp
fwib23HH3mym9Jzxh5Rm9G05JXQ1vqt36ITCPcQijwWa/fGeIT6gZ38tPahznaC+oLs/W9xlMYcZ
IEcQOWgY4icZ90KcnBe0XtDa+sud5qLyWjScj+7w5Ot8btdaa8COiA7xzGGRVbb/XLSwvu8dcAIo
YlYg57bgpMzepx1jqWDLllUIg+9aojhOe6he25JZGaMtdTFhBEUTAwBh/A73hLyRQkyhPRZjJyXY
3P4kZvBZQYxmzbqWWQi47KHFIZvVzhZfU8rLSa6DXsYrHeloEn6k28l7U2oJH1i4uJkMGdjefWSU
hJUJ7JsL5c6Q3RVsGL1b5vE62Bgf5rRQ254pOigEnDRbVn0CtwVuof6Mbk10J4hMGLyNmzjkPMYW
IjcUBLTzR4NkhC0Fyf9ZhSGZJLCIMOC1g3nBAYzP+5VUqdhLkBbTSUWBbvHBbqhX7tiPIoLwZEb1
dfW4PnteBlqN7ZOWqCzWblwORr7J/r8ZLfcGxF+npCF5cz5h1+yVhdxyQKXb78QXWRzKBQv3cTsP
Vj9jEn5YIVML9258AZwEHTJXA4xnhnhtsmP0HXjh29AJbs0JvQWfmzcLndLHPYTcuRJ1gRcwr6n/
QeISZReD76BB0L1TogSxVg3xXy932MyFOp9tF4bUYbV/9tfcUMvLL1+D/gQ6Gr+pLKO1JNwGPuUJ
MfOc9RU3Sa+//fGPyGR7gFXdskcA8qqPNqbOZpXntyGeNwHiLXqEJGHBVVGs6RyQX99VedyKahQQ
8g9R1Rdb6+Uq2IZTynNLNiIfhboZUrEAd36CWYYyLX/zTIa74MeMFiGUIWO23EZYG+eA/fDM2YQ/
D0aVZO2eY1FG1eAjsVskQkRM8+rTpUsZoMv2WJ1EaEyNlhZi7A8lAOXdJG6NHKqdQm0fziA4CdTA
blyXZons9qmq0rnpPL46BRAfqGjvYJSw4FzNzzvOmS6NV97WQUfR4urEuJQG6fYFaT3BGlUgg+Jh
EdK42UFpPdpidUz3w71YZbh9ippkWuonhb4Y8r1FG2hye2JlfLIUJVOVXvNcY0QIo9iys+rV5mtG
CnfZycvuWmvMGZJZT6Ls+IWmgnZyGzWRyIn3R/jB+5ET8NlEvsLWKfbka9I0FIwPCLyoa2rnYaKm
pjWMuLaNA10rMjWgkHt7sptGTqTOeDi6p/6Fdk0ZV6VHN0W0cJLZ/xaO8kpBvnAY4WcvrU7P4X53
DNreLjKeBZpX1aSL2LDYA81qlTawksFH2vKjhWpspFx+BNCbzNctyXqowVAIWUptWSDk3AvrC4yd
Vcum9717IwHA4sUb6fX3zJBk6loosX8KbW/ysRimE3H3MdeBz9GqdvhScR0mF5YolCRjicbf9OVT
haevM8ANq7G/UaCMq4gyqI4u24NZDysPb9J6ruglhDnGDcOTQrI7uY31ZyPZvEOkuZbe5nsTmky5
d6IsWeMJENxZQY188ks7JOtbhGNUXk1uQiXaRYUy9H48GBjVm7pmKgsbeV/51AGUNY8TYFStWFJb
b6u47kTJ8NBmc6vGZRtdrhoAJxByVAYWeIZRiZYX7dZQgL18QRsdDo4kEjzHe3JgbgWsKajLXh7I
Ae4a69kuPdgNS1bmZ1Cu2/lqRrIQEjjb1P9cxnCn092ocRvXESnYw4/hEyBxL3osSc+7/gler7kv
QUg376lEaOsWo6WnFpIW9AXWPhMxNOEC7ttgBSIZm+GO1T/bbZAzDTlDMbccvaHiH6Qb5Cvw3dK3
W61XUKIhT7Kd0HD3B6FOHfEYZkS/3GbzuRUKhPlJ2DojeRLqVJymcfGJwgvCEGSKz1qfC3Wg7+Av
ZFyOUxFwU0GPr1OeDHZpPC8Gazc01mfOG7WvT7NpxXUw9lHgc9FiOxjNo2eBzS+q9RoaihIlri90
IhEqxEGEQtAKuEIdesRS7c3HBswzpbkpjdLmm6fLCNrPXtjOqAoX6f5Krgm7MUqbC+MtW8Ol89I6
wVwMvLhYTHLuS3rB++79YHPQmLKs8TZn2dZ6DO0WdibMkBgt69YgLITD8lFB3fpPsjrLfP+tWOaj
TVV6E+PlwshdESAvdBMd0KndkLNKUjYJCjiBUBmG0CCqignC7L8bk2UQ5Xvi/xzHlkXtVn+YiZ2S
Y6Mk4OuS62RZ+JwlFRQcNLZM4bKYzgukhYzUZotgGkV6T45a1dYcsDEFviUXBPeDF+iz2ZDdKIh6
wgbn/17XdgTVB/FVx8UEFgqRLVTU6Csr6IZahQEQ6AB+FeZZksueIXuNSiuNjC5k6ZLnhRFBZkiN
wfmDv8HL0ZxCIYQccm5hEtqhNEGaIIVJPCDXKt/fwmItvTJnbnBgw3VY2f/icRtOFesj5CX23JJv
b0vXbXObrTlfqRlWNFwoQToW0eRgBhQ61vBNuaGCrFDkoImvy24PGkPRkyrQ6UWz9S3FdRBSMBIu
KlO4Vq7BfAcnLC8xPFCxBcHLAPgae3QE8LMVeeL2Z0Qe0wEV+HBVbcYdHVMZB70vAp4/KhE+brrZ
BOVx6bWs6sI0nA5yCfVhykrrphsqa4w1blYwGoDpP26vLvenZCSg1PZ7jUKi/IQ2pI/Zk/O8+wWz
cfmWpbwgr10pHnIeMSftu1tDj2Ezaa8lL2W2iCDgQuX+HMqXW50MF6PXyI+KW01evxm9UTkSJ8kV
5oILasWYAQu9XDxpawtgJX9PalP8YmH0O8be8CdCC2fxPiPb3CB9q3BuC2fYjRMCBfUwFMWX/0Vl
16+hWdcYglsGqUZqQNwEAo7uKOnIKXLTrsoSMQKGRrMbwJ6wHYQLO/+okAtFN6XhxJUXQHLH9sKd
2KJko28inB5gW/DVMCwkLFt0ri83F4Fkj3upYJ0GFO8H5gDXyTFCZAvKerx8nNAZCrG9iV/K2hLO
2K73rRiiMVcBROKF0pzMFl+0Ujykn7vgXB3N4dXoRlqIQdmr5V0xrDVfEZB/drTcDDy4MND2B4WF
s+PfkukHoR+9O/aOGwdKNDOZ2xJreuSgWUBflgO9TkmxNWhb/qVuT8WVEg3FmJNb5SOTyirODEVQ
jAOSb5gzUijXdAq1D4mTOWTxKY/bDs1qO9gf8DDSlPfguTRnpXB5WFD/i0CeFnqlhVj7c5Pq/T7L
J1MeO6FqLAbMvEQodW7bfjp/cst/Jybl68bal9QXtDoUHdvbMnaQqZpfWVq2+NBeVjb7jHFVgbP+
wfXoBQXEjWLSMimu1nByILbqMDHGAhwK7upW3WRkxHC16zMIhzs9uX4dxSUQfruTGnUqSyEVxXhU
QXr7cXWQiIpW62RnxHvZ+vb8bWTLMslUrJj6h8ijmwjrdEpFs4J+4sZ4WID9nMHKvG7bvmoIqNz4
0UdlnlIWvFkWhnJtsbGzW69vKO4dYRUoTmm5561Ka8wCyoGOwsLyBv0Xv9uEwohCc85u82XguCD7
+WkXPIHDVemhRNdzAfYEZa7ztPe2FJGaJQ/xpfG65fjpQoyf3GeHRm2qI6rOxU8fqkdma61QBZjt
T2SUcoo13bDJrCjMJFkfPkWUZ0yadGPmzFIqyIiUa3zqjVoEPmTQEktacjXpVnZQMORWRz2Nss4W
ZQoj3bhXwMhxtM2xuBK6w1huI0sWtsf3O93MufGD9OgRbFl7dVAkudVhb9UuJ31nHA45UqoxSJ1J
dP6I4y5FSrfYAxiYptkGY1uQD/WT4AvyrZKxJLXOsrg9XPb2bnoL/7rkpAjtF+dwHQl/kePZeMuq
OHQFTw8IyFSRbFGbY9DE699KcdgOzKi6lsA3m1wzk5uI4gsy9mFpEhCn8r24mcXPAtifcJ0LjTl2
mmiFTraUxsREKzkCk6pRH49FWNES3E7lXbyWAoeiWzWOuILDEVf3JCbYegjczvqhXDc8pPz/RK4A
VONs4x9m/3kIpDEHh10GVqqOhG8oeroG/9VmEyRg5mQhOBfK9TiW18UeU/zvSt/pkNT7ZttEGvqL
bi5FGrKgaIOlqm/iT0LPdhcwaMl/x5tp3c+Ed11XisVkJjbh5tA+oiXO0MT6dpwx/kLRzANMngAm
SubDIoWdaZAPINI2wiK9CucMJ3ZDFojwAnnLdf6PPrez6uAHLvNGQ6Tfg/tEx3CZXZFB/hG1ro45
hLpO/4a2u9DJeIpF552Vi5jPyC/RgZw939wJnlY/biL3L5MK86GLzN20DPdDD0SNmRQFeTazn+K3
RDbKSNV6cjBNXGyQzztsJo6/lWjVGcTWhfMMLZEzkYYKMAjvNxbScrNspeyc4GeE5xCkiZ23VEcc
q9HsHgFzzA3ZOONechj/IEFIz7ofee7P4E/4U9W9GmcBDk+bmnGNxVqJYlW35yaXE2/CaIRoMBVw
SUn7hJRk90lLhrXbxfWnOnKGSPqZervmYoHWlwV5oRRXWX/+La/BxVHh+SrGLwv2D7zV/YUYjxNR
jDiV+rirwhWsChY9gl4TMY+Rc7Mcw3kbPjhf864uX4H/4+sI0nFKqTMyTImTTULy2wyW6TMSr7wn
OPHmwLH2NeCzEQgqlUiW9hLvnY7OG7LEdQlVsVw3UK64NfX2PBVNYCq5g7YCTS8HXf/il2oZjxKK
+i89TMaFH4pAHGf+V9TGvSAgXEm0kI4qJZH5iAHFgShrVxoUPTRUCNqaLaOg0swgv4gSEixXjCgd
GLTeDidS9bhdAc77I2tykjEyFmX/m7jV+Kt6rYvvi1HptCuXxu3ex/JXaTDvr5e5pdN/qZm4+WBi
ZSn+UOQtXHoO1lxgq6zjSShE+S0ddfYi1VgfM6uBWgPJcRFdfqNQMrYCf6odgDMePq2ya1nSb2yY
MHYk9VnBurMrVRF9MEoyQhUYfGS9fu1Sme8RNmSuCxKErCUiz/rIeMMj/JTOC2i62KDtF43JsSZM
5k5R6tBfvKdGwL84OxElaBJ1STTK3hDqES8Zc1S+i3/8Jh4ChKy98n77eGNB6xLANmrfx09JH85P
8iCfVx/i6hdU44nEFqCmmOJrKTKOR0Q0MGhbsZBEnes2omI3GoJPKUG6//N960kDAtwxOrmn/37T
DsLngR2OUVcPum/RGYm2zkJ/ychr+7rqe4vSCkGOEcKmLlOPdGPkkDFOAMF1jdv9CoLGVS9C7KSq
Caeg2ZDIaPBbEHE6UpSRSLbrKi5JtZG2PLh4eJFcBmYSvegqe3uotm4htznQalE2Vk6B22SdqU1+
40bxgaK5kBIs147FRsWWrsbNIlufYkDe0VGcf8ikPph0y1QNYGQXdTLWAQqMZ+ab6UUrDIp6gnh1
Fuf+0ex0aNT8xIbobeVGDMuWirYvRzjsa+tVafjYnA+bkqC9Upx+6izbCWMui/QyIgqQdX14wToO
eSdtpt4rrrFdLJFjfPbKB46mwglZtSc4ZakNajxF7BdgWqFeUDOeSvv2bjWvgcZAQo0scdMIiilp
h7iVjIF8sWkidq+YIB1qbC0tPEGYwuWQPIA5HS2dOX/7hi6U70fHneP69Z0Z2JoOHvAfb4u2VJNl
RwfvYMVbrytBBASjpql7xf7EwkibqrTIvfAXhPAEQdtzeqYJAYsiHBEG8vaank+aad59nplZEqsI
utCOvcpGLCFsEGoJ+vjvDqIAAtOPIb1BGoeyaO3lmkkeXpd2bMkGFxe7HoWlj4qPr5vPyw1xF3Qd
wolFqA2QrAa/XavVTSag5NCANW9t5/q+hRRLuXGyjzPPpBN9EJvbO5531+jkP3Aq6bvvqGI5WOR/
j408D9Xk709NGDvK0e/IOyMvhxVfsFzyoUU868aB/2VB2CDlAy1/tXDlkwMKiISrgR2xp2IHHwiF
gojxuvYEDk0m0StCuMNo6vwoK2hVPHcgnShGfitDtMjL8w7iyo/h8QrtPrVOwqdTYnCRViA5PPye
qD1GsJoXQo3dsH99+yyy8xDFu6bPufoqTkQVeDlFOrVZFh2ZTP3+8W8TQ0PcUc/Uhah+8vwuWyow
1YXIUNgZNnQmJ0qXYWoHGkLZ9WUSWJg+OjqnRT/+NyGr79o4NEvoJrss5h7z042IBSgKkrIhbrGu
HLvD+APZiCepBuWrH2ifuM/CEStrdYU+sC2P7Hlr9Xw/d1G2zJWrpPBQbb7f49ueIYtzjk9LPM35
6kOjQyE1WLuIIyD52+mVHzqEQlR9fir2eaArGpHqXmEVrRHyRWJm6TF4+VywC5b4QQ4VLKVscKvs
Ilfzk/twQzGWI8OSlrM+K5yit1Y21ImJRxcxVheDfSPoJ91/jWva4fqhwRFIBxu6r9UClJlUoMtp
IVoUPpVLAHqzgWarVHoy90k3FRJq5gGC4OyU7WSIwmGmiLchitAU+kZDxKwf9m+FLIkmkWTKkTF0
c01q7d0iK74eAlz8XP3H4OPIr+rAGUoj6BKi50gnFgbVDjySov4QlRvibt3vxViwACFO5DJf44CL
73/DU0xiHqBIMveqwAoQxxKFRZW8HDyfs2RBCBiaI5+TDAks8KPNs8riEGVBk35rD8XSVcVqcLGC
15IhTSKH4BrrK+PDRn8B1n0JY6th+ipDPtK7KOdItlepWI3Us7ZCKh94Hn/hdtRIOFVklLiV4/+W
BUl7eRYsptq6ysAKOINVzH6ImrN9lZAjBcE8UmhI/9PsHBTLJlIi1EGEo/NQMJ76n4dCAxhcp8fY
XBZcYqN8Nu/ikr2FeJfZYirAFCK5Mq6kUlVebmjWnmwULI3pmVw76zG69zMIlliu9agv4/TnObJ3
dsOjJVDWEW+eCJSftB6BVb2+7qGfwoAaSBSev2KQmwEUqK9V5NCI2mqkXtpCiIgwUepiaMcHhaNd
fNUK+Q6o/+4lufHXt2YCKkzChdSPBCjryZF89iiqEX3QPVGyuQPVbc7DZOsc84UtBeJUgo2FlPu3
lr/xsWG9kmNm4gsAo8O6hQ5iZ4E5B/h5q9Fl0YJXnIxJSiPQKATaoaG8AvWEEHLNYHD+N+EUACFV
SeinAfmJnzc+zLS8nXvHbDj5VQztvHOhMdp8tTGg47IQEhGscucAOcgp9fdt88czXPQ5icX7l04E
zIQr2HEfl+hlPNGm3pYXypAkXpEfD3vwU1gFGFvRwmmvtk0Qe5G644GWQjW3Eqwe7qWhPT0QgCsN
qGKcDbPVJr0B1c+6ak9svl5AfBl2lQt5pujPCLNI321SgMIoydGvh99sprR6l7vCxPFYmDkYlILH
StdGx7Y9MAKJdTMFO5k7HTXVqVOEPr5CS3FgzrJG1IFKyBWa4fi//ZHpEfLHO+54cvliRB1h1MzI
2MU/58vl6ejWvWbtNjjJ38j0bbSuEUeGR7V00XxnM3LEZ1/l9h04sg908AJgtOUa77/pEZ0Z8cbR
WToIrWeKqmOIVbfwv3Ehhi4y5TMMfVrA4fUqyclCkguP72f8EuKeZbWfvEJOPjDOQY0jEourjqCW
vphgd4k6CdUxwzexFfJkeVbNhp2joTYLUe2nC6i17g1Pzy3Mb6QJvigqIovtIH4Rb1ax7gf86lK2
IMf0cdBltQtiDznQY9ASTYwsLkzbTjInR+dK/mp/gC1uIIuqsY0biwQ51BX5bYLkp00K6wEBepc5
413etUsBBEdu07orOzxWeVzha33Dqod6EKPgkgJoE3/OYT1dp4uBykdHOOM+KhsDkL4HRi6GHtZB
mvTW73a+uIvEnoAdtQtY9DFmA6NOAIEtqrGLb12zhS+Zoi0Frp6px/FLtMHHOEOsmFpp/sa104NF
XsQQHbRSxx5UlSlAjjen/Hd5HfzpzafA8IeYrVS8j42kXLdCxqpMfClojgIEyP73Nu7d+Q22ZyzG
4P7dnQWUxuQXWdPpQYd7xiAIqiBlBXTc2JCJsEZfr1D8GYBistuPjjAs0d2jwu43m673V8fEdPtr
cibQUzKiq+rfAIMm0opoG3mf+GQYAToKh9ckvXLOQU5jjimR+P96CHPG9Nl+ls8LqR+TRvjZZxNE
dzkZTOVAUKXl9MMxQJgjadB0CZDS1/DS6cwplN/nG0Jj2nwKyW65b6nJ8OO0jQn8pO8glKf//09f
r6UW/MOqRWCGBESpN/fUs4e+4FAztmnQ8fucaFeCzqCgJO57Ht8dtqQbjHg9XmU1NQ6QUTEb4wji
VQjp/DZ0zpAnV3MlTZtKSGvITGCmp2So6rog+FSzP0qP+R+1iZLgWSLB4c3vvvnJ1me7QB/qsPTD
GBbv9IYlCkDLbdSFp+NLw0+dhWdE2uwyt5H5KbVNjDDoJDTJmFBGHq3x3hEt/muptnSTKjOa1igE
t5YcTlQwg87urFMkOQwth7n0wQVkC2rcxAYd4TUluih0jJLLvyVB42mtEabVHRSjpAhdc7V9VdJA
z9jr01G+sNvPW1a99iumwVflNajWDxJLazBWkdwHT6l9MkSW0eiyNTZtfyq2qepv7Rfm/oVO4GdY
CxprtqinxH0BFChHklBF8v9lu4tIu3kQ24ftQxqYjxr/cGwVBvKk/92ySJ0ifcLyMeQaOCSjODfs
ddfI2yQm83Jmk6Zkd0GVZzcqtpdGyO37Y2uYlbeDRbw7mGKFkTYbPO628MFmW6WRl/Pumg6TURWw
BaQoiEE2WLMBeh2iWeuym/B656Hl1aM595n8wfR8Ukn1hioKkM9Ahj44nV+TaIoOXl7nQyZMiAv2
6/o8cU5R6xFSRrWKmDdVqAPKmoLLizLy9iKtWfRWWHY2W2ERR8SM7SSaTz0EDK1ZxP182lF6ONS7
E1KdfKaCK845hRbkWZMwGfKgMSG4yUT9vNUiL9Mh1KnA54uZue+QBbAdM//dlmayl39ETg/Oyr1u
rR35zKg2LgptVXT9q4laY1g7nFq9hR2xNxHhQg4w7+obKwwnkiY6DM/n653P0vtow9FYdK/jsBQ/
c1pDTUaDCfS59JErZp4/cc7u00SMIh98up6XZpbtn9Q/kplpqKSIwfXFKMZboiPud0U3898I89v9
t5y5HUOTS7nsJwPTXehzBVU2skvwz4fBaaF75nHMoKUSmc+EouLbYhSdPLNcnYVcGEuA84CdFD6u
XSES2HjXCiVAvT47j/SVMFoJLDvwMZwsSozvmVxhl2gLwaPzjuLw6/8F0zXjF1HRzeB1N1ROzje1
/UOdluJg9r1u7fX8JO0CvZugH1pHSL57WQ1EwQQSkaxZpC8j+3RrKr4KyoVHmTDg8kE1lXshiK4j
cxYVoXUOFsgyFcH7odMRBP5MzyMiNtTJ/J8GLErpjzIGrEkAnKEHykRNlwaarSssrE5EBUM6cJWz
ddZRIcSbO/ykUdMLy4K+dyfQ5NAbqRmWiyAgpHLfA6ohCQLC7Y6ebLVarcDTkuqhQcuIuW2ELu+k
w49rvSxDOWXjxnV8T6joVZWfmv9QCC4ts61ry/38X0509anAK9kwe12a0WASauy1pJckvE3sh5K/
fYh7r38iSLnEa1d2EKRhCPyzdjqBy3qwWWELkkq6bnL3//cFNECyuaBJyAjk5ImwKe8OGlDC+C6V
gq84peR/f4bj34hhBdD5H4WUgwyqvMMQrKEQJxaXNbBbChR5gtArSLOEAE0sXu39QekznsqHGH+J
E2XTEwCpUFji2uaw5wIkOZmlNaasZqp3Zi0LWeK9lqBZLuYZm1O0iWPAEbw1RnIqAivhaq360tbB
J1B3945AQIrqnhSwt16KALInvM0mbI2rSMj6/2jOhC5epQ2yfGTRJCrC8ze57S74p7Y+ENH2CVWf
tYgzDMZSa73IlDAY92NqDqVJ/n2y7CsRn+xc1B1NGTkA9e8Vm/zTcLRvnQXIenTT8Rd2LjMIieMk
5rSblKolY2XLgXJas96W9uf+iBjCO40zBmsyHi9JFEesGt5fIMpLqYpcTQw1VMMbvhyBDWoBPAVa
63l1RLiT1rL3OL072Iv0FyFO5cgiUR9urde1d8MzvIOE7emOhAUf2XA8G5AdqDA4yX5NKhlPwzMU
8l75rQ8iy0GwHbqUhu1286KGvt0WmUk+Q/jPKuOmZevFOuaTjwvgaCFms3Dt6doG3bcZ5ol1eeP0
Z7ggiT87IEJJ2htL/WlwzHPaS0zrOLM9BI437rUH178LKbvkUa4If8SSvZZH3pERR76Y2xThFqu6
6AxV/3zH1QuA3yoz/IodUx3SFbBBgOfGIsBhlgJeEUcFgJbh+NNIBcLeQlijknwQ7oQacs9/0W/z
upD6+sZTYJEGmdOG+VNr7NremcAw0XqIHAfPHWjA1A/g27u2sDHcpmOYoVWs9jwbG2wO+jxcd3tp
otK9ONd/FB0kMlNWjMMvLRdQopo8DbjOghSyWuj+9NBi0bN0+11zat9TZr742Uvlso6/mpNt87CR
0ORKFsAfPwGcq1OOamTPHme2fpd+2Hr1FqeTSLPXpH1UZs308a64Dp5uAFLmEK6vZNwJT+u/Vf9A
VrRP697X5E0LgD8WRF4j8TqY4dZ8ZbSmfEx9cWAVAbLRS5nJDD/+RItZ/pFhnyIQ3X/MfK6dbts4
yGW11AtWmuTpz8kEoFCKlfea8ENcNcYqEtseLbYpZer1u/DexEIcqFFTMZoC/fNOMHvHz3ysjLug
bbNn6yLLkJHvIKsN9LDuzwgs6PyDDT9WhvvY1steGxxaKA1yYOq1pq2yJ6ES+bda9vz17dtQVXBT
pAA7OUN0/cSx4ZG5PinFK0bX7+WK2U1XNb/P12pCutwg6iWzc0vmR5oucSUAbH8tcFhqOWo8RCRb
kIxPIBKplA2REkCh0zZO6evhm6Sv6519EieLRXLS+xZuMPYWUDXG4+lBU0eu9UsiSJ2TpuG6xgvK
ZAUkGhK/jO5JhtHnV39hV5mNx6x5a45j0A1UnmYRmlIUeqMIobMpFIxradvkveA/eReQfWHhZrBZ
/uKDDMTPKrWs8uil8xJ93Z8Aaa7MZA+8pGCf+bqMgnFyX8rlv5w2+fVVro1BcQ77ioheer6PcrwD
8s2ErZI+4c6mhxPddgMmlT3aT0M3IYMyoE/q4JNlwQnMdCnJ7Axta4l2KTUrjSej8bz1nYobzeEE
RYLJIziAMCrLJU1R6mhthNgZLhkrZiwAS3L5RhFMxvFXiLsofE370rqPKC3LE780R0C+ZyeI/kL/
BTJzXwEAa21XkL7bfWekSheKNkDp0tFKJSeHKFNzqujd7frCzxsu9FLi3ztUZXNMR1j2ivWwlHlD
JPeZa1+yq9VbnzQgZOvZwYetEkabkihnH0CpHdjHs42n278Z6BzOoDq4HBbHFOc/n/EOl9vHFG+c
mkl4zmNvmLholkQBFx67ZaCwBF1977db6R6kzG9lbE6XCR/oZfOg1lfSUGGh1nf5ieHt00idyXC0
cvIJ24DDsAIAOOH0Mvfl6RGEkIQDJ2PIv5XUJvDieWQapRWwxidBLdbYwktow0nD71fah+YRYlRj
+tjl02ZeZm70WkPveLaNgW0lIZG15LTr85ht8ZLSahtzPiCK7xTGHNsPBJ8rrmWK9wmmMpfdQ+Ji
Nd6idGwts3L6u9GVwHN/7DglBzspv1hp+0khh5AbYO7kMhhjrY4PU6DrA3sll5LY5Zxhp4qdW6Qq
zvnyhC45isiZpy330Ok87Fi6J9QyATAgubFcwNWfCP3UF1c5gLD94JRkPna3KS5UGFlfd/CrTT6m
371WOAmUitx0YNev6OgzQvyj93JGog6W2ewmQpNHsHxpB9WBQDKOUrG4GKr6q3dfb5BSdffWrliy
hoy93PUbMNpOXatyGM9nkDjNBvG2qOiw0xmseTqGOFfQ1Jmd0gAHZRN4LCQlOPMDWXbhUIdEaGJJ
ZCAWN/Z9+nWp04/OWEu9Aw/Z9ngVQaSdSfQaf+ZQdZYhUcmmPUPSRWEENlc3+C0HOr/DUJpptrVk
m0OcZE/+l56C/fTbkVBv/eGGQ9l+vtL8t3yfuobP0f5FwqoMCLejWmxUF01J0POTNSerGMM+Aqpu
T38vDpYFyJqLvt75GitrqyExlh7FQEMeDvMVkuxL51cOt5SOuo++X7WIQEblkGISMox3FMQR4PY+
PmgYdvE4WbVNSFOQFUKwTuy7F9AEJjwVYAWocJGZva4iO2j5tWtNbUP0S3Krgjy2Iv6d4XOGTba5
94aH8HjYMClrKpkQxo9AjlnylLIiY0XkO/vusfaxFI7KRAaoqoAvLzVeaHNrlAU4ajw4mnAciioX
zaYacFrG0D1oAKPnSPmyqpTeBzBgkJnb3YTxzmllGNItPnNkR1W3PiNynMud9ZJ6LaP1L7gmIt3V
R0QjB0BUHPEoZ2Pdocu8nIJ2xoJ2ybRYeXQYEf1bfsGEvOQT4jmOEJdNRUCeKKDehSlAgCAE4S2a
I+3L5VMg9A1UDqxYCGSPH28b3Q9Ea9KwStm1Hub0GsJ8REMGzQywyf2TFjI5Z7twxZ0FWXHkeDhw
jqBG8x/PsYBgLO+jmo+mYPcUbEuc1IsxtKno3JCRAy8KArchtv/56QwngGe7Sx89XLJCn8vDlyly
jNyKiBgSOhx/6/RRmWAM9NOVCvLQgwMsOa6bDwnJ7kA7vqUYnczUXSjkNFTm1Or6BGvxOPxXp49i
ACXAm31FMHOITwulUZ7c3H8P9gk/4dKch588GSoGPBVRxcE3OtE6EpOcBUWtL63JvD0QkE2VetQh
NMJGZ1SCoj2CTYoovW3uBE5ApuEv+/gNOZwr8TuyQc7o6xSWbSs0UuD2vMNXd/hlZrjp4qo1AvBP
iwAkJSlvSe6QcN0kRdHPIURTMzmiy1Eg1C/5JvFkUmUOeg1Bcc/c7eQZOu6W17PWffg4DlU08q/Y
FqQwySOScBynUZS/SyMJd0Y2pvKTa6yJF7aQlTi3JxrdBIPVYZiYNtCwWSpjXkLWiY5+WzZEB/5G
2sj2/6uVU9J8ECgnKhv3QFDRMb+hxnOgElXJkF+Hr5pW+QgFk4g3ElCljiwjtLJx2iyKVEJncD4H
IL3SaQkOjQvf3lLnL/iVdjZWiIBFpuEr4oT9o8i7XhIQEkmL70ASnDHr2mXp01SVwt2oE3tb75sv
nBdHZFvQKSs2/gpe5EpbE9Ns3hkBT19CvRwOaHz2KgVGp5yeh93e2t8jvFdgqNpEAgU4mVe7b00o
K3nspcTYSwyj4jkeK4ixt9KV3z4+g9rT+Db3nfUUb29PpTe/GE4gmVgamwWWnNi2xHpZEhI8uFRI
7iUq4pIfAAW7dfuMAXL8oilnV9qOfOs005IVNtjYItCsmgp7FP8wmX9gyecShW9TWc8BG2bDCwcW
O9HqjVz49EZFCMJuRT+cPRer2jW3P8Gc1HRRKagH71riNhvbFibmKVVvlvoO72te1TivIyQ9dEK9
odi87R4BYTvmzev8X/jbmiVZO3sX5QLYSrr5wyY+1VqDXy6PysTXP8H915BwYk/JSNW5A33gDouS
jQQYpojh/8FQRiQZ/NnSZaAETTnYh5TJHeXz0V9Jnm+CFUmH4vPlnBML3m73EQR29i3RnpiXY0js
+hou/vXGl+jQaLn6sMDkVCDASvZ0B3bSNinYBUFybtidfybrHXfIji3X6a8+QR4NKWoXPryDmWXm
j/RLtPCvFH5NLK4o91kfDzdY9owLrxxs09WMzjfGTYgpBqqHO/PxHtjQBl/TBuwaF8ymGPqLq+yF
L/AxTasUFPM72fdgjRamClfi8zyIBD9aA3pnvGW6OxUlIoBj/kNxgRRcbKiC7v9PeIYDJfRjtQKq
XWcptKjSm/q2Q6y6dpwF94DdeyaoJwGQhazgqPTdBQ9I10Jf5FilUweIQgrqd+d0p7V/gVJ91zMO
gg0mmIE9l1CpHkY6PK+fEOWz3QeJ3/PoxHJDlNeNE7T6BqLPp6VRMaBalqpXbDw9q5lQ9VLdcPDV
gvyBjj1TQVFsJxE99q269fxOL74129bjb533ahH1SwMJhrtyEALxfM+uGD95qTplGc3xcCuQGhpA
7TUvnFXKQ3mFRdCgQ4O9+hUa/v0G4Z5oqSCejdQhI898Fypwo92Ymk1KyKg9nUkkHyigtuz/Agaa
LBCryuNDWFEzWljq8IyUmozCvqeDxY026hT1gEH6iWX5BwPLpZYU+hVeoRgvKw6YvLLqvq0qBi3Z
/bGhL/Q5KRuxB0sJpARbqRskDs6aTGoCPZ6Bymseh3nGKSY3PX1GZ9VAAC6moNW8XehgwITA3/wv
eblCQxrxldXqsXLHB5vPIrTQ9yAA9kU6j2w9XNCbSzYTzzzeXEabrRFGxIr+0V7oH0GhfQ8se9qQ
gXW1RtOLmHkeM4mwwg0le63PHDsjyb3OdmpuZGn6CJaFTLPJXuRvnSr1rWj8UG2tZXd/iapkCORk
4/UlFfxrwjr5zVF+PI8atiDAs2pYrWR0pwhUeJ8kQKgVujS4ubOn54jpqmTFwliJaEaMg2mZmdrM
EOlJvnYisSVallWpL9imZXpkUzakBx/1CXdzsr0gEYOkOz3n0F7SmFNnIDUu4ABLk7zonujWoPAA
uqnYyzsozdeDqV8w4p3PypHH4l/bLBLkMtOoHwvLGEZ++yxWpewvhqiBU10Y82pIOceBXFsjVYr6
/VvoAUBEQd3bDYAZCHUx2ZqbnO4VUBjCHNg2aQ2sLzOkLPmd66Rwtc0/BxlYWznSkrAkB9f3ARU9
HLOaqpuggBNwwWbV1+1kklWn2xdMLWa7pbpQkD2/MES52xb97sd9U2kws3drJqFfz5hPDHujj2IG
hGtEBU/iMGDIjMjs0kOlqfm5X3SbE0yNzYkAdBoFpUHHwkhs2N8QamDNyCtq6qRMx5IFH+wqr+2g
YcNNpp8YJwYalB3XigfmF0jDvgByhPw4ET87FacGdrC509EnauZsxhrS3HAoyajed0BGE3d6z9uA
hUIo4jgq2MYmjA0OJyKjv24+rMJUY/tTx86sXJUEFxg7fFOldra7u9xT/J4OhxbW6cthNxWCPDEo
GL0N4LBsj+Bs5lDrk2mtEIR0sGBYRBvm5FuWbhdJ2SWTejKLOwuOy549F2/ceWoq6dizYONfjH54
+6RGJB8IxndEXnz1qS9I4suhtkDcjIjeioPUSL/EZIZxTSzZSeJRyCg6qmYg2AYlRFHunjdQk37M
k8TEMxhZaZmMBNXfSxn0HDtKufWkpx04U8NINGz2d+AaIvpbSGF9NXv+/a/FvUfyrLPGRAqL1dU5
FjRZly+MYiSFgSXnspcY89GaBp/bcT4g6jxGHpmnpF+nihLCnL3sgXYGq+Hy60yY+iLpSUkOA/Lp
w9CaLnKTlUYXznM0jvouRRWKE5OXMrXmKmlvZSPvncsQjiWzv7dE0GXQcOnNiLLRmjU21nzADLpp
2xxehicTfLUuxa6SzMmX6ZE5SvBfiMmbKMIjoX9Rc3o1H8ye/CkCoeF0Zle4ic8MxI5p6f4XCATm
CtUUY9oMSo8UPxcxvA9bbfB8VZjRL7qxJpU2P9Mh2MVVsazO39Xga6wf3vikxoteSjS5ZpbByo/F
21Cw5Be3/SLVDivxPCBhoYhJQsxBnhooAvJENcN57Yk6V9FPOTC+MLydVwgMOHZm/zXtQJ1TK+Jb
MjdUIqunhvcZtNd/991T8TQU6aljNqiOAtDI8RGa8iG8M+1JWGk0Iq8RaKNcZtIqD88KZ5Bdr1U8
uI9FIEZfQFtT76NPmBRaEarfH2unbo5pBneDk0lGd7OaOwU2usK5XPqyrk3/7VUtmgpbPMjQJjqV
iGuIb/ESAOrrL6zhkL4gmWy7h3Y+qV7z0T6bXcW7H+q5r7uOP7cuGvL7PZSt+xTpKUB1xTsVh23m
KvYXHqGo9+YxZMsnIskAYPjnbtptojrMagVMEn1pbAo3N8NKxZsNRJuNabQPsp3iyFIe60XrigfS
DDFTueUvJi+tSN6qkEGg6SGFoZUgEXIQkEXQqe152SrLJG43VbLdjFIg/Ohiuj7czSPgYpj/+wyv
BQ+nslarIF5QKXTUpjLFF7+qQElXjn5RpQPVeusOuVQr6Ew9GUwV1m34S+O3dMiw346qWwmtejz+
Z6V8pAE2LSO3JVVkdH2RjFT1GyBsRvZhkUju89sTU291BkBTIop/MRsfGbT/ZH/IR9ehwOudejoA
NlnAerqEl/N+xw1Mp3Ju5OTpRSKqzXsBMGHkkQea1DfeuTSeMgfeiN4pyMQak9IrDVQgxA/JrbPs
M+Qs9ePgdm5PjzxpAZ1HpIKrpfI0FOaxVPVt/jA1OdQCLSgcpokw42Ib+qwM0+el+F5D2prV5lMG
+4IxBuBDXaHQScW4yiL8KO+yFg6O7yHilggUOrt1XTqKt7Oe8qCflDUfx82zSlrlP+rkrzQt4HtW
D7Baa0zDw0y1GpB5GV6G2utOSJKdPCnSVVuN9l+Dmo/I4Ok6oYyl3wIGxCeJ9hFV5YuXwTUm8Az6
yMmp+f7AVZsBMuPgZzecZt+suItP8q7TQrDsKVoM56rY7zo2dtpSLCvQmHmudPAPwPnKasBfAqjj
e7EgFGGjcNWOBgA6sEMIvPSCk6okR83xOdrvkjwxu1hgVj9ws6OzyuO4iRGjpkFNMSxzzE6t9wST
dJ9JeX9I1cZxiMz35lD7z6rQ0EAlGvIecRuNtJx516A53fA7Sxqqs+rH+WXE9HNcAY1WI44AFtrG
MHSr8Clu/WRWLZYVU2dV0Z95GTsgDw6wgJvMkjXPM7dB6Fu4goxE6qXUghsKnshrgS/0QCpxhP8r
yu3ghJp8B8cn7E1+H92Qvn+pSfmzRxO/1WHXLDqLqURjdl+b54/Z16equof7mWDIrTyvp2QQ/PB6
oOlWH+hlV34ALyaAKUAip5DoUGahTIx2LMi8U19WZaLrr4U9GZWGS+ecuHnWIp7Vob/k7Q9QGMRC
SxXHohDjPHsN0MuQe/nXbuZK3p877VsHAtMO9PhVQtqTArF5A9/02dEJN7vhMdoKycV2ykZzENvw
zZqY6RPuI966vjkPaq5bKoc5wmuW8RerYWWfhIkSF9G/YZbxrg3Nc1uNst0YPNQ5ikyci1ht3vzS
M1xnyBAEBNk/f1IIn9w+QzpUDKoeYaa41RQUziekFApBIoo/FvZtUxHZXy4F7PJ2OJWcl3DYjcNZ
ev/t4xgPoWqhVCcMS8AxvSP+un9HpExrdY1LccxO0j28Lpnc8sz5JkqshMNVe+MmJWR9EHZ6uGqR
PvZblhQfQAylwOBDhhqZjyRJgfbJZOa7VK7HIeeK2JfUqTlnB5334ALmaoopxMRXrY7NyW9Do01a
FZ4huJdnwao5nEszJhGjQOjQG52Sse1io0lUqoPXeP6DbBaGjn67LlX9YWTwr852ko/nO9eI1lyv
Kc8jp/p68bt/0FISy5CCe9IsGRuv1c6EiVMdJJLu1kVIfmxQdJwwbMO+fa7lqWjwMPDyxgDMvdn1
HF38Wq/wZ1WRUxJQKoth6jMqrB7jCaPrZRzmvKrKePcjHh5tJ5IHKB+x8IfBni3hAaQkkONLsM2/
Snj7egIFIIeBaZsCqMQwax/QWEJ/UwwZNupRnZN5ynD6sqqaASkxeetzR8t+mu/8cV8fhGU0dM/9
umE0NTD7AViNMd1iTVpEnNZpt841FMtW+Z65TUANnfuw+mlaznrl4PSK3xb76kxYv3oq+6ofYJBM
qEstuAiYWmGOiiNqSJkN1LaTmNoQQrJjkJGnfYPc20G31rogYKnYRPuMHtH1zFcTT29WjXBMxOHb
nd+LI3Uxp6REV9fL9Ku9lqqEeSB7PfS5I/Fsab0cjfHZMngyA4NXa/naFjOi+Y/tcjDLV2OLGD7f
CTe/tUNHp9ysYA3M/WHX5Hqb5/+v9YuWP5bvOiqMFO0yMhMUTD/pUHdmTQVhHMWmqypRs896HXKN
H3bcWqUzrT8ODL3LUgAnHpACRRNQVEXicShVeYRbtwq0kdZREBGxpHhFKi1SZtGO4gSpzGHw1/yN
oNneqHemLHPTpn7BdUOoTYeLNrnn/7/MRNeTOerGXsPOoo67//d8pHGVHa9sTs6QJlaequ74+Rqa
fdMIGuouLgGZnvkoWKGzCrKmKMqcWsfNE/n4Xo/sPHD6em7jU8PykTZLKy0/SoRD6BatFSseC3oC
3ydMBagGPZWWYjLpDNgxhiNZI0p3InA1JNcYLQKfMDBm60gKWYkEWV0s6dj1kXMAdZfu2+eMwhFl
MnULxxBjEikIjADcNVHZaVaPpMuapXLigJ4o+ukZ553RiI6wjetPuN3hyTFcfXVPgg0eYLw7nK1e
7r8mn56/5gJxM8ayhUQ3wimG3b6yDFJu46AjF5VgYAma+TxsJWya9DzeRcb4eAVJqqbq0RGfS3Zo
Gz22opvNrCM4a92z/sLbUFGmvMawdvn0UHXVWIqkPvXGNMZ1RmR54Qori12md+PCGpNjSoROSB2s
WQORayzUO7yeC9wQ3BwNjynKmJBdMM9I7ocPk5MKAiibF3rZepx6JpJDplGUWmYsTLRgQd0WFJQC
qad9yJcShCSMgiuGxxccXvJe6+fVl6KX+azUOOgRbC+/gRcyIbZCwBVluK95vjjBz3nwEfHpcVPP
PQs5rh4+OrVqtiBo8/5FFVJoVALyNIFLYtgtJUAGXaNbFDpsNpXGHC42tQB0brEoVLUk0KvYkd79
6ej8GNFSToy1wHlLdhVooLe8GxLudGZa88GPLJg82aVp7gAJvNX+jLnI9rR7ghcD4jnmd+qwRXRC
ZDnToG8XhaPnIb8T26M50GplrejVGkD8JXAr7ob3hXsfCt6CLn9dqAzZl2sABKUsoLxevejo4T2t
tZMr5qfiCln3nxhPMHJxyxim+ecADs38+8eJU2Xkok6b8w6k8/kcWxQt+vyOCNKA1FVwW+495jRa
PoJ87nHS8r5BMFZnyqu5UYEgoMchDFRC2J+clg2qtvv+FL8vhuW60oO3xNbPLRnLCVF1kqHYfj/l
hILEHqFkqF3n0BBqcVNTnBkmbQlCCTeu2NObzKV27XDDeuGU7jYC8AmST1spa6VeMGhW1DdGd9u/
ZhCIoa3GFtjM7PfwnLteyKzSTwoinXo9TOTtJpfZCvC6q8ebQNCYlOgjFkR2S8r/+sMBqq5ICGdI
7zxGvdNCDHYY5OEHcEPdqt7QPh3kZbqtMAqqL2iYdlHnuQcfmde3Syjb/KiVdjfrKvd6M5eYV2jh
/k13juenTBHh9ZJUbfvnvylMoKtYoq2swBEa30Y3ZI53B1lykdgVj+hobRrZFdAlZR/IS90/JapL
a+MM666IKWIdifwgs35O2bSG3vbSQl5b1xDg/BlOkbhKekvmubzgwRt+Bdn2/BSz4hvc7B1fYW8K
uNDuQSIjNgmyNv/73lfjkOsyWJjBHRP3oYJWqhxc5MLV3YHadPnswfCFOjLNM7yxl4VXj7jZlhKI
4WfozwTxwXx2Og1LumRcBSQ7nLlJGcAdQ7cqopOUJultNJiKpw8KRQWGHwdJVrktgps3WiLgt9Do
O3B44kdNcOcJSqMq6qbz9QgvNUnVJ/4qPIQFIVnD/gM75HjcUNOV8heig22pT34O1Vca5VLuKsx/
yhvTezR/bl9sbPvCNp9jJycELrrgxPvibZEKdmfMV7L0ovood/Nrc/knW8poIxslM41gyyhzKo0o
bwkSv5khBICT6wQty+TFypwWLq+jRyJEHURgRQy1h0W/5XD2fu9Oq7koGkcMg546198x9K5vEihI
atoZKNydpw6nPrffyRvhSf1D6ts6GN+NQzTB/c1OmHQPKYm5uzYvF7KF/t+/PE5/X8FuPa0TsXq3
hg2dkG0G+I4ub0mwNvTPXHltOTRJrxyH67w2vOlU6JlTdPaE+US7LKHOEJoNH862Ys/USaTLCy2B
KuzDz1oawTK7dyUDUy6YaxfRowRjH3TqdIPHt0Y5OUPsV0tR8/a5lMTWZD8xqR+tW3ye7YHBpDgW
lQKsYI9aIgrpOs7bu2mZbotoa78+W0crdXshFNZKAFa4q5+GoZFggB+lLEN2f3aZ9qZ2rLqw0TJA
BiaJKpY+4vOY7Bm59JtC9CPMgSXpDAlmS9tnl1THheDQoIbDbAbjchFVbbF6xvnU4cy4p0rRPqvV
Vca966/vTM8djXJBL5A+0sfVTPVdfFIDqURtsqF63nO63avLkmGsBoYvidPSmrMaaIafXGCO1J7y
EpHTZecCXQMqo4KbFM4GlbyjixbscIjwIQqPC/PD1Eo5VTtnDORAR9ijmqFhVMMpuoM5DrOQWlfw
oJdNQGJQzeo2dezRGX323hmoEuMPKGnfMz87gZ6abGjPpwauniSS1rn3G5pC1suLcHbtSwIiGaDL
RlPgK19P0aXG6kgICx2snG8NMVM5okQVI1ykTlA9K7wlt5dWr/lDBivboc4xfuh3FOuLmU2ezIAD
VXyez2DDa/pehrRGhlQ9iWr7VRIBiwYEK0dsuxAxALJ8xDMqdGk16hofHdPWFMIQ/sxWAnQr0kVT
LtFKti+oRCS2jPhkjHx48ilXqPpCmuObhWIQmWV5Rb31gCCCSwdVQaja+5GkUwCc35lG5Xy6NQdW
P4Voj16lfYYYd+liHgQTyeACKICBxWVwO4jxS8JoG9HvtOOXC3XXN1kf5Rm5hS9iblFpXv17Gu64
BrorMqNpjPif2b+0t9k2rs2RMtRjIQpn3dW4BCbFj/d4XMvMwEZDOmNEEsCqNEJDBc8TRSGqBOOx
KE5ZaULaiCDaPJkRyrna8yvZk6G0XDGUvmVMeX1hBe2+1P/Jn+Ant3Ykrn+jTkB8Ks/eMsm+Jeg5
LLrdRk8zUhpqyae6+t0ovs6T1jLh+Geg8jqjrRNZ9ykGjq6nJyAAK3PD8Fouj+tz7oBtQV6sy2gQ
O2ZGuj5ZyRJoK52B/KZjvGZPYu3p/OdQmFcejpUPxcHyZee1e+zDirno0dcblePMHX8KlbTpHqBm
gDkP2A3rOsVwo7kRAn3JiHC5EbkR9H5WkQsYMC4uLjW1QM4e5ufrX72VAU7iJwbhrGScS2Cx2Qew
zLxv666a5L3JRQdM8/NO/sKv11YwLiN+YGecdOmtZPhHAxF+UuJrRX3iVXDwEOLfgrRMO8/n+jt1
USclj2BWd8D4dPVbtrKqyd3LIs5TiuO4o6kzzotudAEiiSxG7JBkfnxygGcN7Y0ietv3FDcaBPP0
lJE4ZsBsjP6hBU/tV1SRk20Ne1VbUHWfYC1RBq137NKTChJYr5XKNx/TDkoEq/IfztUDgefQZqZM
WIulsej9BIthfKFXwjAOgT0CJ/dTG4C4xNFZJ1IOmLuZOtuNaVbTNwad75Ex2Cg9QnvYxfViizpy
fktylyA4gq0NwDctj2DJDpeOlIOSIks6qyVIqnAAeU+5PSuXKN9qhlwAb2Co4VvTKyizFwz7DYEd
Ns4E88UiVGA7Up+GalBNeZHb/N3MQQztjMtvD6u2YdxCqrcnqWB3SDUYY7J5FWr3h2heNLuK3Mue
OSgPmo0xDxvLK5XE0dRybsZLghpRTnEMZEP8Y9Te8yLFrK9oEv/R533l6bxUEuTIhIqaxzfw49Zx
QLdzgNhWtEPuDpOjP75FMyzf98UDV6Mh6Ty23fBYuhBsxf5/ESnR5SKGSU97EoT6fJD8c/GV4Gem
w5UPQtxOqBZ2/bT38i3ZDN9DHGKOzIKpG+QCFWG7mz5SuPH2gE4BC/T2ueffIg6sO5ItFAj4PN1v
q5DeuO2hnB+F0SYHjH1EJVc+JL7bcvZCXCrLZ244tVYBcRKzA1VX+QBVhGUqKML3spbFuU4BObPn
112bOf3Bl30+nVDepW0MPDVKv22zkhnzMPIJzvpOS1PsO1mePJ1NXSsCzao9e3xbuX1YqBwKYGOO
tAPnZfz+ejgoXh9EZqi3Q7/tzawdyDTcUOPZrwycMh1sPZIxIeVnGL0gA7/k6JfXWCjuKbZpJW5d
JGCy0X7tNaMR4Oeaik58mSslk2y/OogooabpbMO4X1272KvzkjgEqIHdzCHfth/mvTxx8ulhuUSH
bUK9U9814zsAv31xNbz/lZEUy/CrsJuw95rQHTK1j0++hdXF/A3+2djnpj8VfdSVWUDr/BFTM5I7
JtpxfAVAFlB8OVq4zlSPVcWdkCwpotvT0+loX8K/gUTzX9c6Ush2NynoqbSyZKjyz5uA2Y6zzz8i
F64WN+DV8w85tKxmICACNHQq4zhDkOwRbNIVoWG4smd/JPhKFFrmhklKVyx/NoXkI20yD54+DyTd
35/2Nn7rUEsBmNf48h7S/eqMgD14zrqLLHaP/oxMJFrI6/7Y49ILN7LXj5evsAoqCFAigx0kbLRR
RtOfjj+U0AmwF2vLwAdTNMWbPARbufCKmu6E+H1tt+U3bo9usX6m5GJjYHKsVVNbG19gtXXAnYWf
oI3FkMIDzCSWY8dqM1eetItRIgvNjTO3y+mj+gW3DF/q7lsnKoCvUJBrbwQNS8aZElxHSSiErDtK
j/t+43NItueSwyEciRjRfU2suFi5zDLHB5mfP0EbZ36rp+4q44pY8gSpQ1sFVlpb8qljorwqrAmx
pb/Ich0h0/n9xaBMZ/DWH9Ey6AVDEhuCLpja9KrnOb7qsiLFjVkXI/pyVnIgBxp1zwD0Yhi99s4y
WhqGHWJ9jVk4EZy0bBP9yiCD0bi/for8W/Bb89OHuatmRdqWIEPT/MBX3puLRE0cFS/1RbOmd9uc
8zwAHwQ2AuIZ4INV8Fbv803Zn9+eP9XhY35HMcs0jbdoSfh3tQOXTMtrJFl+j3CnFQMqh0neRpMm
irkFmkTsymnL0gT7fNF3zAh+JHDZfIZs1IXHYZRsxYNGje7KH1pRqiBF3423L8SsN44z9qcR2K+N
vl6wwtkq8JErrfPPu9ZNm94rAhVCr8gesl/F8a5FOYwi9G49sOgUjKsddryhY/Org+RY364wb0nX
JcvOvLr8tPJ3biy13i27xQyWmaHdTw/18zYRXPVpHQMpZYrSJuMVESVY/a2DkBITf7LKvQhtbyiM
mzDzJ4UzMprqivQ+c909FCiiwBqhnZNAeJr9KdON5b8X9s/iyRsmdpd4FGBontwJ5AWs6ktlm+AE
JbgwM50QoT9IijHL8dIXyByjixDJaq/61k9RSdspfbLBUdD0bFNnmtc6cH/+nM6/MTRynn6/sSOi
7qQtfqEG9XJB6O+nAn60mqIN6znEfPOPuAsuXAWJKe9+gKsFmZ634SWoYcK1mAGi0X+YRCZAmKVU
UjLiGk1otoLQB3LrLbv6UaBifhO6IMc37wGkZllqQ7XPG0ohQAHgZde/7GN0KmM45qP38uUHE8zZ
GdVv/ZpeVOY0ds/bPknuWvmNYPVD0zA8QjIOgy18kl1+AxaZZ5MUSMrE3voA5NATdZNfO5A0aqpD
EUEp5mcDgJ48iXywTSnT3C63lNITS+Sph4klasPytXCIjMfpnhC2hMU0bZiam7fb2Ox8SDGmNRTl
GPcseznDEB7Ya/dKXKv42/Ber/6y0Q2u+hHP9mjtFrjWDJ2BA+QCxaKJUN1thKqGI6ThO+uFvHKo
cxZpai8S+ay4PVrNHe3M8CPjVJKdoI7Fu/TgL3UnvpSXpEmV9Lw+QfALc57/nHJPJkRzOBWq2t9m
hPYXHeuQ/sFxU4EK9RGW9aPOz2BIP3TGiu1QGxnRk6+bn7O1nXjpMuft2L5jHtDX3s20CESAZSQj
HPZ4evQ62ujg8xDaftdGvtAanrzoJbqZ2Apoh0AjcMZoO7Ph+tblDCCLcPabe8gaS6jhGmtggzSb
OAFYCSQyH4DmfMBMqCM28CbkjUlLwt8M/mgLZu4eOGDPREEv/KLpUh6cMGnDeLOMVxRTZt6UmUpJ
oa9h1a5RPuBWcVl2AGQKbr0vvj+g/kI6098LQFyObSM3mzAOFRSIEZJ8i/rFWdUXGynGsCWSsECY
7jOiFqrZxRkZraP8HhqSfCMKyZxlsFVYf26n5ruwiMvHnBVjMaqr/b6njiIQSalttLJ3eO1YjW5F
iEP5tUQZxnL2PGOZLLExosKIG67JN9Wrnf4ajPG+FxIo1BcXSXWTBMYLFVDVfo80vcVSdRFBGCwf
5pWd7rbtBfEZcTuY/6liRYd/zs/vOpREAUjKWlahdVfM9Yg9ru6rHpVQYNAgz5F2TRETG+KymOrP
MrNahpzeyyzqKX6SuGxKTHAvXofDJtJlJIKlyWTf0fNLVHLB18DzR+3dJ5t2ej47Ro5A+JALm2xA
8GwVml5tkbcYf8roTnAJqZRlIWlysE1XRr3lamiMvYVsbVwgo6Y3Q3ILiPDL/bin9ZGv/WofSEAN
lx/+2DCQoh1LU/ozjdfpHpVZXilwoZYAYcJLvAiaEohT84yZlOvid7lZUrAtA5saguqaVcFH9hhj
fqs8bw3GdnlW7WNq7Pr1oTQvQ9sTCd6lWR2snRegHqBOslslGjWyCifB70mCr5qBFnH5Eke+gspv
FcIPi+DEEElpF2QrOKigpzCAyStETpF1MHRe2V5ZM/cfgc2tM8AI6uqWhcfnNeI4pnW2JdVFywZk
VUpd9VuQB9GreLVXYf1J/7S1HcATu8kNkyp1oeYrfbjI4w3ZZgIC4u6ytAqxT848bH0jpKGoykPl
C5zHeGbzWbpxp+M5j2NbSxVm5FMFo6UP6zISIYjKYRv1XOJmwDf/VOIGAT+mT/Rsd3YK5JQioRyD
Mx7l/KzfjIPyYsgNdW5Ee+qW0HR3UTGsfo/f+v6lZD3zKzPZHPYqgXPakq2X9PiNQp79tysnGu0T
SV4iYWECbWSo7x484ZVJNfccBIJWYgQsb+/0/Ts+o4BAMiZswofTkQ1s9S57dQMsPUfFYDzsQb7S
LjUwr1m17j2zjqw6+opWL/6q+Pc+TozGVgr4q2gFpaPQTJ+FsLGIuvklt/HbKaYPEL1Lucb1H40/
z7YDlL4EuRRal71XkvY2provfwaH7jkwBUkl5zE92jM/eFrpihkq5kTiuMmyVyBQkbN1bZukCUzu
YsAbOY3Y2kQgxa8ESJeCkkAJGpeUH65ka+hXD7d8snUdpEQ5oHxMGM+K4nk2uVwpP3KGe2IHWPrw
YJp4d/3i3D8aXfFfJ0fC4MRa8NSk6iIwJuMGTetRGkFXZJAoI6xfmBS4Lz+PdaFgd87jxOWxmBVX
Al93y8c6OkxZWRuvd9esqACIufZc5AiiNPvn31fspz+uTaMZHbhIpnAnXnyTSHE98hFAB5UYqZ+R
cNi6/8YY/2TwVadCtDvgtPVCsx64lfX0Cirao6YSXuRJEHIgwa/jMh+pKxiKcEWDTDWg5M+1ocrt
pHvAjvzNQ6JBrbQ9m6FTaziCA8i6AMS8T7FyU2QsOoR2O8Yh8YuBV9WLUcYbhU4y1jlpC/+jc0Im
si9p04BaMTRlvOMOccNoROdJ/GZvIpNnH2RgCRkYEjEWapuNWF21LBsDuXs7/aRNZDr60jWK+5l3
A0h1PGbi4BWTre8i74uf15wO4T71tV+FJVuI3yR4aTyVsyzo5wZz922R52ir8t7ILcmkbs07/ChH
vMi/Nl9KaTPAWOBYfN3j96enTpe/P3kQHrH83QylX1YWQiGx3mzJVj5+wVzrrX56khEAqRySEose
N8VRcrrm1W+u8nq9FXmMjz3bpWn5/KbJ6tAG0h9uj8JAMhwFbfe+atHjzguYg6W1zriIoEJXD+2f
RmQ8PjwW6cVsFr9gkJHUGTj2oMumCPbT8yjnOUuMpmV3gTXQHHrIeKaxD537xaM10MP/zaTtTtq7
+xC0dnYRKDzwDAsDZvlzUzUomaDhYZk7B790tSSsazjO+cD+lzWAJRF5wQ6HLF6v1KlCdQ9zygGK
Fjg4Svht7fjI0mokG2rhLn1pg6JAtZ5w6vgPFVK0stV+/wCyNw1KwGCDAIp/TjRKzGDLStGe8LM/
s4/3o9bwCMOtmUX17UkpS3hY9snFFlCnDM1IdKN0tLm1xICHoPWCiKcmbRiDo469ARoL3f7CzbgF
+Kxta3ZpfQKmFDFSsq2Dfjz3Y+rjhN2JoWAVRVbpHrumenvzAfyX+7zkIM8hdpyXyFjIKo9OmWoo
2frCaDjK6xNeywY162fre80V9666uoIBR02wLUilinTrnPzFTKTKWV8SuDv0XdWCKAbJN/BCACqv
xWFcfZ7bl66LVSxNWeorVegIwRfuKUD5xgnrZtYPPom8FiZ9r6sOIvV9ihn/VCJ40QCO+oho0b4E
ERCHDpc0UFBWbEzetDldLazpHjAt/2j1FlnXmTEcvJgr9scS8RKL673ZHUO/XO2NlWMDSERGqezV
aGSxPq4EI2Tm6onXPbz7uNnyFdXcN6H23HOz/5mkd4PwAKiBfUgW1g1CzHUcef0nNQv/OY0uSJCl
WVy+asw0DXuiH8RP3p8Gc7N89mjHaqQofy4Qv5oPrYwr7e1GQaKlncaxm0l8BLEMg/4DoEdQ3Lk9
dWWSfR1QsSIhyp1LStXiMWglBlBumpUzq8Ks6JVjCc4e7nb+suSzkX1RGf2LCHtSIaeyCw5IwzFP
cMSnLnGRkW0OTKKCVOakFgK9DOknNGotONkNv6gmjrsMhMKN0kHIUpbGkNu6KM7U72zB6YUhLf0J
ydwt5gQ6RyG4t7Q6CMIVsvDOd2cimNUsVB8ywq14+yaOuM8gMrZnAvwqN0KBfvSuPf1pH3HyF0/Q
tgH2xhdbiTXeP55vRXv9CvR+wiUPgHJT4CWG9dEaSA6qEjSrpx76DKRh4XTvzDXoQ7QooPTsIPyg
AKXkK7EaTVD9zskdf1XCblnjFoHi6UMhlO8sY+Xnlc+RkchwFAbth4SLhYe0/fN4uOyzG3jKNaWn
c+BCk4UXwCrBZl+c5l2BZmXwn1i+/xbnDcawpuxuzsqLtyJs3511xyMvNWI+8LsfPfxDoW9lNlj9
gWHYFqq/J7FmQIN+f9ikVZPXB5Vhtua7Uljo6/xBKVmNM0zEADaDj5miuIdRKkXfT0jlCS1o6L+Z
xWarwqTpOhXWCyLWHVhPifixHtt7aWBTZOyNmrCSPzsxF7J4EwOerhD0giSWby5zrHOiDJZ1LCxX
prWTcldS0SZOeHh66MuLBxCj6mMcspb0vRPrJcT6YgLgovj4g5irU3kqistxPFXSqWZ9R0sYbhFB
l3zYsTZaEX4LFv2l7kjE9tR/iDSITLt+ORsOi+1XLyhmlXhywX9M7A732FfpybJgIvO+xOvuYDvg
zVH9ZClvmOoFl9dPBBvmU+Qdof/dnvPI5xhe4pFrdE3L/0AAMdZL/Qwkbk9/Bzj+2fFdcK9M4cTT
VzpvE/K1/sKuMiNkdWhZhFdUy+PTFLz86JQ6t/8aEALHw8pkaLeTQqke1b6Gv0Gy8SalxgNSQ0vh
P0yWTmw9OaXScmhoNOdkZ8JzKCdRDIhpIXg/3Q4EAqE3/bJVVaP7ad5D7WZmf1znsYteuDgt0SFs
Iq8crEpLVvE0TTdsfHXgUFg5NFmYB9QV2zsVWSAFEs4De1UugyO+6OHwE/dE9x0pZ44LVQro2OeF
NWHFg1esiShETHY4PT4W4nry4Z9AwlB3fi5pjozpRn8FP8wFS2Fo63voLgFNY/9BJr5Qp+vjnLZ2
IELSfJw+aPIzTHXEDn1JmYsedMymxAmeK5lCuKmtvKLcYP+ZQIqzJ21M5RLVBYj0MSAOGm7XXX1n
fXSRXDABg2xp0zJS6i5AhDJq4DACt5refwz36g1w/E9Ct/lglp4QPdjE5tYsDzIVAdPOz9vv/NVi
8/RCnUW6bMMJqIjdzp2oS4aSLAnupOV65aA1V4t9FE4BGE/KNiUUfghxXnXjIDbRCiFp0FxL4da6
EK/u1hwCrc8K4wcYGV0w8uxP7glbwcGy44mKBhmrArN3hDszcOrwguwIHN7nSgDEZt27j0WABP7x
VkXURKdpanygq02iOHVQ6rk46GHQkk39zGZdSZJ7G2doPtd5p/PZVCm4oQPNdH/UK6AJAxb8R0AW
zdi2ws5vkJq4gj8a2comAwrXME3QSHrTaiVl0/zg0FzlDSfSid5I18bUfJNTzrmk4LGTaCUCLtVc
sQe/QY8DjRIgQj9YuYfdRDUSvzfF3rRwjj+/RoUqbu3GBsFYQ26HpfpzDKvn/FDkgfMy60k15IhO
cUsOQafKyW461bqob1cjjMZqLHl51B+95MLBiuG/im/HyD7hk5ENoYaqV+pL5tQTmY+hTShjIvdt
mAdIKO3Uzld+xDWKIDzaGHQN8tc+PStMgmgOeRo7uV7w2IRZzi0FyGF1CEj/TX4oK1uaqIEYlG01
y3niEqSVUHq+6QZLVs/JYg6PL71vrKY4NMBfYE8BzCgLEHHe/TtGw64FlAJW0TlYOPr0lGC8b5uZ
ZQbvSymtfUob1J8GRyA3x84mmp8qM6eefNuvtK4GMGyZ2f5xPMRb6hoNxBHBkYcSVUm1+ho/wDa8
7u5iVOcCdwsKYssbXBglHKy/L2C9afQuWZVdN+XUWUXLZI4AQDozuQM2Dp4S7QTlD2j7jxMLz1wl
j6SnI8rD8YeVu0y5yWNChhLufmvq8kG/z6y66M4C39nh7eGjgJxXNGlK5haFHrZndF6hjv+lO3hO
9AgVMK8JDKIxSEXA5j9yVJFCSdayJ1yfrpaw5Vn0k3grXVgTw6/3swtgNr4R22qEYB5kzOPvvZzr
fkJPskRa+pP2EZAmuh0bmDjKL5HcOHAh7JKTksMdCrRghdPaNegSQiWfqR662UJjkhqsyWLeNbqI
UH43DIbS7lNEMMV2KlpKIa+WDA3gOXpwtt2j0V4xnOYFqVyJ2xGVzXes8NLsL9ei8onNhBjhvf7I
KWbrvTPwm6hHTogaQQo5LJ3bvWVIEDKZtELlyXv0aUhcqpZFeNuEfn7XQv8TnwzcEf8mV5Q6GkuO
/Bbh81bbzpu/gddQNpkbGGDZ7pB7w0hu3/3dk2AjIP3coMBSf23uOmS2hYeqEU8oofFJnbs/krB0
tFgRWUSmYbdIa1+cV0nYYbqvTpAm1dWRsuHN5D3+kCwhJscuzR0HUKJvvJNAUHkSuwqhXFfLKgU6
FsvQHf6uAFUQtAAwScomklVOXB2tOg7UASKM3c4MVoBv3jLfk2mR4y9JVbNVbaKigxhgzvRSBmxt
oUtvZkEoGxcPSOBfa/wQeEGamC31Tg91m2gs2G+4FDkZAC5HiVCH71D3u2INzfWIpJoRWWOZTbv5
C9wG+EfN3CRIhS3MnrjPEzY5PZCs7Z7Dsb+OW9CZQyX1SYUJ0Vha8OABRuZbokijCTi2VpL1Et8B
/n3YeFiVjIL6LViy0Tpm49TaZgTlKLuDs24ccQjM0Hg1UPlGc7ajU/LI+279zuzYtCCpK4qpobef
U53XA+zWGbFMHG7AFYoYq/3sfYmz79+vOOsnxZX1N/YKSLnfRDZgRb4gJnYjZMQytStJ2ypdSfJj
Shskx2X1hz67rwyVyXc1G7ewItrYLOpE0G95V8gQ4Ep5rON8tGnTqXTWoxZP4gk1YfbIEs8GsXxY
AStbF53Z83on5UUjKsCUEBLz6pag6em+r2hxjwpWXVgXiQ0+8s2UFFRwsr19Hdz8lq6lK/VKq2dB
NwZndumysqIPFqo7pF8sXh6UKsXs9s4tb6WMLGgIzU6svz7iaqwahESvkRgTmQ9kFhnitRvkVJO2
h1o0LbFkXIsjzjGw7hjB0y2oDPRT8HHHZ+KRAe59C6Xxuman7Q4eYQdg/ZX91wtO3BRLmoINYyz4
1l8zTzqmi3FMwhn6wM49tDvxD418oLkI/komGVFzxHBP3aK2ZbqtUJOAuDDAh4/St0tWv5YzAJbs
f2gaR3Lq2s9BcGmAa0BS/jxX/y6M8ZWk0cSWjoicJgg4iiec9TB4ojoJWPI+3rF385AL7Qm3om6O
A2M/Pgo1NM8yJeQ1jo4ayGla1NlEMGwL5lGtqkSX6GOMEt9iPSqswstD1NZ0DDqUuICcw2Tejk5j
fMRO1O7cRw76QTn1/5DHloNmxt4iQ2d5/ZyFZdGpO0W3ztBSZHj1ztskp7m1ED2xOfC2dyTz4v1N
CVZcjjB2i4TaOD5rdzDue5cBENngUPVKan6sQ+SCINhhaTxie9TEysTa8cpk1pssGQa3SGe1SU0a
9Pq08/uuTcJIYTS2jI8pslgDI0qI2mg8SywLf1zW4QlVrspHmxshzdL2gLljIhdNYGxZE2+V6uak
w9SIbDReP2xHZ+GmS3V3st4z2Edd9WJdLLjhCpdknflxl/2I4/v+8bV6yRQcRp0Brekr1BNMijuV
d1XI+MAhM3jjaXh4EqrO/4PZgDizHbm8yGjV1ZyVzaCO73NJe81HZVeB6BGZWojW5JQPexLgxASL
LQNSTJzCvMaT8ZXiENlHLsSMtb/7M/iCDGfE2XrOPMQuA3rc9gzSykabidTjy+J6xU9Mci1wvjHj
6G09HBwHTQ1LgdD1+MykPYgZv0SExZYv8yOpwA7HctkfqZFnjbRBCyhg3uRYTn6CIKsEYcyTORPS
9Jp//5Fkaj7Bdf73Rb+pKWUGOttk+wT/vqbcgjHkMbpyVGEinerNk1ESZKMMa7ngoxIXNbEWJdET
aCfCqTXOXjCOGrV+pb39eO6Pv00vtkB5K+V9DJ3XkI2XU/qNPBiMFvME2wSdk8qWnMUG36POPjSY
LM+7akyubdnpNMcEzJiEqXniN/LNH3Cp5+fsMM+8GaTQyplHpMUfLgKQ5owszdP5y8ZsSvZA/nLI
W5PY0Jfz5xZJohW0o1JUK0GNxF/ycTjQK4xqyqmRC0Xw0P6yENtVozHwhyIp7f+1l6/+2GNFmh75
Q+Bisz509gk4u5R3wsUrE8UF7UTk/X1TBGvDDQp5YbQUAJwHBfhfL4zSN/p0pgdvfLpbjxiExKS5
PssOfkzVwiMwydzEdh/Eoc+gVZhFN68iGYsqT8eODqaQncAxco2Ibw9BtfjmE+Gd2HUnyfuJcpCA
jZLHCI+qWrSdDnBEM4octvMRrH1r6JAR+/2P/bMW4uV1J5kg9+iWhHB5msALuKy9GXKpyWUXM3Wt
ab+PcUDCNF4AkvXzRz8wKH56zizAg3voiOyDqe8Wxh5pPcfDzCsEjAu0677TYuJeG6sbSugvFbQH
PqkmMxceutM3SFEmCAlUMln7uGc1VZmiFNtjyUUzV1WZ5MrU9/0hJHXS8+BJi97TzsRJ0gQiQoWq
d4XxFJq9QErXQIDB4R37xhG9dzpBftuDTV7uIVf+EEZiPyGyJFZ4M3LwMMwoKDlZGCj+mdfcL+i2
0+mS7jF+D2O6Hz/XbgcJjZMhxEh2cyNjmSaqflCDTHxocD2hAWbDJFjEAbsonKZH46Qfg3bzNe3M
R5Q8Qjz2H1ODwvz5q84YW18cKdGOP08eHH83p/QocRGEfxXyeP6WjbPE/96HAKzAoUZ4pD43OUnI
QKEPmb9PuE3jUktbY/EbDw+cJ052i0McQyU03PrUEoA5CCWl++hBGQ9LaDrbOK5zh1nD7zAAnWtv
gfj5Fa9i6Ig5m8vBSyJVpydCyR8s+EVrYEV5Cp/o73mZic4szfJAViIi/Sc/+jvMzapAIoMAGbtQ
l29FsVsBNirznFfvIK4oqXefhiUWQV47plEyZu33mV+xaAfXdleSHIm+AyRb9N4qsBQGBMh1H3CY
AVbSldnuA5KkE2gVtRMzRIJXHxIH8nmyi4A+MryKWHi9y7DuX8ACIR3NUh35joIx2pOCsbdemngd
W5UYCwHCbvxoIKzCLzX9NYaEo9ej/JJHfLQ6nZGAFV+rNQpDCGO+o0QOpDkrw7vvQz7nEP9oeoft
xcR6XIFxNs3TE7qvku0rNyfEytRAh709XB8tEL0QI3ZyThBnr4vxUkReFIMIlDnBDP/7wQEUq9it
/xPQpbR4+2VLh7RIQx1Lpga7Zg3AAiH9nKgp9FqwG6/9sdsz4RV0odhnV/g8wejE2EYyMwQW5giR
9Pao2Mz46/xKu870CgYcXPKYzwdcmhgzqW8+3/OFNJQ2f4fihCvDMSqGy8kE+TJKJiK0ZED+P1Tb
J57Glb/26VpPsH2k6pT2SqrenfxLOdao7TxpY1U2aobAC8PFXqhkTd43maGERS49fy4p5ONJt8fh
HbBbqTiIEVdTHt4ntUUh8EWQqntKfvj93qohfu3SrCQb2ICVgiINexvC4ayPPjlmsikxF/9sBdw9
yuKX8Jg4yoYc+AOV8EEEQGwowiMeOmY+KE4nQcEe/flUgzAcdbzZ5k9Hi8kyN4ub1NyfPkDP3jda
uFz9DA8oUUcm8iAp6iR5bGAF4epqOzNcRQGSbOXGwFuRnkg3N2sMKmCTw7CrBWHw0N+hdvZtlwgd
kTxtwplnVjDU8Z6peLyXhjFfNMk3/qfJcSMbfbT46MSv4yGqgSIVBazKDzjY5KY8RxO8I7C4Ys02
/XftUOqeyk3qivkvKDZqhPHJOiycmQOQ7E5rrP0/zA5WPjJw6mQNvJQuX90NUuY7kVJoD/Tp8bpr
0Wefg5gUjVru/5zJX+/WoV90aDgiTP4IwcV6eiyYSRdxQCxAAo3rJtLk5oEC78NYrbk7No5ZreSG
GeYNiH33H/wg+jEZ95vqFSeUcij+2atrth78g8VJyDpfeMgQbz5fTEN0a6leQzsEDHt46UvNiqx/
ZfpxGloQR6uECZI4OWZCP2YFmqS02+1GicP5Q4DvKOBp+MOLDrLmYbyoCqEJ6rxuVIqVR7613h6b
WcCUQqurj/xhRkFNa6hC+k4NQXfkn1YEljLDOzCrrmn22eywEFaG5wEGNoKu1IQE+q9BY/a1jMMb
8LAh/omuLuOXbpe5or9brdgjLk8gGIuvBAtBULpVsaXKrW+yPzq7Zmzpy6R+EQyNeyzFrICJB7LU
7YA3rwSHhKpxKxXeb3LANQFLkLTSA0Z2EbZVkWyWQRFZPlzA2lvm+YdoGeZXsNSPO8Ig6ISQ6MIh
oNL39yCeHg3z0dNa232ofZ6hVck477o3tgQb9UqzFwCUVsBopdLiOVwEs50eBH0MkN+odEMaAjnN
HD5u9S4ppYPpGZdymtuGPNfLKfoF+G7eUxV9iHU6PWPkSqYKzYU8WmYV+xuAyX4DTQSdgyUeiVSG
QwHZnazNvNdG6czi+1IC9n6MLoVFcqGa8nYphHU3N1sLza+srx3hSt3cWe1hYTsU+OktPDEJS5S5
PBNMWtF8PvfSTYphmgcn8ndau60b1XZKL6B3EyyFjRmX0L3ktX3zgzbpL20/4USDHaD9lF/B/WOw
6Q/jK4F6SVhwg8lth3OrYVb7emy82X5155of/a+Qk9MRZXtQqqRqchZupN4b+Qicfca01vLpyMze
VjvidcryKtYoP3s55guPzXt0QyEGgBtg3roAd4o8VaIhR9EfwCJ2ZjlNbsh9n2W0Ugqs4+ZjOAuD
aePNzmusGbJPLdFTagxz5YGEkFPavWdR7jDm9sAtGuVSJVcdrIUWV9/fX0SXHgSI0Ml6h0st/MMZ
QxENMeh5FtEkrDI9LLH2PhiFzOyea7H79if1E4Cqv9gsdsX9WEaSoOcXTVfBqnAe89Q54snFO+1W
Q+vwWD12I3Gvig9NxrsBaDKnBWrjB8wKzqM4Q+GPN2UQhUq6GXTgYj4M08IvDhWqiBqJnqHbRwQw
LIe5EoK+POVRvQmqd96JrC50ORY3B8SSA1ii5h/DOVs6mQb65++vHyRDMYY79+y/btsvC9x4cYLl
mLR7HvLD0s0jlEGPulGfKPNmVipOArcS7EBSVgyRZGrlA2twj6Fu+0eKYcr13ZM1y0NLaBhkKUMQ
EjWb7jlqS33+0q2KwABVBlVMYDpzlSrEQYCihGFlMjnnnX8X+W9F4Xv4PQCBNlXYvLmCcgoW8SrQ
jreEcJvvC9tecTBMyH8qRTxWc5nFest7AKjFJV7VzIKSKt0Cf5CFf0ECjhllVvkovRvqcmw3qnJj
wrFoDzRbx03WcELhNZjuKUpYAOFyAdYP+DQ4WygFrnXUtqdOChlNH9dRXi4pDUwaVo2O5hYm7QBn
leDQwaeruqpIHBrPKzmVYR44nkGj8YE1Ujukvhb9FGE8M+Cns7CJdF42iDosOLYYjbqs2tVXiQTi
/IEUubG83YgRyK3nbrDzwP2ozEKxgehSruNNbCCVxu0ks8nJvwSpE4DoZRFtXV1IODj0aXI5fG7A
1MJJ4N4+fqyCZZQhWnlgD6T+YDhYf81/l6+snpn26AmLX6A3kD0XBUZ3yf66/nD33hYbcbS/32a4
4vPlW4J8zSFrig5aJ6hPObmIt0jklDzq4ndnCgkVTk0rK4D/nT1M35ZusT9sQycVHhCW7GmQt41A
om2FuTck5HTCGdU0ucqs7NRcpFmqDKDmOiGSJp1NrtgbgnpPVwoUElKBSIOkLn84qedC8IOjhUvt
zbycmx3XfWxtoB4lJ2HRPfJDlrqvfvRKfIrdjisorCrFZBLWyUT5frtHCbh5TMTBuymPLsjjHCsj
vjl1Yiuxd75bfu1VeGybM0I/gP6ulEKRhmtD/Kt2hkCIdh+QcyQygs1q+UBBUwPs6Ph1Iazwhu1Y
Uzj5q8yoUCgMVXQiavqsOIraMnsK5llRnn80+as1x521XK1UeCBA4cge0wB2/pTa0x2k7spQ2upq
MecE0xxLXr8dvvBSrBWDIY/oCr7Xu5EwERv4zBgTUAmCetxGEGxcSEr4BgtUCrvV4deMLW55/8wP
KXYwbARQETX16JXA31Dn03ecAMDPigj+5Qz5TdhGpwpaxipY7RuG8DhzZYbMPbeINuZmL6PcCJBT
LgFZcAMHbTFNiAN6FegkyGbnMVv0RR8vP9CKqOFJ9bY/J07h3zXfMM65APFNzBKHkfMcFsQkQYZq
NO0vWd6lfFy4szEuLc7seTLJwYnbLgM66RWFrSMFNlXyLceV2B7eXW1VYfDeYPJQh0IeFcVwVr7K
xEq2gwnnYw7XCTtQVbKq17kRxd/c4SM5Iq/DeNc+riq8+X0xzkejjXSP/2/XPWd6EevXVzHPA1f1
TZjJiV1dNcn/ph/zNNfBPP4ZMnYFKKVtLzRi6QiltNfUAXfgicq0pi3iYKhknEQjjfbkPdpRHbpz
ZxvplGtNGneGIg1KGY59KlSOouA+/k8SMI9NItk5Pp1cfqzKkFhhyUK4hgcj6iOVwm3xyNDKtkPd
vNZeuUXv/HQOT9CvRCdeGkZHe5uptG/TZTxdgrWhE2tv1UZL35/D0Afj6c01fW/iSqr3GXuFQVrX
ZlV2mSvxzdhMLQuQdX3KQy15B70fT4NuArkKPoNZGC1JMGAhxao5PxzM3CVnV9nut3VgwTxj8Ij+
AuNCGqUxh+qSXT35DEGPwA7+Bov0TVbHRjq0UBYl4fyzORnA/AYbv30YnBwViL2eI/3dA3hxM3YH
eeTSlVDDXjr7CPwUwtw558JvdwTj4TQqJ3bf4g6SWBvFcAnAck8h2VxJ3rQGE7lneKJ6YjcVlH/a
Nre2NPIbCiAE7ca4LpBrfILUTvGXV5SxvzUSuYeyU4fg6vL0zookrZXqBgPPhd0+kxVmtCcYFXGO
iPAgCagOCnb1XZK7SvEbETMkyqMWhc0/qwXPpVOGDevNogLoHYHFa7T3sgfxM5BvCWJsMsz06MkU
OG5WKWHMD6P+Q6fO7Hray+gw5KMwQy/5+fth+wCgyTRoBti5975DaIXd2m97zDbQzm1QgOWgRvWQ
2y/CMFnsFga31hPd6pL7gfODfldA6n8z6/gFQkyoI/JQKrEGmszCA7rlZd9ilYhhzZcbrceCg+0I
cRXXt8uHKA1tIUerVSQwMKV+Tqd21JjBp0NIM2eaE1Ja0gSKaH2MPA3CBAIy63w3t1XOxK2Y2xTa
V6ZZOHRFJ0SfgpPQe5Mz5O6u77KCmwh72eRgDh824YPNJOkoQSph62SL5Nh3ECguKJvcnhDWudFZ
frUevqycdbCYnBqQDnOGySM1jkM4pRrw9YjVaMjno+zR5hhusql4MZfKsBMo3uIXZkR/slpTC3Xf
SiDWzAC7bDb3g+8BJK+dCHZNOy1l7HCSVvSSSSY/R1+Z/+FiQV8Evko7Z/sFfLtKdthXJT0zDJ+a
KGwwbYBrkzK0bVCE5cBuO9SZqX2qny6POKgqM70zz8IGTGYiisIXommLo1s//KEronRKkkjucmtO
v1S0RDhCLrpbo4oopclXTxv3GiBusNShFQpwEuIwczCvEb7tXX8heDyhgMBJQ6dj0pQ5tRJTPmWR
LWog/dTTaVOtC4NbVZwNfLtzJlDjxo8nNLi2R9XiN9tBjMM/AhHWEcCpnUmB69mNnGdGUvFwmhYr
bXG17uiScrzleZd6DwJrNEdlkyDb3rAITjKfOltiSXhjS//m8+S0dTIgonZkoWsDUM90MxB5F0uP
UGoJga1ZXbRwGirsgGiOnAqUa6OPjlv/GijhfRaG45ydL325IF5xnpotYgvJXwNQVcnhrYQKVEQY
PylHoKcJd5eciOJi4+GlqYa8quOVQ5s1NZwWbbHBD0PMGykyj4pfZUVBtnhDcvoyupLAne5AkrA+
tzwzxuFpo53UO/bSAxI0dyD0FOef7Rc7XpEHZvNO6DctK6dxrFQixsiA4ifCtl5fKlTJjAhsRulf
gDlx3lBKI/diS5bs70BKVQR1UR5dWwXngq5wQ07HCLl0468prj+kHThFBNuVvVjEVxd8Ee+gwruT
59Z17TBA/TyTTyR38EV3okOJ4ISGKQRj63DoRPa039Hv+pMrzFtsqljtv+jDuQU1mibZLeJli9dt
egaMryrfrz82DQWEKKOvmhO689o/RIuTjFVxZ38DDEf4o++cLhhS3Cp1pl64yD3VGsrQs0WIXyYQ
kzNeRgGknNAKYV2JSCyM6uV3c8h1nQfYA6d1rvWIzV3uM/f4faoLA771lI5J2Mua2V9s5230IzzX
SV7/3m2CXot159x9UqDVZe4s0Gs3Dd3vCEppOxusN2JZuIEHz5dneh6bbEw8/iD8HTSS6kfjOhq1
5/lIMgvSx5dY+8xivSBo1sXSVQHpbGUx1/24ce9wll0L6HGnkyKin3ITFoZp1/9HQjWrKaXkRHHn
esWxDISi/UjqYS6wUyY5CmBwu3UY8CmgDP0tG7xLIU11H6sLkcIU/WEPE+KAP+nM9c4NKDzNo17u
5QNYR/VnPj6VdtD0fa8yS2VoInOBgvYUXMw7s+ZoCsCyAIqETlyd+PKHPaSIILgDwtIgSEr4LR0k
+GBUYTgCr+wN8PIn7HvVLknVw+wsT8sWxRb02FlMzMnyiJF/W+wp/crgoIwmmPvadse2Qa4rMRW9
lee6gBX3eW4tAWYFDB5ZARqqX5Aw5aTVOXl2Odz+uPWThOrzfe25xCZ0q7xCVJYr2haPyXD2A2BI
fN7Ov6vQp6rnZXtYnDExuPVSRaLOcVVTux/dmWX9k0GfpwbVO4LusCWxfNiy7gEeULVRc6O/VW0w
+cIN4lCc4vWRBAdwuQNaKQSYAf9qxrllnMCeU/LNabr7/B1sHOFhwaUzdOAZywtmeDogfhWAn3zG
fv0nRVCTuPzVhiTGFmU595uc2+taliOarT0qS6UsaY/h7FThLpKsvf2qTSUtdpIl8+33XaSRsqxO
3Zemw2aGuRuhL42c4BqZGTVccr+Wir+rmm1tVr+r03yyE/kq4RC7D/oEyTX2Pj9vN0WsyBMOW3ii
tTyefONjW2t1L78gAY30P0oUtCBzMOfmAQozmKliFoBRRn6KgiL2pDD1pXy8YS6QefA9ABHj78lh
+EvdnEeLndJN74EXLylisvNahb+IllHoz3MvrqkTSzHO7Ymb126X1maGyhpqpz3KBG5jGHQC/lcj
1rHzr0IOHvypqOtWi+Jedrjb8nggbnrOm+kk/TF4Du0sVTOU4MHjbJqrW64PuiDmsVDyb9GTYoeX
Z9ChN+/6Y2BM2HzdQ36YCYE18vZOnJlqzyzF+qi+HfC0nHlfpqmSFMoHj1cv2893RLRlWejkGa/p
74pw72pGTWcuti6Ugi+U5cU5fqroBtfnifmDNRPPzqpBMv48LoYDiIaOv4Ab1769w5pQp6UxRX0x
3E8ZddPEEOXz4LHC78lPDRiS56wWcRE0VKQrHO/5ABQLAl2m4dyHRr0Kg1RHtG/947DSBuKgXRwe
A/1JCJCe5alku2t7tlRJ6TYoHdLJFwa2OE0qlHsX0Vllbqvg1l8PX4M3npfw43QGbJsl3WoCjc+V
UZbVM/MbXaA1zF7D43bOXtnTB/Z1mFYlu44OhpJrkRrRXkZBS/lnjXb72Tg9Kbf6EkjIVnjVICtq
fxBLti9W5BVZ012REICTBrcPzzB0zQ4B1i8eXWOkmXKbkqK1UFKGHer0XFXuxNp7FvFbAT89g2sP
dINQ5ZYasSPPmHV25smGgwCQ0loREkZUR6Mp9vseDe9yyzVBueO4zEaWrSAV9z5GpKyPwngIYxt/
detqHgcFlGhIyDu8/bACb2tkUAOejTMmTQfaXHVnZL4v3l5SgPGcf71uvri4nA797Dg5BiT4ggkK
AGNKKqtI3sgzHXlqnon/98XlrYUhSQKAKAvWG+Bs0x5gFa3EuQy9+8F6y1e3JoCTgQWWs6JZqVE3
zPn0j8trpFOSq12npYnbZLfIoI/JyQA0mzHKJp6F03NPN0XMHxT3Kz1qAgstDRSyWzP+opIptrJI
oiCIac1DD8eQm468BvYUkX6BRQFg/468auJyqUaLe1h0b8gUk+qXTRJbMklpajf9c2fK7OjfQJsa
4rdHAMVSg+JGpP2qEnR86jSlAkdgPDFnVsupCk+jxtLBnhRXMmT/QH5oS6ReQ8wWA1jPWxXHqEcD
UKxP6Em5Fg33UJKJceY+BcfXb/iB3q84+dtYZdNR66R3V7kJrjWZWXtiiKuDeSTGHxRkN9i3/nnf
E1c3xmn7aTU3i24g08e5ADCsYFVAQZobMCFjetUmf1SM7Sc/YXKE/v+AZv/1ntaFExAbXE/GeV5J
SF1rniay3yX7GHXPIo43cQiwdPVfcdEsyr10FE6ruVlQUQ5S6JFGVh4z9eZ78YDn5ewmxxLEuVYk
LltZXK+kSjr5YTUPI+/4nl9l63/g55+8KdAVb9gHSX/FmeA+3TNRTGsy1YxiXDUfwemAkoK4/P+p
dQjS17bNeNSVWzQPHrY+kq5EWpvEXc7eAIQbsVEQmf+5AldmTQdgaBZ4F06hz8ON5l9PO20qTEix
ZEtea1Fx1v8xYFXl+27ANYoy7g5IwFuVRlD9KnRO0DPaj7QE2fe3aAwMpmGvb6fkIVfo9RiqoVWk
QorrXqL/LzxX2SZhJXajJLLu39wNtNZ+omP8BYqyO4me90ZBP9wxqcT7EyFL1f+3KJd89HzsxmR3
6/3VKro6WambVSTU6oKXMQAEVN2cuUOieEWlxdDRw9+V+z9nmoFWLoQl481B4voSSgOpA8Lbkqdp
vUHG8U3JxSuxQd+ENckp4fAMhSD1B19h35izyIg1wbwfMrEbjTFVnQWrC1HvylDx04ZmfVYBiIqp
nL0mCGsYhs+JebTY0rVxd7zLWdT7TM/DNVQpY3lWmY4V0CFlZgxataFGhCCRKYgmybcC2YTBnAUo
vBdqunGjw1svd4yDdttoiZcdA4vm89qc9C1/xdi17epslHP7F8gRi+8dYjHCv3b3U9WEeDfc2NIE
bsNsthAu56XTxNYOqcHBHisvJNfqab3KJAzijrqofnThAedElaJBUmx71ZvkU5ZMGqs2igFR22+d
BIqRIrSArMz6IiR8EdsGvAKyKJIQAz9vVHTz8O8LElqd8MZiKeuUjsT99B0KSH77rZBUhlqXfUbk
bJbcEOwrHVubpxrZmrQ/MFFEjawh6S+VMev6c1iP9zSXSSogrD2RG2lK6iHkEVJ2mVbjeznuik5G
I1GPN7ZggHi8y41vdbjjftzqij/C/dCZxpktNC0Blm6GXrXkJtq3mX8nPz0M8XugbmrUBLbhigmw
JzzBgEI711REuiKeyv/YT/QOl7AmlrDdUVp3YWT2y1225zBUHnky7Ch17pwhfioBWjz10hU7kQuY
2wQ2ZCVbrNu/JAcOUDPdJNDeFSEHrhC8BwdWtTwitZ6kl82yw68uQ7mzepMnVybTfZ24Bc99xf1K
Bb5Q0JRYkRhgsuBhnp+o1rk4pNQUmA6lq70WCJSyclYWmGYsTFM6F6aFVyNMAto4YjJWIugu/4fO
cIk8JsEDOehRDdriKSasqCYvBdsDKGRt7IaS66orMawzyM8ajJaIojxKrqzxghXdk+hRzWUBMnnE
owap98i0ShbdDphkgZObkEqekBC3zT8Bwwx3bSA9ABIt6YOT/Q0KRrRjTHCSEDctDcEqr/uKI8Gv
BtTSQEAin2Fkyu0wffXRjdjKCMDCS9ktmbVf5Y/C7uVLH8o0TfryC0ufZzA9IfYEGX+kA/0SJTn0
GB+aIYgppTFBJ2DzpX1MPCj2ysS7N6kfq8nASO/r6ukZS9G6e2hTOeLdWOkcFzLHyPzZGRXVhlI0
4dhUeOdaj4TfvimelIsG9kWpbd5DjZlbtO/xB71Ouwqjquuu6nFPCTJu9TJbrm2kQFYfQ6NhkdiO
J4kzJCgBnmRHXCmsOC7SAI8CgvT1uNRR5S99CLttpX4jheAdMLJyYmbY4haeZReoQkjyJ3JywFUb
6hJIMZCjdaJJEwwMpBzAEo3lDAf1ryECLzeAhPvJgrdnfVqfIJji3gqaa7GmZ0yTD5RkcGjvLlDr
eI6ZSZxhuKMX7nsbuJsgAeVCVniVXAdi9Bx42TEbXrXMPnyZx67S0msPYB94qZ+qrgn2uQ7BU3VT
WGBkQHxL3a2EEBty/Gzxz8caS+KmWXhk6hmX2S+wKMG/F4kyYWJDLFQSWbrAKSuK2ipY4lMieFtd
hMBOaoTrdp7wD6hAkRz3HYO8X4Vr9KcZ6j5rTKPWczioZKgTPKlpvFyJjpO+M0qq078XI3bcyoRC
N4y2o0svttLTjzd3+p1d494CXXUPpEP6r0oROUO4oWHkhfwBTnJs0YjT4vEUOSln9HTT86EoVR1n
VooTvPVktQ/eeYV5ZSr7Stw3No3QA5v9ApQsobtRfunkhMH2kXPMFhjCBmXCnothTcCugbfxG5kb
h3Vn5/7ikfY2WsXc0tMo7mwlhnqy/hFSdgglVKqam8GwPppqRZ77AJrTSRaBdVJJ2Y12Ad19m4bR
/QgkPS+WfTg/d8j20qk/PsoZL3CbP/vcFbYlnwAvSSvqpvP9E5xe0YbTZpJ9KxSTTDQBN0nI/W5V
NZI0QkITMDtPexZmu67Lcbm5/UFyVyhb06j6p+h1/UK43zFupY4vtEVYL6go1bw6QPSd3GcuGVVP
tkiGREE2Zz1JiwarV6NWEEdMH7zM6+Hx/sCoEnR6ddTDzIluIckmjefPQKfTGPz+1ALT6YFXB56+
P4C5iVKgQP1gVtQQD4zTbf6YrByogS5CUK0Weh1zv24x8QyfT1U0JlwL9DVFGks36iLJAHQIZeHL
mqVSaK6a5Whn1+1B7zfN0PCxmawW8znOcPoYKmdnuLShH+C+OsPlTWKRK6PVEIYXPOxAJqVYIDtR
VBFff+OxQ9H1P6llSQIxzZzUVTcjGKNK6Gy2i82YANzxWgek5iJ+B+MWkyCvqfmIsDsvKTABQI7Z
i0zJ2juq2IXSB36oQG8q7u+pAfW83Rui87u43pSxYKMcUhAI0nDqNuxON6gVtnh5eVCcFdcjBKWg
8+HAaGHWUh83OZIEHID4m7kfd6oImdtoU25j7Sy3fEeOSGZrWgg3E5DhXIxCsq56/KdUP2Fn1mCa
ntpYzS5J6KSpRD4ouPU+lGz5QV0PFp+b5567rtJgOavKk6z8OKamcNM1U26zI5+7txpoXuqY6r3o
I4iQbDu+8raqBO8z8agxurOcT89F0TLrN8xogU5R5gvLNNbMXk5Q2WZZ7XmLJ0oTR53eoqHitIaj
wLDt3T7DFpxhdXE5nPHYcZXPQPb3wZxV1gcpi4B3eiQ8UtDSw6SySufYT54gyvM2XQKgFvlvwcKw
1XFx25HZ2em4KOUYZAxBIPiV6L+tqEiT0rdBAKGyTO/qLueGhlCgOyAg2VF9tuygJKrYYk0MSWAF
9vWr7s5WCPFf43tLOhz9emSjPomk2+eNEEhpLUVZNc/YWY+hV0oi6JqknxFT8QmFS9sSJ9Pr2bvP
mNeZn1y9zAVYLvyFWSqU3Y0xbDcghVv67xexMnNWP2yoZQst8cjRPeiodVJdZ5ePuAZWjqi8GSXo
p4VXmeKepnxpAvENL3MvF7gQz2DDWx6BiJKC6peqRN7VWp8tMqLSBo+1GkvPn13JC0YGv56DxjID
eR+nulIt4L1KqPtXfZU5Q1Uj+WW2ri5acqthUjI3eUFOsYLfpFTOcnSugYNVe8fHoHWw+UtXWecy
zHTVL/XAY9wstl4jduKR6Q2wYLRgLHg2XyqUcxRRj2Zvycwau492zxv7/AokEWEszzQGXaIxYMG/
OgJEP/UJWUXxJBSIdOOqY3LSZcpJ2EGMLPgem9quZAQfca6U/vDb5gLXXNHmRoN8GA8Yyyl4S96f
fC/tOvKgUJ5IYk1oWM44QUCPuZCiKr1Zd5KHfvmouUAwO9ElHbAgd/Nrt84D6Vv4uCtU+y3XzJeB
WqLBboqTONEM2YciwNR3SO37P77FrvFM4DDyB9d2Q/vy1lxDSJ8lbcFsNLzWwNOq3REFLRjzX8Xh
AYQVmBnFfMN1Fc+cp42XFhZYK0OML7NKdaKvQp8olcAZu6g2c5cbM+xfrhsZGnvVa4S7XRB3JT97
fFZm5LGwG4HGIOaEWYPbRdGTqrrwJ7nFWic3RreIOj73fxHlTE0teYirk4wo/P2uEKJRg8HrM1UZ
saaZnhXawX8Wlwv3MpSCFJ3SA89QQlgqo+TJOuGZ20ZiayhR4Kddfh9MgpzXBSHsmCCHZXtQ3OtO
OFlw7aZKStJP/rcAohyRxftnUBdBk4ROY6tUD321ajvt9NERd9D/fWBddCdgScKosVmg7By38VEs
WSiZ1m6H3T5fTM0f+qjDDg+KOMWn90ezFl/AQ2Bcnwe66pNsXJYUFfjWN18aQTiGME5uLmUQ3j3T
krlwgJ/MD4TzprBAKhJYd6IoQJ1wiuCDidjipr9PKZCWlmGBV9yz8NA6EUEjUM0VT0VATcHiS9/Z
c+lgCQ5dJkzaIeTxxEYOxUYArYdjc+8v4gM21HnTmdM9qMm5v57l5l+I4PpqFlt4yBxci4tQHm8b
NMAHeUeIuT2b/mRNnjwfl+Bknh/nJdlbcYiY9DAoCDXHh/DcLzM/3gPt3yyDIG0HGF6h5e4UV33p
ZNL+pN0w+kvkstNqjoeGx4HiaRyrg6nK8jIYX6U3j/DVnHF8oTj7OTwn4KX787Su/jIEYssWpvvH
30St2P0gWdFADWzC3mYXhs3SGe7cbKsaWuQVfeIUtaR7XjZ6qRJUncbnAXJ70/oPjzUnso88YXp0
QvcJirJUwfVHi0EFAjfMsxvWwM+gd3RnLWK21ZgkiMib0YaG79oku7YHgounDneIDRY2agI27ODV
MoZrRfuOQralI+IflpvuFUnPlIZDreR0acrYWoEL9tDAdp1QndlHrIU3F6coqc3DSMYfebBVPl3W
jkkvC3PJP/KxjGyCzNeN9IuF4Glj4/TeHwy2i6mIy2hW268/gqJmNX7LBjq34hQUuX35ewQ0fBpX
j5tqRVpKCxFbVPF6EnI2MEJCz13Rii/vLZjmRJQL0MerThqSoeroChF6tqDGBT2vt0IYj09xQGPl
430mmMZNslJ78oxqpD7liTjFrg7uyCvwCk/MxId61Tcfc+haF3FJh5sqkoJYm9DYy1QdSlYQLIM2
BgtpRjmEbCRoFvW86eeUdJb0IwK5OE+SYJkqZnvuaN18QEmCxe+0zEWkk2y5k9t0okph55dp6UTm
ISrBPmy+Pi48zevRS4wDrGZhH+4LM2vXptVkcREE6sZhrm503uXwBjs7xa+I/XtgN8oJUs6Q3mWm
enViX94KJvsuxEGc5jOXPpnwbVgr2yEZG7vDKIGMqyIKc3C+4ejtOlZx7TLp0DQcbE3IyNJ3cpZD
89aI8cSHFg3sih6HElffvOO2C72i04gWp1bxxYj5kbsGzn3QRDAyWhuuVoW7hf38XmOZECPPG09O
EM/5cBBOsQOLj9PZc45uLFs9MHAy57uLTbtQKZrXSbX9cFw5rrFl5DjtKygWZja7qpEHDqwHB2B9
yW9C3uO3axaeqUTI4xJrLw5YnZYl8UR4if1W2OKdbRVbZc0SIW0nkJDhbv4DsaBhNBx4Ls4r5/aH
88roxTEg+JpgB6RYXqOck41Yb3B2eiLVD8UbeFMQLliDjTH6Prh0lEtederU6oGvyRhfVsYET8yz
yiw/Puef2AGDhfw1k3o26giAUeiER46sDSnNNcctycl5wxzXCQpFrb66CoSaZlpzT2x1P4peSolF
LLTNUkLX0KtKwDboNWy4lOa0hgQANVOVZ6lBWJi5/1w/Z3ZPtuJbfORinYeMUTkBuPUzwKlKD0y9
DCLcTI9IXHdtIw1zxU+mLpKyMogRzsJrLnX0+FTHf9qigP+qJZ5K/fuCODZExZ2BMdsHSOXBzsDr
huhXrjw+hCbm76zP4NXix6ysZ1/+4yI+egL2OW6N0QRSxwo8xa15GtAuIq8VekAPFPa+Pb398R/9
uYvy82xot4Pv1VtInhLmgm6694SD2SMpSvKtsPo5bvcPlX8fWhnMLinQMUvwVEqdHWNtinbUFkEl
0rqlp8Iy/g1KR7E0TD+2jrZCQAEVXtEph1hi4OYjHnjaaMaE+4XBBYQxiQv+aTobBpeQRh+yu8ax
yyGkYq1qd29BMrpkwcvD6h/voTOPqQkme2N2ZB8sOR6KXvPL/qjRpAbAiJh/HUWcrUYaaQa06W3u
aRftEDF96qtuz9ZESKhEbjdjDPU54QGlhr9SXLBP8i0KdnoRF/HYYTtr6TbFZssuVIsKPljK+hX5
X8Bi+5gKp+2G9MMBTOO5h/31ErCGoSVlvuwrOMlzXSLxzxHRaYNJrgasX7ayXH8dN1ZqoLaXjRgC
XaI+2zJp+O7auNdoteSYOt6x96sRDB3/nvCN2+DYgOg8RqN9SylegEhFza2ppp8Cn6F1QWb7PsYc
qjYfNMnB//IundnP4uW18sTrpjubYE/H4ydLk+MJmBEsb/kZig1H1EqywtAszD1eKEuoQBUhGZ0P
xpLvD8gxgZmDjpQCHqvwXI66grHR1EaBdGmOWvW7h40Hknuv+CBO4WQEfqdebcLFiAAfu0Jeqaux
BdfCo8CcWzFTWoKqbWnz48s6Ai2BN1EtStPbgC0zhoDdpfCiV5+CkbCLOu/12g/B4D4wluRz8HsE
lksVG0aIQPW1Vm/UTQNCCwd7NvZDcS8YgBGnKIT9RAUBbxx+xQ1TY91pTPomK2thKFQfeYJqNdNr
74wwUwJA+/L5y6kfN75oiOHqEGdPRM5V7cdgkjgtsadNvHCvQjJ3s5UkUkNIBsi98fshWJlRW4LY
W7O7RqId1zXoGXiIBlfLG97g4VowG7+sJs6hOgAj2I8YqMDt6y2ColPr8dyfNOCrdOzUkXbYr+fl
TlqiesfmhZtTbQe+g9WVngz4XIH+cbyiUhlH/m53CvKmgy4wcCvFi6mbgnyRvNPfYKI1BFXrSSrX
RGfUwPCLJTmo1grahGI78cC846oD8XmQYTRgkmFQwg8zq8W4PiN3arolEYmbYAdUeop0JtIaJ4Pp
4yF8x8bdX/o1k0NIYjB83oQYZglxuNKNqDXRSJXyw/vAUQgklbDfQhWpLvu1g5PzacryCBgho8J4
PhBP0VHaA+w9nYOUWZjiLTfnXBSVCgQNCvjI/NLfrtmp7xXMFkkJXrXHFevpa6j3nq/tknsnMx22
PjR47F/oVUSVLFd98ZvtM9XTUEZ2cH6agipiUGrGM7bl8EDJJwFIss5Va70slXind4FjKZ5bhgl8
T3vnfUY7RiVF2py9C59d61aiycKviH8NyHeZE9PGV5IO6vfQwBNOVK+BKbidHPOQ16jJtS2t8/c9
8fQhG1e3IJnQo3Jy9cUDyO31esYRe4ia9+8DURyj4IHkW+qtS5tlSj2aLc+ZBYnPJbkzI1sNFArh
Zo6CKZV1YdOO9GSVrRMWHtCN/wf8+WS19MrCCSJR/IjOZ5lUKQwCYLqsGm2NAfRJBsl6AHrGVUyG
XN00iBgRHTG/fmRv3ZXGeDmqK9kreuxourthqwTEm0qOBPhxvUzqqfDrtAuMSXWoE4JwnYekxZXD
fOO3BLelQ9xbxslRJGYwbCASZ7O2YgJz/yLKO+OrInnX9eQYyoNuqUf5o5KhMR4VKz22TlalY4QW
/tm5cvE5b81JO24pcLkKPIE+b5L8odaNUkASkk99i8KFh9mtvNmWeP+DflkwHT8Rbqb4nr+s7Wb6
jgpXbjt1RVZItmZ9JXuXGGCiWbbDb1gkA+pzARdivKORzbuTyYXKypXkUefVEKTe0RaR+7cMspLg
YaU/FmxntfEXkhksxDUFCpwTvgf9BOybjUnZbNX9q61Xi7iYIXxRPa/Naa5DF13DlJvAzoMaGG21
5DPE/ACnjxvQ1ExHOHEdAAv9ErPW9z0O9zNUKgIJVav0Z6ZZhck3Ubw1JlEOChchvBNTvSint2ip
+NZ2o0hSsjkKs83NLvv8wL5/bXGvdvkYHuSBKU6+t7k7WIJgv7UZz/qsQGh1xm3qY9Kq/0yugv7w
B5W3w4mkBvIyRbIVlTsNiZdm2dXRuadcw7e/oOf+6hesWogN7sEj29tcUnww423T2Jl4hEr9xeie
ojkBTDIrHEyxoSkrBCNifUrfEU4+h4sQth+tMLqJwaGVs8P65VVZ+3H2NUTkypMiEguQD+ih7tLY
u6qsd03GLtU8CgjPQPVe41u/r7hCH8rH3KXHL0Bc0iliIbpr8WXfxpPNUbqQRb9zA2aor3xIr6Ro
C93DGFWWvu1XDPjIP3OH8ciZ6hOOw4v3r2YpAriuEEZzSoCo+1JO/yvKYaEMeL7O2TcNGANqWrS+
dBCHybVOwc2p540cn9tlM0veZnEm2tZz3W6QAi9PXw/4p83wfqC4oMcIbQe4KHyxUgHxWmi/17Sq
CwjY3v6C/XQ53aIgSgKjXoh8PcIjAd++5USnQghU34AumJz+1oy6zf3xsoljPLs2bHFnHk8BVvu/
/WAFHXbcpoqv2HaQablzHTjGZF/ElDrwm7AosCPClmMot3NCuUBqb1onKDTAUKdHHtpACImYlB7P
epJrRGosla5kcMI8kaFr3RUIluOJKHJ/vs2dGlDFtVWZzZK4N5gU6hwMZkki3LPabnMgUPFsi0LL
2nuX9f1EOjbc8yiDHrtVIInqM+c9GYlIRqDRtAjPwR9yOQ+TOzAcVcSqk4WnWH6KwXUmZ1f/Y6Jr
GRoBmVpgX1sbWKx/eLbJPj+mrQ4Si2zeRu+EWJOO2n79lAPw92RvoK0vJh4DuSSu1GmLoSdC53iI
P/wgfoVUkgpT4TM1T+1sokX11HcBs6YnEKXE6BURhKQos+oPLb70x7D2Lex2+KFdOGCcoWib3MFf
QcLPM/Ge6WaUUE2SuBwHbP2MlzwRDTkQoXTENXXWVgt3mL1vKAzbxo4rBY7G6E8CcwntyhuZhaes
8vo5oqAGt2o2KqRe0MrxiVwqrBEaynUran9E7+z+arcQDYUebwNK2l9C37jfEcHXS05DDuiDjuLi
8t0WitZXrH9ixoZvhv92F94Z2OFxfJme63vhyDWBRl0tzlzY3fuTo1ZvAyKZd3VNYp8SZ+AQ0JSQ
Z8qogv3bZ8TN2XZJDCCRMpoH1orTkNAfkMIUcSKb4mLc3HD/5k4WvQmMkNmwKvu1/WH2Z7Bv6Bfq
ajUgSbIAXLRMRp4JoMNzkSJCz1JdIoNGlqrVnmiZOf0irSsUTzFq3C2YURylS/CuCiJ24Qgdw46t
vDhtfzNTef7GVZHzkGtIfOml78mXstQV58PNn98z8NyqVicGkCSXIxSriyEGU8KeT9G3E9tw7Gsr
V+JPDRbocIdqbRGrCcfUEVHkA7owo3tvHiXu3fDgj8vKR7f1LIxZh7+QYB4ATuW0v+3Kl8J2t7P3
WmKBPszmkimdSIirMNAhhrTAbbxS8iYZcGXoFt2aFg9psqszLRk3KkU7QxKjuwzHVmuNHtrvmq7d
lUWwJY060aFHU8bPCKYXIG8oBKBtxI3haS13tSZz/vXyQab9fHhv7iVVsG8f4q5JBq9lMYokXWDF
8O9SSKn/U0I2DH2VHxnQCi5uMWXo1RmBxrsgSYwhAvp+p2esqEPh6CVss1Zr7LGApQxqmIpGblOy
OX95y2U9E021Njwg1o3O1kT9BYSpGWZ4q2G2X1xUH5uPPuXrfI1hNe+1C44twEU7E6B7u5C6E/Gm
PJ+QmU4fiwCo7SzSpC8BnLCOg01cxb+8sXq3tpiTgFa8pvmR9yAA++WpTdwhrLTuCZdsMclmyW1L
kc0InVqj2Dd7g3lIi1t53HlrZgJ1BAnUyAWMFkbg4jY1E9LljBMaLk3whZqq6dv/6YYCaChTRS5X
LBstJp7ZjYEaaKnU60psDkThQlaSpFwZY8+3M+oydzgdW/5QMw5/GztJSciM4XNZknHUNiJrJ7ho
qrAbYbXlzJgqpdA6Y/8mOmwOWZgDKTo1dq/k7MMlRx0z5PDIsW8S3iBmITPLX1HCWyiTujShEb32
Tg6GESdDzOqFyO+zeUu6feCwVOIbflvoEOGFFus+8gXo5qW75dVhsdni4hLbqwYa/hT1DC2UWrTX
YpEP4LtWYBHrvqw4b8GYWIIYCC7+gb7jwk3/PdiXwU1KfRbzIRH42tikXAvPd3LuiC79BoGs917n
/N54+X/lul/2I8YjOAiic+6gAlx9x3396iOqS4OAILgkOR0C3TGdlgKHtSVDtCFkj2sSg5tKJCaY
QUOsyr71jdQpVu0udao+MZPO3+hSCy1Xg7vKErUpriD5o9WDIZuKuokUj8RJXRhe+Niw3zfxUGrs
VCg6h0wXeO5YQhqKPPXsr1fxRFofNL7hMHem9QCQrRhbs61L8qSq+qQTsTM/0AFAg7Knvjgu1+l4
DhxnfPixWJf1iqbYO+W1TEwfr9Dlem+kYno9HNbbxGp640EssZu5pWsyNR2vc2eOyfjVXU86ffz0
n2kgjkWf8KR5feG7ZB6Yacjb6err717P0qDqrBiX1d56pDfS6tDRDbemkcZFgoKxIvWq0A70Js6G
it7TUHdn+2bwM4f8j15BOhDBxwYQVXV95zMvh6z6SUVeIhFadsG3Rj6sQeahZBGs1CvwGEPNug8t
fJPezGN6hpyBAixqxLpTWtZNPE/IFDAv+Ug23Qgb1txSm+Qbsk1VbMNVdgATV4qOa6bb2gb4kI3w
4tkW7tGloLCPjhqX0hSMdx+V+C5Dgu017xQqkHo43eHfKkAcLbIyDUkPmxfkm+fmdQnM/itb4rRQ
b+zpNn9b5OG52milAuF7GljIEIi3rlB5OjGrK1mgGv4g/PAl6L6QZgFBBisSWrQheHRKt+Hm+y4k
6zgvWpyUs7du7Uj1toW4+PaiMetj7RtYbDso5f5gB5TOb2eJ8B+Yg9SHeWcPLl/BUEf54K4SSX79
vjGdxH70X8tK/HOyXRr4CYqw+YLgRz7dFookbeRiYtCDaZKNHLv5vSQDVuwO01f72e2CUnAi9qyB
FlN/lYjb9jVYfwfmm572CaJ0ix07a590mGU50CYsLgIYmTSMRcw0X2LjynnQSItInw83hTBZMVvh
jy45b66r6YxX3Vx4a0ojvB0YRuH7RHJWvEHmfXTj0Kke2nc/0S5n+Kjig28FoPPGXHxEM2YLmvam
wXgczFfPWIQRli6y/IC+NLEBPu1dsnGoCZo0cBfTGyrbfEO0KLCMVjE1K+SvW/dlKUAnuTWDKkqt
4eCQoEj9NDUq5AvmUKHL+NOxJ6VegUUlzJQHxxRBPQfW1gsChLHH9opIecds8pk7BuwA3zhxkgLn
+FticU+Z8J/VBeP8+leFUVJ5n/hqgWaaOEF/Px6R5V4WSlHBc6tdS/+XI9D/lKKL3CTGdthU+zD/
C2KIzxAtz2N2xMJVWobmBeSBWCavE7B6K2/rC+WeUP5Y91am2lMKM3Gk47SJ1f6Zt32aL7STWVur
wYRPt1iXPDgIUy+Zhdd5VCJFgTeVm34y+8fGufgJvo/ecHDDarWTiM7sCSliXJjgRLA7yT0JRHgw
YYBs8mKzAZAJ4cW22t67TqD0MxQ+dCoolQ2vKbXAdmETFMlBdZ6Kq+c8//AtuHL088eq+e5p/CPt
WSCth5T8YhO4iBJEUrovJm9Xc+qGzFyAPG3pAdkGsEUDcLsD7uLqShEfPSoaUkjkM5qMiWFLB9Cq
gDzTxg5j0q2PuMoplVMeA657cpj9+ue/aLUz1Smkgn6Uf2/nVSXyWS24qt75rKYnHPL2lXX6rqRE
bcX/8thQKlUfIhHAdLF3po+BYjcLY+PIEU0bviFlV252/FFdum0MAUN/lZuF9KsNT/aMW3m90uxe
r5wAAXKFonyEPUkiPu7oog7eCnOeRKImJvuxp5ZdZ9/i41VTD0Mv/dpPhT7+byAPA0FQpGwVFxG0
vAhsUJsKN5IvDCjxVLgUWKJMnGqS7LUosTz9AwUhKw8ockx4y8Pd61dSmW4THXczhPsB/DZXdQ69
8AaNkK6WqVF31XYYQyJktYOUOjlRjvKdHOIQGXXGN12T8vfehSul1nWJ8XlqzZkebaDDRaWlo+Lt
DKKJv7y3q+l2XfDeDNF2/uE6y9t5TtjK/wCmyxfNHuA4NXiAflja1ogIMo7xSwc+c4iJzuuAjF8t
XfL++nbMSe7A21eUWGGMeRb+AXUFzddeFAiIsv2Zw6oLKdTCo1gdhfeTAH3PMjIF213iO+OUkHwt
O4kUuW4qkZmalQ+iov/oNEudubv95GQldOuO8W6nrG/ASV2xuDKI+zxsQVb1RpxVPy9psjrLh0sV
5QnD/1yptgJYQyyPjuSockzeW16SNGJ4KhsMcve2jrJpJvN+CPUXHBSHGaXYyTbAkFBb4som3CsE
sZlUE4tRlvTn8zuE5ghooEWbsMXmdK0NKJuw152EUcgfaHhNLOxSWSkSMrwD5OZv3fOt01xI6dMf
YtXTufXjzp9K2P271x0ykAQxMkPCVjP/Wg3NXYmmkI0kWKnfHf6InCbNoiQh3JtDAnDWlNbMZ7U9
Na09vk75+/mTCgnS8i2eA7RQuQO+n+1w8OI9PI62vrau9HxcKQo0yoTj1WdE/pnxfdk+1fhldMHp
p384P3GKSSHMffuWPWqq+ftbr99+xu5cExfSSB+VbMC3kLtfQLgeBjXBvi4ErXomR8QVk+LqvtuW
Faghk5NQjPNSpF4d5zA/nXAFl5j/gTcqK1EWqkPcwQ/V6BW9XRwYI+dABdRGoMNnPs6hSTLPhznv
J+31DVuaGt98CkyVsBUNu7DaxuEGUswR03lAP7wKx4e/1ebGW2wsZftuKP9mlRrOH6tiaIsOORqC
4G/8nlehPHEfpZ4hDl4kAZu7mP6alicf2Ve9EhFJcKczFy0lKxBjRJ+1f6iw/1sRUeOM66ysmk1a
WfsGdmXKxIGgQJiRGZ4zXX27gflTCosXbOBDrcEdEIwyJoGcc5kn1uYAym7dYrnGGIPhQxYUBiTF
/K8KOK1AYIPYIqQTDu9U2orxI+fY81qHBeT9cIGA+X0G39Y3YmNYt/B70ccZNlrnMNhuK+kXoSwx
Ysnu38a44fbLO8/XHTV6Kl60GGgYZG5qLcrbsJnaxZCNfybL//bfZA697UVWOSFwug6M+7vQzqs/
OcC7mdQVAP7bs8TvKL9TwoYiCFX9wIkPNm8+co+bUqT1QEHRfqPNda4cXbyqRfQTHtQEiADdqm1l
oQx2k0IkMSzjl9WgAw6b6no7aXR/2RJj3+45rGdTWgIH1TcUBluyvA322iGEquPtBzwCFmd3azsr
dQjjE9upMnB/VW8DeLZ9z7+I7w5pZGRrMOKJMs1Y2T4c6ZpO0kyMUo1Teta1TMGVolj4SPtLZVs1
zH5aZ/437wsDbyO0rkIXJ4p40yE6p+nedhneywes1fSK/HEq1GbvYtgzpsWy/8YpjHkLdmr3Iu3K
8CPhPY7bHNDaL4vMTEP5alGG1hWwWimz0GY2FYJKe92Jq3SZwngKn8gM4RFGwIpvVegDcFLN+0+O
pCVgIwvww05fJHkQt3vDN6sobkve2XNFiPGWfz7/gPhwZZUbkrimalYjakS07w7TQqel8XyucQWy
+oLvqa4rMpYpIYOH6L7tGluDLaLqg7xUDLy9G8Awl6sTMSPw5XSb8cGPt/U5NZhup2+I8s7e17pT
ULwUHuOc2FdUUQ4ctpGbMmnGCo5MtAfmbZHOwSaxzYzui9Ak1xKHEjOqxUTMHa2LYi5qONCI4GXQ
PpyQHqM8xkQLZA2GeGq9AttmlpZrT+GFJx3Gnj9ejM1KKKULgX1A1QgSNsDDu1nP+C0eQeAyOzrL
3r0fHR7uSEKOb0EEaxg3GaP7i1rOyxMFRRSwEOnqNWr/3YIayh7QFcTsznXPW6B6f8cq9EnX4apL
o1TOM2oMLlwBP23ZLtex0yA8YTq+cOxfJexJ9MqpRjiPUG4qlOZxLSF1zPwCJB1Glzxo4BoHnahk
LSoFu5IrQixeVhyL8s7tmXsmDn+bYDd0pkOaV8zOd+m7FliyuY6S1LesDH9e8CShkjva+HOH+BVf
EGhiIFTyPcioIUWkZ+XGQsNDGC6QEy7//mbH8do4KDMELT0ip/ptCtevkk1wlnvtPNexVpX/p7uE
0us9BDsVPLHY1edw6/5+zO63XYlktGjrCvIYSaSpbDg/DWadAbG/hA2C4TTBvAUyH5iQScpYnp0g
N1L2KSzkIZaYN5AA8DYrqb9ty/jsz5bxZFpUngqNLVif0m1jdPUA/1qX523cWCZliwMrXOf60qVv
4BP3OFMa7JduZXIVZzPUnSHN00D3ktM0taYwoMaESd13QXTpGEc+aLfSLE9XhBldDSPEsizvPJ1c
tIwZV8S/5O6FeXl17P2uzIDxnf+abeQ4I9uYMb/B218TrfLho/f2TrWyH6jPK/y3hbwRStOGA3zX
VHWDNuaTCxmArGzLU5JHCl685SOVvD4LYv2L3XkFITZKskoD/CaO3Gbza467VCPej85uwocc8YcM
yGOn7/a8XldJ8k2Mjq2Fd3466Gxs9+u2ebJU7N5e9p2U241KV0r11eK/MPMhLSD998pNt5sA8w35
vZfOn9K7T3/fVI7wu9dW8vz++tbEZIWyg5cTUaNf98FwLTyeHagwNBgU7RYC9Y1y0BgDKWrh1jyC
YBHwDtw9pLzxz/dMEaQMFWPLfL3Jp55yI4N5Fotv0ila6Wr7oBu+2nMfxkNyd1ZONxk4acNUBafi
rWy23Flpb+rIvQFMLb3VxsowwwaRn4pHhLtfeymEYEtBCGqjfvyeMOmTLTCbWz3ATELhISBCY9LQ
iGukSU1zpcut4uzeAEp1fDY5gRpnnuKA57JdnvZWDvYGnJFmIpXT+NZGsgOK2+Omh46as5yL+Luf
Z5I3Dzn9gkqyrh+KvcZfB3oJ+uPSIUopLcvqn+nhjJW+rG7PhxOa3y9nKb+N7vEolK9GPOSym9lZ
fpeP2Dd3bbLho8KOyCOJHf0g6I954H71atRq+9PUGv2ubkM1Z71ltbO4BEn5RccqR4pyhPlNN+B8
6CGgxYuaxI2ebZS2K0Cpz77PlHp+xySm8L28W5i4+a9+6YrtcmJvtI2slfIuWiimzyXpEVE8NYLy
aIP3iDwNO3QVRTdHI4cJpNbct5XQmYWLQ9IoTF9jjLVWmqrGeraRtdT4JgvmE1zHOhRoO4AFBWOT
lyDFBYTu8NUXxNjUl510LXGBwXAZQ99Z/N/GieqKcCbkOjlJxGCh9psw5ytguu41APYXzkr+euFi
XJJf9+VjA/BiPamplXCgguEHDNih8uWFB+JMSI07g6R3c9DutHMywUsYRwdJxLO3daw3GH9wp1H7
if0opFmOlbN/4eSf/z394Lgc2R6RwFBPP8BSPme86kasH4ozSmTUXtV3/XQM49pLTXpVTeLKJyb+
iGuf32DIEZearjKalWUnyBnxCwzJimESzjx8WKK7u6OcvpTmPswtwSnXhiNJx8stIohpJaEzFpED
rYGWJCiQNnHlyWSwBjIqaacqiewqAhGiYL0gs993eRqY7E4pFz7Pu0+PVpIg5HMYiDOTA7EH6pbQ
wPM1wuQaft2sCNAGqjC7u7FE01axtu/tDtzLEOaQYPZJhlfn2x5Um8cbL9gDHvEH/ttzCZVCB0WQ
adwRSHslsoVl3YzjujTmBncgTjs9IjQOMMkTzTFZ0kcS5E6z1uE7sE4XJUuLJFF+/lpSE3KLzHcz
UnOooaMfDmGaQ8e7QVhM4er39rH1LkGMh7Uxdutt3OFx//cGcUuhhyRGEGUrZVkJF/LhjUNd8ODt
qM/KAd0fOxt6APL3vBaPn0h03q0kbVk6HD7V29mgtP9epfywObcDzl+k9/m4SbOpff1OnBcVn9mi
9lZqV+byFiqsfIbuQ53ZveLnldhFcAXck6eJeye6mJZf8nW4aIz+6JO4fCbijmt7jffTwP5s5+Yx
TMjIW4Di087BYuP4fRRWkpqtrg3y/Dq06u9kPrWa/WHB6lfe0TnJyPejDosG43Sq3P6YTF8LkYeR
XFriwpJPiDVDjV3Gc4ZE5NFGeB/suPyDpUrH2uCtqXXm6KiK11/WdF5gV88VILqga1XMJXoVzv2p
Czz/ybtgyZSUczv2MtGSFfPg4t2AekPbeqaeQ1vVCsQaomiZEMNcafAd7+3Mgj0E3lMhvKGdtHoU
Z/Wfa9JgtnWp8d3fZVhECzcdMcSL0DMugWhVa3rsqlb7JI6G0HAlcYDvZwjL908GxWwVUePQhQYV
ArfWTO8c/hM41bB/PZAlPk0ipAb1zL7h4sdpzl44fwFQyO+9evFuseC//5Ku/cD4qFCLUyomeGN6
v2UBGEVZYbSRKh3AC0SpChpgM9FotJOmesPhxfNjq2Wjb0/m8Xionq/kbYYmgGFjGoe6zesNS/5z
rBN7l7W9+yb3dToL1FdP12mA5WpPWzZvDnZpXubdp++iF87jY8f0EOSc3hlyoxynUGjw4udLw8e/
PWjvo2HhFU70s+h9FiKndW+kvL8dyv65Lh7VIvWMS6CuK7W7eZAwlUkoyYPdwuj+v87WlP22Cs1g
EJNeZPlEddvNlr4IjFFocPPfpKyTBykEUz9X2MmLL7CB1LIvIoi06gqIFU1M1zeVa7dbD7Ujtdvg
D5/SccR8QAgGrzRxpI68k5FMWZ98bvTszYBJFtMyhIVAs7AkdjWSaF/BjSoxrP7a2yAMw867/1kC
PjlXOw6HdY97vf68bX7HS3ExlFg3OuYIbeObL5+8/ZjP+prfnzYwCCYNpnduhe2BkEnP6XyQXHli
lTZg4/UUYw4FjwqA44020rpOj1HI4Ph/I1+5evm3qyjPDmnT78kJjBHqzwG3bGVtTohsGtfrt0WO
LDnrAgOM/8tAARalhqXz/r81WyXtY+oDQjTkZE4E1R8L/msf6WuryZv9jBk2ePTfHjc3b+jZ4lan
SSY6gJRdzyayXSO6LY0nDESCNN8oIHrjcXdLMQoiudtRXU8E9/31nFv1eP1BLyVFu4M+6WYBPIQF
Ne+gwpIDlhhqLUf/zTwbgX5TzPZNCm6OBc5V4zfMTA1SW/Bu2E/dwhNTu4CKVLzFNO/lD7LAIsUG
Hs+tGyc8bAd8a+jPx7PZqc9PEKqBWhD3V4qWG5NzdsY0w5ehSC4cDZpSziUeTENIol709/A6E2qn
MqOjO4i/yAKG0Qz1bQI7rNVWLTSH3P+d9RxmOwgaOaxE4+dwcWV6h7OY4Vd0441Fhi45yx1CZGEg
pfQHyUP2mZLQjxhJ7Y3gyXHEuwDUmY3Cb5E1lvBIuBouGf2mQCh1l7QMT9b/uHO3rlK6DD+zml0Q
2EKcvMqUq2Bzq9C382CS3PHGFj6D58+Qbjchv/kDRPKUBSryOr5tp3sWHtmKOrGFvbi1+6CWtk3T
y9v9XXDwk0PU5CncWzh9bXuQ/7XJXMHVfPw4yOtNBdAFpZYuWS0DjOrPS8fmrg1GAdW/Dk7wpzoj
GdahU1B/CCl9OGDyE/H5njBKbAWwi9rHi9FMmYT12mj1XgJiSCqYBK00IJ/9tfDpqgmP86YJ9KXc
3jauNtiYY9pFeXXbtmwsts8FrroINPbgszt7z4w23DmTYzyflbPHKHQ4gt7fAS7dpAcWuBkmHOLD
AV2WMnnFfeatMipIXyD6J+9wkAqcl1NvSx3nL3Ytz1tKTb7zTfoy4GJgfigwvPYXYtnI5naxj1lM
vYuVo1oUR3GsR/R+Xyoqy9kSFBznLRVKAIIDl0BBMh1salMVT691sJP3GZpdVJBMrWWDaoQv/BiV
TTGQx13wxHg7YdJvDP2wk8IY1/iQ2MxwgmAR7JSpnSWwHMAIeEYqODd60dLHojjmZxrJjjuBzT/Q
DJ5D2A2t5/ELUDhSDNbJBpoS1ibNOYtZxfQ408w27+kmxifzwzrLNiDxG/2k9cTnMsbIHF8lYN29
QCDKMuFw3bWuqrx8WxXf7zr/YUsrUW6pmW+Dj9yWDIOYRCgG1+UgEOsPRMEHwHMnVPCyuyWVKyu5
X8ZyiCjdqDQR+8kpKUwZxbYdSQo0AhidzrejlkK8ZhFbMJHbR4j6dOVhVhvLuor2EI+/NqDtbBkF
qm345F4hXXqCdLBvIuj4juaaxH6PFugLwEoZVx/G4EcKrfmQ7VrC0Gr9ALKy0+6OajEjLYeGxIWL
sSqQQl6OL9db5PIMXxm/69XAQvPccvpyDinepa/0vozhlbgLdFptGO8bZ26tt5sX29vHF4x4WO4j
oXv0GMhZmr3mmWSHBeQim0j7syU67wkK8zRdNUQdcCYOIsWHHwM+JS8b16g9dqKgImT3kBxW0j3G
7+o7RaQUxgYsbPSejcQKHnZLtO5svJSwsllpKmRymsdX03PHKmWZUVVim+EGt5PA19H2HQBgoHu2
YG6HrplES3dujoLMDY2k5EKQB4BlPbsLjU8Bza28rRpfjQHxKvPZ7K36vspK4M5p4zhIAposu3fA
ik9V6ulv44PN2BLc0CVuHfiCZN2A3wn+Oh+yP364lmhYbUUyCkqhmCXnDyCNqEBdKI+tMVi/d1Tm
3evjqHfMlnR6Nrvkx731mfgvBm0/LJRprxjiA/cx9GP4/kRVsbIGilp5DcOUfqXY5bgFN/s99dOl
k675cqhWbj20GZ7+v6FItelSpwwfwgbie/MbZH5S1cxLL6I2oXmFfEcKeA4mZGOZctQIwKSZD5m4
e2O/vlpxNqNNzIof1envPRMCsB4G+8a1SFnZmTPXv9JClCaTcZl7ksOkVpvvR90e1HGUWFEAxVOY
o70OAmQ+nFvSguv2CGQIAJvgMqN7BKD/53hpF5eCpD+dnQw6qmFdLGy2Ju5ZRUOytoxBq9YSceTR
A6kD39wbsiSKYxoas8cNga89oqWVGEwJzwWNbV3N4as3+yPrBUScf/tBqmKXgtwtF4d7VRaISqXS
fdZo/McLGnKR1uiKROTJzm4P3sqvBLFhvIhRtja2JNQnOgl4JN07ABYt/mfwcyAuF0M1aITm0C+y
SOTpODKQBrNnbATr1u2dGtiFZj887c5PvFDotNzNZGqr9bDdHnVGU77O9aLIwrKnt/guQTBk2EEq
gq9gAOL95uGFdKoNnxlfd66o5PTtVaD4op2qijI34yj9QB9dxU+wO81E9k8dg5YwKqLVvX8gxgwY
B2N6eCWyaSGLuWPWg32fzbtw5rUdTeo8sgHcasYxfe/+QEBQSUc3lIFKF6Zt/cm0aNrUd2hAYBpC
I0As8ml2DiMbhj5oJr/B77SXzaakVTi9ireC4tVlkTDtF0uCaYhM0u0MGg7/GnWQXYeCo/KZgIh2
qrricuWPFHlHMU8gocoLfH1mY9qkdCxiar1APm4wQQUji7bubuFFrjQzQeJE2NHSFdzooss1puOc
hbwv7QtNCNUo0Eg2pEMNll8FXjE6sdeEPFOTEZtYF0duGMtpUKvom2S2KeDcl+t9EvCi/usHUzYK
A+B4pbVTYSHc5tFSQj9HApTCMyoq1q1mE7WvbQponLpc3HLwFCIK+E9IQHOSxEg7LY9EUqTGtHZ4
82TgUKTGtGXnLPPN1ml52MWit9toCS9B5SEnJY/btJMjVucMv7DKsY305c0lQhNSap2s2uYoQ1/J
rwmUvm8mHPj7AL5ABEjeNae6ylWzbTjFESN19RjokkGF5w6+WzHAD8qplnCCZt2vythKwxPTv8YD
5o+2tS9mYm4GOBW8UbmB3It0Mh5/4EE10GP/On+52sPT65FbObb81MY71IUIKn8TQSfI6kEpzUNU
U45Vcqo/hZysLGfj0wuM/1KitBBm56Z6ZY3uU7bAcplHGsWnuN9GCJ4FGdEuKx4mA0ccVQakOlBw
O7iin6eQ1PjgIJ6kVauiuP66L5C0DOUTOFxKt0e4jMB3cknZFymoFL1f5lhVdDbrufunrreOEDd3
IsiAGNANIKPtvTpab8usU6eXljxlVG5WQRJFPvVVYBEtwHphRpz2NeZGL63RX/vRtcaFMr+fl0iY
ZEuwopkbDjom1J7/bvkRQeG+ZT/7XSAur39QTvxdRl852qqHifMlRound3mL4JifhzRhPnF9QsDT
VcPpYyDtMLzIbyPpbOrpb7ls9DeywRRwdjMicTkU8/RMTWuYYW0GgoYECkpmVZO65wq6yccP+B2K
dsTOoMocxGydDvZHZE3PYKrCIUmlW8f8ZZwTGIV3xRCBQJQscpMjxfQV0MMkNZSQPI7cXuGgcaGX
w3gRM5hpmuc8rNtClB4w1m4d9/SOtlm2o+dSBLeAwodcC0Gcv0sC18SPHN4TjeTzbd95CMzokdAJ
vG8tMvqTgO2LpnI7OAPdrttw0r4vAyjWdl1+5ju5Gv/8G8To2MO9m/sUH/pwRZDDCld/hUSFs9cE
+2YuYDQqwLqAo20OAJGA90q396M87+IXK0XINKJJ3IwajmCm1SxnOiqLD8tQp3kgTV1rEgRK9UTK
Jz/fGvewdiCP3pbz0LGtjqrlgmztgF5dRpmU+VSMioJuLTdBR54XoPdMY398KO4fRrdg8fRpqNvx
w5JxuF7f2kx5IVMtvAZx0wIn/LDepZyZqmFsXmkA/D00MEjs8tl/KDppUJPxYy2Hz8xbfr8ewYQN
9aBP/mEl2SE4MLCC0g2YiebwgBFKev73FOQI86qxLxO7bm2/EFI4zFNUW+vH7LQkzcGHU57ZzM3l
Zwj9K210OwmTMnvoaUnXiLVWWHYo5FCp8QoChbW93oryhth8k5sZWsV5IwhJEvCcAdvTMZ0EvkA/
661Qnw05Y+ezOLgi65M8mPCpRdiITdkKbyK/C4GF/fmwd9w97pvSzuRvkJ3HQe6lHPUiR5hPDw3H
DB0z0+4sqPpYYFI+gm3Ct97yKOn1lmMfFEt8u78gImq74kxuENC7aaI7H+r5qdjFnP+CjJVak+OV
cOF/jd3d4jYVpGyth85/ztnnM5Hlvgf8tyFFkbp4803cWw5yOO7u68H/IeK82iaZ3mUTZr1fM/kt
G3SysGj449pOv8ArQzedmSb0g8ssTl420UXcU5Ciq6KZj+OdrHil07dTQh0yHyTOyBzm+r4ul8RF
rhk+9RVZTHxsk3AciV17xGveJIoSXl3psNZ46JmWWCLBdM9SBt/lnvPTyhg5/njflGlEArHJn+wD
5BC5wCws412MMUNaRZMvvnCvrfhtJ+VSorh2ywCksJVrPBhYRoN7qXwYFdjy5nA3mmWdWbdKqEpA
oasmXKAPK6Li30/NIHCQf0+tP05qitC6zbXiAevsBFovszBkD2YL5RJqqdMBQOuBoVlobgJWD6sP
JJYCXec5pRJxZyWM7cxkdou47T1ZDfN9doL0RxC3+RDOjc0aT5mUy29VsxMw/jfs8LHOttJ6KAgV
0jU3QKtWgNlultr0SLbHQF6Zd1qgArGnPOYVN54J5wEhPlh3ecRP1qe7X+HmTkoZ8lu5esO0KfIY
9a+r6taOVir9q5d91lu0bdkCi6Cb7vBVWVhf7eHNy841tlJZeLdeP4Hx35sqpnjoDNLNvCHvgAnA
tZkvHizI4+6nHr5CJd58y2Xe6xdf5zlNG9rA3l37SMH88UUxt7mzasbUc+A34qVJzb1zy/U7FZrw
CdXfcxNm2vh7a0DtnW98AfIP1G71StFgvRzBwYrAmkmVy8+ZtBHmY8GxPPIz2nK2g0RfDPhezMRC
DxFU7nd9cc4sEdHJQ34ajk1pkEsJIXWL/oZCzKAdmG+PhyHrS82yTOyY9OZHRF58h7rYct8wHhYu
xLQKbC1bdq+hTymN6MlmTzwMEIU/wSfEVK+D6yQhxyYD3S/DvZwnMFet0ZMxzeCsIXtCRQwP1uwx
eKx5lfKKiTRNICS7wfxXfCpJcqnxK+j+PdiRnNjKi2HFz018EfuK8kCjMy/5vkQYddnmvZz8U+5j
y1pqv6uKtq8PWOz6gEVhDZfIyNx0+jvHzmQ1CQrClv299uLCALikNDfHF/8iQpliaIH8ybhv723b
I40yNlDL3Cy1bdjs+rEPvs0hp/pESo0DcN30dkopxIp0lNaLQlCll8OiwFDhxbPTOiUOYmG0iI/F
EjjNIytpuVtufXCdN7XiNP4brC0XG+uKySwFDiwVej2AYwLflbTnKXuEUr1heFQdyCAur5b8pkVS
iySfwptWDDSjHTkEPl5+5SnyxXoW1Qcx301sl6CTc75ovZ3ouanPIfZfOhJEU06Dq8WzIAwe6qX6
XuGmO10nt6ZmuaaGEFBU1/5NvbO7iKfegaKBPgtf/TiNMa85iRkkbjcW2jxcIKU6dNhFqxvrjO6e
JlZv4NwH/jUIeKfu8Ur3vJzii+vqYNIEYIxcTP8XfUBADula1MwmOob60DltqVFbGmdID/qrbLPz
0bUh3rGmk8+CUFUNzVgy9yBrU0+NBnebXoO7+1BSCbydcmEc9l9Qei5rviH4nIb++sZO38hz2GJk
LVzbaIykviFUnS1OPzTLGkbA+JwsEjjfX0qwO/EXi4SldUnkrjO9Bm2lbfuZCZgjFukr+f39hbzf
h0TgxY7IV1a8fn4GBaLPjGvoOUkKbqKOXmtVykG2C1UKYMPmI/FQ7cbC9xlrMb8ZX+WABa22V7d8
74AdrE++02XG8IEWcdbYvU8rWh7Hl1IPdKHW3mN+Ds+/JI7JHNvUyB4e5TpPWcdc2QBwBKUfI3hJ
RdfJ4QvGHQ0tKaraYRBs02O8mCGGWd4bR2sZ3cijb0vYlWUT0mbsCy5uobc3jSBRaQfqf/G795L/
yOhNwubdxvoQKG6pwDQK9NzlNPS6CZdMQNuNYtJQoncxxqW4XKvpwNhdgFYze0RC5bmkj7wO3jwA
/qLv/IXk/i1h9cNbOtcp3zJ6d8ImQt91YJboIvtaG2V0Tx+nCcxq7nN2HGB2Od+jGLK+pw/rfVFG
hH9BuxKtBMCwDJ/OJP6IuRILKKQEXRYgfaH+MVRac3nbf+P9SK7mrcb+IhF0Cxuj8NFm7NrYZUXq
8GPNu8aCdgAb8X3AFSEPdT5REnLfCoVsvkX1RNKcX0mUaeJcdsuUOpWapeTXXbissh9d0wnrdYAc
41l0LFT5GCGaROrkXNss/A+DE+8glSzuz77PcWlY8ivWfF4xSeSzm1YjsCGEuWfUCGl2G6FpZE4E
uIj1d62H1NXfzf3KI05xuL7xD2ONAlXYxxlaOA1xFS/oYvrUzW+VpUUC71Z/WvRsdl3UJ4OuJhAL
q5JAyx/kBj8053C/ZgeuSSytIfuolwPOxgNpkg6Vab4fh4a7rfXkaW1e8Me7BbydSoZjqRVAbpJk
ku/wMLBTjkK5Bzo+6cm4zyFoJyf/XUkS9Beala5dfxC28Z+LJOafbtnUdpeOIKCzfn/RhYZO55HJ
Wk32rsIgECRWyasimVlm3thUUswGCW5wFbxO0WrSTj2mmGoRXvouwiCQQGN7r4v4eUNBpYbzWph0
5QwUtBQ57fXrPwAirDaVq9cKY1eHzgwZRRaqpxFuT3IRAFVX1XnjmOpgnb6jVEVvzr8zYE4EceGi
5DhOc/M3H5yYdQZ9CBq4yRo3uXNNZ1tY70irbeGQ+oi3phM/y2NJ0iAHNOfCipEj9Bc9eRefWiIX
3GLPMUYINeBsoVBggpJlQ72B4VL6677amPlO9DsuLa1CpC5YTD2OqLGOAIw6Kk5v17V5XdlbafCM
+Ybgj0QF3URbzNtaCO1lAXeMNAVo3qrMHe/vX8IHQ2g15R7xAD3wmcUlJaTQLH1yEeZ257BE4y3l
4NVf+2/gjTElSwm1vlLm26HeS/V+kP+qApboUPNXkm5s2iqayx+HIiDlQ9X99qWf0LZ2etzRFn27
1MTt2FCTLu6gbO13lntdlXhptHU8OPG0mf6rU8+s1c7cOEBGwoQ1lMEE+ZI2qN+TNQ9ub4CmbbNQ
esEnq0OHazC7nc+GY1FaRZUt95CeJcEm3CWwcx7Tjk9cB9mCVDcJYNxQizVgsqdyzImtmfLVIYVl
3SvrrTD/MdZRjmNHlFZKtjKT1yYZubHlf0W6PfNCNkX4CytgMudWNxICYUt8GsNfjbUWo5UOnP8C
XYKIrYdn4/0itU+JNFV3E/KxSnkfuZ7wMkHVMCkiCaWG7GoBif67qPSIOt9SCeC66/PWrpGyaUGC
WaNeVfZf9LbaEOZKcxl6h7U2S6TW+SW8aKQUsgIHHCFVybJ6j0DTQVm54+9avFmJCNy2Wy67/Lhb
h3G1qNYSmpcFrblXy5kiH9dK451B0fjgimV16mlQ+149N2CXGXgFBZkSkBYUZbWhvIt35lPx54em
z1w4z6VJ66g+mOwIfVDDKaVvqNsOb6Uu/6hIzV1CBWvr5Ww4Nw1RYp2jJ/p00bPF9Eobs7OtDRuG
HqwkGe58L3XV4CO/lcIGdMWH/YFtXjRhfTtCxnLg0dJWPw9qNwUFUuATaDzP1gvQygVI2393/wHi
ev05lNipG2g47KVvvhoX8sxbGt5c2tlFjL1sblv5VMOvHITiFOg0wnaNirRJw9sUN9T4HNhE+8SV
CUjrOB1G67jxPxgtmB3fkrCm4ErrKFX8UZAc4DWVNbVgVO0v5p2eqh0CIfShOuuv83ZJxLM971tq
+C93guY6rUO7BAxvFPjkxUR3lTqa/yHOfdw6xNPy5o0TFzb1jCDh6+kpTr87cjp50iLchZcSagoK
olyyJP0NAoy/0zMbLyM9RvLSWePwcjdF6QwsNK01Sc6VpafzmyY/t0HTqsZwn+GkamQOxt9DWBlC
ClzQo77NpNkuly1TkgpCf6ZdP74HH5qv7L4jt3uOHFfkWu5GIL4fBsE25CKsGEiFOyj4yVXw/FrP
YSfr73Qfn4RzWi91FaXF3QupR5/Hr4a+4nsq6upklKKea/4QRXiS5d1xHmgrJ+BKogYwbzx53Pqe
wwyAYBwnzXKlmfDmI06lP3eZzkaQ5L+BD5zMTd6EofMouT7HkGkghyO2irm6Ti7LQHhNWu8jdc/1
v1DjRLcgNzN+t8N6g2tApOWOS4HqDn4ZrrvL4oU2u3GgLzUPxiKorlhky2O0i8NJR+fNpAO+mK+t
IJOxcoqQ694iOQmx5wosTqQmKrq00Lj3JHZ1V/7OGH9zroIqXXcUwSV6/eNIVeaPZVvgwwjvQiz3
3kp/sVXy+Gaylf9bS2OMm4weplLcTCXBNq0NlUjGL70mrnd/KP9SLtCmdxxztBokKBvvZcnQi6ow
xdXnlIBauz5Hj98lyzRJhgtDGMTtqQSF3g4FQRAY8HoT8vt+hF6cyyGtsoVVch6DhwETi6gp5YnW
qOwahaNdxzUojG9bKYrXU8KWta4b30ggAT6yRuX+e9M2w5lfCyk2pGTckrfnsJIsxVSsybqh9Myr
utsQqrh2DtwkjV9m33pa5e6hwNdmpGmDILdbUoIlc59qGiv7D1hmFvW3KtMmKG0cwC32c66PnmMo
Y2rMavIX/Sw/1ouLS/5FmfuhHQphZnaEx99TUMX4ldIC/GPbdG8RqMpphGNL9iwaBUaySrsOYyJV
f4YwfVIhjed9JaHmBDF/NMOkok5UfBrYVy7AtQXmyAFSPVa9a2uHiPZr98o81zS+FU7i25tp39QC
qxNqKF0d0Q/1Q0zQP2a5ON5LmJ2p/4RqHdus5IAS/I6XA80LtVJ1JkFM8kmkINOsKr4sYanXJPWy
Z1mdPv3bF7jLzONCTCNl7UVnolBruBVgCL8L1YhJzw8RUekUfBKTRzlrBejlBVzbpU6ZPnqaQvw0
SgIvOBuREYSvL3b4jZ176RfTCuf2Jc2ieLj5hlYQ8tuVqkv7qKygp2jEEKFNFLrQ1uwnwNTTy73e
FfaZizhShXlVGx739JZZuHFVTIDZAMUQEsufcWxL31p7hrUi2RFJpLNoxDHozLMnodo9NZPY26lv
NXUeaGSrUu3oc/Z6GAhyfaTEeeGeqL4qd1XKacP9J9Qm1aT58RoyEBp6SBgCMBJxX7E/AQmQJYD1
O7jhUK9j/BQYIhavEA4RuKCWlC/RV02hdAXOqB90cqi+9C6LzFkxGRNdJyk5on86egOtecc5Xdlz
HAW2uHiHbns7+lWnnCWqJ1m21PkhXDr+gDjUm8upgVzuNWjhEXjkVM/CQyTqCpw2f6AV3Axtinbs
EWvOhbzeUobPeSB5UEIPmAgU7gHzp5RjOssTVNkJ12/VdL/VlOdVHMr8ezPKp6FtWZQfAmu/HY71
VJ5Jra/ZKD89GeUzg7I+wBuDggnVKhVMJGXZvgSLt/gHw5VJiNTvQTyIAnofsecTprWeLilQ4+Rm
kFy9+Ja9bGK0CeAPLQy5N/0t6zpyY7nmCIY7hbLpimHxetb8Xt48Zr+l+u6EKzwCdvMAWk+xGlkd
k9hbXU82IYjF/0IMY/iFcvjcX6l4xE8dlAP2jxyO4btjBheMpq2sH3WVSLqkscg4FMYWzHYWfoQr
ZjMW30rb7Xc8DLDZbUvCJZsdaSfr9VqJ3WN2ZQTtBvDEIlT1nsbNaBG5IN9Vcg30R+uLWOys6+gb
TnPdTErt80+1PI0qIkdpDkIA/1BNVcMtZBdH65jYHB9FxTlyzBTIGYaBnkN0bd/xxmhFVtQEYuec
VS3T/pkd33ITK5vuDCfJ7lduQ1ZD9hImz/xB/VqaljEc+FE4RnA1KmSO1/YKMOZfxK7544JNngcS
2QZdSZ2VlMf0Ouwy1VX2FDeD2GNG2nctxk03DByHG4JZls5v1EvrAX+aGtl47OZGN/2at4+hLa+M
p/XuqwTJ4Ot6Pk50wBLsfG9MzK7841AlVneLpNeZm1xNq447M1DZ/H/AIc/HA74AljAolpWmpsoY
TtmIwCbiHAGz+vhAywXRWzAwjRnwmDznNndFIuyJEymUNUgpKno5ijDgvxStAJgKep0Ao+PL7YLV
5M/bOQiVSkg34gSoQr8KI1GU/rWVkUnziq++6h2kVYU3hmcRVmqG+Rpy4ZAMVEDgv1diCh0MOOqT
Aw+HnQK++fyph/4W/6VVIoBvA3t9cQ5ewLiOCEBaO8+M78KjOp0td/9iPp6AhPWIvWk1uSGyxTg1
a/ZWzGSNYkVklkQeao2Zd2SKo34gMGHVKcWDS3g+oClaKLfbV1RUZR5OZftF2D6MB9Syu0UkhQpt
f/g4MSk2bjYe/+xEmZtLxCgwXt08QUQ9cl11VD7MIw7qK5G3q/ayj+oZKbfYT5i9G2B0xvYFK4ri
LRcfvepn9kHNMSljEdeAo7CEwdhS4UgnuZTTDMFUGc2tsEYhaAX/BLfHIl3y/f5Zu6jByDs0M4BT
sysJUJYjciyy7glo/HHXMTtessaVDj0GXRVJDcPZ88TCWt0zBltSl2oLtfdAihy/61hKMEUoZYeU
sxq6SkCF3wn78sBHviq/ZVfw4BiCCcMpB6VlBm6bataq8qLOmGsVbgqlLRzp1Aq/U9/Y6BAdTetr
4cMAyo4e8Y7LGzhj9A02WFtjCd2h33E5LSEov3i0mOwIuyy1JPLuT6BLYjDWixLuX1AKnsiY0x/W
74v3GflOMJW9vnh4+0VwbJqYo5o5UBF3sZlZOLaeuH9b4J9wwRxKmh18bvjvAtcF60hZgyIEzTrr
UQs+5lIO0ZVvprRnXXQVuD3Dn9031wiwQ3DS9unHup7nZVbKgidAtReRFUvt1nx7UyfvJkzflq8E
Sal5wmNDyTJo2/LjZBKe8W9scnTTq1l/Fuv9QyAPmDgZRD929cZg6gEzTDADIDIRoToG5DJcUPnv
UusAJR2BvSpgi0UC3DgajU0UeylMhPDwkkgRAyAQ2jdOqccKRHUXnYfdAJaKZwPBIBhSLcM80Zvu
qFoVO0t0rUBdpXuqb6jAQPPGYn4LB5W9OU/Y+V94MLycd4W12HZwon0G37Qg1ABv15oohZQMJhLq
T4yu3SaC5cQyra7bh2l2qFQcX6VV89GH92Zc65vQKGTdbvHmPabG1yD5x7PT+4Hwx/zvd6jBIFiE
RZCGPM0DizEPk9cSb7vXIeN3oGbtjLMGtquq2TYge26bzuz65dVQdR0kkqLY339Qd0SIOCNar022
t2HQ3Eu3Kgr7gwDL7jpLsn9Oa7UM6jZjo5uTXmatWvJrGCdCrNmIn90wipCqG5e7/xRg8sqpeEjP
9Jm673Zm46amOt6Wvw2ZERN59KYaIO4Kmv7+IniEc3FqXoB4T1/5LJV47ewEjyQbSKXmqhZGuex5
5q7QC3X+U+m0PIh+/0Lx1ETnI6JJ4ySMB806c02IB7QLd4Av4cj1uuR/1N5BURMnYCixhH+1hyEV
rRGfP4zqz1dulkylruHqE7c+Y/vVd+1m5xU7kMmDvl/8JVofNhb0uuXEfepXx8O5OQ0/4E1QXf4t
OMSZotRo6alp0d81Vt/nBLzZ25ie2K+BhVI8n8ZgmFOlJarDrSh6JVIprd2/2Wbyi4GT5NLYBNPm
Cy2Y9D87pJCLkjBOZOk3KyREIhFt0hx1vIymtIcJlXfVJjjwyPOviJZHdi7U+TTVyDNyxBhewEuq
8vkmLUDNimxX9xOTfTkGztnXzqxz8yYkSvGGHsOCgtIdQne6AhvSTuOijiTJdUC87uoRBILrtA40
cJVLnkH5vn3CwzukuzeyVmJ5UBehpcXURWJVXkv5IpV8tMa7odbjYQ4M/fETaLX3Pws8OBe9sFjy
e1Owso1EGh4792jtIaIioZfUbBVt+w1dmHrd6N/25EbuKRVKZ0CmIkgAX58N6jwlmWxMlBUFh1uH
0gUaSvzPsZ/kvQiuiEUAekZCzM3fubIlmfqdS5n/dyplxogrB8OwRlnFLAHGSr+vgqvCq1NR7K1O
O1xOaUL0xv6IUXZGj3jFnZNZd55/rPNVZTIKJ0gRz37idPEMtjAyXGgc5EHUbcyYptS4zyE4JUK6
fJ4/36HSDEibniWXVGbWpD8pY3vUUJRHVf7tUioS+/To+KHx5A3r2zByYOUU75ahvE0PiBa+9b1d
2wlPLDv3cEoUYbwecoDaGg5J1IbvppJnQzD4ULQqgLUHPJEmMm8cN8Hl5IfppmluJvHYGL6w6HDS
F5oxn6XPLUEWH2TKusdDOA2/2KWtHpsE/t71JChJcPtypBzmsBNgUw9Gn8/T49a3UVK2wCTfr8ZL
ZrmOcQz0Ml9YwIid3nwujOLwnFbg2gE7X1ydyTsl5PNTPHR7sqd/6EiNFoEDQgNWJOclnioYZT6f
r/rFCTfyMNTOgQ5fZD1J3w+yRsOLj9usySOtNPF2y+IqzFJFkpq6EHy6gZkhSIV9dWcfLToDsBwL
nR4GO7IWqHBCfti3dLjVkpHXeDTUKc2hApNWK3gzpW5/hqyL8nDy3Y9OMq6OdjfgZlNWb2BRj7FG
P2lCmUuHiX7rtuOVH9lt+NLs86TEdSk+Q7Qp9jGNfXC0nq5Fc/tkp7JD1NBEINDBTuGh9U2r8vlc
97GUnLqKQMkSlowSCpqrTNFEMvvt2ChablYHZbG/Tuz9JVmNdWsfjJkxKEcdb81l5jfgs8Y5LgDW
iPBRaEFrHJIoJI7U4Xu8pMGYcP5xdGN6bCuzVaQJBpoTyT7tRitIwz+3kJCsABrOtk2xFoYrMCRI
MS4Z6je+j4MkGFYRrG2scOs7HC+yCdT2v1E9wguDQ6O44khH8ZKkdyL7/+vvdUjsNctYVfrm6jUP
3hAbcp3oOKWilyOgXRwz+RiF63gJqEpwZuxXjkoAFIh9ZwwoeL1pf4kGj8zGYeaOF1EIziRfvrCP
OgEb/C4RxK5DUx3ogOGL1Lhong8+wuKNL3hb84hQA15KTlhieTFUS4dP8zlOzEMJ/NsaSwYgbMAw
vNMSa5a7k9XJcd31ROj0WiGc7BuEIi3JMN2bExdZy/IGnaFm/zWS03GtPmpTLGNfhTkOGBwMS0nq
/gEYgT5F3DaYS+hPhvPsS5mwWIbkGd9PbGEPOA/emb2VU6kY/pcJwWiDFvUTb5Jb1IlNPhTEQSt4
TswlJ4yiNHd5c6uf4l5ID02Lvb7uh+Q0M36lWOkium568VlRfsXxJ2cLz8FFb4toK3tr576Ar6vN
Gj2IzEgKoiKaEr80ImMzcytPZZ2H1jPSftoUDSYiNlHbXq8oCyknRtj7eqigmR4sdRe0ZkFb7OpG
dftOeaaC8+FtymT8mIQe2jcue9LVdoHonlcG1zyD7uyC9EIQHL/aTaMrAlhsKd+4rnHd8HzyEFO/
sus0UIYluP4eaG8vO+wWoPb+LUEg9/Hvh/b7LgCtP4LqH5Fx8uOExH20PNnZRou1sHy+qyUrCcwJ
oVxa9ToCD/Qvt9Xndq+pcTsYGmC683kl/qc2Jic1zFOhxulnlCHIlytQGtuphfDCiZXzXoR2/hSE
t+t+nwIW5kaCdLr2K6jsR4/RENTcsbBZ+UZ1tvCzYB3AFAEfqat4/Ql+UKMWIR+X8bk8kPivZ6qB
gLPJ45ZQUZuV3Pi3aRyYw8E220jGqXASbLBL8EpBudlvUagBYzoW07XO0XGbVN2J0oG1lBB/0tYz
d6F2xoZxqJIPZtofECc5Clsk8uq2C3r5UON1pJaM/eO6gy7NzX5CxIKJ+81wXJUHo1667MZgWJUZ
ggUy6mE2S2OrbVMwk619BgcNbx7CuS1xDrhwz6TWegyEb/YRVZPlm9Q+PVBt5rqIUhhJGkn4e5dy
u+0MDoTnhMc7mjZAnSBEWrCi+Ecd1Ii0Jxv3tIjT7Vi1mCB+DiOGcL2cn5ym+a6OPiKy6gScrvIh
B5n7il5AIfMk42UyxLYK5SooGPkpiEHBkmWtCGHVwW1FLZa+CgJMgqyGEbgMQRq/aOSY4R1WKFh4
9SesovVnzRWjiG5bc+82L1z+2DmY7QKQu+1ObIXg5f0JevertllM6KO3nzvq4BqnKdAc16QhBz2I
TA8CQCDaB3OjDC7ZhZCXarlNmt62CWRHGZ9W71VpaYMjuV/c1nmDeWVJS/wu1OkCRVLlf8eLSYwy
8yd/W6T1EF0Ks1gxnphaxvGrp7OStDZVKnOSucxj2sOatWDUSAWCI8TL0fqSBx5vCpIIaTx5tBic
znx3yDDOFCaB8mNRpVR50uqQdaFL1wnjofqo4U5U/mYkBOrDtv5ecAhhq9eKglU241izlc4tUofx
MR1Rsvi2qOq9ZpTfB3dcYxZs1vCNR7elDHr04x47VuiZ/N76mJUGM5JlDg1OPJwmBiETTgiANOiS
d6xOa6YNFvbEmec7X6d43k4OiVoch917V0V+8PTFt9XaxHRHOhrkVXPR5jTb4tb2A0Detyw7B9SW
owwoMQg/WsYScnqcbVrNutzXRgF5ilL0tomA4XU8lVb8nqf56lxpl+40wpWsyJlbDps+4Ngf0ssg
jv0ox1YZsWKvoBpzxRirw5WoKA4RFkSlXsg1wVJlGaU+uC88Ydv0G7B2iMSIV4cZ5ELaEnLnV91E
wu2YFwPiw3sjPFETJjdRMJLIu4gSZBfM34IjP/KlqrWu5S/URctn2eHM/MtaxMAZb1MCeqesYJkF
dXi5pBp/Sb3/5Fnw+pszjhCk8/RbvujOWV4c0/oT6RN16WNEJekt81u714ITGZ6qmbHeeG45zAhs
wGZooumxdExw2TNcExziSPWkWv0GXuNlAHk4SkQ8RkcoFXYe9OpGzvjsxGUGaSGX33apdfE74TGJ
I3Gy3c/1KKsJXGRCU2cTpvUIHvDXgrFNRNEgTAJNgv2fCiywZOCMN6JSwy28MefUPjsCUFRjo4H8
O72esEUlaYDN38TqEaHl/y4Vs8KQF1xUbXPdDBBxoIa9VXaW7AlbfrKXTRMIRcjmFAQIh3TFSbZl
Xe2AiDpp7gTsImCov7Yw/onWwrbzgxVCBPjFMYB8tESBspK5Ij75Ph8PZvemSP7+UbvXLgXLinDE
qKv+2uTJMcnui+r11++LO453If6kk50C1xr0pPYhzLmN1QJiSVTN83DMLqRMS+F2C5DhacQ5Vvfw
VBJmsDPPcxKq08+6VfN7SIHcn3Q9kYyZ6RmOsEMOGFappdN5lvLmOtQtSRfljBu6K2cJ1gE6uCkC
x+ixlmUBxBpekCaO+gFXClRIb+QdfHdpQN9yAcgDeaZJoJ6Y+L5wYUdlrQcEnNDQkSdL1OSwsLym
DGnlWFn9KXlilH4I8nGSMok/CLgTr/VjzydRnEkF5vm9wlzWFLSmlRP8cSpvxw8LXlnlTeY9Q4hV
WIHXnB5lTxpTKqIHo4YOWdWbtafT82nPV7ANeIyd58xjMbJ/NA81wcFhJ+eNIZoYYd4CJz6258ak
SBAWDDp4v+zd5Rdq5OwCKqILLkhp4yo5arKfRiYYe+U6kUlYoztPDPFaJh+Da/uFnYS8sFzl0N6m
2X42GAjv+v+6A0c1Hf8BIj/nZRnsK1Ziut3Q4ZDxzX8+O/R1BnokuSqOnwpV/Bghn8ksfE8igmFy
8xtguMnJJk9c/LILViVoYVhs2yr8NpumnnH+sJrFWY9qpm1jChiWk3CQ2AygcfrSYl0HdcnMlAYp
M3npxtlamZ3bKGzNNa01p04nhCmBQW6agCQhgCNmwl1sRmrH63zo2sdyKly+dE7+Tc7NMqocaZzx
cCILw+9f/z4gVsjOKcNHbbl202kJcmWI6FGy2nbMFLybzhEOCC4epOlYTSErXftyH3DJEc4MQ+lP
6tnpMjuykrJIAnyRlRA9Y3bmASaJRU6/vAcEqTum2681EswOTSGlZ11bfV4wcRpGIHaB5xNYLcRQ
9oOciB0RkIFj25mMremCIrn7kf87vrvlf1+X4Qaz5J8sGGF4MAyx1aVbdL0DUVJ14hjSfrmo3dm6
BL7hq2rnQ3j5I3y0qB7i5TkLBJcmKSROWndeHWRc1ybeCmHNuIGIGXhTqUklletlP2scEyTZQvjC
QDECjTs38+Bmucxe1qUxaRuLGv+OQGZ7fUKguv5FgobEFkAvJX+wjyJlqB8to/Pa9Z1OOqpoF99l
kWiMZNiVj4uQ4vJcifwXh1WJAYu9Xq5+P401OvyV4BvIOvnecg5fUzuSt+9nQYJsmXOfuI3j25LT
QzYmY7iB+uJheFaVzHk427WAXEkdY4//BXFsQmpsngQRiUgSvQjB9qGG7HDSV/SgXJGwIPrdh903
WdhZ1lv1JZ6bYFpdt8p5rAsS4BubQFD3vlgafXowh7HMeh80JLssmZoAdau6V2Qcd4oZop4lfoI+
EATb0xz+L5JI59K4Z3f0uDYRuEF70s4JyTVh+9eUPAvMzNmWsNS3qO1/q8P+vn6WEf10nbT/yPxA
atNAemegoxW/Ma5Jp3z4m+2I3wi1OWa4eQs5F41KMe3m8aEUWuqGnjBx8BvUXcLx/tjDu0CgYaqP
kGTkhVNdYCN0o1YwlvCjqC17rcGOppXuiCUApwKi7QXLAh+bwCJSB8NAEctgsQbhFrPYaTwPn3xq
ShEfPR7WPQc7WMoL6mSUtLLdHJWW0aD0VAoEoC8GzC8KKFUbsLi1bTIOmowIqo/pSEDB2NUYdAKm
5y77+MSKdnXCMwk7yVyaUzQl9bmC0x98/c4zWS3yxgPnrChYwCnZaHkqCzSW7563gJm4Z2fIv9om
SXXH/bKsDDIpfp5yH4sQ2F38pQza4oqr2gscC1tZ93k8+ov4dSw6osoq42OccJHsEktP9IDIXx8+
MfEkTbo3rggOpTP8hJsMBBGa9f2KibPCSmJGJYh73jgGXnBfIx+X6SBW5XsFSfQJ+JpUXh9PGL3Z
dsCXAx/r2z3Jm5mWo3V5Ztzf+ZoNNQbhC230GxVLZD/mF4XZviFzmA5pYbnCrf2ugpfQ/lRdf2pn
vxwxBmUEnf8cJLv/Jr/6XCJklpqHz930Fe+RzImjWZ9lKAqmeN12K8eYYk7Q7PtC7L9alO+B0//O
jGH63r+wYSz19ofJTDhJvJt5YNk99eiBJpQZPEG+W4JqGQNDZu8F7a3FMWCsyKRKVSTTVpLCklYk
Edw38pZVI5xFEl81NgRuzYNNk43G9Kp2s4Yb+zVoKyBaNzvTTslXRRvv/3E8YuGkxDQFhe1aGZ+K
yhlAWsdgxZQwjc+CVD625xW1zj1GSLR0T0qz1m8wsbyE58AyoIiWeVmWw4q2asOQoXsDw+DrbY7w
OwB6/pFSeUM4VKVq3wTMyqOqm+3lA92a9S1iBP8PTLXhqpPeNFzT4mI4eYrHVXavveATycH84Knv
KHGITnDk7Kb7Ni3ern9GoobqWRjNUZC9+eEoac+Yeue8/NY/z3vdbv/xhacN0ZwV275Nfd0NgQiC
N1L1rUk7xd65w2Q/5k/tHE/B8c9HTewgQ82EvMrG/3Vieg3cXahHI98aGPIDoclGCKFJgYmFdboI
NbPyIih/x1VnMz6PHKSfnT0yizfUhykpTS680jgIcYPmEMGo4EuNS3hSbchwIUSIrIENaVfLPIqc
rAk9zA8yDHDYcJaPQiopqbZH79nZuS1pT+HEnhldQW/z
`protect end_protected
