`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50720)
`protect data_block
T8eXMOMZ3vQ5kabRtfbYvJf/cN5gYhiOANqBRUqUXcT87qHn2xKyQkyxFjCDFj71GJXb9+EIx30s
Je+MPFjuEHhPlDe2IBLkmSDOtyK55k+gDyOkGPn0Kv634Sh372cO0rpe6donsoYHNsTu1bar+wU6
KRr2KcKipw53ACKySxDCmV56i9dhagEp+EQm3WcOsR4SiN8Za28VmfusGxOwQ4npYKRLCBgmACyT
K4/hDbBgG/iFUUIB5HQU2pMvhJeGGbRw6Q8jaVv5pkB77UfswVDd8DSDN33tto5rbyuE9Cud7pv9
Uvh/vBgWeX1ILHrFWybMrdktEUX5c90/2z4pf1dOENnv97S4hNmF2uNloAUoRPH9tKGATwkoG8xx
2ATPhpkMr7c+g43k8EAgm9Ioa87WC8FyQ15P45q5QsQ/0nQh9GA4vQgcyDkJuAszl81LNfwfbvK8
Ma8VfOKqMbT97Ay7sj+Mkodggts9d1h/y5J88CexfJ7leqxATqC0Ilg0CjBz8BFV73eO4tgC4FNi
j13tUv1tRUSJYfAlu1glLynTv6gTQi3uJrC/D7h0Uwcs4cBEF9aq9Ui6ZlMG+6rdTQDBnuVuId2n
us2bnpG97RzvDcFsgGRoEmaSkTLVygNuMw/JX+S3qh1Q5YOzCGdHLreb/bFFUNO3nDrGe9TSUGCA
yQ+GuRf8X96f+lFUci1cL5X/RSexEzTdZU5bkZJ2zirnqELgAkNFX6RixXSNDYiiR1LZIIQI226z
xKrQAku+a2eGTV65NMujHef5XufOIbVtvPbQX+gPSmFAoR6p+KYK3dX2cMNfxsLigm4m2mn+oDmT
lxxKL6HERY1ToeL2Y0FMzIHBEKadDLujAHSit2h0sbBtgoQ+5532klOMse3fsz/HryhK4ZTVKf2z
JiciteSk16+2NH1VKj16iJTuSNjbVYCWyOxZ63NuuVuByABmr9DDer/eB2LECIsb1U9Hr8L5Njke
JGioVaRUuIVO5BHowDyAddzOGX0mdiCaoceVlsdVo/4rjwHFKW10E2yB5fSaOZrSWXkl5v5ZYOYb
lwyp99bY3+3yhcdsSnszFWFOC5dFJp1GmNLOeUvA0uZ8Fkhze9tvPVeee54wSSa2JbHq6aMcLg2H
GnYSFybvPLOAfiJqxp1qoEppmDp/358Y6t/rEnkX4iFkM10SrpTw3e9Vd6bpsdwAz4xP1/lBTBxx
C3T3cAzbXiaRW7wGCHs4eZuJp1yTgZ7V8+DCiu7ld5ogMdx+XQrxbmPZN3FwOJXuQY9RKtThvB1n
Y+9SWaT5ZMSW2a0KgdGg4p5gWukcoNPZIzF1JZ8hVvokkO/gasiBDqh+wZ2bvvJ+0Z90NvcmZbVV
QQgmWwmiPyTBXcp2Fz28QnSP55rIvO8amDkK1ViMHzcUfX77MhFoIdbLoCrGCYHyCT/m3TZZAo/u
PVl+PZHOP+Cj2AwbrgSBfjrOWUrRITeQpB2Ziy7XhS98xUc7aNiYVlYM3xTZGlWRvjqojuuZHBlF
GKlWI4HKxHiQi0y4+1Hlt8aq6xT3SQHD3QfWBerW70UBjQm3c5w154ByinspuRqjrKzDQ46OCdwu
wXEAOy/li+i9gi9ZkIb4WxJD90abNlp2+XPkwzB1MaPTGTnG5vK9BEnnUeaiNbY5/DOjHi5nEUv5
/TEgWwqrQiHVxkCayx4L/YoXj7e3MIBFLIlPOsA5kGsJvxIGXJY2J5wAyb2nvOMABxgE6MACr1/8
917UpN52TaMSxet6iwzHFZpgQMJ1JTkjMAawomuMveZ1oMg+hGKNIOQ1YvjH/oS1fu/WlBUTM3j3
NGQaBvzSl4SI80aBbJ5Jrhex8qKmzE14rtDQBaXjPWfMS9GuojhpH9FdvxSsTnEDN1greE6X4Uq/
85eodXfNPQoazHzvyhnpZBnWqkeA71ybpwrrb6XYP5isX3isLvD3dSX17rcFhJFwaMFkYlFviuII
qAWv7OLv3cXVCkBfOeebKRdDzpoiWzFGYOO/eensutMsPZZntmdqwgOnRQmbZLih8S8sK7nplSnQ
MMu6hp4IV+6iy5PCGRgu8IvHWlJ9Z/5K9LqphQt/L5D2WPHM39K7DVJaitVk8LSfh2zS1XNo+2mf
7nZTxZTCTLx7QVprrIdpmwP5zRY+I07gNCwLD3fJcD7r+B91ypnqsNdtIO/NcGjqKpT/AUiL3tVs
M7mgMScNGe2wTSU0m3yGyxQXKXeKp4vOz89Hmu+7bf+T7BNZYETxlGs8C7it8fEYcIA8Hd57MePt
SyRoiq90dn1G7TF/nxrf+EnQYJGPB7wVw/WiwRJxpll5IeSqfboTfGYIOYwvmDsGK6cznE5xsQ/c
hrU0eVRSPyRA8T+uqvYpbf20V6GiPKxeMgbRbHJl4l7Dl/DzdlQZJBxKzc+Dy7GlZ43NLuzxVvNA
RAGWizYn2MeLhO0THIhtkwlVP6ss9KOxVfIfBiiuHcOTutQ+pywgbXOq9DchRm4EXf5l8hvQg6uX
eymjf4okJAmhVyeXfonihGhv6QKYqJYesMgEV1SVdZ+HQDY39WODb0bV5LFuKWG+l6o+2unLSsyI
aZyM47CGYJWyJkjVBoWtUv0gN5EsqxG0PuoRNz3W01dvqeeXKdSWMK7BOX8aeCwZYE5KaVRARo5W
ZDm60oWoRSmUX047qEzE4xe2gWVgOvdVyL2iYM77oK1g/uiXG+X9qTn3bPM7PBzzHC0nGVmy66PD
nY60hyv2W1J2jUCRBxERP7tLtZWEtj3k0jQtY/DDsLzb4TmjxXGn3qnjji6fflGQ3Pgo0TaZMISH
zz/qDsGS1iiRhz0DxGdSmUq4kZIxGXbmUBs52dR8AZtskmcUDdh015ZHjDtHILn7jK1PfbvIdn39
wncXDg9F/6kPU1ZacnQMHPT1iATauzYmnYkP6XKM/ODG+q84TboaKOU8vaoQBne1gM3E9Wmx1Nfw
lsbtNnkzg+1/YFj41lltSvRK35Dc9px2HJXWD6xXKRDOpQ2ulcN6cns4FKvh85q34i7fuqpPyxMf
AUrJvUFswl/Q+vp0ACJ+8ETg5S/aAKKPiUVeMHJ1VHxP9L799H6vG9lUvr1xiO72yHuVq4FPpszq
bSywCy5UfmBzhFgo/b2hGD9BdzZXEsiqjjjNEllYV01tqJjh/c8OyeHA2YQai1XDer9SuoEW7dnq
87cCsF24hMqB54jTXh58qjofSAN+EHhO23Map6CwV+FWf/bGOV7vRJYj7G2NeKp2DVB2ogqOSDfQ
qBGAYv39T+A4/aEKwMAiTYmf6uk4zU+tCIFjDTmMc2f/3XoTcfeyt7PAU3QOEC21wThIHwl/FQex
uyKcyOHokFvPCPW4GNQcE363hJON8I6CwvEctZj0Fug+beuWKIvhBoarlA8qCALCcHLPwGNprDwj
TauaJCDksDV3ad4JTSFy9KlCtL/yo5Y3+1OrLeB8PD3dp5n+RNOm0ngVz0bKqmXYQJRU7iH7dxDf
HvqR0LYUZzg/f1FKvrD6ngTKCZlgPQccsSbL86wPHNlrIUADOjN98S0oT19taG2gwM9LFjIj59Dm
9QKwNqqAR/fxht5+ip7GmrZGmZQ2wNZstEzEFtXhcVYECYPfS1xkqUZNlq6KbIwSwMp0+4bYeY2v
EYiJlncaXSrHxnDxCxi6g9iAM+ZZu+xYqlL0tyRGE4dD1B9Isw1MBFUZpHvpfhIA6TqFD/0DLymc
+OIrHy9VnNzNJNqd+Y7RjTEd4taOh0BbPmDukYbXg3H3UjPTXSRSFVKH5JZl42QdN9eO8HeNa5p0
K4Bq6lMT8wGZF2f3JD5njXEnZeTFolVrUmpPvpQq493F4wNBASAM6Ogwbn+hqKQ3EmNtnbfB5fM6
njGPCM/vGmrBssktxWnrAadBWmADPN0DUi2iT7muNRuMgF6sVfDu4D19WcAvAbhw8NkEBWs1Y0fx
oxeZnj/SQbqnw7aGMklPXFHl2fQ1Xr5Nvh5laQky80Xc7SWDf5rcT+gutJ+2+dln3F177wK+yJ0E
IFgRjX0YPU2xmfM+tO9GRctGu7pMZOYL4ULtrEnKqEzgbCmgZOAw0IwbWcR7rlzH7OjErWEhjLOC
W1lZ6kLgW3+JKIEcAJM+Kr2ctMVm7YUOCQHnDcXwQuoloEZ4JCI/e17Pb4iKcvtQ37ecfOfb3CxX
pcG8p3Q93t9DakidtbzpIxrgyVbp7WS2E26Rk2C2nOKVhMAfiXcKJoFu63Pys8UpLdAkRYGkzzOr
si+lHf1GLrAH3PNbAq3EIZvont59b7JmN6bUv5WwiXa8faPV3unsWF9I3vG/40SOHQ5ALAzyH4Tn
DRZ6xamj4NG7DqAaOgtjximZRETIgEZFDjdrxJYzSQ6hyK5/HKqeWDjfPC4ttM9cqltfMlhwkICD
DSbEdzjmM0NynqPkZpZvFoej12cxGfhoZHoha+fEIAotWCDt+Z+3/GFe4T0YfuEG1RsztA/LTR6I
VxBvjBNAkXqlpg3h15oyqGntXAd0REQD4f2T7WrNexxiA2q0SrEwp+VRHSb/+FB6SHpCAaGFUNhR
EgKhhMOAqw24lRs9uy53OyP8+7w7F1GqtofgsPA9yeuhAIQtHXpeTV6vr1fTQt4yK4jAxP0qoM3I
QMBYsQMI1/Cn04ZukcUCp/Jl04TGjygWkKV8aj4AWkN1qQzGkHQTsjaE0H/P/J2AIOo5rH9AFZ05
Z2i2Z0dTVeeL/lMOixMhnPpdV9YuyPSm6ejGLXKUNDwn1V4aSlDf4O8nfaXWyoyzDBHWL7ZLtmsi
2wIBtj21Nz286LNAlRvEyXdnE7aPJUODQdN/wLRIMnki5lQ7oR8rAvpqpFg3V0LVsbql/si5OyqU
MI4mVUvJzNMMAuUxF/euRiLlXjNTJdh43m4RoMfKaXo2j3oNIzujvvxUOe6BPYJo8CZfQMr24Qup
6tXJlbFeFgtLKVebLqmDUFsSU5BgBwibaw9b+lW/nTW3lRW2HuhMs9B78xILN04of1/nzfd8Av0S
SrcJmhLQTv4kE79v91H7X0OresYFcMZpUVKY16RKaJHjEg8b92nYYLtjRSFqt+7Kn0C0Wrv5zrHG
9i0VEgJ119R5lhcgUwMRUZBVLMZSNr83pz8X4gqLmBh+S8sd0CBP7hb+3AMMM2zM/cuI5lTKeoQF
HvGxGwrFODPHyvn+NrsjSrYPp7VtHDlp0K5tfQYokjUNiJ0gPmtW8yYshK3m3fVmv0Qu3U46qsc5
3wR6AP64bjpAnUaMoK5boimMi2Z+Hmqe9eJt1ncRUD+NF1D8s3FeVBCoEKmws1B68ZZLvA24LRYS
U0X/a4udujKQoL7HdCK21ZKSzpOUy7TkZGvDW8h1WKB3NW+oXD9iRiHp0VqbIaUdbHz986lJKOB2
Zg1rjnLrDZZHCxhL7+maCOEWynrEiwDtPSZ8ImSGLVVN84Vju5ZkrPBSkwbk3rVC/7ItVD8rcLva
xrdyeZ3FK1X3FjZ74Zt/1YChqlaAa2wYUWVkWkIcJAHGstCxVunSq1XQfjenBWAmOqJg/G68DJDe
384/V6N4tSWXLM1xLvzZFNFKX4n1sw75xjhsbozmF4mL+/kUFVvZCZIB9R7gc84trg7s4k3nvWYy
nz7WnuCWag1HUo0x5xWHT2xuJez1sdoFcBnL6wPw1sv33ZnaKiPSc5uwOY6ucFbRT54KgMBklQON
8K+DAGEKZGp3NRAY59hYULR/+rR5/Ioh9sqMODFt+QUqu2xt7adZz7YqDztLbqWTf5wqeywuBoNt
UDqRENsPtfqHof9aaXN+Mq/lSDzGRI3uJH+nD6rRa0Uuo9lAU994M1K/AFqtBqyypiYVLngx4kDC
KRWBWMfYG3LYD1U+fbcfOGQRN3lQWoFtcPt9gB3qfDjuKTdR4U8DH4h/nsTtqHO3UbTcYoZx9KXD
o6P3ZTHzBKGbDjgPow/UWk2SQu3XKcOw86C+4vBMYOs/rPhPYd9QQs8jFAxLmGf888KcWTwNR6qt
H08h4gQeIxBdhxp0r1BjvX67CiEe9DXwg8wunkYbT0t1l+Nz00h9X//IXGHZUl5qG+egY5RCupJE
zR6AEVoQWHlCp2nfM8YpYjC8AfJRzUNwEhXn3yDtIuAX7vwbh996F5MNJU99raEvOBmgFW/wR8Qv
5WJTh05XtSIjcQ5HLtGBuhpzni73TU2uzN+w9tkMUCc03r1KTOCwkOj/lAy8qVeqdKRCTy8s42J/
yTbIMb2dnvLuT3VJdwVEeMmW9xh+Xrbjtfabv3xQU+Nrfknk1Xs4hhkXxbzkb0Y/9rOc0E97NooZ
dmn/EXA2ql4f3tBYKbbzeYCNczdYnOv2H/8m5qyGIxkwAvZUBLlYTVIMegYfcoMmq4DZOzMff6Wg
OFfvxJCDrnvD+AL2lvcg6NbBAYQNXm47oXwdiD9+C7bLVyrCiG+1lyYaXr6WwoFRq093JoVIByaC
K85cOtKBKBwskBDbH4GVCSMdgomZ36lj4sV4Ck9Yi3x55+aHsRZPbTsjiZaC4MDb2dnslLshf9fU
tdKenMh2RMoEnAyHSF6zYtT+Dc43eVdIR+uHjOtG7Yp8+En0DUfGaywfF32TtDBq3oJOXKGzbSiI
wEY4QCzJ+S2laJC9Y7mcDnwvYm/y2l9w0+aQSf3CM4LHGCC+5CeBmIYUlIOzkC9ja6CrDzvRGQ0j
gC9QqF5PdJPyyOe/Q0/hPI82Lh9WbGyHBxNU40R8bgu2eTbakAqOYCArIm/E83O8ExZxwIbsAY/u
h61voR11ksDuw2dMk71VR3I/BZiWTjm3a2QSP2ZOrdHkErQfwaxVSLCNJD8sHCrDN1lfHiJ5b2Y8
f8yWt+aG3R2fiGu+5W2r239IchtUIFf0z2Bc6u4rDtdeU8533CGlrabBaCdSL3BQkK3VdylgyUbj
qLVx5bqb4LX2IIdkaGQdHDxzEgGP1xb4T6qzC6qoqZCpXyK3YInfgcP44GslPlky61zs63Vmk33Z
Fj1y0OMUe08+4+XGLewlv5gNdLdP1NcZibXM3p0ss+YwbTIa86bMaw9q5cytsSnN7Wa8Mv4brDDM
E5lSOQhOGTGB+oGMisI3Q00L3PmT2Ghrx5ci+9QhQu9U0h5jW+w7j56Px+TgIJWH5TbGbgojlcx6
bS/FGmA68jVTKN/9IHeJfd6aBgNKFhfSXhdqCxxdp/ej7uM4HnK5Ah9KnFNvV9PURaEyRDCBR5j4
Xtx1DPoza3w0oBWiaWr5yDd9ZA8DJYGY8hnhcvAfi8nEEpJ+53pPV73pVjXcUrBneM2BdHJNnql5
8BvhtinTqdeV8VOwnlSa37++1RMOpSRhBPB8eiVYTs04HC+eqfz+4cAnM6hYfbk8lkC/pmHQB/nn
OB6LwQYH7R9JXw5b6ms7/uTe7R9u70FwjM4jSt+TSeebg1YX/RBr3+qnuf+j5ampTr1FY6BqgUIY
UJ6+96ncC/jwdE77RpLO1a33iRoNlVE7QbiM9dVRoK3nhUak+r+OvXKYSrqQpGDHOMlmc5rjgOye
njzm0zehEet/9sHKss+9UiUL+g5kfxXOZgkuOtTcFzH+11bLPbrTzOcIFnwofsaQaur9pw2rOc5a
cG30dcKoD8AHnnhuR4DtLEl4woQVeJNG1evJ2D8cFpBwql55lBLrfLms9vHNCwqRlQBSQl/Z5Vje
qFh7bDSzVtwjlNhV9aDs1WV/knrw7T4kuid58uSXcVjp5Fwa2fISwZ+8BlQx3ehTXjHoOho0nXSC
i3wG28NDqtf1+fbKwGYWlvB+Euo5QUFOoTzO14dFkxAQnVMyd3o1Oab9LvXOWyaL1ltjkEmw5L1W
OoPeT46y5Im04qn+OWFf7Ws2tpJVQmCdEpcJRgwxUtANK85+b5+jSg2VvD6EqBblQ0lFg94PKTht
QeXQnyVZWJ2/dDGhH+4uhzdqT2nG8Ed1Xi4Y7m3E7RQ+Gnju3g1CLWHx85mfvSJC2NihI1Slvm03
jlcz4fWcKtYnfM4QMpTj3IzYR2JXZGA/cP8fi8mI+5mjOI/B002kObCgbbA0XZfILku3HJ7pFFme
Q7/yNVn7MKQr5ZRq4fU4+RLCjUAOaN6+9Wen4WGN0djKHT9qv49m5pJ3P6CfGUumCdI+nq7CGIeR
k+b+qYKgufZS3VraVWi4Nr4bidvqUbfIAYedcImvzXkv28jSG93ncnAZU3FmA+3BOyFUTKQJidmD
qjtPBmYv3MyZDKny/gwJuy0IYdShZ6/BgpfalFvicopWwSGKkOP4Ox21AcYHN6QoOGfGvSYpVYFn
A5s4c/gfC9tbWhRz0ZWxNKQZsEzlw160fZfq+VAYt0wUVjr1GfKf9W3toQS2w0FxJfcVsKDQd/L3
1ulbiFO+o2JTeKNE3nmQyOqyOxUpeiixmbdT23RPlfSOn9uO5nwt04MxycB+fY5+bi6riO7xR7O1
EIjcLCI5YAQOyxbiodfxivrfIcbp0BVYXH8+mf+Q4psMNQTcMmamPWhFvJpCReX3gMCBsL9KAqvt
XkqpN4NlmKf9jtDTQuErE1JB2GaXkuT9QcdirsmouE7dXuXuO/qgPIr3GVoI5efW6vESSsIEnVJx
hrDQJfLhw67S96e4PiuOzPq6IifuulGt7mYPuof0TcYXBjqSdXt0EOwbYppMbneCVmmB2tEbGpI5
2O4b6znTEQ3gA3olk6vaW2W1lWI0gB6RSV83fj38BcZdp1Pj2r07PkPxOvMLxyjjPbJ4AKj2mfTr
PovcatXCWJ75gtcZwsEbokdWxZujP2bT8DUJhFJdLQq3BzopPR0DVvEEplNkfK0jynD4lsQNjALS
4oDDpCbrP8SvoiMyqY5M0b4dPXnM86ZLbIu+9mlE78Ykrb3zZBUqxLFBWiW4ZOtlswSKYH0cFfip
QryGMWzJzSnY2GmURUYYwfEgiU50ychD7tw7qek85v5BEguDPZSHSatEAn/25eDySOGBlIH94QZV
z5LQ6AXn75zY3ykakcwhSnZzR+akFgL0NqMGiG2ace9lj3O4XgVNYZy+lU86TCyO5neYdnj2tJoG
1ejxdeHenh+lIvm0irQS7rVQBr0oBYkVPkfNKLU7kkohDRqyjqfzLh4K/6ZIEb9ajmFoz0DgxA7h
qpE7M50wCHlSidVfVEGlBzyUKFh8YdDAG1pudel7uVBqCQBOHPwNchXcGbHfII3fac+CH5ojGMy9
nVlWETpCv0bJrHRyzKeJWmaIrK+uMjtwwGjpNY8g+1I/hQlJCYLD5mPDUyve2YgTFCRnZuLHlawB
9cFb12bNn2NcddmbdnUmfnUFIAkMGv/Ex9YgN5T5okfZ7JSnvKpWvhvG8MwR2T5hvYEY7hYi2xtD
JkKhlbLPnlUxUmFLbjKZwP/2JkGWq94nEYksmQewof5wgGPgUxhNAhq4tFZc5UuqR0//Mea1HNgD
+iUTAclcDoj8gP9gOlIuRgqRF9QrwgFN3u4Ll0hL0xhmxxxrstVpj2Z6BtVqXJ8lxJ8Ga0NQ3wtm
BPXRn238d88GIPO8m4IeocT0Z9ExVzJvoAMCJBylI3RuhzUAsJJWPXmG0XQWKyHfokQ3XZFJO7ij
orCRVVHzR9M9UwDdIEglgAfIxC8ubAjL/m3ruGLotnoFC8BNsTo3P9+we8YoA3UXGHmIjTSeceQa
axMlmAnl/jFw9FWZW2b/A5dvRCwNYi/3rburHm/IE9l6uB3ICXZ6ubp6fPzaWgOGPNMXPpNk0p0m
VuiTApdvqc8Zrp9G5E9oMQCCgWKMnxK/Hpjl34XpMAWpSuDsJ+yAgJ3LASGSvHtNULkCFOcT3K2H
78FZ0PWGY0mHC0Kxl+uvAVJblKSU8+/p9mthkJz5oZbY5RYDItcQzpmuAV2zipQ9Q+hKl9xeOZfr
3FCxVp1BdObEH4yI/Uual+4DBLUb5oFYW0ABd3Q2F0Fmr+Gtt8mkvudDzE/wa0j+c6Yrd2suwdzu
4AockvHVEq6CfiLPKJIAjIrx9PfhlzsuUiKg9tW8bq9lKPRveuox+BKoHddJ55raTp4IWZWj9Zex
Jd5MQlhN7E2IB1RrvBWpOv5iYoDZvyq/LY0wqJtOWEoVvMQ1Y0bwMHdid26guzHh258LX751x22F
DSSQ8EXeu85zUAQKJdtfmVdeUpXRhDDuW8F98r252pdz6773cPT0IasBtK238okWsRoo0Lei2Vnj
x7XYQIqC2RgBtjtkqhTKBi8aTHm1v5T3xAlDeXB0LpSyNZUnlW5LTN+439yWxIw/C8B1t8t9CwUg
GJZiRiThRh5aprDV4h0XkQ8qmG5jNfxU403adynvPM56gAmOgdvIfxEINUR42PJv9vywZXj6HKRd
o8l3VEHAEbMLvGVWoha2Emm3PZm4bPjXBu++bpCdGRIwIVZ9Jm+lnBU5dAl//ehsioGhOs0KqeFO
2GQ8PO4ehhMe0/mXehGAPQ/W37BieQQWhIy62P+8R8VS4uJabaCscRaRObmc/e1d16pAer63IGUm
Cs+UpPm4wzof/wvH6n7W2CXnoJUpL7iPuvgHeGvswKZyNnj/DTHU1LjTCeOyV34uNZJvrm+dUPqB
i5XSzS/u2JuAvv4ylPPjWRpWLvQOy5w4cUT/SfBlQveELb8SDZ6QCrfw2I5ZGiFckVbdC5t4ba2D
m38YBKYQC7r04SNMmVTAnehR+HuI4QFqTYvRjmCTbwYy4E+KLcMHVLIRKH1HrwbqaTEP/1yMhdNO
araW3jJ3u4d4jvZPDK4obhigKUxFksKaOOgRQBqpRjDRm4MmCK3c36ga5JqSQhJdl4AotzJ8tHI5
C11tFAPLFRWSY0WGNLT5krJUig+rYoLLMrCs3lUzxTrlAQXZ+HoFmJ0wwESYg9vhclk8zdHkBHoi
k+b+JcISw6GJYU4NYmEhFWCaPHZj9E6Ru4lzbu4SwvqWhFDfJAM524o0D+0SjFFgYqNxynKRYRk9
/hMvRAguNUyDyqKIj2vIFTAh+sOvWUgHXmaZCpoTS9FyszUeIFOA6n+GpW30cZ75Ab1PyJylJUyy
lSjVJk+LUtP/8nMsOnTolVxZRrAZiAw0Bxi7eheCthPZThTMi9pQVh4hE/GS23VsKakmP6yZKFkl
XjjY7DPFvcDA0IqBjYxqIboy0pUbLbiYW4Y2EDNO1zYLLJtTizxQ0aN3ijc7oENVHgx9oH+oGGnU
JtKEJ9h+YEd5jT7zldEfIzzS/rFdSuACZNz5Jacaf/ipi1S5a0SXEuYdTyFjHj6igaxqoxPjlXrI
7S4PcH1yB9iQbVvuW/dYVEWxR61AcYPH097K4Q9pbJYcQyi8G2nuJflTIFTj6fxIBD9jx8Tn4Dm3
ZcXfiMID2o4zb7v739LcxaNHhvWuOLrx6PWhD+GxHe5D2vzYTQmQM0i/2JbQqHZOGyomjBehPpuU
jX9Q23/il5JDeN0kXV/yxb3DEpe80Y8qkngisEwAAQQrspgJQYDw9ttoZ0F52sMhFw88g47dHnq/
hjgdsuef7A7fRoaYzqHySVivjKZJYKACq0vKVvX8YBCBMU04nu1SMuhFud569P9aKyqR1AfybDOL
ItooLizysNeWs8RDRO++xrwtAiRUW539VqfpUZgR7V0sF5nxRKYlOHWT1kpOzEbALhyX6B3q1cOx
vlyPXpfKUO2IApavqXhO6xwqMjPSZc5opcHkDlGSoCEZcRZUFKkSCS0w/h4GsclcBehi5NqCvmGE
lr2NMURMp05mMEqHRkod/Sfu8YODAXGJp79HaIp2eLLKbtMe6jKKLMJKy/YyMNVVX0FTZweguj39
JdCotJN61GCk/kyNJH06XB9s5s6uC5qQyB+yV/6Blu4e/D3gR0sH1/CajuxoE0phbT+2ZRbsnrK7
fsfkactPeQvorz9db2R6L4WjPt1j43MHeSwW+wPTMrRvvjAR6UPzHdfxgLymwNK0dY5uaeoRAeGX
XDNC00eMFX5xVFZdgECzph5Vx8Ddb/eWmhLutA5fEykc+DvUqK6jFRS7XkdME/CI2glwq6mrjy08
reAw2T4tPXaEA67Bo/7Su3YwR5HLjKG1/mIwjR7gGPNQtsL+JIyAZQneu2Ptn/a4BxY7pM2sx236
CUydeMfNLc6Qxy6nYw9qEBcccTMqVgNo5/wnN45qTX2VhKE4rIDFvsPjVqUG1ol9MTgCzxKtMYZt
9cqM5fxH+zMzt7ICy0O7Z7fY4NBtcTUo/fguz0/obC5oLVkS0eZ3p7Q/WJ6ZESBkf21w5vyMFHhG
Xgl1L2EEYMS7PvguZA4/FglnKcCv8vwweTk0OftBS0sGYtRYGT7gN1DxDw5mGw/oMHTItn4mUNEo
ZVd7oqDhxFkLzM3qV16QzrcdmcCaLkjoIYmKaIWEMf32T+FfsLl0iiP17LDz+4BFtcRr3KRwTELZ
bVYc65tc1vJ/9QBkbu1P9DXks8HNFC/2VUzad7LJmd24YtDdNFXSLc76fKeBNl90GbK/xZbRq902
ay3tSHf7l4vE6tlcsNwRPPqMy8qFSPXtyCPtOK4y6P0MMTtOg7Mp6sG1e9HP9r2X0XF8Gyt1RoKL
tj0bWM/YMhaJ9zlqC1HxIvYFWWvXr6vvwUiEWJEa8eZl1X9bUUVEZ52IOt23aYjrcRwLYSt/fWJb
PTaWRxrwTdWArMxW9hrsnHodo8adi8YgZ70f3IY6CIywHSwxtG+wW/DNSP4rXB1+jYdlSHbf5M2F
4ETLZk5f3Np4V2sZBq7zEp0Zz+IHLJlonvKbOn3FCWlI/kWmgtT6r3ko9DpVln4Zklc+byEW/RqJ
1fnc4FBdGz6ILMF4impwS/fiaCWfsPWRzhA9QsdD6Bz7E+EyFgiSVvvP56Dluvr71rVkFgwqarkt
EdtqbTknv1qruvTUiBz5MgnpGzzxRlhHTKohvEk5gLrNXIbtZGeebo5pyF3jTkp4HNke/XShthRJ
ajtLfo48i8SjD241p0OpYSE+bBVb7mKOJZdyx3sr+JjTmk0YxKQJWFYGPeQthJPczsiK8sYhniHq
zzwUwb7FBzleHi93LbmNaiMlImDUsv3ONczlA5KPoQtnH6UB/tw2otANDLfOifWQp7JLNsydKEN+
CoVie+TGMJAobaJW56XifdNMHyOR9a7iuJdh/VeLdWRYUeVQpny24mPKfskb2qqtF+zzICt78AMk
Zvm0ZUcCOl+m9zGfwE9CcuSNejesQHgTiJPi6Z+5KFIJfz127RUqLwM2XHWUUdvoIVyCn554TsYm
gLv7lyDzRnBw8dbIC7wNDF4wBCj35yuu7H7rW8B4haKuWyIYtSUCKtWBxqB0GxhMVRcdAHke4lDQ
pRXVMXv3KCcKSNempyk+CJnOkZUB1UTfcS9p9y9IlgOIJnAJcEcAG4FkhD/1QnBFe16w/WUmFcgq
eRmH7nENnoKysBmgY7J894uuoqbM4Zh8n//Nos2OLCQdE4aYBd5MsHnIfq6dvZeb+5V2Nyxj31MP
Jcv4VYu7cIN4faG5WE3KlAOVHvnfxgPXeHjKe/ZVwQLEQWTt4AG4bTqtEMAeXIUnmmGrw155sqHf
kuTrcXMGg5JmGlnNxnw3jvRLzusgw5sctTjH3yjuQmEsxNJUaHqYfpk80QtFmqfBhZkM7RoH/w8b
EWMBLKLEZPN0HuFZfcKeaM6+2DkvoEwVoabDjQGpmbLnyF9CqzXuUoFltbtUZGR041VfdVGs47X7
5ylFYqtljwhuG4eTSGLNVtilkwNI/Hh/PsIT5j0eUNuPRmpwUA3PThCIvHvNJ8odlqL5Vm3b4CUz
WMelzqfliP0W1qzPj2gLnwJOvobKj4R3gqezrTzH50j9vTGuIZbl3qEl4Za/etcHMMZWnI2cd0Y2
X3K0fbhpNuUW+s0btO67uXS758nRXVvk5f2RDQ9jzXc87MjkO3JEBMbuowPo0SDgytufcxSvGAqW
xnnAX4bP4GX9gJBBMfCTjXDNpXA6eBRSdxi/79oUhnAOuTITsRh1bO+6anLfckplFV4t23TkuchY
wTXlm3oTXqHRGQK8jaD039Yl1Hm/uK39ZoWLq9tRW9baLVL4zd+O6CjhxvJKasBY9qpnzUZwlLFK
61Dp7zR+RyQhZs0FPy2MNcbvpcIW7zpAKcRiPO/h5P06CryjyEu6Hxz+NbnGQUo2ss9SXmHvcUAX
DfWkoIuuM1ITpHoGiLIbLtDeeQntheR8MAITgNb6v1hDanJ0w3iqKf3Z6nY9aRyyVGaxBQ7xgT0U
FX3Dk/eFpTCKjSiQxqQxPu6ZEaH1bEesIlBKdrbhQQ68b2bMHJpFpD9GXSuknmzYqNZeySigNzak
bG8jJBEP2TWsYTYNqVzx6VJCbH+wpAIBmLL4JVDqSA94dC1lwnEHhT3UNOXgSdjdeVpmooBBjijh
pfaw6KQLZnBeumgJ3hqiRXB4x1S7WVbpNfHRF+M0SgJ5z137q4Sx8ldM5qMVe04PLTgpVF0SQpxy
ST6jzeRcatucgVPxL21JAjGeAMBZkB2TA55DInSIW01fApcYQkMsX6B305hozRUaSS0h9Fo0rmnP
K8U+Dom6Nvk/vxDKETsEATcN5/+qiyKjX9xI2TEr0EEK2b2Nl2r+Xn/HI8sAF3qF32X62McH0ik6
Oa9rCHGZaBaxvZ9silVVP5mpPBCqH7Zsz9TLHhviyzXfxJtkg5pTnsyCkqWg6HgMjYC0NLJjz1Oc
2GDYt7p4m0DL6hvoQhas1PKcKdpXrNJS1d3FWkNdkhmd3cOLW1PeeLH8mCPTmSqfe5BNXfbEG9fC
0hFc4qSxpZnEcr00O+19us7Bk4FmoDH3g6m8Cszw+u2kCvWOcaM/7Mm0dtdtdzXkPuPnvRal+mUe
BNqKjxNHosnF5pENEZjkgNJWi6ycMgaVGZhfOiGXUwmNkZEKd0MXkQXm1mAWnQV0hKKJ6xRem6Ap
iJXgbnW6F2QgxXfcKxkuDkZ3j3gUCJvIXZMxr7gvAEuFhvgHiajRV3Ggkm5BMW0eFAnkhbPrqfsE
L/apBeKCLpYeqIoxAk/aag1Tn9jZNOLGe3N/MLcBZM1sBg6KvzwktKInjxJ9lZENZBg9BY4sA5oO
52fkWqUTdqcfs2B9BjvGZg/kXbo0xDdPcQNoQaVTYj1i6s+ByQSM1xxHF8OTKkd82+2AK4XKk0kJ
IZFGmbUAmc/2oOvabFjd1X4pzXKDBKdn1TxAeF+5h8+9EP0g0WENTvzH2cu1VivChuG144hWndU7
JnDlyIt7/KDew8EXVm/YIzxLW3V9MbqVd6sVX6DbUn17Ct4aqJ7Tnsp5nP8mw2JKb/6zt9QPfxDZ
luHOK8kMEe3lFtsGxiZxxOB4lpXeJambIxqziUuIaG0kCyY5hP+TdKXjMjDh1f/AWTskbtqi4vc2
TI0JH6S/GayGIwUh1Oa19M3eHG77qj4eqKoxJlASAp9uoMRNufQLhy0MEoIcS4LmAB6It2642eVz
aTaNp4Gx3GTBtkrVZMv1Ym/1Zb+qNrkjjKmZDW1Tkg12LSxIQKVsVZ2o9WMEr8uo8P7augBdKZEN
lRVqMjXwYBQ6kpSeCB5C2K2+JVCIaQq92NTFzeaThqAwP55c+DN0YtmtsML3AIPHSAxa/pg7vkwg
QXDPEu3uP60vtoL82vFoaxUSPBbG7LsXj0gRFJsTUumvCp5ui3Muau4RV4zDtN2HntzcL71COpVu
ZYcTUHm2G8+31pw/etEvYOa66MLHH5aTKxzAtrOIQrWdPS7unQ8xefKAs8xqpgKs6du5DAHQFK2x
DhTEqcbLx5sMI2+JC67cUDFddbePVJ5x1UqnF0UwDlbaesrqXAROTHf8Rbnpyn+Ej1CMS3SwdX8h
NDGoCjIe1RPh7oLIrV0Y55gQu0iQdLwcvS/lq81mL+7AASyvWl6biMpoXq9ogk6kFSp6YfI1KPxa
SIQiRLhB5UTLI/dXrnrGNNHlLizAJYGZm6UTKc7fOL93KpT6sp8h5aBGFBDmmNgwObV2pORBBRez
yp9YQfQPihfUugnVw4qNILL16sq8xFaRmEXet3o1wkDExZHQf9woqSMt+qKoZeaSej4ziC/wOtdz
HIVH48WRLmSyaMwMbg1OS6xvDT3YqX64OSpCYEP2Uhy7WVa8VlgkhyyXBK9dJ/cJ1gGCbwl8wsGm
b0gdmcO7xR+sg4pNuKGHf/kukw4lHJRNSyD6ZPafS6sHYaqUg7AUaTBfW1pWiDZjOX2WKO4U7Jrt
c2F3vhXv6jh7FQrbdcSf7Ld12pd2eydYKolh6eEoRlBOQQZHmYRGnmrJ/JfRKjWxynch4z1Z2x4K
dreeWIkns6npRcOaoIGhCND2AJpzlj/6RmgLoTwgHE0JSSJkrxpCZ5EmvuXkw2IEaN/GnCn4oCCw
3429arQ26yQfJqlefJIxjtBnjGasI4zYCExD+bAz36IJNtuQh3lCvwLgoNL/rNPH+gMvq8Cr5KmK
nG2rERp/icr4xYLc8OsCr9GV94Jn1kbGMbk3OKHAEhIfgwOqwHk3SetYOoO55rQhwr+W9kpSSzrf
o0SGo22VbMqTYBz/6+nZlzk9ouLIMlMiqsItZ+f1kVhHSb0W4fDV/7NDog/pySoP5oifd9oumxKP
CXUr1gB9YimzKVIqkpudpiYPCbpeotmHxEz47Uv4LF+AZsdJz00obOf/e38tagDL/SyWdF10xvVj
vrm8gASgThxHo8xxO27Qb6fkICMtu9vEPniSvc6wowwp3kFJwi5ubdQMVoZPGihMtpGMYfRb+uin
Pjv9ApwNVaBGRYNdSG3tbVn8BKQsI+4UDoy0DXUKbNiY61yP4+6RA661DhOtBj5FuXvQZy/7D0SJ
U325HG/j2BaNFKGSSs+fzaTq2VqEb6trb+loQjONnQ977T/2PvXOANGTxglm9piUYYvZ+Rr+PfyV
lUgjvTd5TzJt+wKEtfDFbGXF23tKfrzV34nO/Br0XgfJANdUfY9hjE6kkeevq4pNEJYW+ptQlAw+
6GBH2A0ezu2UCtArPNJNyAiUYfgYmmJV3ZiKEYOV/TwcoLy0OYvNrmB6gddSOQwli2Jvf87x0hfC
j9MVk3LuZ7OC4zQyocsdq8QgDW1PHw0FG6jPb677kGKIcDw/KQwcqnAFzMtW43GTcmwhYIUH/Gov
QUqCobCCPW1Jxx0QRh2tjLdGPZ0hCzJcV9Xn3TCsygo2y8E8OzBlcmrNVUpUEpVMzJWrvaQrnVr6
xcn1XT9lfc4tYpyAfoMtR7TSQNSU+vr1E70JVyyq+5JTDAyJLeqrV+hEui1nR7fp6Fb2NpeuVD4N
HygcJL733mXUCW6uAvtxB4DeROWRYaKzIOtD3xhXgafh6rTuTW1SmxCJiVvhOPIzzYv5aMrurhuc
1W2WbEKCwsCGgisfyK9OOBsYlc3pfV8L18t35eQ8j+FP64bUpknngwJAdONzAL5+ja2rNM+NDFeH
fauGW+pKoevzSjLntasOYdS+W6lzXZMtCtPJDklu8xkZDa5bjkqJlnss/+/DbywUh3GBmDRyZ2PK
LB0R0ti1ioDtEGs/u0hGaPKq96N4GXARsiGZWEXMGEg59FE1AU4YFxSvNUB4iNHdSwMnUtvch1eT
Au5gBnOFZ6vohgueZJ1ytALdN85DIlCLvdX3u6ENh5el2cvgcdO0SZ0PEHXO0fFPP8gIoA3TUQgm
kYucvPHkj61+rMw2WeARBzUKwU3STfkSu4nTu1QvTwl1kS6AfEobaofy6M9nvBQnzebCNVXwb5Fj
v8hN7P80L0wfyjOheerDd98eVad1/5ib3JDtZMOIidymUlP48ExkT4Uc5kUzgHembwIVJPUK8GOs
cDF3zstbt/81V0lwAK/6ipu2dw7vKpXGg+BBdUaUbd20Qe6L0H2fO0Z2RRpw5mIK3VM01lvmsJS/
cOkBJLNBRO3DkMUVDlu2UM0em8yI+Jau2n/OhWy6Nvre67OsBlLl2twOVfb+3CNGiXjpYTcKZaxR
l930zy0qNdVVbgHK5zEduF5F8Dmsb4FOPFaaXrvhLGljzLisqDIDSKdzWq7//Dq3iaWVlTxyHvvN
bly/ZW85R69807zyS/ftWxIm4VARQuzdaQpsOBrgJtFxvi3NfqxEAJbpGi6/B0im5CN8jsPgFlSW
/A2NyHPS4v2noXfHA7vsUYH/wTQ0ugBzqb+NLvmmemEdPavgAJbf6PTEBs5fG/etB8/lolPR3B8m
w+/JQakzM9NS+23UzSSOh10eHjS3SGJhC0/KbszLxCSfh1d3qtrlU968xrnnOMdFhHxxqiH8+tyS
dsFSo1COT4J+/kv/ym3dsTSrTNxjieYCeg6y5fD8AaEEWS/SDfOJbJRXCk2SUzERy18taLQaoYiT
CfYFfrjOunvOW+4wFP1dwnhAVzjZi2EDcoE8Olqbqnq0dbKS9YFbM8WtMBQDUVNw50wVpq+5DFa9
/03mXP+g457KyUa3EUkBPfrJ+gmFUe8gTc8N5ga4HQ0sQRzuJY0ADWExPHjaKgGa4gt4n0OZJGBZ
+DbUGLar9qz3kGZrRDaw56t6zEt8VxLUvZMnQnBqcnFxFnhqLdr/g14RsXVRUK+Y2gkr3UmKqgSy
y3KsORosj98RnChzrCy6jMK+ZfQrgyW9aydOucQkzkn9irs8NoSH/Q+Ht3wIlDO368kQsbftcCqA
b5cUAoJVjKDndPOlNMT4bRhAd6qHufoy/T7RODw9vcEerKoQRHmugdyf/5Vv7mASzUI1qdYUrWw/
LQSsKyJ1AD/XKMp8bU3PAv96J1ixUDbTDz599frQth5EwxOmPv5wf5tJBuHOPQaP7hJK6iGaROZG
rq9cLHN9kjeZsX607iWIwbzRWtniyk629+soy2kOOuz3GewjTIMTBel/N2Z/Ngl4OOdfiufuJtJe
Y0+xMLNYBdeOKSmNjt1nZI8coCLkZti2myBNJ4YlNfgV/vTxBPYyj78v3oa/6HZsdt37on4aMxK9
hStBOsAewJGhwDpNh4q3/kMejEcs7wd+/TS6fteJKCZQaAOkkhN+vVgE20g7yb0EPOiNAPZJkO2F
MvyUgfmcWNLqJjGRIBgvdr/d6iSB6/cLzwyBldn+sTnLIsT1ODl3Ae2beEJF+nnZXb7R3JgXHFCj
c2h98QIhWgDmbFXexi4nsagOH8Own49UrvKJZRkpS8MB+SA2OExpMbimtbPlGWIaGoM7//mDfGeo
htecKjapAvxzvArpcvU7JzmBAuDwIO1ooKhsRa1o+uLrzqK8+f/TgPRF49xlb0jRwKzcQ54H82N/
xIysQyHD99QR/kiBp9OMKA/F6ohfZKDXuE+nSfhUFbf5jWgwRPUpiKyIeooyLo7SmanqlBCoJhZY
bKineFgwDMOpX/CbhVE64icuVwHKc5K29eGg4erZ2hg3Yjp6XXp8nuw8IKjwBa9GnB5mI9Scp5HR
JOXx9XQF+zfMHuteasIX21h02ZKjmrIS+hmncmQNWzCI23o2C1l2jU4RzCnNhvoOXkHPhfAYqVzh
aabfIkTrI0hwN1hwNQ4POs1W7LeDIYZ8ZkAAy456bX40rafj6OT/C0J4A13ZUE7lx8b8x5TWVhNs
s0YyYCGa49gDuCQlMEawVipHUWpeAx8gU6XzjZK6Hu9aeb5d/JrpNZQbRJB+HScQUqU7BTAtCE2k
zMFXwfAozbXuQtMHD6HuUEMrB8NSY3WpbtLp/G2oE6/R9S1z2bDQPJ20r+bRDsmrOm6DlHLlezeQ
/jIGzbktSGEoT/cuOuJT1IdH/7GEwKaWA/t6xqcc8BwC17VpCCx/eQtP/syVIfyVrdAzuQ+gkZWb
w/xnrd18eHE2o1b4V1x5VTtNHUMCdsBWy83OW02jOeCxvmeqyMk6d6lpkY7aWTa918HbpzGIv30n
GiRsFBy/SY6XtpTPwf3lvGmadnn5fpOv5X3CuHGzjC+JNjH1NYELMDCfR5791HMe228mExKHiYUr
ad9IK8SfXGseAY7gcSeOSIYRzRgA+Jabe4c+Xc8TPGnkXCF1im6dH/7SuqkCBBJquTKLs3Pn0g4X
HUTxi3BEB639Sn4ibT6A4sxKc61qLw3dNBGYcHqit2eW7T55gg4buwtH4JXQ4vNQQWrzkCHCOMiL
DwiUzVOmZdLFe/FeLcbfiCQZGh43srkbVpGvKwEbHocJCKlkDby2I8YJLNZnwtYpsKO4f4i++IHp
3LZpJ6QjOLMUPXeYMOdbCNTCuFUfU44yVBZF6OJ6UzkIZtG/PN6dzLUskltP3qJJerOo+ZZvq3Na
Xpusv3nUk776orraeEeAqDmuQFbnAQ/WQ1ddY8koTyyt3l/uJO0laFADHdEeda4L3FF2TtB/UUKj
hCHOcS5pZUWkpLbpSo2Zipkl8YTLsrLhtZK8EkPD/aoSeUtq0UlvdZz7skQ/3ct8uOUQsDhezeRw
v8hF+Hb6NNUwMwZBB/hmMPLTg0IyN1BGZ7EL5H4Nr+zBnmKIjUoUOJgsaLQv7SdjGBvTx1hkMm5I
41avgasDWpqkShge5txXzlpXc63cxOg7sLvCH0RhQJkkk99Cjt4Q3wPSjp1G5lQspO9raAJ86rLH
bztrAiK+of9IbVuREW2FaGQyYvRK909erelG9sYGTvB0UWCAMWjYsOhlahYyvrqkHmvlLE3bPZ0U
ihu6WqP+bKhZLgQJurFjcF9KxLppZthOB7v8r7mJ36a7LXevK1ddI0TBmiNrHvc8jCVGp0DSlZlv
f5AeXY/9fcOlXP2YLBNMK9fO7bMGYLrnsBjIjxAHwxBwz1DEZLMmIf4CG3huGYXhUDPxzw5aSP4S
NRlS22rsCYSkrjgAlWnCF+og0/Rreaikldd1E7KfEoX6A7NpI2wxobn08yzI1r4p/lYXRjXNBnCs
SWvFaOVat6VNq89Q9MKlug6B0HOVd+Bj8EtKcBU1crj3rFkSJLlzX7FefbfeIzOgxUNmzQ0/ENQ9
kgJ2O75T8B0zVPymMREiPMrWF8EJbpBVpYv5k9hb5i6aiFQm4ARRl38gIpmb9O9x8b37b+FZTQ5s
k0QGB6Y1KtYzy8+CzD5TWsSmbd1U5YYKDif4+m5n7mZPbBswD0EUxLaFz05QpRT3oEZMdEhWoy+M
C5I1EfrYlotKj1dV4ZxgR8C74i4o5NmY4KoEz91tHSW5UbNnOuz+gngTHkY4PpQgoLfrBdsDnY1F
rCCI0cEzpXhIIS1NN+cllmc9z4Gzup2F48CHfDt9jqWAWmHTvNbi3/XtmUpg3+5ywv+gf174zt29
5SAqwrXsFOi3fuNDQ6199tRvpwaHsW7c2PwhDYYmsj+KkaKs0Ksig41UFZuN2YZ8AK/jusaDZpM4
+6KhWzuS+WFfMY+0+uFS6DDLk9bmQehA+sp6GS/x/rx5luX35UxsKuojy8GopfQmiN8She/NPTGw
21UinEaB6pe0NaL5eyA6uDtvn3yP8APCzpaUEAUVdgN4EDGFpNVZzysyZxZIOZ5dCDqxoZPY8eh5
KleU1lrXEvSSqA8DNbJswMkfF5ImjZ7CQw+SiQ9YxumSzfEyr+kf3wzcWcnDMPXtNkXR44c/puO9
0amimjaP/QakZBYDSY54EqyjjP3xBzJuT2e0+ZK8queBak8csZ1rvFK92lKwNLsF/lT+x5L49YaR
cWl83urLA8HHdsS6V9ILXMhyaomGLgGb7o6X+u5M2tV54vfMVoA4ck+zteytbycunIt38MhKwYtJ
dfOcz9cNGBeKkc9j3+I3CVclo841n2GCwI1/i2pSehYq/uNWDWAZA3ThgH05B2fj1QAOUmcJu+IF
TSuRK1/S3q92pORwzTKf7mjjNuptc4QARJNRKbGc5RNo77020OE0D6Z3vuSSnFXnmXa4Yy2J+tJ6
SMoUlZJL3exLhqNyhKPiVA9WEJUkDV+ei14/PAumdCr3QH4xGkd9tyYH4t0IwXW/w/i0YFEBjZIv
o9eqizq9FSbJhqk9H7XKBzrH8jDxU5IyvJT/hRaCzpw7glL1mNZI6KW9+0WCdncg1SqfRMcxUmFa
GIfisAKvG9uZMlAxf7dyhMC2HFM/Gbpw6Uptv1toKPtdn4+xHttkkWix7IfHD87Zkkl6f2K9+w7O
/agqfn9RYz+7A2HGw5XvGHy2IxI/ytpZA4SgTi63y8Wq8XGQ7wM6FUuvc2h9qx4y/C80ba9wulp0
hQlLuw0qWZn11IaPZqEXW5OeUIGrQPwKzEhiyd4Aep9bylYlJr/nRt3uLGJdhzOG+Je4NJUDGr5k
3f+1moHTyeR786mIirXULqP8AD7Og7Z9DZLIT/Ew9eR9vo7JbHRcsbwLuM0UY2DvfITP/yGPg3tn
pW4gZIKlsbhSNjbs5XNVa84AGMFW7vSHFWY7GBg3YmS69QH17BRDfCVuhdxvWYLgni2cz0h/rM4H
RYGuFEc8s0tqSfcyrxC8Zodzf3aSPAWSJCIce2187SmJVdw4+gkQuuLObGt8DIkeX0+FLJHWASYt
4phHMVlwrYN9MXnMoRbl3IBvkuLv6T8nFWZrc5Dw/IyyXPJ+PvKb3lW4C4Vk75KOhr5wYTjTYaR/
F77IFatIaAqum6LbDTfR1LYuSMan9mIVr7HuYItSNWS6FuBCuG3GjfUM3tm81tBJdT9mmVkUfoiE
EIp2IgED8ZW5ldQTtyth9SrSjpsUWx2KY2cBZwJp0gP/UnTO4qWauMfKURC+nUUSpKA/5Bf/8y8k
e42MGkFPtekEgjUgmoxnUMHOP+xpBJiX4hbmd0VdzAyGgep84BCHKP5n9vABu0R0kUtALbRD8hOb
M2tgBNMquR7tGSIqgzYuy422loD+gxU9UD8r4M9TbBMmJbPBRX4lryBHCWR8UDvO/977ad5kc+w9
0pHq9ZU7LtleVFBcS15kcQ+hfl5VaqPN5TRtmmsuEPyaXvlm16IisRzXJUzeX6DKemt1/tq4bkyP
Y5nAg2i63HRZeON2qObfq/4/uoyzbOVxz1u8hZL351Vfw2JAdSN6y/Gs/9MLtqS0Qbio5wTCrhPe
7U09vNxzDWSHEJBzQXyzOPlcWI0bgt90myf9bI6gqQjB22/r4O67NXjZAZi1/HJyK3UhWi93GRhr
O9IEcy3VSwwq5YyfaWl3kCIPKbW9MVww0iuQEkzBApBlKGdDqVNPXr/iC71RC44I6yIIIhhX8O/s
KgZvw3PkGJYTvIWU0sHLu06aSEqioDgpT321qlVQ8e4YbvFJ/aEOnDbYYK8pmB5ZxP5z8+JN3/70
3FYmbYr+ORiH0nbOjZ89gIrdui4ejHUnavYkv4BQJyVBzNB89cidU5X25rPNL1F5S2AZcsxBfqBg
rwAoMAcreDmPWDkwHt5BPFctLolH8iUL7Z7ZPxWIOInZvg7bgVd1y0CPyahao/6QU/SyJPicCX4w
nLNaYRiYlnmmKUjrILtl8tbHA8TWyqv0AOWNJs+ORxxGZBMMt7gVDm95t0Wfkl/+TNIkoix/kTe9
8FykPSJvnGTdPh/VMsS66mjp/xRSLK4NgyeUidTQFfHTgDZGzRV25Z1oXe5wHpaJWxJ1b5ZJ3vNk
qFyCeyyYQvA95ZrO5AYDkujfi8uiOX49H4/QTGNBZfYtJY7NFhy0bFve1wfuuyzFhpCunT2bq9TU
d854oM2EAKquaOp3pYD6bRJeAMHAgaIkEu4Y4U7xC/PqrPwHm6V3JJk/yrNUi0IGNdw0lJINUzVF
PEGeRMGXsaUjQtqo7cejMa/8VkmhsdfV48IVP5dLmVSQ8HUMGOJKzGM7LnIl3P3exFyyDtZc9+a1
IGb+bfy5mDDBH0vfdNCeGUHU0o3z6Mj5zoN/ZwXJt7vLjsnDg7dUvX/E1vZDCQFdbwlIWnV8lKmL
ytNj/ZrIhMi8Xum09xYofcEEAZAt4gREyxEZ6iMh1v0LDelgPJnj7h76+4NAsCU8OMZCP3541nYe
EZEnhOWFwLD68MGxqf9xE/Ur+pCRtiiueXSxqjVeqxccQKmEVCblvuamLxiNJdyq4glYnegT8VGv
ihWITGW52/gU9gYUgyium2YK+TR/va9bD3+B8afI4rWbHTBLNlwDMkCR6yJrQctTZz+v3srkkCK7
b19pCOzp4Ab84W4d6MBND1RxgCUlC3eF50j8aW0UzY+bNaMdZqD5ullqC/F6UPfWAwFNsJWdltRf
bIBxLgdF/vuIOf4gsgfh/1mMpCEPOCYRfqjM4uIzOxNv9UKqzGwcjE9tK0i6qIQ+s4tuZdpBb8Bd
mcgZta3dCiNovkv/cL+2hrCtn2bcVbO77ahYMOCwcjcsmpHfku69iqzXVu2s6fB16naxYdkJRmHi
ERF88W8444q9Ei1egtc/FYyVB5Rqu+QjGsKKbf6xUl6Jmv6fNv+oLsh6AcMZI8hGTMhDAgiCSCLA
bEs/NEeSwOVVAVIVUtyrjSKOJWqb9RwzwBiF+J12GePVJDZn0tU1SpZerlVswJSKHB9WCGTRct2n
TUdNsBaJJ+EbSWFpUvfcIk2HpTNjIz0SrnFDLIL9P1anWi3gcJk1IsZpLigioS6MO2fRYpYytm4u
hqKGa/6Daka1oMtRuS8CR38y02n3oFqOqO8D7vo2p9JLo0NegX9IGtZ6VvZB7FwnYByI2wyo+IQR
edmKX2bk3YOrYnpl1wQ0Y3bKUUTGOyxT9a11FS2M5NoVdtut4kFXm/ILiW7gAaBFJAD9B6hG7N/h
H71HIUwRE0aLc/99MvzamryuKdrYg2lEhJN40cDNO+BeatvpIcslFUk9jndNEy+Fgaf4RhKuk1mV
6Plz2ir6IRYIUFe7jsSimGN21+T8hyu0bxBzAon271P28HOj7ULhlaal1yJ4fK8/Y8Uuvl9xqF+C
/4aWQy2xgSCExEu+5A9104otDpJARNEnuBKDb4hXJUEBfXvmso3mMRhE3xMVIpAtR5TQnktc7sE1
gHZq/8pv0BuEc6DXrObtmb9LlXvxmRgLKOqUtat6yxBB2kG9KtjNOXu+abetjY8fIcpDO+3/5oN/
9il4fSdqVQrmXoRAtm/KQ7baB9npZi7F26H+rgE85i9BUFDejfZjiaivGCGVl0c5g/FsuN8CQ6G4
P96gF04ylJF2N9IJ9SvajXW58Yk46qvvHZdjgDLUoOf9EozZ1ppXAHeHYenwFoCj4vcNyVGLpZjg
GpZstrFxS/JYdEkFU6aArbn4oFx7eMMmX8P07WO2eL1ViqSgpMCkUikNvuq0u7tCJtrXEMHc4k0N
i5hwrDCrptZGOKFMSng6alJ1513JzEYIY1CVDx+rWs7n//dLGNPDwExGcZ53XtHStkcklvGSCUWD
S1bJqHrVFjpuTRIsDg8G/5FPzbwx5E+s4gD2xfn7erzIvqcdsjZJwhwoXIsLyfpB2ZAnidRWa98l
5rYOeq9ngcCU7hfe+8HetvN7zN4C+Nmyl8eoHY6WBRBE9bWRszQKis5fKXIRUC+5islwa+rSK/oE
XRIS3BbI1bhJep+NVvxCpLld+CQLJQYx/xeQcnyNJtKDPKJesTGs9M2Jqxdo7sbXh3f7AphKWq29
9xRANCU+ua0LmZlPttJ+XVEk8oVUmrNGMaBY5cZFUFquRNthVfy7aDL0Rrtn71wmH2AkV66jGgy+
mzVzz0HVAl1xHvLSZL6Xj6eUhxLx+D+mUB/1BU67UvS67CRSpOTcvzU1CljDHsHS3Gt2fxzBEwfR
r/KTAru1LiXvXMzXfIX9jykU2LsSpGUyV4bb1GaLwW7Rqcxzb9Bp7iXUTmmzsmELGyqkFfrJXKdk
/xDCwnaE7vbAJFED4n2zin4EHAVA2K6qPqq6YPno9ruw/Aq6+U2eUuolrR5JA4ypUnp0VzmoD0AI
VGtEi2DyvMXaG6hXTpQyFch2K/WLaCdKXl1kCGIxL8UmNaZBxFeMdv6k1eiZq/pFG/rXqIbPuFbr
ntIW74hm7bpNbGtDByO6Mp1pg/IcCPV0AdAD0XFghFQYg789WsCVGW1MoQNSymIkuBl201VRy0UF
HIKT/jiW29WY4SOrvakZoLPsVsQDKxF4FrZoiCBkK32Ejv8/l3TQkOlv1fLhu8SsCEOuOBz8RnXH
G0ErppdogrGfzuOm/sft/ZHshKStsoqXE5cxqEG2Xrllqcew18wtZATXEp2nX3VBJMStQGJCfmU4
FNuL+FpaKToAuZyaKwsjSUKmHBrthd9e+VEVQFNq0m2IrGKUQDE/BZRO0FEYNOPXuh5duXnHESkj
lM5OXLQrwP5q26qzpNzURhWTsxswJIe+nRgE63wiJJ9mtxy4yDExDoGwvFtDKeV33rSxa1sIX8WJ
8PsRfB3oBipDNQ/mc/6hHktM7VSLbdug+F6C3tgpOJs1JWVsB3r654CweZ3UiaChr7WTOWmthTmp
cYQa7Pb/J6cjD6i2zmCBaRibBfUVEuqAh23Qkc3QqL59U7gtPfCCLgm+DuYka4Xi1+mvNxljoIqx
7yKDlgc57RT3T0kZ3ZT0yDVGvkmo0YyXFDqZHWFeN6ymgfTN3WejEJRb3h/MyCz+azE5uEFkwWGE
GtgJBBvBDZlfindLmTc78M42tqSjaVtUdzadZ2uicr3bAOVYO2qAJSOxTj4mMjO71nVUHTEJTuXQ
wuK9pSq+8TiJU0dlvTSWIwaj5T1smN+2Mb1eBio6tOSQuyTRjRtGaK+jNNvjfWpKPNMtB9ZZycFY
FRiUWs0LqoVCZzuO21WM1gZ5H87cFyyhFIqDN+3/1feJ1BrzvEwTtiIYnre+QD5qxjH2zUUBZllj
qGB3YbzGijv/LED3qZU9hPFDCleLLmt1ULktZXYO1T3pXoJlTCHQ0OBEsPtSxAc3eANtrTxKmioR
P1VN87oD/gEhlTcEBKMyKvl6yPYiHCafSDEPDP5cEil65K3PuSWeUT+RIAIT4IfenxvR+vOcReDH
kXC3DZCnVNzb5wAQsAGDtFKdIJefOb/s/9Gttp7nfuhUsBwE8ksNbF/12fQKkKx2C6EGYGeriewz
LL0X47tzrzXJhTbFYLjBtG2xK2U5sIufzFsXmhoHmL1p9nj6mM3CxFhreJFlw9cOI8+mi64j1y63
FTwRZElNW0Wi00HaG1jMWS/hfxy/F2IEcMzehpQV37MNIi9dvTzi9qzADhO0hHsGm4eHCRYaCHpm
+3MFo4oudzTm0jAXn7TWOXm4ooY8RBd8znh3ChhrZ7J5X+laWZ+REaA3MXo0H4DclRTbaoygrvC8
P98fkzBjBKfUPL8O6M8fnaZ3bKRozzGrbWIprdrDzwQCDg/sd+hfCoRoi6iALHK1uyqdIsdPYVi5
Zl2YDygk6msM+IIK+k7B2DRR726dMWIXbsBp/pArc6ODuTwSKcIb9umAvoBKX+gQ0mILtjlxpkSi
qhOqd44y4pjcnnC4TR1rdRmblR9toteFvpSGzBrBqQ75myiTzCy9Z5bRxLln4csr8PwVimMR0qdR
EGsmLa8Q7dBB7OBqFtFGE+oJYTQyrEXbj2B9BRPvok17ULkMSov2OO2TN7KH+Kj5qIMqn4OHvMR0
MYiUREA54UZjOtMrhoIA4QjlFVKq+1E4peE1WOmXWgT2VkEM2Sq7hrdJcZeDzv4rL1Zcrbl1V15g
6j1yvYGfOvgRbLcfUroPi8VUwhnEkNthh6xk9L+LUmXtoh0dMMIWekDQq+r62tqZjfjMS+/v+Nmw
UkXVyTZmBLMnd0P2GnFBt6T6YYCPdcfrf/+bFJiVNAJX3YaBPRajIijaQVBbaE8ekdU5zXrcOs0f
zY5PIn3ncCxR/hHoERgQa6w+RkMbTfNxcd5DH+oO1tE6p/iXHrzfbho7AGj7RKrKABR/WuECAqB1
xL2GB/4/5ZvNdxpqnHjVuzWPQaifIeWK2zqvymyaAsRvi1s4DuqEchyhhbZzQGqmfjSZWo/6P7H8
J/xbiGjfUlkrzFwVFdD4EfNT5KoEXXKGiL7mFWqpSTmw9GqNflEJM0uXOnx0wMEHEVvFwxWPDFD9
KffYUMTtsx6wsPdk3vvHTE/PTHvhLIQrqj74KLSSrXHlNIRUdS1hzcoWF9rtH6AiWaKde9xQvIWK
0dYVXSdY2XxQe8fhWebXGryaF5s4yUnmZWvdM91W3ZSZ1DL3VuY1YizGDOUKZIMQbBotBdClJmcC
fuZqIt6Iy5nqoPYNk2K+30SUPpETnwzr3GICOPpVb5j4iatYCUrdgI3nMI1iVWU2/X30Z81QxV6x
ml7rn5gmos8sLky/9dKmlqr8ONyEhUCuSgDoOASBdb+1Yrala3HfqQL3yvioXeF+XlcEOoXSYI2V
Ya23/FZUFFZ9QbESg+/fMPNwjLyTTZ45yy6bS2ePpRs8kmdZMWaVAaovizbXiRwYa6J3oDrFR42A
PnGlL8Hx8LR4rISqYzZNe2JkByv5mmGQFn5YI2XyIaZ1dOFgdBuGjHpkPMoCcs6DzsJbbiBLhKtD
sMRG+mPLpfkHuhknnrm5MS1GnfODgzhiF9Tael2NrePqhugsbBwQFjzDwCYaC33ZaswxPfbXpexO
BkriPzGnmyhWEikTURzsH+IDRkMdARI1mND8GwQBPe6y42dgcOpJr5efNpYMRLojKzUzieU4XNdt
d3uiU6JniJ4wP4QRA3oz6Ire5BH+0nY2mbcMm09S9L/jY3WdOTDn1Q9WczRJqBqc+KqWgltqNZdg
beiOzxSK43J3Ef92/Z18wxcvMPYsi8RKIPLWY9C+RWa4HYrGp/FRMcW9NYE+ljidx74v7qwlOFUj
ny7bGdIUbj2WDB0cCywYHM7NiJeMid+mnCHgfXEDPHmASo90rV5HhZoprHFfq3Emx8WZTvwS2Oub
LGmbS6LiFU+EAyDG9EAdMn4O45ATlqXxA7wSq/Db+ErkK58mxu/DZqu5bnBJZ4C56ytS4607n7CZ
VQsQmNNAYFAj4+YZ67SDXtZ2oZTlGQfJ004EaEJCSOrqITLLuwUIW8SmWetlzupjXDPpGSoi0VGF
00T9VveRl1KtGlca3kiCf3nwdv2cp8/rVclk9gMDzUVX4L0iZYmB3mMZYaj5lod1TQGjpGNfZemT
bGzEyFEDFNfHrY6zjVA0GnkqWzSC1Q/92S5as6cqCW4xBQ38+IvbyiNlQDvdYdU/hGMjS2OjSj0G
8utkWws3RHftIgtvAM1uXbmDNzeyPH3nJjSUfbZGiCXcZDEyNctTzf4JXfmXyjhzyiuelCYQdQlv
DKJ1cTsmUsUHw5XajW47eXESmIIz/Z8t65LqrubLzPyXyMr6P5bh4IzMs2Kh7+Atp0IODyZgtdse
umkgBaJJ4/j7mw5zWOCYDqzX29Td1vFnVnZwOw5GPHjCte+oAiTaeToEBpoKssYd8/9Yjqk/HUI6
1x5ynLYCYfg6fkbqNCDrUdQySW9nhjyFZwDtANsX3c0neuLtZq0GRDdeWL7mSpO2PoWzEkTWyUio
bNpp5nKLRFgxSmZ5HPomKkK76hIbkFUSrkJNU7lnSmIjtKRXhzBQHh0eCT0uOC6gWSzoPSsUHBqx
W/lrleTlCB6df7JfjYeMJwx2250KmyK2sh09KUoZEiSvhyqfsc+1CW6+BpekfaND2BeuPmBhUHd9
a+vgFCBjofXn5ttIk3FJL6eH170Mfn13gguwSbxrI050Q+xWJOtXDoh5CghDsBbHIwJpew0EPkJJ
3MNxuDGni9HfROH0Bj1qW/U6nlYEBike4H7zK7wIZT4bR/qkmen1AtbjHg9VLiyVhYCuSTg64aS+
17lR1Am162Lrix3VFz1iETho10h5PEXwB4xdBthigI1ceWWX4V4I7U+1ZXYCbenzB3vU7A7vKS5B
7J28Yvv6yvNc1g4ejP6bzS3UZ5Y2FhkqPyE/stOpHKHJqfVaQ97jsfpD+QScurBbwbi//L0Pt8s1
UYtJG5HYvKig0oLbk9tuAH85iwEhA5iD0g0QTcYmxKGVWxKJAzboBhfsVEOGHtuSKyebsrXwfsd/
73rlUvp9tGTr0fahLZrze8QUcU8njH53HF2X6jxEaB3p7Bl/jtcrSbdBr9lTl6uI2+xI0xmV6dLp
A/JihuPURWd8PHGgHV5PTFJWWs8G2OzPvhmgOypz9pyDxdVHv97/AkzvcSB4c2IzzmVPncFrhD6Y
DGijACKWlvEljuRn1WgYuHyGeYliXznfcE8xfrmNqu/J2eON7phiFaHJFlvuawfRjrq8upeVvxmo
ajh+AxhaAAkOpHCvFznTr+MFv/ShDTS8CeRJd0b1QzcJU2hdWa+VwutPvYm6lCuVcU0BMv/bEPB7
+kyxo3ggW/vzh/Ld4/rjjCLQIVfVrun3ONZ+2Em0zcTGaqirxJz69838b+RILmFSVvpcDbtLfgxu
ckIVFHLfMSOgXxQB/4ynYJCpsA8RVYSDa60kqEShmsKKDDsfFEaiRJttjijIlyNj/igJoaQULteA
xamhZH6G417hvdbN0uz+cnDHBbBe80Q0i5GwTdFUqtkNlbYwRzisX/WXNROY2phBa8NwLw5eeIJx
/A1tDMXKA2tnmGC1s6anGSWAa2zp9CjRtauHDlVuQMLrwjIOhaYRIWQIv3XV+KFN+fbJPSDr7yiM
VBDvymz4m9kjfwFg7r8nVMJ9QMHrp8gku/7wKVkaAfnTFud2BJ9kUpnVKxw6VYPiiCnHlUSpczxy
QIWfEVoql6ZRTpzOpV8iyRbvPGUqMdMSnuE5CGl5f6JOYnaI8wJOPDnMWhlF0o38psBv0HtXh4G4
f4xJ4KT5/9hkhgZlim9j/gQmLksg7tYiASE3sF9CKsVpIUU//TEFPscpVobM2v3Isi9RbNXZCwbu
/BsuQztVOB3cBioMEkHddddagd8jvQU0RWxhnczcjzmh2hGnt/9anQz+/3d4YpE/8DZu+rY8SuSB
buGqTIRwcaKddO/sVnlrxYxQlf/fIr3l0jMY9ObzlJlao6sth3p0kggrMvvhgEFSe16PBJ3euP5+
iDzd9XXdc42theE/z2GcHgqAD7cDd9nTf03om7NG2t8moyUA1v1cSUNaIGFrajItLzBmmfXN/spE
dGcFOzEWRMD76MzRXHQTohpRX0/cawwYivg8ROkp90zWWQHujrrXL9b7dkFW6nsJXDL74xqHaVKM
nLZaCbHNFPRaAzF+glg96CwYhdAXUcomTuBohr7UWSLfgIiSfTY/5u6NGClnbGYiytgNRpWrPsb/
W65im7QWdW2b8V8t1T99WIhNQ8IeolN4roy7Fid76O20LjS43oskyj+Z8BAAWaQU8mTsWBlF9mR6
oQLmTBn2BEIVcuAHhYJ4T3p9K7bgV7hymZf4yOyY9xdVBponQLSLS3ZKxGwf0QUieWRtf5U5g/+Z
gjq2GG21mhi1DCml9hQTokh/HdrBH9U+KN/zx584iKS+Wf7aRdBZv9yxV/g9xmtc4nH1HL8mnZo5
dyHEr9MvThsEfRCrd8oRUX+zpIGO35LMZpPJ+N1sDlvm+dg5V50TNX3kCl//EGNfI1Z4SBSK86TS
bh2HAvr79yydouJ81nbJzKUuCCDEAsDdH7nQPFSuwEUr8xrODio0BouGF/zi9Y8rY++vefsFLek9
MQyIkcBYMjE1L/kZIs89J0xUZn+6vEif2BiJ+BwH/WlTyvKamnoQYnsltuxUt4Flf/Gqxhr/oskU
KK+OsuWbeSjoU/3h73hI2ILecD8QMizHQUmTvWiU3k8zh/W1iA/FyXWn3TL3fvfl123UISUA/7B5
anur2ylTX9UquADmnuIbEBpZDoeAyvI1eosl2vf1UwzFLkntfqPPyrbM8wrb/AYZm9GySezeLcH1
VKUROuJLBCn8f4vfF0EkGHrxE+RuL58jnFZ8GUDfVuqlcHMdNpUxhEHAb5e57lgbgf0o3ixoSMAb
L0moN0nJOAG9e+PxzUrNaQOwWpunMuuYpDlJCoktSt+gpU91CROEeJQ3RQoJlqKzGVBE7H++Dbu7
crL7XuLqxYGYoKZKRQe9TfyP9YVyyb7SxzuixtXWzSyWll4hCrclM+vpk6F2JpeiWIv2I22T3B5y
eyag1MHXTp8/mwZbOrA6u8PyXuS+q44isHdvpXpWCiOJntep+sYF3I7rhyUPd0hM4PR/YllQ5/yc
Ks25NWdx+HcPflJohuAh/0tiUzPDxZ3XJTbSMYzE0qzfJ8FcWXPh4mmrF80ZzJwIfD/YqFmTNxzr
eEcqlhTVWEh0N9drdN6t301ceGkJuXLLbhALRyVruSkSZqB6X3+/1pXgp3mxzVB5iJx1JcePS6D4
57U4ReH1tcLlBa8Z6h4vEw8i3oJwGuV2Uzhxv7waFFcSTbvNH3EOKUyW6ghYIent68af4X5/udZa
1AGYh6BW7JAC7ZRCOQo/LJiKbDydIsB6fj+Zh+HPav4uTFGIAurmyVNoiiN46WeRPZ3PE3nxiMZx
Y0PNZmEMc4v+iRJaWFwHGtFQtanSDuMAHTAE/1/QxBVk3bBmN/gxlJmgCulYgWXeGvMiohP0yKo0
93+ONCCAuj8od43aLZe89LwKUs0VtRFDy6j9ARqeiOnskJOew41TYdFWKJswsI/nr1NtB04AG+Ha
5Dpx9V8byYT2ZSwjVY6cm4tIDHXqjibJQPRHKJnq8s2E0ikjFHqaSt5Hg0ukD4/NvYL3ipJkipDa
52LnMMcBo01fgFInCDNbNjimUX0jA/3DLgFxgPwlGxdxjaMLxzGMasFTkbs1T3833TtBXfchg7Bm
/ih7KFMP1U6QRlAQZfqfHGYAoVbNMIHQ5y6GXwz704aArE1tyjoges/j4iUqCgHB89VTYMwB3MKk
pYi544YRThhh3KyiVafMsPBjGDssYGGGy6du92Cda2c0MxZBw5B/3a7065n/zu1OflG7UmWpRGaY
Vszl0iCDhhKIea84bn2RUzKueyYx6WKI1Pw+x59vEHAas5IhbzpI5CrDF+BNpk9ii9o+E9N7Cd9+
k0iQaeUdiA8NHGBzS3NoiaUCV8FvNeUL4oSGbGz2g0xKaCY1MeJ89K7XkdyAAIHQ08GhEN6UYTL0
6rUIeh8rP8TWdiiBD4oX81gxruqtABJQdsevRDRaq5WJ1trjq4RVfo6eVzRTCZbZ1QdyVwb9blaz
c02+IDYnYsZZXdM+26C/HmfAAnTgFseJ7UJLRKwi8JXZ9gi64NVaEqhcWrQUeSN1UwvDVk5/m6JI
5JyQjg/+pLkHtaVVSoikM9uYfFJnAkNtsW75NacG45yzxQwlP+N1wsLfjyvp9juOwymJYP2SlyJ/
zaR+4wZUYN6WW86yXUk7J9fXUTBN3QkpFItTu1MPS+NsybQGC/BsYd6l8FlDWkYrxtA6jKOAdhn4
XbMvbtFxxja2i4fWj3aL2dfpl0I+QLyt989y1ln+E6Ne7S89H0eo2kfsB+XFkPdrpRV3qiD9+mat
al9wa0Shj5cmKQBEWOfpzXdBcE0L+gR0fPwInQeztIA4GOdbY1nBDpr2hopDnCEMRAw0G/JKdqga
I7YijK/3Ev7zvcd8QigZXe3dtMjRC/yci8oB9if5IMZ4GtLwIjsVvAo74+xB+OAyoy1A/QwRiSXr
+VS/0Tj+6CiaZ65KBXza6fpZrMwI5RRfzreH6ETZZZ6BKBLRlKDFWTvmoSSsMFIyPbB8lIML6sz2
zZF78wedoI63G+5LITpmpVpFOqe4obPVn0reI9ZscMUc+zgvq1aQHx7v3JFPTNC+zvwyowbAIwEo
KRdXu8iwRKlL5y/UJIKeuKHTa2Tr8iUinY5Q3HTr7I2+vumtvyF0D+uS2o+154siXZhUuifdBNQO
jCSgcwBAurVrGDJZl8tBd16Kk4obfnnl8Y9SJEIMqBPhqPm25WVwg8tCtR9OqGT08MKNh03Ae2z5
W8rIGwRuMKKuTYRLtm6ACu0cQfbWByIH/q8fNdCdAZx3s87VM4tRoLtpmPeScyrezaH+mPKD2DzJ
3yzInm1X3f2jFbYBU0l7LBCdkVDJJuwG6GpM2HIwtaJAvxyBNsRmOEe54601wwEDPCgFftZzMqXu
A60wTRurE7v0K22/moi8IY6bttdpX1vyCw6s1bNR+EbiK4X0qcCjGtV0EwIOd0NsG2UdBc2PofcE
9JAcR9PcG3bYWQ2Il/8doVCqRJcN0/K+V4Dgz3KsWWSp/U82cdicF7tGMmCT2aZZ30wnlQQD3zdn
FNx//rf8KJopxmPHiXvm+X0astpEJdf96V4Zu+DsDW7JGnJqKE1YofdeSorHXtZA41jyPh9vACjq
skXk8gLxaLLihKNj55ElMzvIfZwUli98h9+Epwl/LAHo+5wrfPrWYTjS3xDWU+ajamy78SI5J7gX
plI9vYNSgC0J0oitASTsY78NQZrU+QS3UGJNyrmatikciwokjjktVERwex6Lw/2qy9CL3KMwrFD4
ws96SFP7ylm03DJbyjDEcpnUzvZDtuJ5BGCYWq4gwwxT5/XT4Q8oUBNdlU7RsFbwMp4r1NwiqZps
/Aiym9O0SyhQmxGafWuIG95WRvXJiekbeaaFtwwiZgkaq/B/ey+9BwRogSjp4coT1uBgeo7W0trE
DXN2Z3YnkhWBA6KHJjYBTrWsygdb8zhFk6VGYo5ahDDfW/binDl+jdHuRUm/uOfWnLCuB7jdT26n
HsB8N9q/lBDoEEk7Sl9tCJKqSc4wNPXuAkJ3uZujgcDDRrS43PPhHB2eu1+Sq7fUfHb5GK3bLqVv
h4hjHVMnz4n7gBdCC4dS8G8MHN8Rf43qQCEh0pRSXxx99WZi7GMjOdubxVD4/0W2Z/v/HF6xJawQ
NxWvSb6bBvlY8uTzwKc5QIGi4aDk1OMf/eDcPKs2L9Tvc7szu3a+ANSmfuJMavreAn4PtKzKcuRv
+d57isrUOkhFQvuTk/iljes19MSKS6in7hKAI1dMD2Arwq4GeMkBwS5mC/Kb4H8xOGW7WSW1jd9U
Tp1T6zVvhEs3Q/vUQ10zfw7g+Lgp4RVbKAQAtCA5757v8gjz3rngsChkH1w4uKQQ1x2VrjortCOu
F5HtjFpreWMpdihPvgphOMcf6tYAPuz/YMn1RO0PoiiFulhLMJ/LCAFCuaGSkkXpjiyClS10mHxX
7dOzGP4H6ZJZyGluB7bjbP+rj2afOgmjevZ14M5G1SidRCgv5PZgXUFmPZYqEPsgwD/yBJQAYJWv
Qyzdt2RJPUDbtwI50xrr6h53vl6xA2AV89iL3fwwat7wzcQY7N0XpGXnR3thEiRZoVIuKbTgxFCC
QHiwnlcsUaNxNPIG251Z47JuoJa5y1iYZTm4PQ/81T7cStF+u7twX4hjSg8RwSqskO+Y/HJZ2hlK
3uS3HsF1UiEdUQDLJJEOgr0R7Il+Lfo3MdJvJRltl26AVXnOPl0nVgE7ElOOTs8mz+5NsePJp+wc
LS4+D9I3cIC7dHNLyxm11UYdc871qsi3FoRCI0KzBdY+pVh1R2v6bSo5ZkDwRzDThXvVow56LJRw
xY6WtO2iOFfRYqEUeepEhdTXcdCMmdxr5130T4m6g1JmaWyWzNxNbgUXuBUk6Xm97Zgnni6CyFcA
l5oUrKa4WoZNZBnv0Nw7dPu5GBavGNHjbY6H2JUdEM+KSBIDy61z4S0e1zzcHSDp1u34xB/EtlUh
X4777gCSwbpzUCpvoz3pOOmdrJ9xYJlWSK4Ri1sPPkK7dpGNIlojCbjC013TIPtzckwXMQjMN4Vq
hspe5xed/a8x74GGsLHIVWB00PaM878IYkE+lnNBIZ6vNCnTfpQNKkZI3Lmdx2YRNVi80KbjloPd
jLYAV2H8sYS1eUVxVuh4rXUdBKvZT5z/YoA8z5P1IT7bW0KN8gNctCLQBVZx6GWrUCh8cNL2tLYT
5p7FuJOdvZdeK7BbzC/b5UaNYETb52ZP5qh+72qbyf4DHPmOGqOVJZyWZmM5TbBbpYJ1/tZGvLnn
ij8YS5F08/Uq1RSP/TU2bkcgfDhClB0qd3UtOsXY+c/zHkXUU+URoWT6XjBhulvX3GsNMhvw2b/2
zQyoy+jiwmULAzkhZ29wcz2izspT7iyR4kBTXCW/YVIlPJfGhEjp25zQhzvODG7ZPy1ftanS9jJp
WGlqhVKDB0rzyUMVFunZf6lP0GO5o6e9o3ZZPKW6HL/xYWGEtT8n8BZf8canYXr5PcPB6cZy6U8X
q3ULkAX5TMNCHkQ19Z7EM84ML0gRatpPu2o3vvBpWJYe4vjETChRbRaMnuHOab2Abk7EMHEKNZt9
Rd1XwCxId9M1sY4T6ihMhVTttJdCVJEPatFNCSDjnCTSjgqOzwf+J8oFpUYLHzlmqqZvM8OT2oxh
8U8BX/8r+LbELz+t+mfRLrWMtyjsb/9WFcoIVQcBm/TARmOYGurwFFyd7l9M6FjDRj9tbHEcCs5Z
cGbpjCACMT7DlVTuufVLiZe0VWnNo8bvp3H22TlFRzay1iMqvCH5yYUC6YaLgk9onjNsIIlrNSBF
DZaKsEHsQLA31Qgcdzxtw2SEoyjxiOS842kQlAqdD1q0g/J9LrpRjVIZArKPq/5eDrotNozClEnF
Ms+icsv8oLK5UiHBPxKBk4RX1rAd54sFdB1a+BHp4PvAVfMBNb5NXqYH7tkrogWjdnUbil4jQMn5
Da/f6svZ1/1xTZJujFgruimYR+Y5XOX2Lq5mVzIgv1IZxZ90j6rtl2rpDmwA94DOC77ePWKwRd+T
e2j3uLTH07oJS+F7LMF7syQ8WIEu5UaMHk40E09EzWCGTtAQi58JHEfTERo9sOsYgyI7NbQGWp/D
rZcFhOk/gZ1cWgVbtHY/HScJyujhetDsYp9RtvPlGrARBFbwIeeI8wsIWot7Qtad90cKvdhG1arB
0MqjCXWua6+kAcOC4OL8xxOYUu9D//qlJdB5drzzRIjiV1YtIsPL6Ww9G97CQ97SSK5ruOsZBShA
S04bRPC2wf5qKSOztXVv8GPZ9DfKWVVf4qztwyU0kOLfMRlhcgKiX/VVNfEvfIjrFf+/YSVCTmtk
50fM5aclmVWotqL3VkriAd7D9wQKxTwrfhfNfcgkVJraGajKusKx5kWiFEdjpo7bvnj0IQhzSYLA
mPU9kpHeDvqa0Ll8xqVZ+oRXOsVdNpZMX9IEVaBNHvyH+jWPpYHDm/RLSlIPb9PoXCnxGAEc4xEb
tJDz2Su6oFTC5B8/VDWc7R0nYvC7HKrxESHmAp/I3LQs0veM991Rmnvyu2vQwwFHvrhwZvyP1aio
19NuE92ionX/PpK4i2B9j78fbDnJ4JWq9+KI9yz0jIslQNpF6YhhV8CL4cFRqb8vcRPO1pfNVySI
dwMdxesg6etRZorbagj5pLytCzwSctqgvuAj7LPlmyDnLHMxQmYln/4c1u+kFGC5Tdct39gnZF4U
akXJBC2Z4s9BTapKl/x9dx00P+fvRhD6/2ipsHLmVC+GB3ZEDEPjxWMVRN7UZ/8Zx36Xul0DCEPg
Vw5nnJONymmSzuC7FevPEc3AJU1uAjmGjXym71CIBiyYP+PaUSdDVn7PNXwQjrvPpTDrpBffwY7Y
RLpxqAMB5YG+DXcxN2CTh2gw1ll6bRRrcsDBU8KsKG8RbNcr95IhiP+TjtNw3NK+maJs4bSdbD4l
IqpikWDANzdDQ/nF4Mg9B43ImsPujJu5v1J/gPrkDz/ZeMxRbySru1PJzvS9f7dVYCXVRkjYApGt
oPcrFTkgTMJqtPYJzNBLyRlI/CCRCJ1bl98NNcZNNYuQImtex8aAk/FsCCow3lFDSt3bioP0cq2F
ZjbALrtU4nlUj8FT7rvSpwOAI+r2PC8qmB/NzLyVUNCocd8QsbpQlTPg0+EgycEBs44uExet0J0z
wXonYrVrNITTPS7mz5OcQXYV7R0owlffOIl4emRLZv5zNowdBzOLuvLs/lzWKoiKBZiGYfOaJE3k
fB1ekCNlpj/dbsMIw2oVvaiXJMsI4pFgPBaUmvfwfhrOL2RF1zcUoIrjzpz+4fQFu0AWsb1JqOMx
EBteNhqccXjUhQioLkWUo5y84qcW7bzqLe3zJ/RobU/JjUXv7FNZgjTP7kF6pbcj48Q5cTaa3mBH
rNNGspxv2mmJ+jbCby9+HUWpR1Is04bP5iGRhKR3sl3/0Tb+ZKNMTnJBQGumCAuXgMMMoE9cWfpY
dZpFWXq9zZNC6BLkn+6+tf/CUxR1U02IJmAf655i+8xI3z79XOK6W9xPsu7tajMSYegzzVRwSLBu
Yn6GP0xLk5K1B/Q1k5inXDn4oD+sceANiPOgjkMNkRD0a3j0TEO64cHBKgjDPvMXGvq3WfIS+z4k
JDg/NozgEMhvz8YlhG3UmHnzAH00R3/SXlim+BjNgCc3F1iqJKnxwuKnlrS+dMfI6evEMfh2Xc5n
9m7lEzLtNCp/dxkKWQBxUWmPFxPa63484ewcAcRV1wBtJbagEzGh/xHx9EK/nd9GPV4zLLkVLo5x
DiFEOHkzdmeOSGB3GfWYeLjBmWFB1UFB4yp1ze192AOb1jWqh+0t4naiU0KaY7dUcQWFSUQRIalm
llT3oB+iNfgiUysXdlwl498N6PjUZ7ZRWL5DJb3dO/Uz2jhiyFGVbLUI7h6ned0SjJli6BEOXJFn
BU0Yfj3EnBP8Tyb0PLbfLAldE8Hx2PHBZE6PxQAWGc6dAuCSheZURLz8IfkAvjw1hYQ3NO5tJX7N
Hd4A2rlpHZq7mmW7kOnHICEvnvwsH51enkVQCjMRcK/eieJGiO2O9wRKjcMI82lkJzn0EiXfVnzn
n4e9VQElcJsED+/P7wPxueEADR1I/EQaDl9xX+EEzE+YGqixPrRJorBNujgaFErMT9SaNqLOzSBs
dVPZxRP3WHYpxu9W86BnjMb8uwimLtaaUI9dnzu5knFDuRKMH4sxdk5ZCycdzh5xoSVKlO3bw6AC
OLtSPga7lKsvfim15NeVdlJ/G0zquaEaqb6cCGOcA3RVSob06DYQMh3RhKBD4G0P1K81xb7ouklk
Dqe3NACr2p6Ztyf2luK2mBZCOzh4G2bE90gbuHJKFCCqLNfCPtAVHIGkjrD6mRcyqMCEFT7uJLnI
lB0N1KtnBRaGJEX0CxsZOBey2FGJIJymOFYWoSghonGOAKXZcTbrzobGsXCUPOtFUXainv5H75RV
jXiOD145eTx/Ck/45ma0AmCMMc849+GdBiVn0eee5T96aW9vJXeyQ4ISQOwnO4U8NwXmySTOAr1A
VBi3+oM1tFg3ic8/Z0ku5hixjuynVO/4JLwXmNCxHASFytvT8CWHalkXZwha50NB810Npjyv9AHU
f0sivcCnA92H5g9EYZTx6bX5x+A2iNI4ZPTjLbRGdBGRoIiI0NJ35IxPFBA5GkRTAdXCu904MFhH
O+Bq8Gqv62WtOiHarpLsPEM7cJjCvsjll1eY3TErv7h6Q3j/Ye/hFPicV210Hn0w/C98RSwNYavW
/hLzajrBDCk/m/wlY10KGwbYrXfLlj+D7tVLrGKRfgnlb9YlCbk3pD8F3J6W8ipuCw7Tl6B6blAQ
TVzidUZnaHSETOUubTLufM9SAbKFSZAABmqXGybabpnNDDwcaBaBiScZEZ+YBWVyMhyaJ5U5edf+
V782x7rTQymzajOBI5oMlD/+3CJqasb30u57GZE77dAP4ci+b08oSKLKCOI2ZUzKcR155J/MFqBz
hOZAb0k+iF6qn2eKt6Ccm4iHpXYbWHxZRfqE2xb1C1OpgYLv1Bsp0uPABiS4GB1JQqTbm5SSNsyl
3H1TBjbr+ODTAX0pQbPbARjC1jJEvRmULsdyIX0tnuSsQOluN+i8tkje3CkHUqt/E3cd+mTVSpVz
Iy7o/ZJCbWTlyMH3ZDWz5wfnnQsAFZhqDvalR5u4fph/t333ut+JD+PYrgb3T9IWW1cc9B879fhv
qGHH+v1M5myRmTWnOSUU+UuCu5D03slt1OVeHGECvPJLXhz3+dY2d5m8WzQ+wUQM/MGQHKaqWYif
Vu9S7J9YhD9a6SZzjS4HId6aD8mM0C3z6sLJirnyzT14jv87zJoVYIB0LiMVWB0VIv+XWdz43+SC
RheyiDQXc9wys4sQcblIh+aN7MV2HfTCruvyORBcKFmvPWiWUGacumtHHRYQCYHbksSG90HIssan
Sak2HkvKt+qLkA/Lz/yRfrw2HMy1tuR2N4ZMo5mkuXj66oBowL3Ucc0066WHfuOhm4zj60Q2ZbbL
ejip2YsVKkoRopR33SZeEGyxmnahW6Npfa6nSDtEqW0cayjroW7k0tfKsMhCIpeAloVDY53YTzWN
YvYRSGnSWEwq9GrXcaF7ft7fKb1GM7OUMzzC8wnTJvkEJCt83GtbyI/y727kIXt6XSXxPipj/qNf
B8EeaaJgZqe3SFWL1bGuX07mXSpNa2eK4zl8P/BroqXiP4YHctaCX4iT7AyaM7ei5/U9c1Bc3q80
1aTk0Ogjmnzg0Z8N2+dwrOLgqfgb9EqJjcA2C5TECuDxeIk2G0kgYjQRU33toXsvDmWaXwXnhNy9
gKybfTES24sIvO7r0ZlMy0Q8bgB3Ir5GGfIpBs5vKsFVB2euFjt7wcfi1c/5HMHxz1JXzEWgWI1R
cRGj8wojG/80i6pOp9Fw7VV2+dSRZyTkoojqTjf3BAoRUMtRD7zMvyI310pFOqCiBExL2zAodWqJ
G+SuZl9oFkbU5+N4yLRvBVnyHZJtyAjJqFkyne81CYFhwaLEDaHGLEOmkIBzMqOvtxQKIRHBIY10
2nOhkiDxFRP0m3bk/JNe88L51a94I5XjKgRCqVXnb+lzMxO+wgkbRHdgdPsnJfdig5OHDUnGjkok
CBCEKMcI6tR8V+zpKGFt6z8u+GH0ECwRZQQwgFEMCFlLRAAmiCb6x+iQ/NqZhuuuT0Qjk6qQhcgQ
cVte/FGnA7s+Bv5frVWRJ/aaP/6/Iy321G4ZjG2gYfIG2BHwI7/o76wBF3tNqmmve0xfi3Kydn3E
N0I0BqHx0Gt6VUkFSn+YTUMk39JxHoUv46NdFYdps3CkvSAxX3oXeGwbueAL1H/N1gBgOcskiJJc
piBmLe1oTNCITMmqQmWVpjR84FLthBRk52CvadUYcpX2g/a++bTvkCPgTUpWe4N8Nd8scIwTJ/9e
H+zKBG5MTvrEACHekPcyaM3Pmdf00VxBhUJI/EO6tBLUwFuNlEqBE0hyP9B5+AEGNN9NAYcaO3Do
2opXPsjyYu4MWARX6PCI5BXmvpO7MQVkP2Tb2upbfiGfpbzwU7RluAc2336S2o1sxJz+WtSbUQjh
Eb6NDVzcpfOSpLhFb4RfeNagzg7WGc/a49XNlQEVIW2YSsMwTGf3UP0CUpuX7grvktvSQDwE1EYl
/MPRJnO1Vy0LIw4F3Rt0yxR1dqOWNHdtJbjjD9OlFwPwybHvnhhXo5cmIIoIMeSSnCWw+Yydz3/h
jIHm2Fyi4A+L1DldhPYhMJ7gPm8hX/kadxxYOKOWk+kB1kVcobT8uGpzSP004nnuGS0u70ZYptEa
QEgojs+/553Y/Ado/MIoAfvQ7S9CVLuopjfjzPZbTQWF3sMTh9R/99d2N/QlDSSqOcLB4FhaQ7Vg
j3fGgsLdipZWBpdr5G2L01ZjlW/KWGaxsuCLJmW5WL2hrxA/JUPF6HWSaozI560t8xW+QFm5rcuj
z32Mav0+Qso51lFgS+SUzyrOlGpEskQ0N5csSU/eQLDsXIYtDqCuqdAPNFEs6DrezqBSYik0r/u1
3zV5VcZkxvbXlm6ghhQ2Anyuh9dqc4QnYU6zjCmicYlQnWNadpmSeibsln9yYq03rqMCOPJlJ/og
UU0cp3hHNBgEOPvZoAWhC8xUJON9sKPx+HzYfQ/B+72Yagkfu3jTaWHGsQJsfa88pjImDJ4vjhb4
Ilu/Ntfllp7VeqhkMFC2n64qX5FIurE535WuhgQ+lkzG5BJj+OZCUelm76MwuZKNK2KSKiYIIKeh
Q0A3LD1dR1/wiosfS7o29r25pgnxvXIY2tZ9pv1KjtB+eQWYY2FNCN4Im5pC+960hQLDswTAWBah
4o3Zg1zD6WKLcUdhwM2cI4rnn1xjr8Q2aaePWi5RG7InrX8pLEf4M+LUJru3bm4f4hYIHnbYBPJU
wLqZ6eux0P40VGYAthuVGlpUIOevIi3rDoz+sDTZ/iH+8MW496nunrGFknnYLvVaebOHUuu1oI6q
1k+0YLpUkEBKjX/9ladFV22dKDjFvdG5eJ2JvH79o4mWRfuzZAXDxsiPdoCcTEmqNLKnMNArwiZn
YpM3y9jDEM7QAweeam2tatAHHO6/Jo9CdGW574hB0vtxWCxSPlo3BXCZCTpvohyCVRYAv7arx1zc
OmDxdJLcZvUEMdnuN5XIAHdVk/NKT0PENZaVghlzv5HdVVO2LwkPJ/dBqBAfMAWnRMw0EAa0J6hA
hSpk1h6iOPOovA5bAiO4ScS++8yyT3BREimJsb2d2Bzu35/vMb2jSKwcA8IjPcy0lkaU6fIiAJ8h
0CE83PFWfiVm9Y/ehPYmF011WviDwmA+shhbuWvc9vEU/qWn8d2SeZ/V/XXsiUWGw3/qCGyGyzjS
hE6zn4GCr0r/LY9glSXv2w0NkJj4RC1vqnRzk3pKICGDLYUv5SVq8V5paHbsCfgC5Vdg2JB5IuCZ
6Nd/Ta5qR5ETh01PGEAMoGECSl5FmleRSUYpTHM+7E8XcEZ/i4BHsA2NTQqw1e32XHWKznwWnUVB
4FuQ13KzYlL1+mfo3wHp8OgMKmSphjL2ePlHEyhcOcC7pvFhOjUH2D7tgxykfvEFwD3lxkQRU9g8
ayNF9AcWoMzm9aXBvnTihs4Ln1tGK9VzXmY1s+3Gmbew/JTScnD0PRrd5MG0oJe6MFXe6DWhbyJ3
lZwPcBh24puUBRqLVg8fVaeBes+Rr4MtP9vL16y/HxpDW7t1UC6NPQsjY8bnSt6B507vxgWiPsSx
iwmiKayjcQyWbpEGL3FsFQGk4wNbPhCa8irmSNriE9T6V6ik59BxcTBgSNlOEz4PQFAHAbRtzDRv
Yx4fyGXrz8VMnnr64GAqBS04OYONwyQJbtYHjMxTapPsE+krBtBLch5ZHG3KyKM2aIs+FQjx5O92
IkwA4i4U+Kvokbfp8FmFAD9MgX13aaiux2vRh0RsDotZbgDcCfpLJgMndisqoRQE6LAEA6SKPApB
Eu6BkhMffmrCDQJagHtJ2T8X9J3y/93tRBGLWcIdFTVFGqJAioy5eAtFjYYCmkQMRmVRHxiqspkA
K/Qegi9E728nq5Y9HIQ9I6QXV+FOJ/PG55vP2Dx+B+MSR7EQ9E8FyssIWgYReIN9etAN7wscgcrB
Ly9vA3t7qWzBAGZ5XeMBQTCOjvaGCzn93xg2n6QGLnFn1imhUZZGCdfu3HVxh1nKHhQTSjRgODgu
8m8ikGuLBSeTjta65ERZP9M8cTr51MzWHF9Rv/jq4GocG5xgVQjDPNCtX78gJXSm/EmOPVeeZMr4
k8Y1scVvo79+lqZ22/z3g9tl2QtIDll++VwnAemLj1T72LS7ysuKzeAknlwBmaKid6lqn112fjqx
4v9D0XcWgup67YnDLwVl2ksTsEaYwrABOl5vXaib8EHllIeqKZ12QKyHhnFBV+0xWpzZfAMSmOL6
ob6o4sn1ppkaUBLjk3/01s5J7n7/mB8Q/2ks8V5OzNR+sZVJyQc3kalwdnQ+KJqeWJr5wb8JQDV7
lsCYOC40etBEpMXCaA0vAgvNaTvgXqvvnuRipWjuTJ6kNhrrsZfCMeSApnZs5kB4J0wRnRlPFibR
oyz365cL9wAPFME96Cam0NAFMpAHeyUtdwySxoxcL9Tx5GyX3Vf4vqC7wRbCl1agV0Xeb2XY81RR
wmXwUOR/HKOoG+JgQbfm/xrWwq8vpbSu/N2B2FEis4DEsoSXt47aOZWxvdsFzxyXZPoHoCdq/CHD
JJEghVrWk1WKBHN+oGJb/jj29gx5KFtPNZXqZxE0Huv4ag+2lvkA+pitIvfd7tq3Cqy7xoLxL8oj
rO8sERa2j4hFTwPl7Mv1LRIhy40qDFxFhywVZxH+4vHP4b3ZsbzdkBA8JVXRx/5H2UiEZ8UZnZ0N
esxl21V67YzSREmdL2ph4hss6kg1F7DUcy1GdtA0VqQ3sEiO6oj69Neq5U6t2oGLnCjanVx6JQDo
iqUj3VMIfnZC6Nqan6yW8DeVHooDDmqxRZ7zcS506Ozgb/gkwRUj79eOrtkjrNv239XO00o9Y9k2
8t0F7gUWEIFJ7MvFzgB50ceQ9xkJbyfYe4mxVM8ileRj3GjM1u1gUjSXd3fgUghzfw1oJ1Owrvbv
Sv72K32KkSg47IKOHhhLxrVvTkNYFjQScX9oCSwDSjotElhqQrEqSFssv+SrQnIJupc1fDfbqNt/
qPZrSFI8NSaSe3YM4TTac/rUOgM/oVOHLs29TWD+3RmF+KcTYUOqE5XBUVnMmVMmiJUlWM3mBD3u
tR9I4YtPOi5bOdrpeeLEq1iwmdPYUDrafmKmL7hzg0y0TydaFKfQxRMvHLha5c6UOGzjm6HvyUSL
7sxflK2MWpS6I4EAK33gnH17brtE/s/JFQu0ZdiXoHJNssIT02/KNlDgcfMCsGA+KXauPw3mUKJX
PJ5dZzypikfYuArz7nx2fcmEknhed5EpWoscbnkPe5zuIMJbqDbovOG57BQM4lM2PthdrGcCoFFL
bf4mXhoS3sAR7kFyHmi0ejODsdgiRHipO2gFYDnwwM1rRhxqJijJdNzs/1vMiYCT5r4UJ5w3qQPe
FttomOIMwZg/PGeUDvzZQKz2Qo23hJCGBlvOhuqxRclIw5hsIR8y5R1KIsuteWO2Rdr55bwll+zb
/DFSAgczT/9KznQWa35Bt/5x8sSptnT7zXTckYf8Bm8x6RiBzmhfi9uGJe+0sZI4yMCHBOuHqHfE
wl1Rrw24ajb4XgNeAc2xuADHnixfrw+HmO2WOQ4YgEiMXslDn5kSSPUR3/zmZIEuHYs4SiVWSJDa
EWHzxwdHGgu+3zwndGEkdDHpkHVu0piEv5DwZe0SDhZdLmDKa57YnSV/hvkCBTPMu8UBTJwQP7ME
tCpXngE8UBv+rYwp617oTeCbvVGbMC3g3vI2NGNNsnsiKXPvElVtO4eXTF7BdgYqxEhuJGbeXY0T
Po3Ob/uXwmSOI9lTC57q9Z5ldG+R/j6THUQDuJtINUBgUptBR3Vmts4R15Y1BmoMhacn0DMMI8Es
A/d7JABfYXAajTW3LvkWRIkRJJUdS45xrd6fkSuE4wPP7+WqyQEpts6phvVc6vVZXrzm1WxW45B+
SIxXXDzH2wwsM4sHgNCzrb9kT7IGBRxsvaPFgKYQ0285zftKM2kjwqVBu2zvxGkkClcZQUwRylJE
Kg1+bx+C8IatDD2CpBmY0wxY5pck43q5hDp4uYpfWk3O5RGdYQiiIwrhbPH2U8kHAYP/LMSiy7Ss
x7Ru7My5VFMbAHf3/kQRn19ZMfYtVsN2tHHNobpAiKm4VrptdQtKn05FWVzyCYairF6qUH0wiGMA
ie7+2KXtbv9I8PbdayL0sPuyjQ7kdgdq++kc7vIogDDy8YDRDaNSKtcxIW0NXVcZbZvdV7CxCSNL
DWMnQhH2R/Dthwnp2B73dxezIk2yAvr62LxNTH+f1TssJRfIkJlNKanuaXo3FGvhz1dJPLXA3GOB
g1NoKa5xv5mMD/Cr+GVi7LV71GJmZ5cSa09p+1T6yVxtsVC/XBeTJq5MyP36pS/xUgQJE1XzHIYh
C9ke5ez09uJTVFwwq78/ejogkVq4q6/vGO+fVlXwbuo/Xsn4VRetSL9jEkckvpd26xZIBdlGy3Ir
wMeh8GXij8WVHNxeu+2sg1W3SG+67IgfgFAFA2gThty0KOviWZ7y+tCh8Y5cJED5EAhjnjmdGOR4
OtM2pvUz5S7jMrpS7g0+Cc/eoZf/9dM9HI08SqhlqhXrgsSRunTmALm0QjT9iVqoGBnEpz8EQNlD
35dBCg5Be2ph51tkEw7ALZIpGod57B/eVgHUSB82F+Vb54S7Gyorw3WJETZyTj1Zar7akpT/Coa6
L1G432B6S9MCXnKaQI2BjSh4nPfaXv7S6sY0nk9loOJHujWFhikWlVtrQ1pyRFwvrDYLYlQvSDN6
6xfbHYrBIJcQOQ5n3zHRKBKxN5skLNrlWumibMbwTsE7WRHXpmQH/vlM3mV59MBeZfL4M6jnzyr0
7JnGsRM0irygwt09+YiHuVndEoEpORL6+XVybhMchoZlOhQQieXeyKbWbm/0R2Xxj/hJyMmkLwjo
nkNKvMaUzaUDWXgKFn6xtkw0ROB2s75FOPbnKCUpbVLDnBvCOSBHrezvdXHYds2g7lSoeyJoJpjt
K+dPB6zyDMWItM/1YrAyy5CmDYO/3nfTJYgWAdMxXnoy5Xo7QTzOYHjL7/TXqoh2L0m+qlVcwy9v
3RnzZrMUNCJR97UJoi4rU9X9/4iz8i0zQ5faephKgmvh20SSHUyt9JMdvTGVxPQpOsF5JxhvqoQj
SiLbUV0U27WRZrMp+8Z19NCUhd2DwRshjs6Iz2Tuos7SGIm0dKRzOj4Tk7MM1Jor1GFZBvMOMCoi
XEboGlwl7wTWj4JK9bcCtWDA5ZNUrvVNW3TG2Dk7ktr0Eiiy8qIt6dfC+H142mn3EyxLmBYIKlDa
1DsA/36KPEz5Ym6ZEJTsANVuUeVJn/F24G1/Y7MCeMz6sqkKIfsI7nb/KmwroLell68KKEPo3/20
qbUVM+5esn/4D+Mm0qGJ+/ZeWa2Phcf9UDT1Iru3sOixhZHrVu9WCAsLoPeBXy6Nu/t5fb/yt6y9
g9zVH5siUhF7Wy2vs3MWvNXZO4UGAmZos2/G4byRrGN6uNIuY017TxoMkBBeEwcu285R3IHxPaUG
CbBdhcxbP/WMSJYRQFqh9MxkrckiU+x6zh7ollcvaUQQIrvNOJ/Q8vIDX2yXDwQ6gKl89RuvEP3I
94Icr5OfH4Od23T+TGzNnFibrDNiTGYnZCec5/5Q1idg7CesckzaFovdVcHd5dvf4jixf5wODFs6
P0yriuQ+ntH96rnyiZUTcLndrH9mPoCx1X3QkI2ML838HGLgZgti/OY2+52+WVSZDkacix/hSzik
MUJeeqS80Wgsy6qORuTKjxz9e2nxb/y44trdVfU4vT2MxoMf0eMmgKJk0szvo4f38cPV2m9NfP36
ld3uHVF1DcmRigFKf5ef0mIkJnFBjIZfmqQXJmynSyRABvBuoixLkVKmmAFEFT1slhhqZNbdY6+g
8twbHcBmKSsJe0LtW6Hav06b2EO6AUVunUScwoyfVUqexkZY2SU4f9LRiE6rQ1gu+uzWPy74OX8e
lEfIYeCDfGk1gs2XtpBD3/bSIwCVIEDP67lnsg9O21039WUDBD2M4E8ZYgfErmWYackJrNWmxveC
0Mvkz0+s2q0bVAftyiqoScpK+VEml+lu4upzIamKAEc8KYQ8tqIe5PpFGRbXnR47SAUBB5cu6Doh
tcIjmCrkVnFrSMb8bj1agc5XHtB9GTzjj0qiekAxC+RfVVDrLmiezgO0Nc/8HqQi7NSdv2e/7HDV
fGN5NJr59uLhsDerhLFBjdOOd0r3ECU9hgccqlyLKJxvT0bLlErQ2rD6I5X0p/bQwwLJ25QTg2Pw
EIkedQwiC2HoCBgVXAC8ZzvNgEraqpnehb3m5UQx0TQLKxk8lS2KTb9xRaE00+xvoCGi9/r/00MM
oonhpH+3QMzH0WxVE0oxmUyGTHaHC3ipMs0wx01uvUycdIXnIPq5mBbceF7RduihC59KG3KK1SZi
ox78KKPTEK4Yd/eRPhBhVMGZDoFzzJXY6wtSJcCVmmsY0nTUKYY4/jlcTXSOkJ11tq2kkE6kRV4+
ka3CFD/RhRfh3wFBT2TFjFsQl/kAUmgvixRik4g/NRw2q/a8HkoJ68CMse+HjlmiBjwNZsl7Fmhb
5mFaQbbeDGsiqwMB3ugMKXl/BiaY+DM7oeSynaZxqzSFZ9kJY9r2nP2Y8QtN+77hYIePwwbBC84Z
2OnGSEdr90kuEYVzfVPYfeIt7l/WvZ1ltF++5gG9/pjrmeSiN1GlWSP4NVNPvOiGWEPDTmMDKs2F
uGbhwQWd1lDCxX3SExIKVjjJd3v5TFErulwg7S5gbcY1d6NPIfOSLRVg3Q5XqUiRVPjpYhwN3Clb
dFhPkPVv1RXuIzH5I+GFWZkPZYtgmUhD2M1fztdMzfO146AGsTAQyFrl0Ax98BsFwpRgKMdh9sxJ
kPu4G2zHz2mGk3F33mtih0BwRzhZ3paESE5WCNPvltBG2A5pli8Xwzf9Pt5ehyAfWAdPf2VFNVDC
URp2sua84aBoejUh9/kFbihgJDBa3ogNjK0et+Jl9KPcQLFV3KhtmzMFfXA8dWrFiYfsP/9xFpD7
iK0tAyMK5jm5rUROfDUbR/19dQIUmD6TfQ1E6mqUGeaXNlhBt5jNMK8m8Oagr8Jj2PQ+FVhZ2HwU
Sk8q9DLzpbMffqRVm5Bam+xdsBiLJFU1CaoZHA6mKLKuwmBQlTbsTFtjdz6urDctuowAUEckjT5L
wBF65GoZAQsvSzqglhsz/J407h/vP2LjfHo5yP7BhA1SMKwScidbm5Dnv+ywuRQO6vtBGBIwQCvm
59NKOkZW01tAIoZMR2IZGwHv71ptgQRYlZvvmAIH8Ecm8b23IOCHz6zroKaVgLDbbCDkdY1qxyMh
mVZ2g43hnaTMw98PfYSWI1Pu25gCIcccB8thrsjR1eiEhpKHk3gjxeOKRohLehn+BD723k11nhwj
z19qDJPZpquqc6EBnovR9PJLKiJ/pi01tfBKLRM+WRU/WlDEnwt9jpb0aICEM8sc052L08MY1U1S
vtS5oDA9DNvTig4woBdYAFJITFxmfe2frMMiKeoN4GaPspKaXRiby81iIPMnny9d5+nkj5dTPirS
/yioAMC4ImXzB86+ikHI3DCHwwitEHGdP0IkXujvfPlIRhSSbkFGdPwuseuJEIe7KNCUysCatQiC
z7UkQ6qJFUKgoQItD/xpH5EeoYGkb7O9LT8pI2byKalJTjeyMw6s9rzr0ViNKaCFw5VRaj6vVtug
cXWn92rsjiA2sxN75ovitKSPTGH/vumtLuWymd28q7pBGM25YYBHjiRt3t7PHnOYKN9UHFaJ0/b/
Eo7VVJt0f4NmWh6B6q6bXYfj8nfrmjmge+hOhtiBwtvd26uwxGHhV2+fgTOdoCl9pROU69iJS7Te
SUCI71FLdXJYvr5exKq3Af5+hpWLdqCr3VHBn1c39opb8Vcqf6muWn2l9uLwKCeOtJ3bBV8WDtbz
37u8Oi4VFOyz0JmGaXLINofNtFXg54KqcCJl51c2zlD8VGiTW59uLzXrm6NobwuDowX7vb5oHHNt
svbbwlSPchu0FkwqbeR0iCokCCmrPtJ1Z6qM8MLUewtamSH61FCFQ6EwGWldGX/wCLtdpdQoOsXc
5A4BbgFC7VBabZRW0sNaOvDeIyaOBWTEtJITAWiBuDN4z9ojra46qJ99DRqLZYjvkeTo3rtyrK+J
QvNkzF6iOvNtqBwMrBaunCPCLpo3YTlnsgEkfcoaxhI7I7MVmLDaqohJmf4TGf4alrcDtiaiP3uS
Hyq5ZFASgfxpst+YlNz/rSwa3HMXxspMX9HaU/PI3/fdqBfeGCxRSA3Wthmont75vvkWmdI4cVYR
aBGgDA7VfMEd5GuktIjcvWe8fpRF5qtOrb7NzwcZ52Bf9VpU3vkm6xYLSjZVl9uEdE9BcYvj51VG
TkggvLp7uXZWpxfgKfzYIVj5cPiCed5Gp6/Xm+AP+yY5Sz7YtI/vxzOnO4QmcWJ2AUHKiX1jip6O
KRriDITuuhen1n6TD7ursIiVVvI6tlfpZaCyh3YzwW6KdMnJPuTtoO1+34lkfvugIkcrCdl9WEYT
sW+ZDq9CioGRIVygaUqJD4h4IbXEPgpJzRWEAyqmc5j6viHlivRK09G4CfxcZUZVYWB2vZn5yRrA
/KJiyIqZYHukdQzwYhx3OuTxm9M4cNBl/B4ihbEkHkY9d9K3/jR05DlU2txse3NryveAvSJFThjk
+19geIpn+pwiBZwKrnCNeIy/hZSVRu0SEazXIhElg70XhUTp1B5y1+oeVtDJaKZ+uf6Ii6vnKdjW
gFy+8AUQ4b/+Cwh8ygpm0bQhtawmvkAIP8S5M1oyTw2oyJl1c2zeBI4dvUQHnZZZ74oIr8E267lF
Abk5ngflBUKgQsKTGmhr9nEfgZTHC349WTZMqIGBgqkzjv30b1Z5HvfJ5frMtU2H/nvktpjUDtVd
qNwW5WllrVG7oyX6j/nOpOSxupcUnXMEEUWYou5ZOO4tldQFdwbNDndcsTyhWfR9GhGE8n3lanj3
sl1t16m2mf07GECSycOCbhqcH1AzV1KigbausqTbTqVBeXYZNxxVFHIwjjEI/qIFX4kSVohAUih1
dUYehdXDZOJvLhJdsCYcPsm7zSmkZo9CgAJthwCohgv53rQhpeMdJRbY6oGKWMTVxaScYwWViDUA
7mAPOvELzHbvfbne7tJxzhQJ2EI+wWrDIt6b4GZUd9W80eG8AUdwczG0egPdzMcPUgLAwvFI7s/8
WXD4ZLInkLPtpKTekMVMWiKpN6CR7DpBhIJZ/KRC+aOLUusC9x2l8JfAaDiopsvuetZ4hOhOTVMj
n0+vqEfa5eX/Cn317NicKFVmspNrWIPR8VR8gAS77XiJfONua6c+QRoQgmBsq+mVEvIMlRDdyHHb
9pu2tpSYfUopzvpwMP6o5Hz9q6dgARs1irMUI804/qrsOLOpFIqjgN9TtXSQJKR1gXoshU8apUap
r4MrZ49lraC2F3m04PV1EmZd3o/cCvlYrSD7xXTZh8qk4DbAEx6SNwef73YmRJzCuFXZzbrMATB0
yog5OJAvXfH+tGKnKHkO7kLkZ5tQ91v+Bo5OQemccwBRyuv6WQ/F8XEzx4021MYRVKBcXfXrP/WT
8WidmwQVDzocJ2ekfIcOW3YXz2XOdKqDAGY007RI+2bCkBheSbHB3kyu145Fg1dXp/EKcGGZZ+5o
Nb2pSCiPny2fCTadvaAyIx7MLninQHO3sAR7EaHA1fLRxIUriCGaQ9ONG/EPqLmazV/xZkpVep4a
2/RxP/5RIu9fWhxmCW+Ug1sYLEakSUxMMUs6Po7B0YR40H+MjZSDm3rPzthuK0h3bMwYUjFqKr7/
wzd0jepbhUpaa3JzeYSWAygQlWq2mfhTe+Rp6GwqUuCG4hqlK8YUofYlZob1pAHGXOjWE+Vuw4OE
oU8w9sIHR6oUPiTwAWpVbeJMlrInlomB14YiimCCHauUXMYdVMW/omFxHjNc32uFRVFhP9ydtRYa
SVVBWeksoD/EkfNvkzC8j3Pg5u0A00wpIUSMSj+rZ+f+vilURSPsGzxb9zaJxLKjvOqO4oPbZf0y
7NOe+Z23EkvrMhZqjsy/6R4/NDvG5pyiG5tPHF1VbkK2i8sXe1yfsSJKvwtVuiuDr2W3wDemqaGk
DB+3nQjn3jueWC/xqzqfpZlzSfv1VzcXv4iFx6ni30pgnPjKyuLvKX65D5d+6vB960P6du6S/scJ
ljbxO4WPsBgGd/Z2gc4kkrmITodBega8uGPrGTikKsbwZEpr2yq4rMxMHZYu+dZr8SyGIqFObxHY
g8R66GY0K2VmgeGyzfG2B+3Muppjkime4Ih3mdrg1doxLpcsddH12XNM3B6oljj3bWrhTaM0OjTD
47KP2unWQoVUkQbvkJeimZTiuDrx1N4nwqG0I+/+IjHTwTCl9q5tFjQgl1GEGman4uR8Oay0IlxF
VPwA/u9qPgdzsjqXvgktNmoyX1k57RN4Pr0sOMv+lf8ITQYHpJe0y7racX06HzaKk8B3dHTp4Obh
+lYqC71pDV3SQzVmKq/aZfik3DYWoyD9ON2Ap/gOubkuTLuIXPGBKw2bWyYqHp/1ezoRYeqVfPsy
K0HicJZVQmBVU9IPbShMS19SZC6OWhrmxpuwnSnUzhuauMRcWIbmFrSL2lpwNBxBkODlNOiey20T
KujptA3T00w1ABGXY9Qd+vSheGr0n21CSTCR4EMEpZf7+OsqybhuOGZFmKKfbOXjA4wFtrL6cYMw
IwIm/vZOtm2VMl1P751BBF5wXUzBq686tBh5Vyf2VdJJkmj/m8V6E2hqMYVWzMzZHetyvO5cR1zX
2LfqjyG8cLGVyVByK+rEG/hdqKZd3UFd+JT5pHO1mwVQumUIWF3FwpGnwrXu5+J7uASlYNhRj6yZ
fF5gSATCTBVf4JvkqNlZ3SCsKP+9zXKJccUIWI2+NaMTzlg0qOTbGwaaUurbcZxYJ864l/+4Tglu
bo7usnGq/RQrNbJtgwyRsjxTs0a711upYn7tGY9feG0uxRzrh6sC/S690AIVseRUYlunbtjjMu07
ivVQocbGNbySfcD6CF9tx0Az5LzD7DQQb8RhdyWvRp4Aw2MjxO2WBpx37ipIuFwIwRJDm8bH2slA
CPKAeD7pwSvZwY83/Dnw/2dxPC4Vqp115/jGFY6BiUVMbFjdptUBHlQhTbO0PKIaERNFGACrYkMK
xRUfKkwPGfTWFQ9mEyAuIW8gUKFZvmXgx/V4C0iS01gjF8OCkbQlDhRQ3TR13LO0MJ6CAdtEgG/r
PZtbiEmu2RgvGkDzxhNvQ1OyfLNoavNRxnjyKDr3zY+aY/3GwqYVRBSQfSieYEyLb47/u/+qDgar
yDYST3TOYe+b2wqApBHqnBzBrBGO1mYiC8ybBjCnugjIbX7SPuhtumaG1omFRW4OVGKs33ZHC+Qt
xq0tIRpag62WKBn7E5WOSv2ZxKE4eJeN3BvjJiv4W91T5Oc8yw/2+P2b7DHSSzX1wO4y4GlViF0X
HGBBDvQRBFmYet6MUuHSSSViojVHlBu9EPWpGZvTdO1YbUX1Uzvurxm3qn6A1ie8WshQaW29nUcP
sVcBmNMFa00EurP2RglB5Pbey4Pnc06E7KeY6a0EgrvRwBpeeH9u8Zepz8grpG6Fmqxw+SNzqpVH
w45prTz0KDMIFH3icq3+dcwsJ0ErP6Wjlhz8+fbTeE5J/mJQBbIedL87tvO9GzR90tiAdsy/xIdG
+JHLGc6urSNHTYkPy2J5eZoG1tzGVn9NzjS+pE9qyj4wQ7kCk/3XK2a2P9AcO2bKddS7OTFVAuzm
6N+1PsSLzMlf8VrVMF49jP2BrX9gEA8qTIxBh9nL/+SRO+JhUyZbJ1dFKGgASEp4rWi6jodaZmNT
juA87Zbl8oPKKfR1X09ImeVlbH/QDTcrq52adzPyjdX9CpeWoCE/M3u5in0wktzvkxxg8Rq+26dk
mbCwcMgBk0/FmUmJsH3DWxR2OpNlv0qyxacD650aw97lOXnyF+VHpzmxh/jXlCZvWALIg4al8JxR
hR4/H/lRdHe2dekkhMyMl2H3P0HY/jtUhj7eD9fjg5YdsU+Du6rlaTiFbm/eJzEkmhlHw+EUbizo
llMEDifWS1IIXTNYMDQFCJShFBIQ9DQY7m80AkduA+VZvlvV2FRROS1IF3xogmZuMF9HWmAOcTIG
ZHA1g8wVIXrtBjThbcraX8XD9VXpG8EcQcb4IGfDx+XPG5StVggjYjLJv0RiK46BO97ebUrBpFYR
nTjN9ng923kOIDnVJNz+bd7rhnJwCSzFqpF+rND4P5ExB908bj0ZJXf5a1NIrJNIB2hhLI6ctDNZ
yV8aN3c0cTsEaWqWJgXjXx//UyWt7TFVjYWIxNklkPsZTskKgHz+rtj6ZjrioA5cdpwqtdwNMeVy
+kbczukES0sOimYB/XOsWZHI6+C6iZ7xVVFfSj2Rx4Wc9g+Tq775/ZrCEI911rlmalsmmRqGoi6E
jlLldtDg+6ewbRDrwptDocEEL+VOHBFfjJDxRlRw4xPkpWHpf2I/cgSLQrsJclopyVRnkbTWK1Vt
q4RPXV31zR/W2nGZoqAT1aMe0tOlMAYFmBgEsJ1Jwf1t8VuviyBrvsHS+qAPEzlMz7LrdkzqfCu6
plAFOL13IHlgeoBmTPZBL/zPGMak6LF1h5W8S/kKQQgm0+CSqept25xfSICw5nQ/SRJiEJ9smY4J
E2FHc3LWhGF6wvrpnSyvTmYxmcDuBfJY/TZefCH1dTXeyUUCG4xb2zdu4vnyW2cw3Oiw0ET/YGw0
oS3q6eQNvITbp/MyXKa6wP1r/Kxx2QqJSnljYmhZMydlwDE3tsoZFMkRVhujjbabkZbltWc2ok3T
hdHtGuIIdyY0hgZV/jBuHf6DaiMhbr/6fDzmDmTFzTBCxtddjfLEAtF2tEvjlq67/guSKQtIBeI8
NqRhKJ3ocymsQ31thyj6ZM/Fo0Ko8AbstlQCoqjZg+1Jq8qb0yLJ0nIfyzCvAf6xa1X18+ch5AK4
VyR4i/GIkA5TpjVuJ01Uiu6k9XTW4OgbUVyxiwDv2E1jAk804C9arf+PEtV7Foe8apMMaxI+btDj
zVMCZMPiD+J4ySqorY8UGuOM/SXyO4bD3rN2HIreWarPmvZQtS7q2rV/W5x4ryDzdsySJl3JimT1
hMAxRBqyC/1nNgT3kBpu3o69SOg9gfqQHdUrrD4OsSlZwou9PI16PM6eFVae3nGMSq+IWY/P9s9D
rkL19c6jd45Pl04/HuM+re8OkPaQXUj9amdJjWGGW8dsVlNwselyeOjqVqqRS02WLJmE9sSKdBMt
rCKe2ZEtgifSrT29BLUQRsQkdo2oOnZ456uk8JyTwpT7tX8WKfyCw7GLkoTk5GexI3robzGg9wCO
XHvJjzu7ttxSdHOSdrAAhL3fILTyiTfOYnyZBW0RAsc/MzuFWr9rXqPRCcEaBzI1HMpsFOSilmln
skLhj3+sXrAvtIKpnTIjp3MZ16W141FAr4u36+NQFTTefvNtgAHN4cB+P2juPkZd1IEgmQMAESoa
K0nmVC/vsvq50VnjpbBNjkR51YVe2BuMNsLQ3DMVyPBIBK12Y5iqnarK/bOpQSxTRuqI58bTuVab
t2nYa9Wvf9a2gn1Vm4pPu9ISrKaKRYFpsh1e8SB4O6WwHZZWGeA6IZ8lXy+hNHAJHzVgqD+/2yN4
WiCRPDv5O0LeJHN9c4dW2yxeCbGogNjCt+Eg4OESU63xdPXWk86E6Nor6pm2gMm7AUw+wfoS50lN
n+dYw6CE5PEZvIfHBk/8PnsiNOSj4mEb1TJJmElFIy//z2Mu5BwZtcVfP3hufa0QqHCc2etO4VvQ
wK5vG8nkzQtZSOVHxxcKwF9CbYUlEzwW2sX+ZXNjEnMaPAgNkvQBODvFYPObPDJiwKHOKZbd/cse
Kdmic5cLiTRuTV1DxQGYfobk5IZ9wWWR2VWXVOvfcd8m+nwCLfRJu6hDtS9Kd+wbI861sqn0OpIN
q5m1MK8+hRtDx1nFhahpxe+2XQ/Lc4uYK7pyWJl24uHPHpKkTS6WnB/McV4+Ne7bdxDWKfAZmERz
Fax/ZyJ+NGpfey7ARAlsSvHv1RzsBghLqTszzeLdKi3eDgrBm8fHicd6RJV0QeAorVCuzMKNN38P
RH+/k0AeyT/n5NMmvAmLXu1rAK2JGrsUAsfdBfZIjW1Hnl6/i89VusSFE0ud57SFT6q3yp8BPTV0
LTTcp3ef2w6RrL3l9sNW+e4/MrFzwfEke42ZaSBYhkn2hV8t+tyFwE9QWu43kFHw5XruszcMerge
iyNhkNm/8YYZp+sJY6bi346oI4dzQKzgS3Sw649yepAWVQn/W/HMyi5meqCOtRmynaxm7Ka5QqEk
zPh0Mq1wOQEn7wsTi+mhM0YSIlYZNLN8mm2Y0YyZJJ7F0+0Lh/r1Sdz6EQKITHFYWcXm+15I5gNq
rpc0KT1y5ihdhFjelJIhOndkCZB6LHiGjxx/dt/fUyHftRVX/E0ZOx6bZD06RPE9czAU5wlSjXJt
bpqGVymq98nLDyFeJfHP4shM2qXGEsEHmgGcZWCLrBzpUFbzUwhJjrToctQIlNz6rrgndp3zQXrv
xPJ3nipKlAnTJpky8wITZbrKocGiaeaUGyFzP1cdBooTCrGBq5aSnJ0+AweAA43pBSR/zFijV8/8
zK5NlJRXdZWdPF+SIZBZqC+7u9ieR262Of5t0TKkyxcK1XYyBCzqATOqrO9IFdkukXZMANKLFUPE
VyzHC3Z5+/9rFLWzl2piLjeHk/f3iJk1Iy42hPMVWQWzgL+e2VcqU0YT0P58MR3b5mXQrPWzO5s9
5j9Wy1Vvwx0wEJarlvGPSE/U/6hKWCuJOu5b36tWBnefk6KkDTQ7wXZHpomc0jZkd8TEQhtfaffY
611lRSwi3vS4UwAdkmUkvxccbzyI1zfCwybPGV5YadO9R7pKnnOv1eM4SflEERCog5Ss5HR60A9c
/FIIVxDtqsoZqI847lI2uKkfryeu87v/uPe7dmGmpeuzAH22cu7WKnnDWiOm/ZUz3QFYe4TqgbzP
NtizfTuH+9wtEQEpnRe47z8q2dDhWhoRtaeo9z19fwGwkCEMB1lEeY8CY5rRr5T10saSqEHI3TSn
371e+kFCXYiFc9/CfX0BIQh+NfcBB16CuvJLE7lRD65ShV5P7J8e9ICv1Lk3M9q8n1QpZg6vQpYh
AgexX2y02uOS8xuWFyxuqzY0Ra/dFOWJ9DfjXHOFrTz1HYBEOjuAfmShhuL1/RHM7e2ULwMUc5jt
Ql5T/8fyMoIO3LJX1WInZtq3bXBNozBqa5KOeNAye1wX8/6yEESd6m2COI3D2zQSBSsg9xhCJETx
yzeAH8dDRgnHyzoPcZRlVYrqI5QoJsidh7QSBEkJguW+PVDooO0wDC2309G3imdSkjYDNu8UpMgo
IAprj03YtC/vl5DJomxele65Sz3FcSHoR8qTC8ifLg/i5s4V3e/3FhYUj1isjpNPwRSr1Nhwit6F
xBE8Fqg2OQRJJjIhf7KgSHOpyFef8IW4kp1d06++YrXsf1iXF+urpGhkg45nlknQx0fSS2D0RQUZ
1V2ZXYuQk12RLR/5YwV8//rrv0lqd247yYDtLqqi4gXAcu/DDHlJYhoIs3KIRXfyxx6mR3U/iPYJ
/wwrYJWOwqcfWkQ+qYhCHUOq/gbvxwpLLKDMYn21qyLBPmftttQkXweHOeYO6zYghTVKXxlFEh5u
gfQRO4OfW9GoQK3F+XOjuJ7JXU8giA4YtYS+4FqSW/bRW5m7nWx+lyEBsfTmVKO1FpkxoDl1jkwN
/zV5U+pY0ffPWJygaJkN2rGYSdhx55OCtT4Xa+0DDVXvPDTNQgsHe7Qtz6FEac9dg+FP8OsH215d
/Qz64Jua2cxFeIZhEzlcniMhgf85cOtexJyJxEsW5H6mfc7qknjVj641q2QsGnIgE0VfXSo3PClQ
ZcDLC7zFyuBQ6oD3niVscHwa+A3FUUJQS78weV6PBPk0DPnIScnkdJzWeBNmIBuU9mbCqsRa4uiU
q8wQIQlsOkK5agGFfgd59PNvPr3se52ueoIBBdUHIWPNjTBWMoo+qVsaI+kx7snZIgxzh8pX29B8
hwaPvgVzMzLwWWd6Orzs7T6FsbAfox+cCpw+zQos4hCDxI3c2g+a0lPuoGryfZZt2hjBdALXThDx
0iE2mSS2l8CccbobOKbO1CMTfgoe8oyXst+Z6g3JEzJ34JFWPWlSHWzEaRfersXu/5s/Yx6YvdTW
53++optthRVbfpJCz/77wV8zCTqKT7/qZ9hsmPB0IbNUhKfbv0VWWQkgCTP3bt01sDMC7OEsASjQ
I3cijy/+fczWG7pHi68bIU42VFHu+yhx+NjEuraZl4tPYQlIqWC6T+vF5b2W0r6iaHjrr7CRNym0
ITu4xCDnjt/PEK++pnL8oSmMxTdbHVIRylRhzF+ml6j51nUqOWWrDc8JqZbLSyK8fCH5ejFVdubV
vtlnjLuFwMiHh2qN7u+fpzYgqlAqQTAfU+ZX1FoB7RrI6ZLSDynVszQUtSl+tkNZ9lCdkeiVHruf
xpgBnk4dGRVEyX6I/1HwJQ6Xt+1Bf9FxrCbxZAndVjUV0KXFsThrMEGF1L3VnfgEMI9wVs2wok9B
GJrG9kwSDgu741lOIenuiLckNckBT4vEhEujNn1KRVCBCQiZ61Y/yDk5UFj0OHa1MIevmmz6TQPQ
swbXIWFjhLqFyLegVwUNJ+fPKbzW7en3/0/df0w8PwUP3AKvCbEZLriIQ5Tc990Zqr9ccF5nyj0Z
/g3ESAw7rXLhbj1SjqHtrBoqym/oxkE40vmQSnUJsbYN0mZakopIAPmDCivOUDSRwwVmZDYh2kXI
NLjjIAvBuZf1DPcifmsao6MULDJS/VhR4POBNtZ2CWNYJxmXVphgkuAj2af1O9scXSqj/q/3cBhH
dVvXQkHas36ZushYUfGKGD3waZWLvY/g7hbbqEnWw3p02o9CxAumAvjVHUFNoUH/nDpn/qQ6AiPd
goCR9ntaM4CUq3hi0XJ5UfB+b7OjJDYzR814gcycOpt5idvjYB5dn/j+EmSyeAQ+jPDAtA0ZXXNN
LuBl4qxTMOUN8uhOfYPsorLUcbQEmQRTw4J4YW66wllFXaPMG3lMHU1QHdz/JRpsGwAdnjbbCRQn
C8iIDxQvhG7zywnuFSufrRx930PJQotqLHAx/fiiOozCg1BBn7BxPBIVBbkGt2dKgSiDSDc7or4p
jVc2ES020t4+dKzb5TjR7bw9XHwFccxrfui2zU9K4ZtGtScx1bwqUNwt7jS7Jyc7AcZE+VCfjWgX
6P0qXbqIUBy81qo637QX1jiUVG5hxd5tcV/jthnUG3eLyccbbfncgMRNH6V4IsjnTIYGAAorouO5
aX2MVJnsoV+XI9GNu67gAT2qZqlyx6VDJmDTR6PYycuKuHEFA5y5ipU3F3IotQKt8KK4OWbLwPwG
t6WWtwjQDiAS3SJ+PKljZQMZI7DikG7On2yCZ5hRwozvFR40H8sTcc0RGawHLD1c+5zjSywtjZqu
qquuqM1Wo+Ws5IaLW4i01wrJHWNap/GZBaPTI/c4EtHYuxC+mqgwk1ILCii8rIlR7YraM7Q+FCxG
wXAJef+Xqb2kX/vJ6weEdzKkB5vtd9RX6SjD/esy5gOa5ZxiWJmmsVdo4sDeYl716Oco20L+XkSi
KBstExYysfrkk2QtVbVVZI+KXEdYwxYFGmebXN3w1e/iL37qet/VK8yUboKyH+IX/0qAqFWf4ky7
5NFIxqpTXJA2X+cNphZv0mh69r82Roz/q1i77/R6uvJdQFLeIGZiAfkmCwglRC52+MZZpgcOpJeL
rluCa74bjyqv4UiTwSKiueB0eX9IpIaKhOBB82MgzMwzVI/5USb8EAjCdJxOmuPjYPjfA0qjEXkJ
+9iZBjqp1R1PcLNP1p3q6J66WCIvGfiBIE7b3jUvOMFKFpGT3cpK++7upHUdQ2yqbd/PjU4gYOFF
6twqmtS55LJa1jJ08Z0xCnuDzmtu44m+f2+7QMh3h/AR3NvK85JgNE/PlwWtO/0sjvVhcarCR2Jf
BrB5r9Z8RBgTq6vUXdRzSbl6Qjjsb+zw3bGTWIw0Erf8LiC+NPq0SIcm5RbRqJ6ZB850Otuhf6UY
VoCoah/p1Au9wtn3SuuWru6MtQvMcmlVVKaBMnofZKdvTXSfwBBGPYn2FICFk/+5gngf4fppPNGm
+h/+O1BTNxGZzmhgTljSyn1COG6Cn2bZBXdYXaJytpFAY4Sp5ezRqeKQz4sG+AP4G1uJp4SpRK6s
q/JqwfBsKRyReRaTjOoJpGuwGlHLdzplLw3/ZCmPSxkYpC/UZ3jl1qfkQb8hH8WHxg4J2nZYxQxb
zYUW2xmeuzJrdGWp2joW1awCL3+UXgHnaYxIxl5SFgBjmpb/oqcrPOXecpUvtjV36I0udKRV7ypT
ZXSn8RBPmBMMpN1s7JcZN1aV6nzRTAFWFOa3KcNacf1LlT49iPdXWD1KLuO7gNavosS2aubdXlhz
HRKYQ8Af1DYpd0QTdcOJhsrpH87bWqrComWtm1kyzu6MPzUckrfFMowWAU9R/DY7DnuPMUwZFAnI
l/S7uCLFuq8e/N0fxeru4zXwYF5Uw+s8xHSlIHthu7/27kUTQxg7wpE2Ta8L2/BfroUR0SA/RINO
QF/MqOSD6R/5zFI3GVpHYp8UGg6Gvrb5EmoWdbuNvjLlp1o6G/osSr0S/kKR984H2U5wjBYSWCjA
nYHaFuORfWo6mo0qovexC4w68Q+ZHTauuFg8dMJTRr4A7gAXjz92ZH9Q4rw8L3KpkSWUfa/eEkv4
ydWD40LnhAzSKRmL9ZtgvXwnFJivTdjYAGyVvBWPbz50fzk+mVLdUvsOdgz/bihf8sOXanF7qXaG
TVIpGVABxN8dlZ6HKvIl4RKFaf9aDNgzs4je2WsFRj8phC1ANEngoWzaQTj8gk9snpkeYFTqx3Ml
B56nxBpjy/fOFzaAST462MgpIk2Fu6eu9IFjJbxn+kAhPUYPinsC51ZK6LwGvJbX5vQRnasqsBj3
JoRaIr+Zx+NoqUpREeRjFJoIkx4DvcOxW6RV8hwO5xuPSQJsvmaIcwx477E9W/mFykGWlPYZ/SYe
irHshXgx1ekakUM8eWlQ6v15hOir1XfXaFkJ/Xbs3JjDh3/TOIUFS8o4Tjoj7PUE9Skzx1gqab4G
DBiLf6AJAyzgBPeOWFQU3UjyxmHRdlwUOm5yhsAQUzn0FYVyAdGkaYam0JivQd5CE60qEsTSqfCI
7cgyrf554CDWH/2pR7Jm1O/HCgWJx90CE5AhRXiR5/FiLJN0k6IxpllSuRDK4GThge0CXyeKO1PJ
X0SErpnydArk95goWzyEiWkcujbbwkvkNHKPiQYUKHvFCxI07gvDg22/T8HFjFGDFn0TKaBULXGO
uncn9gHyoCuD/WPg7qy7HGmdBOeiaZnusYSqQ7enzVu3zar/zQiyqqK6Q+q7JUqG3VjSFAia0W95
thAVIWaXhzYqK+qY5ZmuO2Q4luynjv0DiuFiyLmjDs7VJsS6EvnZsxb9qcGWHrj1rwutG7hee9ON
iPsTb4AmX2jvqU186zvMUojI0DRMbu9wCpV91Jo4NoZydoONq+12aTd8ijhMHbye7Quw/IHJL6ri
28zra1CJh6m9cNduLHzdThjYZCLABnjDQgDcqhHxU+2+Uofwi1UINfwffamjw61EUYb83dbdrQcU
vJrCOFipxGEDVzuFh+awr7pE87bOKlYEouctHnU3mXNSsr2HhBfYMK7c1GrCtIXCLoNd8WpkjUBb
EEL+qN/XA7JDIkXPQyGdZso0800o7BGgEq5lBuH4Jue5gmsns9luXApdflkspCPePQK43nUz6ism
ouDR8I54IKB0FlVi6bnfzCTHpS/q/iAvtHIPvARUDXKFfaJZrazmiiF1a+V1O5fqGqC7qt9sklDv
3M7LMkv/9mxACfcx7sAgDgu72eWpIv09ncb+JjOddmEugUV+JKD5MsxmW5JyLXjoI9DwX7casXnT
6nadvhXtR9mNtrywF0F6faW2rnQTtGyXgxffwOGpF4uaawiAkEG6fxT6U+Uf8K9GAQKhp0ovSOnh
9yF5QChUTo+1pUbFjriT5rUjUDliwHN0TrK4vn43mQXY+E8Fw4l6DWrw4XFjnvYXoIp72YfUkidw
piiNnLMZbeXLtFufnuQKdV8iIP+LKx6wMFvI6w+qXcVTAbqrb/Hmc9GK8LNQHBTJUBuh8t/uTtDk
PeZq4qLF/rMq0jBGnuP5kH290agQZQ6mnLGvduzwsQ9pJzfRi4+NNVQKuzsEZ1U90ZYjjRMzDYaX
KG25x3ELO1h+RDqYWxi6hK9qTyiFB3UEjs0S8P89D8PxMXOlBqUwjmQTIWH1p1E31ZvUb2Zngbos
HDyE4uCJciTtDBkN+v3QrDr0Tjva3tD3mxw7q178aa/gV3PyMiK1ZuDAi8oVtJ49AEEoYMrLjJkS
k8SRp8r4iJonvK9MKWLVeJB79gs5ZcNKfM/9RCGTCmcfHI14Lvl6PtOQAnC0bnWcrefUHUetK0e2
+NmJad+ojKjuQZJGz8kIYvMdkafdRSBN6iQzqmIkSQqRFx21KyXPBiPTnBwxlRpxs5ugNz8iYke/
ZtbTDppKnX73O61Hb1LFcycW8vD8P/nVwYPotB1ofROWrRQt4WwYfiT5wPWCEqNn7C6hNOHNk0Dy
ENAI3vWQrab4Hx33fskEgkS+aXLkabW5LMfY8AqgvoCn9tLFvowbfTsy2cZF9QvSW1daKFQ5BSL8
uPCtEdbWPPy2DJi7wOrLGShojAUOFQKjdknBaGVqKAhxR++Nf6hRrSQrHP9DEIkUJS09OFcizQVW
hlNM3NrLqXUCc8rGB5CXtJVGzIpHO0m2Ra5L2/sMpoLHchzzqXRGQSigk6V7GwP55RC+HdPOWTEt
IBg6h4UOK1ekznweVOpXHA6kChXTGfoLuj5l3mQzThGvRf9IMJQiBpRgLWSgaQD4x7FFTCIH2ZXP
AFbGreDzygDcUIrZDoLde0AaUfAFTalteCJbkZD1q81G4ZnTeEZial1x2P+/pGnkhV1+alawhBLh
o2FPqIqtxYzcyQkhdZukorZnDE8aWuPXNUBFS7RAJ4WrWhNW2lsetkujvDFrHfg3uyn+erbv7DZA
yoe3KRumm9OSh0bnhMnv0NQA4+0EHEdNkfOwd3EjUIDj+/IbDR3BMPQFWtHUg797v/4lVPbOhaeu
9Bt3XltCOb/4cJOujWZX7uAGLUml9mRn5eTMn89ip7yGcYayNeEBLsosjtZg7KirQAotCdIq5aff
lPdWItRFUpKJpabjroIMCmS/NIuTFb1MX1xS+Ol7Y+S+DEvszFo1Ft5AGIiJnzAabQd+PeZXTlbC
MOfStrOm7WcGWCu0cRV2iQ9pF4IEgaV1fuIvaxO6h2A3+2sRK1TU7wY1k8fTc79/asqW83sU4pUE
tg7NdysYFe8zS940rXXgpUO4SFe7ltFpzJDGMEIxEWWW09Q3aaMZfG3DUsfoztGFeMW/EJrvhs+G
D8BO2YJa/p2fQySLy6wXeMcnl5pXehm1clO335Y2r6Bb3Z5vOCWDZDbuvUep9giL+C9UVqOx8WAh
L4FCyjW91jBFUkfrK5muffEHqMcxEUOFWWcSDSoN2gi1Iul7fMEG1fKBQOsd8s4fNe9Fs6DTvJMA
ariGvjP/S/K5QEhxLUjHXdmwyNkKWRoQow0zWRoBsDmD0VkXb8dPGFQYk+ZTA0QU1gsieGX1At3L
QoHp3bpgUUO4NnfwLlnUl9JoHtbcIEPP3Jyh/GtBE7maCYxDMYxOnMWUOWsqE0ehevytPs5wMLC7
G1ezJiDAj8f7NkaC3fzY+E5wzcCggDvSDjbydXoIqb3nS8L1yxjdsf7vF+kHck6mo1FF1LpiVQFb
HDrJTCFSqyjRvhA25Ejt2Hib1BuZn08fjOTywviv8iL28Cpo3tx2nRKqTdHrdZX8cko3IDwbG8VH
RZpre6hiv8Z9btpAPQ1bXKSoa0JzGzCfI2E69bMORk/Hex5p1YsjJz6VYfy0bKTMSRcifkbgyUFJ
AOvDAqXlKKwh6c/chSPvNqfoG4kwxlCpcJt7+H/4PJXbOLh8BGvwpK6GknHoMNjgXulcdynLBqgM
yXsmLg2bd/stgdcm8A/HvJrESg6MI/1HSxVQfMsdf4HIoBUYhid6xINoa7rEN6couO/b7Xk5kkMD
wXmzaFuYsEK9aLX478Ax5hxZGlfL6oWLo5eCSewp/CW3gg+UrqSKHjnqdTFelueVt7bOslweWH3x
gHA4JoYSORek2Huk+gxhbdQu3d9ZIxzORLBvf55+pfzLfwt4ouAtA2Cv+cnme4ZI2gAsnHuEaaOl
7zzKd1znmo0RS1qRZLwGCLXxoyLZcA6PMLNUZcwZU8mB6lwWsC9sbftErnG4WpOCyiQsfm03SaKj
zYKWaOIER0ItMjkNWnYChJKmQk7tjrrz8Ct/nuHUZHigQ39S65FYlcJrnRVziNnqS6Rrxazd7YOr
NSI9y2PGkq4IKp1XaK+n16PgNE3l7CTfIpdj7yJGxLAdnZxDXNcIH0Ze7P/Bi0k16dIYpDEdXKuk
i+Po1JNRYxTifUbF6qjv2Fsefq+1JbqxZYKwTzKhIQAeTx8bvW3OW/BhrEqC/P6N1DOgZ5hQFRON
C85n0kc+OjG+4DONyxc3mDUt72sAVncnAXTQSed3pSau6xPNQmzUVKxhg4aXG9iJZTBAuksvoHGb
RohQ4UTfhDDqh8n2aUVpgdPCrkSSUdYAPzKn2c+hYuPMg8UDhbI7nfU4e/gJviKd/ZntqkjDjYHE
mXVRyODn5XPeqBQJYMUamZTR0JCjKK5z6Rgju3zXDz5SloIxxBlibatHem0pO1RU+17Dp7KP1vbk
DNzUNQtbj+jGYUa9QdoakxpGLaMGTIR10iugbSX6X/YFQQHIOIv/yYCSoD0PRvQGCANBHD1dmJs+
d9ujmufwR7SVaNUlAmS6SOr2t9P/Enw6bKrC2C7o84h6Ak2+tLiZqYrOEspvNwbMb9XaMe/y0yOt
Zr/97Kz7+4rdqocc5FH7iM4jtNsy03f5Ip9V6j+Lt5inDVuLtWqbpEN0etdkvaAEhw2m0lwSSN5T
qTQAEuJv6q8AbUKUBJ31XXszJofitHkYY2MUutP8ltz5zF/4bnsRhc9rOZx2rOim7A287OWB5/20
X/tvmRSJbPKqECIAxSoOmPii+H+EI9v7WW0oMw2VnQHk+kU8oXbgDyDQLXudCBwoY5xuvWaNW2d9
ZXtVKN/TUFFj83RNRytVtpyaAajnP0yD6SZyeuLshfbIwgjNFEEfwYEcmkuYshMVwXkLEaTkcx6D
RZky61MeTx8E2NR0Rf1nueKgLbqG7vhURvk5ut9laW5JWHeO35ush1YkVTRLD1JQuRUJt0U0SBx6
1N2Eg4CJCjaAkTW15Uxi9FdkZuV0OOYRwce5hLLhObvDgdwSx3nGPARiYBEYRWZHn7blfcCaC+zA
x59mOPdj83nQvQgMCieOs8i1cR4Y9PkBGv2/cuRKKoMUQlkICTd51NBmpK9f2Vcc3rr/SYa7FLMe
OgvpIHYqkpWqvF4O+Q8c82ppiKPp2DcgwVPNfs3gDDLEm1/1i2AwNtuew6B2ZO6SN229e0s5TNox
XluU8gnu7XrOhwUlYO6RvTZllscXRn5lgiBNLyYXkjffuLYhKxigS7zWOOPq6xpERfRJwMjjak6N
xQL3RrGS0gT509TOzZ7GGiOW14YYmLx1BXqQw9LRQQdpTIniSndDLSpLR2otaDqJ9WHoGxazKUE6
uPYgahqj34rAt545LcEsAo3NFSYx5ZFVd481FiWE9YY6xjYcQuVlflaUnNSOMvc0UMESWgpWsV/h
euDOWdHkfAYsog+LQuqTBJCVsQxPfAi0VluHyKAzXv6z+Rgq30YFWE1sRxay4xQwPl1wZ8UX9lmY
bh0cWzOiCxBk5KwQbexLhPLP508N/fxF9kO7Z8GPkOv5r0R4y1/B98HvFSZ26P6g03Wp5XmPcKlp
tZYPvZkXPyfDSqJaEvCh25CcdfefUPz3AFB4lnzUfomdKXz49nMQ5BDogMTu95EmPeULQPjZJopV
/tk3qe8Llv9HQNIxiDAQtjPiA3aTFaHZ4BBZGd+5Xe5HGy+sigIq3fYFjBRb6KTvWIDdlhLT3ZpS
pBXJWG1787buE653m7B+Qkd+IwYJCFW/58mn2+wwCHAvD0Xh7sdlSN/fcMqPZIm4bbevcDA+iCcP
HK69Eg6pjnU+cstHR+N0Wah09URHPXgygma/fYWDUdHWKbKIiukKgYQZLG96RVQU/lPRg9RLy2ZG
psCfSSmE2X722yZv88HloWYziIzODR7Br3q5Z5kXaf7vZaTrx5BhdBG2/9TKTLybexhfBPciSzGe
//XyWADaPYQ3Ct1dM90OXck5AmKz1/xaIdUbVXgpUVDW0Gi+d0scMY9RkKly39EomAh8LyAHaNvg
aDXkMbPQeodTcozbUM/RqzEzthuxw0gohb3hXtqS5a54ABDxJF78mYibXnrDYIgHpkmmBn4b255d
YadwOUB3htDTf6pQ8SEIRcpB6fVs1vwyTO95idEBgYeyQBIegpFxkZYCO46gCI+vkZiE16taOLNd
Q5txbOzQuIENX+y92QDfso2OG017NF+mqwKQipgzxC+vaNjYRrPZavXrJ0G0qfjaqhbbvpU544UR
4rwm5dKRLMWtBMRqTIIpvyiVsRKRLTQ+4ilG0xi4QK3VnTYRTrfdXnlyXX2Uk9PFCQfLMj5VdBXR
XyE6Su+TPW7a2LzjC02I+pEB+qg44DXazbR0VGfUe84SMG5KMQrZElJBxu9A01C5hHr+wjbdsIk4
J8MB8Y93AlmZ5umUdfSmzTXaFh4jSKx9U+JiYGR6aLGUVQAb7wxU7IbsgTZiSx/hM44JijodtW9a
LDWmj4eEby/7buYDVizYYhSY63wJI3IQ0+nkp2LdTMoV026pslU5JCpAVnVsqmVPF98vZb7++pQy
C9xly5TgT25YV1jlQUwRyVJDbEvqGrYRz0dsDyfRK3Bgjc5rxOr3KvL6aZjmd63ZF2u5sflStb2m
D0BUapT5Et6dg0hm7odbn8TC6UhTUPHQ1FXUHF5qc0y011jZYK0TF0sFm/MaOJ7347oDaOimGWOT
AxkSF1Xuc947QRecV12mYMGSbc2UuqvOFgm8SkSWOiDllVf/RQ8Hp8SMKUzfW+BXiKUbIjOVrdRQ
0ey9KVoTTFG/Q681eQ0ukQbG4t2TKVo7jDHmeCYmvDGLIu5lSDyVpakjH7w4DWwksEovYknRCTU6
OiZP1DIMJzCFl7L7m7PnikmM3ZqcrLm0v7yA/SGohshnKUzPHxyKkMABpiwLtMoP5gLD+mm6KgOR
OJT0/ElrJnQkJEw6GGrbT8Ff4VTV5hlZfLWBFFSDSSgfSpbKpByRCFpBHJLBqbf7jZPuXYIWfCb3
eyI69MkITawenicWyh17jaMFTH1cuqeHXiX2ibamBhOj3BqUGWIY9gVTqExp338wkCHIB9tt0byE
edQ/67dsglEXBS8f5hpeDX4Zm/k7w1GTW6dCrlKp4FiiudVOtaWcinMYfNoYE9zrnXJFu/EVrmbV
EdscN8oASwqSpLMXr3ALN2Oh6pMG3ff1scfp4EyRMM4B70it5lYhnpH9UK0tRAjuyQ+2tehkLMF3
3d5kLUOeO70Q42X5/ML2gP0g0SQ4wOQX/m/SZd5eSCazI6CweaPzvQkJjkRlXWiW9u0OLUelTwb1
P2ZDSeYvkmgvSpFpdQGtP7mcl+SV6wYCGo/hAzHZTQ+//RdDmdzhfznvvOglA7/0xJxyYfbu4GDk
OCn7hZpx9YgaB155vzNjMZFGXmQQKF0eqiWXYgM3sB96kM7V9WvPqVZPpDMw+Vxl2TXz29bSd+uG
Vty8kso9bCRu6jBx2p3+QvzAYwI6C31PLHmRH5F1NUVixOgRzVpeaneh7FKUGu6Hq7wiMRfAXq3S
/njND2hXI69MG7OMd9NZ8XypZ9HtcZSM8xnP86bprws6v65jDiERJt40STpES/56Io4dT2BIUkXS
0wO2rGObqAmZK3GXwvE9II4/5tKRMhHEXqMIoJ6aoPUUF5BdWe83+K7ZMrygva5jcJD+cBDqvFK5
IFnZrBWErGTrBWdJSwYYI/mlFncILf7rPRjrz0EZNaEIaQREPsZUYjlEiM0Pw5vWjEomBMmeZaGd
khvOWXQaibexJRjtWjgMN85kobIU/7rqmdTE1S1TLsi68BNc7PqH4ypzjjBEKFM=
`protect end_protected
