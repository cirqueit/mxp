XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i"*'�[*���Xn�Z>;�V������\���L��(O~� �ڜ�Ց�0n�U#a�9��%�~*�r`���q�Q��
�����o��Z�E0uZ��)��;-P�e�l���G�-�QX��B���=sf%~���e��:o	^�sg�Ψ4��0��7e���C:��y��?�a�^2g��`����,�@��zH1�[��+���t�ׁj4oe��ǒ�	��P��~e�a�6%��np�J�߉-�T5w��"h�H�QQr���4:B�5׮Ē�U�2�����z��V��n_��
}��`,7�h[9Ek�T�1й"Y���i��K�B=l�ؓN,�=���DKW*>	ǎ�X]�#�o����-�>d��F��t�>�����Bᯀ$���/�X�~�n�����.o�r�-M�|w��Z�[+�lrb��~��10Ȣ��7O��W�z+�ߢ�%�m�`\Й#��U� Wof#�o�yc��Os�����˄©��wc���'q��Jn ˑ΍v6ل~�X.1�/d�/=k�6�;���+��Mz��ojn��b6���9��t��[�i��m�� .h�҉m�����O�$:��N���B�-8z�	Y��5vMYI�%=n z�y���-�@0z�y�r̚aZ�GO
�X'{J�v��^n���n��kƭ\��}/�5Y��%����"�D����[�`8�c�V��i)��\�#���힕���yn���<$�+o�X.��GU-
4�~���d��q�o�� �K�NXlxVHYEB     400     1d0�[�2��8���D������;�M�@f�w�PH]��^iT��䗓M`��T��p}+�:o������ݔڝ��ˇ�JL<GS6QQ)�@\-�R���i~{V((�\ԃ*�����f�'{
e�D|�M���\�w�6�[|,�F��P��;��כ�7I�o���3��0�|�<l$��4I��q�Q5:�S�?��goa_fM͘a�9dV���55 ��d��)�8�{��'�n�u��m"�"�L�lX�3�K����ό�(�?)���*�����1x��E{U����u1�ؑ�
�

��;Az��ZB.8�}�l�탇��Q���B��r0-�3�����c-]�}�R�8����)=%w`����h�C�
^t��[�c��i��`�x�-2���t�Jq�
Nja��xGa��������1J}�},F���Ԧ����"���9]1������v���ՖMw��XlxVHYEB     400     110��䳞 6�KJK��fz+����јFU�UA�>��/M��b����]�)� ��`�wF���`�,��e�X�M�L�F��=�G��v4�v�a�ۥ�զe�-A���~�Y<�Z�e�N"�����^�O�UYb�[a,5�靷,���Y�k�^���L����<l��R�����:�֞�ζ٨8 ��kw���/U�ṋǰ����������u��&rΫF��}��m�j����mGY�$b�T�� )�KnUd��>S�}�[eU!�I�c��$:�XlxVHYEB     400      f0�)��ŋ�o�k���>�g��Ւx��1Ȭs��%�YFG���q���-�{�:�����\��h����n1�|H��'S.i�6�**�R�y����ZRz�-��%����4�G+�R�z���"�,
uڔ��悘l���.��*���x�Z*W(K�/�,�r���&5�����N<9���[D��}u���ߗi�
��$�5:�U4�L�J��Ha���}GF�IɤO���%�����{:�XlxVHYEB     400      b0���X���pKco�Of���8��'�e�jn�;(�lb���� ���{�r�\�ߧ�o����dO��@����]�j���	#_᩟ҟ����iSuŕYz��4ف"�Zeç*མ�f�4�|C�.9	<�K�+��;dYJRC�[.�����#�x�5��f��ag���ez����XlxVHYEB     400      d0G`+D4�zH��#z��0�����a^�t�o��ٷ?fO�hb b�SJ�ʑe���M{]�S@���]p_$B%Ki1�t:%�Y	�v�$K¶{bO���϶��<O���7]JM���C��φT�LI�JJ�qX�,J=[|�.�)��le͋��d�%LH�*0��8�D���o�����(��/�kq���F���cR���"=��3XlxVHYEB     400      d0;.ŵ��Q,a^KbXPN�:m��K5:m�zL��"�F�m��X�b����wyBW�G����K!|!f���:�$|S6L�\�n|�D�45h�"�y�l8���'d��OVG$^1��X�G݀U�ݻ5�{@Km�qI�x�ÁQ:�6b��>	yZ�G�Ab�5��<����ϴM�"ׇ�{
�1� ��z'dr�o��O�XlxVHYEB     400     120��T~�=�je::��A��G�0 |��f��@�'�F!oFE<]u�ֻ�y�G1��@8��'�T�SM����'v�T��k��-eZ�;�QyU��;�� ��_5P��T�h�^��s�%2�+�k���M�r�Scm����֟-��d-�+`��l=|[Z�5�7��s�F�+cik���᝙�E���BtK���5JsGHB�sA
��\	0��3�7�+r/�۽Q(|6ቓڡ��l�(���Z�-�1`[��{#�ʭ�P�Ud������'1i�=��c�A���A�R�XlxVHYEB     400      b00Ɗ�h�t3�iVxnio����
��09ޘʤਥ!�{k�M�$�_���,a�4Mh�������ry���]���Y`����¯7�N�@A���BL3Oi��L��,��������j����5�w�hK��O��d!�������cj٭7A��M-��?�1�K�z&��XlxVHYEB     400      a0{�f�)+{�*f�b*2H�H�\?�������|d�yZa*yڋ����>�	�gF�\*�&�.&�u�)޶��aD�Xq����|�F�P9�TF%��_�w�A����#r�.�~K��#Eb��#5����%�?{ M�*�䭘%�����6����H�>XlxVHYEB     400      d0k��+ݍ�,�<�9N�:�Ђ���^N�E4�gI5:�6��_�&,+�-�o���mM�?~!W�4:Q�ƥ�b�G�<5�/<��ը�L��u)�\�8�3?��ev5��)@~�Ո��%5.P��37% �gY�ts�sfȭjM��e�f���G&]_qM��B��#�V�U��=�il��GQb�C�1%�Et�/����f�6-z(�;XlxVHYEB     400     180DX
�a��b8����i��W�O���~ǽf�2F���-��J����~sg6��H���^>�t�'���}ݹ8z]�>OM?� ��ͧ��ypb��< ��]�H��F��ŵ��<�x�c�%&��N\;;]qH>H U R�3�6_�<m&}�u��+�V�,��wo�ܔ��u�
�T��x�#�5�t%N[�g��$|u
.���\)�Y���m�l�+N^3�U��C�s�ܛ\j�C�`��@���<��+ӥE��L_;��WLm�8���\�"瀒��uQ��OG�e�s]#����D6!')��\���m�+o�X��{y1cU����ճ��F���2G;���W&�v	��N�������D�X�*f]��DV#�=�XlxVHYEB     400     130��3����D��X�v����_����7�^���Ŧ7<I���b�CZ-3�a�\?����.s�<�rj�_/F�F:��'x��%��N|����>:sJ�@�Ǆߟ�o���A7�Q�x����υz +�ϦH��>ܐ�H9���۟H�'��Қ-t;l	�ҧ�'-A�9 36=�1�|��`�`xf��3�}���y4���dƁА{�$�M<lHT����HU�NO7�`E�I���oQϓs�v�cΩ	��~�0���҃Ӑ >VC�!z���(���F�2o���&z�!��!����XlxVHYEB     400     110��<�rY��F�9q.�W~ޠh�,��Gx�kI����D�u��O��s��/9������Ϗ7;��m,A2��ϗY����� �QG��TOah��� &��8��!(Y���H��x��v@Cf�^�.�}ؾ��2��oC�Y����1�Q>9��f|��B#�8���d���Ǖ�s�l.�0G����V��{רH{��~�(��=d�X�	�� �*`7��ť,���`��4Y�^�@]��(�H1�qç���)̳�ͩ~��u��ijXlxVHYEB     400     190@O⩪�p�1hv��g����ٜP��9��X�}��X�.�u:W��{�sG���X\�}n�9�!X������)<���;����u�]�N�S�B&���k$3V��=m�l��{���T�&��w�B 4Ԣ'�-��o����M�)�S�X��rɊO�c(�%�?��֚D>�VP�ʄt�Q���n��X4է���EuFz�Ԯ�ѳU��e���J�dMC�����1�+W���s+��Q�o3�KI��u�m�ׁ��TN�jƈ�:�S˅��o�ɀX�xPȪ�1s*�fBU��/@&_���z�ю��'�[��9N�Ǡ��S9g�?j��R�5}����3��6��~�E�������	�~-�kiY4�_Xg���	B
G���<�x�Ȥ9\XlxVHYEB     400     110�\�P��U��;A.x%̭k��>�!���ר|X˥�@���*���?3(��	 ߷�_��1	�X�k/���G������0#7��F�T�wh�)�7n �����\.��Ȓa%�����w(�th#A���Q��y	E�k�n��,��[����Y�4]Б�l(v��E�S��]���I�$ͽ�T��Ts�p��˼���8�?,ms��b�{C�/IW~���&�኶%S9Oxy��0Cj��Q�����P9Uir+l���uF�?�XlxVHYEB     400     110�@G���`���u�C�ݿ��Ӌ�M7+�Yu0K�G�Z��M���9��TM��\5��ƣ���4*դ���e���WV� G�%s�vKA���O>���4T��4����)��ʾI��cE��	�'w9��"^j�1�:|�]�&_��v3��{�)Ţg���ܧ�=�;y<��&���K��ǜV�����A�'	���uV��i/�n_Ӆ�[A�į���i3�M�s��l���I~q�$�"��zt���Ō����!�@4%���h=�[��'�Og�XlxVHYEB     400     110���A�
��zx)��5kg��n� ��ż�m�y���}�� ��������:��O6��uYR�������b�^H�
,�ᓥ#(�
�R\����'t$�7t�z���|Z"�����q�=KGD�	�� �'#�_\�=�o���3*�4�d��Kf`P�·�^�CfifӇe0П4`ݦԂ��%Ld����ڌ�@�&=B,5w��~�����/�[T�-����Ou��w�Em,hi6y�B�٩Q_�|Hs C^� @�N����V��IXlxVHYEB     400     100�s�Mδv��G����S/.�,��U�2���B�5���YXDb�т4��� �M���sf�w7F���dZ�Ŀc��f��m/����5��l�r��6��}����6���"w���/��4S74�j5�$�}�3ǮL�?���\5LF'o�B4Pr%�.��mLN�h����ƅ�%+�I��Rd/\����As1�l�����U���&}�x<�F^��N�!e�P�T����,S��{�&�?!q&5�.J1�Y�Ƽ��.XlxVHYEB     400      d0�0|6��빵5pCHW8J��w�@��a��2��:���?
x�Y��vQ�=t)I��t�ɉ�DҌ�A3��|M�j�����ivǤ}�����	�;<�Í�~'ITe����?>���@ڤR��܄�v<���W��)���Y����s�/��2�g5����ߡ��F�g6��j>\ˡНӯZ^��Q�Z���>�#�;�Ƴ��aXlxVHYEB     400      d0U��ȉj42'9�����"I�~xo*9�u��3M���B�\W��_k� n&�BHR&g7��z/W�\1+�.��a�r00?�
���y���:��@1�d�9�cT.+�4���ﻶ��(����b6�.���*�����0�3�����] I~��&�᜾9�rql�g�[�$}�4��E2�����On��E�o��"]��v2h|��D�-Og�.{XlxVHYEB     400      f0��,N�D�w�P\�0y��� 'ѭiФ�V}L��� B��@��KM�^�9�?�*��c�%M�2~����.��K��ms�:ee��4�u�S*&�!|�J�hgC����'��1� %r��� c�H�K���a{f 
j���I��������Ѩ�Ń\Vٸ��G�k��x�{
��sfd}_A�[M�
��?�C<���6�>q[�����;x��C�%�?ڊ�o��Y��XlxVHYEB     400     160M�֕���,�q'k�L��n��������֜!���.v~�ٿ>b`�Š�l�;�f ��"X�Rڋ*�]���Kz�Da�R��^?@s_��F�݂�Y���xb%+RP�*Xn�!Ju�`�Zi���].�$���P{Nς$�rԜ]��]wǔ{h���'�8��{m^��b�)�X2���t���:Аp�bPbr�������Z�o���Ĺ��U��5R��.pQ��o���1t��<P{�Yg���Eތ��� ��C�1B�"D��X��|���^#x��W'�d��ˣ�̌�1�6ӏꁧ��}Vh��ή?�<��PL&�E���So���}*�w���U��l]��1QBXlxVHYEB     400     1504�0Ym�"	Ɏ@F�U��Rl]��c����_ W�f��3~�0/]��)[��Q#z���)���8bڳ�Q�5)�-+A �z{{ɢ'_�S�2�q˒��ǃN��ɮR�ޑ��>㈁�t��:��������5���|^��\&�MdB��|a��r?k�E]�(��	߀���2�y(�ͪq�N��<z�98����l�ݍ��B�ދ�Bp����;���ܡ{�˲�5=�Z�b��j/RZfQ�#{V����}�X}��Q�a������d���������AY���\�ZFzA,,�B4��!��'T��d����fD\I�`\Dm7F�XlxVHYEB     400     100e���FJk�!r"=+�������il�4��!�P(���`ʇ�	�w<�tOa�PXGw4��D\@NS ��چ���������j�@t�Q��r���a����x1��[	]T��+k�{e�yg�n=�q�Z"�$�?Y���i[�~�Ш�b,�t� ��e�<\0�ak�ԧ3�p}"<�tOn]e����wOV�-�#��p����n���+16�\�s�|���i�DAj���"�I�7L:��N͎��XlxVHYEB     400     140�S�Ģ�C�]����:*�����7X�ǩ������Ŵ�a7a���z$��ſ�����Tu|�" �)lW�"i�rjk.�4
D�M�!'i)�a�7����K��E�a��\��HS�''�9rprk#����	��7�����hW��aZӢ'IL�=��̝Ո�goF���y����*�{@4�݋*���z�6��0њ�j��o��G.mCU�����e^�h!"��� 1��(zX�̺1�C���;!8��ufFOI�y$^�,�|F��b>Lޜ�ԃ[%MڐyZ���r��M���{���M���'_2���1���_�S5[WXlxVHYEB     400     140�o��ς�.�;�b�a��-1#�́�"�rִTV�) �c��0-�)�QrB��q6�����������+�d���V��	�+��
�/B熶��ށ��-!co�|aN���A~�/R�y�yG"ԇ~_���������3p� �s�4��N<��1�D�2W�i�Ǫ���/4�q�O'������z��S-� ����u���qK��
�Ӂ8�vS^����Z��8kЉ����arN'���>'/�|�# 8�[ٮX���f����\K�E�5�#�=
n��:B<���M�.�.�<�\d\T������XlxVHYEB     400     130����]��3J��Pdq��/�7y ����'ԕ�fBז�|��|�Î*lFx!
�Vn�H�2��d�4���U�������B���b��T���)!s��%��c�M��ҽ��nm`6���{�������2�^ކ���A���7�ip_B!|J���1�x~@Q�\�� n������0Y��/���+@t�"�2�����K���_]R�(#{dpȋ�rv�+��
�poʬM4��L�I;���I�Z��X�G�Pr~ez?�D�&c��kk��tX�_�%���8.��f�I^��XlxVHYEB     400     120{^�^�֋�^���d����=�w����Dv�C�� h���Rt��ٶ��u[�� �������#;t�ˈp�[v2�{�k�"w;��$��5�r�2W4�C�k���?��'lO+�u��_�����+���W��N�k+P���.��?��ˮD{���y��WaݚG/Eä�/hN��_�M���?��W���~�Q���u�����?|/"o��m�k�߿�`�W�fF��!ҾO�m�4���G�N��F+X��F��ނ*~[zKe���f��XlxVHYEB     400      c0|��z˹^m�!�G���6�#��Ӫ��{y��κ�0�z�R����\��Z��X��0Ym��ΊK�����#X�鴑4#����/�4�en��Z��ag�8J>P�D��}����6Oj��9���0�P-~�������V�_6�;$����H�,@U�۠B����S���z�2F�z�[�{�k�r��XlxVHYEB     400     120���n�&L��gܳ(��>]���l��Q�1,��eM0p�tF-����hg��I�h���C�N$��\n�MpM����D e��}ԟ�9�d)�αϾ�8�&t�#K���?׺n�q�M׊p��8s�A�K�p;릈O��p��$d6H���E���IJ�hxGͼ%��U����:%�-�I��y	7�v[]�v|I6Ք���|�ޮ
G���@����=���I����!�Cʁ�_`e�5z㢁u#�'/JUzNJ"p���N^�;�P��$��ī��,� �П��XlxVHYEB     400     120Ȭ?�'_��?jij{��lN𕗡�����m�����u-_�F�W���~�_CU��{u�A1�+���H�5�e��-+P᪯�Jt�:����ǡu����/4��d�y�&Tќ

Z,�0$���u畘 0�輴�w�W�p`cFQdO�K������`6��&8�����,�`>+2	�>솰7T��xMӲ��`�Ý@�<q��Xh,�+#O0t_��$g�X����:!����u����@5<�>-!���g5_jo���خM�B�XlxVHYEB     400      c0Dv$�;���F�+�(v��ð�Y�#B�)�b�De0Sa��l�V�zM̞)�d����\J�7���^4�jy�&��4 $�W�zMM
�l�	�+Q��pm���x��9x'Z_+�ڥȘ1����+Y�"B����������,Z�GI��ۮ~�U��a!��\#�c�9&�C��}@�`&�P�XlxVHYEB     400     120m�ُT��S�c�>#�ɑ�D"U � Ho`X( ��(u�`�h.�+|z��v^�SA#������tВ`ߛb[,Z�XY6K�.O���.�z�$�nn릙��}/���V��|��@Ɛ��}\�:���V�<E`n��%Ä?gQՅ�S!���� �#�����+�9�u�;ӗ��.���R�l��Sᶠ|�����'Z���r%"���w5�-�z�_�״�\!�$D\�dL�bv�T8%E�B״o"]mY���&:�=��n-�ÕւǍXlxVHYEB     400      f0��''�1�<[`���+o$�-a�"ɥ C��U�K��oay�_�&�E�/�5�L5�6��L�����|�+B�g��`��&��oI>e�l�����"�uyp�؀���	=��#S��]�T��֮!��#.iF�����|��$B��bx�I&��&� �u�H��D3�i������(�"�D��6Re��V$�)��M�/Ɇ�ٻ���훖Ǚ^r�.?��rIc_�V'p�#FXlxVHYEB     400     110I�V��I!��fN釥Z��ҫ-��q��Z�%��Ĝ>/zzG��v��_Љ�GO�b��|1����x�9K�O�]T�3.�W��L�sKá�����۵*2��J3�F]b�9�K����+܅�W�O3��R7�~�6��8���#��L�|J������`w\�ϝ�l��-.�3����Z�q��R���\q���i�'�����:e�Ծaf˟qB=V���l28����[����?ѱ��-��U=`j��#� lU���M�\L�XlxVHYEB     400     120性r���r�׳rZJ����#��v�/
��">� ���ȹ'��|S�Ʈ\K%���ڍ�a���F9�@��Gۯ�Ã9��Y�%��y�@Y�)�Nb��
�Jʡ��~t.�Z��	��.�s��JNHlb�XYx6�w����z�+�>uSA��*�/J�N��l�Jӆ���}u�"�d�P��.٬0�Ĳ�ǖj���I�i+"\���4���9����J�M70ȕ�?ܮ���Q>���ϵ����ay4���1ӇjtT�fl�:'�.�6:<u�0��XlxVHYEB     400     120� ��x�J�\5��\��4���e����[}��͋H�8�zg�/�������JlHٽ�Ǚ=o�4YJ��_�|[~�G�zk~�����B\K���!^Di�̖ັ�	��$a ���Y�;�y��J'�z�&�G�６5J:L�-��Y� E�*����5���r]D����>�u���`tB�$��_sgQHP��6!��ՙ�3}4��G��9.
��>+0���ۏ�M%�u_JQQP����4k˅F�"j�2z	N�w)��Y3��Q !�����bʆ�\�XlxVHYEB     400      f0��q0`{��>s�"�,&\�&C�J�v�;����t��/��Q���~Xr*���Z
j�/`�S8��vZtu@A����G:�y���*�v�ϔ����QM�Bj=a�@���x���J�c��{��<5�A��kA���3���_ֱ҈ŵv�yd��7���-tV�Ö�tҤ1/|��B�6E'�M@�列��:w���Aژ���i,r1?���=ch���
����t���	����WBXlxVHYEB     400     130L�����<���&���9�������ۀ��Ԙ5_T��G�,s.��t{�b\�EH��d�ս����'��rҔ�l��P�L�-C3�Tn�1�`�
���ͅ�ȩݓ�eV�M����(w�b�3c�9��+t�}�]&: �� ��sP��t�ӁQ=4��}��C�DR�dls˄�����c[������ע㠭����L4v���)UZ�_�=�"H�ʦ�+��ɹ����H����;��I����q'�-��M�Dn��� �r��[$��[]��=��@a�U_���}�P��XlxVHYEB     400      f04ި6F��s�3F�u�%EXM-�j\O��
��Tc��;��UhiM�'���[�f>U������o�<tS�j�e}�q�{�8��B����|�j��K|��y���Κݏ2^e��fIl?K�nAի��������L�?-�����d�.������h��t���t�sj*;c�М:4̺��5k�i5��i�?Y0EVGQA�D�N��	���m��V9N"�6���XlxVHYEB     400     150���u��><?�\u3k�D����x�T�O���P���Y��Ľ�پM�XLQ�q��� Դ�ϝ6ev�� _�J$	��'�t�� �)Ld<iAV}��r���,E%i��R�}�;���X�`��ԈE�e����8_;-(�*�\~y�⢾�.>�W��ÛI�ÒÒ�C�\Ilv����k�o`� TE���h4��Ҋ�����!�YRHS��i�.����Ȋ�Q�ꑷ���4�2�B���\��4��z���D�I�&� �%��\<-E(E	O�`.�9ӆd�5j�,(e�	Њ�Q!����q(}4F#�n�]�Z�H#(k�Vļ�{�P�XlxVHYEB     400      c0c����p���x��/+4dU�d��������j[+C�Z$�m4������\�����Y����ɑ 	�w�x���Pz�cwe��"1�����׉��i� pø��BEI�]~�vo����A�6c�o��uM�p��q�8�l�1 �x�`���B"�|ΐ��?�iH�M���JT����6XlxVHYEB     400     150}F�t����t���{���?�<�s��?@FV��w�r!�m��(Bz0��(��$VVL�#��0k��ws� ��qAL	
#��1q$��\a{X��8��.�
�JZ�������5S?��g�&*��E�1Z�N5�}5�#׻f�r�X���]}lS����j|^�=�#K�Z[80?xiv7�$�&9�#E�ؚ�Pꙣr}�h���`r*�W�1�m�a����%�]���*���7-��.]�k����h����Y�$��^�z�n�Ȯ/�/��%�n �4�$l�5&4��N�2Y��E��?IָbR�,����k��G	��^oy���7�V����XlxVHYEB     400     140�q�V�"�r���v< �+>>F�ý�&��Q~��F��|X��ٓ"���5�k����@m�Ӄ__���j�.��g�Bi��?��'u1��H,ټj�r�*T�M��!�;v�kˮ���E���r�*mN*I���jR��#r�ѝ����C�)�*x��=Ɏ� �ut}rXH�e�����y�Q3���+�R@�8��Q�CQrĽ��+R�P_i���(>� n@�Y\VM���<3���;�!�Q�Ja�n)�C�"����t���N�@�&��Q7�� �t^�%��j���-6�j6W����AܫSέ=XlxVHYEB     400     100[�菈�4�ER���;׈u-��o���U�9���-i>��1�6o�{��W���kF�B��G�
��"�tз�I(�}����u!+2�zNKb���䉃�	�Q���M��(740x���=���ǚǎ�'�K�s����̂巕��x�w!s��k'k�Iߤ�����8H��u�O���]���@�N��J�	�eP�=p�AU㦘��b�~�-�.��0	���@c\r�[�W�����M�|����/%�ԟ6OqXlxVHYEB     400      c0絾�7S��U����ۜNu�j	�#��q�;��dN��+P���Kq�K+|�U׉p�x%��k�ݫ,�Se��Ȫ��h�
b*�h�GjO�������(��)+�~@�aL%8�2mG﵅��HT�G���S��J�D�]VQ�LT���T�,���n�m���[t���O����u�̾��O�ėIB�O���~9�b�XlxVHYEB     400     100���=������Y"���h��hE�PԷÊ�6EvDJ;|�� /#������Z�=�Z>���W��ZB�	��e9Ch�h qb�3����pciQ%"�e)O��\ ����X%ڕC�}�B��EMz�V]��-C�<����;+k�9�L�>�}e6� u�mo
ym���hj�
��,�������y��.`�\8%�8q�JZ�72\���3�;e�Փ'6~�.��(&�qVk)�A]�ѹ>�tH ���XlxVHYEB     400     110�w��Mִj����NR�"%�.J�`�6��,'���o-W4=��T�8���f���HȬh�fO^F�H�����"����ox,ل��p_3���.�}m��	�+&���-�ߵ��	\Rw�K�s�Z�$��D��i0� ��K�~����l�C.U���5_�(mw���謩Ṷ>�����=�R=5�[Xg{;��� I��]E�����]T�0~]/�#��o^@�m����Ñ��R�zմ�� ���;_���Al%��G錐����XlxVHYEB     400      a0�r��@&&��g������%���+#&2o��Q/�����|^"a�xbS�~�G&�e]e�j��q��3��Nu����Gߴ*~O��/1P@i獹�P����-��)݂(��L���·((j0��w��Rsy��Rς�����8�u,ڏǇ~�8d�-����XlxVHYEB     400      e0I(N�Xk὇���ԩ#I���D���Qt:8��PŰ*��>a�������(��Pe�~�U¤�y�{�=
���#�,K�گ0p�I,l��b�sE��q���q}nA@S+0(�^�>�IKY�NS�SL��YE�,y�X��I����s�5����a�!��3٥ӛ��_�IARIm� �w1��:7�̑;4���?����+	.i��7��3�����
v�XlxVHYEB     400     1a0 K����vri�?a��̡@m�m�D�m��i]�.���ɚx����;�"�Ӎ�0V�<���:�v�������5y�#�/�u��2<�ʑ�ɪ�G)3
��;�eF�?['Ŵch�RCz	��l��[���KMDA'�g�8aܕ�e;�*;�Wg-�v�z���u�{ֿ;'��Ҟ~6r	#%����l��uT����Q�xDQ\�/qR51Ǟ�∺�{�J���L�̌�k�sc����»� �y[	]*Ѳ6�F�P�ܷ�t
��T�c��z+���{�O?d�Za�-�_�!�����NK�}��!��BJ��$Ls/�Iz�f^�}�Y��vz:�C�>���~m|����#�Ⱦ���{l�Ӡ1֏������o���/�a(��P�_��3G��>�m�2��3������XlxVHYEB     400     150�!���auΧY�z�%_R����]�~�=�}CM=l-����U8o�T������v�� j�f�ɌxU8��[6 |�Dqn��G�
>:��`����팱��q�f7@�p�g6иB�"؈�;I�����*E��!��P��c���c�Q�!E��J���gt6�]�6̸Ń20=�_��il�ʔ��2���2�)��uW�N��hE��� b�0�[+<��s��Q���Yu}��Ĭ>.��0|�cc����k��D$�	�|X��pa�6S�מ:_����P`�Ne&�v�(T�}��R�vޠ*��c�k�7b��/�f���I�XlxVHYEB     400     120�%Ǉafg�Ҍ��:#y�U����l����c�@����Z���vO�����)�sKO�^Di6�t�?(}���� �M���&$�R�BܔAu�q4�_�(%WE:Z-��U�b�7�ؓIV�U��g��3�����F�mj���ߴ��"����������kj PΟ�_�����#Pj��}E�κ�mU9�g��V-��8��l԰8��֥X#|q<-�f�w�z�Nh�WY�O"�6j��b���,��""���)���^�U^+�H�����9!�A��g��]	T��XlxVHYEB     400     1d0��:d  zk]U��"� @s��f�-oo/J�W��/�����	(t�ro��'W��Q��p�[ߩ��:�u&j;�����d`���؆n문4d����pnXa0;�����YmA����CTfɸ�E�O��<+�5�*���Ֆ�_�*,Y);F1ȥ*w��~��) _�����Z<�Sl���gF�AqNY��bs��.]D���O2$���!����` �'T�t�K��oJ��/O'�,IaܡUx��A��l�E@l��4�Ϫ�2��8� a�n���ӊ���k�����1-u����BAӽtN�0�-���.�/�H�*�����Ry�.��o,]��\ %����[�20���6+zs�C�l]��g'���-�F�<�{:T(����В���k=HQM�V
�b��i��d~W�>�a�p���x)�������fz} �{�^�K�o��V�?�>�mXlxVHYEB     400     120RS�+�i}t�ŇrP�J-"x��6�0#�D&���$x��?��fS�O(���+�jpOE��` x���NT6k����B�����c>����o�I8�HA4�����z��{'���,L�ٛ�a�5͕s����p�*�����SGQ����5K�4BT����-]7�Y32�v=���6�+�r���pP�|w�E�]�X8X�x��mo`���O\�U$5�f}�:N�D��[�0D_Ǭ��؉�9��N�9��L>��r�(d����@g�I�=g_�G2�P�-% [XlxVHYEB     400     100W��:�-;[H��d$�2�� ����tS[g���f�s\$��)���BF���p��0���-Y�h��c%�_:���)�?�����	�ݛ(q��������c�$I��6���C=�$(�V��ʿc�ة�z�:�����4��p(���$���<�F��o�I�mP ����0��[�5Bi���˲	^a&�&���XS{�9X��*�m֙��3�V���i�&�ļy5��9U��u�>�XlxVHYEB     400     110�/y�4WKY�?k���bSn�0~��?C����������!����i��
��|'��5���#捜������@L����a42bZQz	�[�E�[9���9J�!WBQ��@5�j������p�ƗVu��"�F_�S�i��������^�x���K(�鋔�*HA�G��.m���fN4��cB��+g�aJV�#�l��w^�L�v����mɵF��Qm���"*���a��D
��|
�-�j�����[�2'jZ���1��ǉTXlxVHYEB     400      d0#�Q���϶W@��ti�ĶHN]6Ѣ3�q&���\/�럭���{�tfe�<�#KG'�ڱ�Ⅵ|a�
"'{�/�>*\�fԺ��1���v�Xm���g�҄?��M�S�׵��(\��|��:9e�o�P�49|DES��C���SԒ��b�euc��A�(��ʿ�7�v,<s�F��V�e̼��O'��+�G�;GXlxVHYEB     400     100��.����3w�e�[vp�!�]�=\�3���A�d������CAGe�}}Լ�ʚX�:>� >)O�䁏��"vT�~�}��>�\�gWٳ�3�� �'�GcI��[���L&0�7e�E�H�?�+�K����"B�G�M�v��j�0A��.�-�R���G�b������
q�b�n�a��@_���5i�$��NkRm܀@}����U����P<���-҄�,�
�Lo�Yh|�v�}ez�2C�|�r�XlxVHYEB     400     130n�H]#Eg̨jx����T�~$���vq�[��g*y���A�@�"����x5�r��}N�C���Y×H�+7��<�X��b���.h ��T��h�	��?��:z��Q@�����:[��U]m�hY���CI�����Z��0@R��r.�94A��`^��|�͚����RF��1Bw��y�KqdI���[J"�҄���E
P �� `���&A�tK>
Gum��-U�Sٍ>ms3#TXn0��%B���-����r*�sԸ������ʬ�����`l��y����G�L�1 f$#�XlxVHYEB     400     120����B��J��mq�?>` Ū��L*]^�8r�}�$jg�7����ڐ=ª �,e�H�٘i7�>R�y����i��Rn5����H��縰ܧ�^Ay+N���	�PG&�����K֤~��[�9���[,!�f`�j�;Ɛ�i>�r,3`0P�i���Q����Y�[�ɦј|>�����򹿸GnQp����X�r�;�R_FC��l�8�:���5��:�W��,)6��۾d�\ׇ�Ei?�������*˖ne�a�y}hp�N3��g8��f�<8XlxVHYEB     400     150@JʧN��n�qOw&}���?�OV�.~b�6DXbr�饡d�v���g��y�7R�3)����DI�_&�[i�ؤ#�Pv�6���B���*���#�l��]w��A�:ً=)�P�:��r��_Tյ���%jT�D�*�%	��-l�$4�����>���%~�wd�ꯤL�3�2Q��H�E��Gq�ze�C%�')�@�A{�H+Q�'�����╁�N^����*��RX>}����^-��[���~�p]kơ��U.E�9�\,`���ć��X=���|�\�\��$\dy��yVN�@1��4��.#w�̙ڠ��0dt�E*��5�0XlxVHYEB     400     110h�b#�<e!����ҹpb�-��,P�=��Zo^I	u�X��T���4�i��We^���:n9����M�.�|g����]�x�x�o�%ʨ �IP����Yୃy�u�b]�'�Dz����a��X8P@�_h�2�J¦�T�2b4ǆj��)1,ˠn=7��# "�>���K1Q��ʰ�i�$SC蓱��%M��4��+�u��T���0�����)J���ͯl&88�<��Q�2ǰI�o�E�X��,�V
H ā��"�#�XXlxVHYEB     400     110�0X:O2o�WL3�����jRPo?3XT>ס�˅��f�P-�e�u~�p:�@?�>��ok��d7�'�>Xw� �~���,����߄$(��`����D!��-5'Gh�w�­�3� ����i�#�~�2Ӟ^�dT�,"�����x-�g�h�;�� J��M�/��J�^�K�j�ƥf����	}D�fp����e�6�*h=��h�|͐��G��B�v���?+B���t��L�|	�M�,_�U���]���|��������yiq�jXlxVHYEB     400     120���n?D�X��߱�d]
3���x�m�nzsJ���K,�A߁�	�;�7k㇀��'���ݰpH�]M֑qZ�7��V�9�q�Ek7>X����SJ�$	�P��% Tuo�Wž�b�g�
"����SV�?{�i;%omɂ:f11N�G��yec�FyU�H>�XM�C,Z�FT
9��{�2�ӵ�M�s����!���Fԣ��f��M��d�{�$N;K׃�7��qm�wÒ�t�p(v�I�j�@�/W1�m�Q'��I}^��� �dX�\���$H$Â{����XlxVHYEB     400     100���xqG@y���ܺa�]S�4�F�i_�*�{�$9��w��P�U�n��'0�6wR
	�}�z������a���a�C0ҼXB����Ud{��
k�l�9n�
��zzN�_?�V�9̼Q9~�"m[�*��.��8�A���\�Rl� ����c�_#�&g8z�t��v����g�|nOnnZ�U䫳Ri߷/���D@�;�u����s��HВ��0�I�����B�F����NFq�����xOS��!��kXlxVHYEB     400      f06��M��	e��Pf����g�<��*���Mõ}���l��m�dVY�{��0�w2E)�\6�������b���9�H��=�w�
�?�����	�NE�X� I��i�fT$��Pؽ��Q&P#���>~+H��R�M�<gs�z��LߕЦ�O�#U��<XB��Cl�F.G��ף�p����&��?��'��4�NyM�b>%5>Lt"qY��ԤPR�)�w|��{XlxVHYEB     400     120��D	�+B��˵Npx����%�^��y�hYV�%�ǫ������,�fWgk��m#���n+����#�����3���Uփ=:$D4�@���I$�O�G�Z��=y�˸-���D��s����ݺ6��I�����u���#�y24T8U��L��d�P��h�Yڤ��h���p�'�C�x `��R�<�rR���=�R����J㲁�p\�L*��&�'~3��rqr�������EHi��f��2Z��ʡ� ��z*�%�Ȯ��E�.?T�P)���ψ%XlxVHYEB     400     110��X��\�Z�}w	��s�_�6��V�*���ɤ�b!���ZЗVKB�k�4v�/p4��`k����9��T$G��Lη@�0�N$g t� ����,3��Ռ��7Kn\����g~�1�t�z>4C������]Pw�'�� �EN���Y�UAǭ�|=P����7��ty�f�HϰѢs�Z|�D)ca���Z ��ڛ�b�S��bo)(U<�y�?�p�at��x��A��2�bѝ�L��fV�r?��l9ʺ5�K��SI�XlxVHYEB     400     120�{"s�Q�!O���%r�R?�V(�������D���_vX S����⛖f1�J)��+6�huhv��d0��Ād��|�C䚁]k���b��� y�i=������#=;��H�*p?K�����x�Fy������:5�n|� �R�/�(�b'�J�Y�R��EǠȱ�ò�
%GP6��ho��ЏXE���4]'�UbB6��$V
Si�G/�rx�i��}�c��y�e2�z���:R&�����=ga0	_�&?T�}e_2[L�� �i�1KXlxVHYEB     400     140&?4� ��;?<L�)�S0�l\ޅ���Ás���@�/H;J$�:���4����~ڤJ��.�WR��f�V�9�rPjj0���@f<����b=hN��w��;����7�|��ݺ(�Ҟ�3<eѳ{�+����9�'U���!1 �)�W9�����?�4�xB@T�	3M���3���y����y\��w$���۫�W���R�Y�_ԭ	�� ��P�����	��(���#s�����;b8ɠ�C�̨��K��>_���%x1�sSn��(n y�H���j{ۏX��2 �	~B'h
_(0\��\��!�-�@����f�s��"4XlxVHYEB     400     140yf�O���ޜ�Y	7��d�W�%���JX=7�$�[H��n���hQ��6U����\ �;���	eS�zAz��4����k�gN�����16a$?|u|�Ld�ŲGDGG�#D'h�P�X�p-��!rk�w��d����j�����te|2���F:.���2FƸ_N��n�L	 U�2[�aQ<�*���N䟽�\\qe�z-GY�[;с��\�o9�]9��)oؘ/�d� T���f���w���q ��ǎ-�jr]��潾qcW�P/��4Q.4��w�>D�9�s������ڟ��}]�4�t�I��A�oSXlxVHYEB     400      e0���U�茣���w|��`��;t=�s�$�o���c���TM�slM��������6u�iZ������Z��vZ=��v�
ı9��>�c#��ď��NNFodP��N�wAdO�'w<f�s�ָ��wwT7~D�1c�ECm�.hi&�1]p��;��~�fe��[�0\���B|�JW��a(7</l��)?a1���U�)�8P�[��:�L��:u�� ��XlxVHYEB     400     1406t�{J�� ����՚vQ��Z?\>O�X+��?}��@��e�4���Q�yn+��#^�[©����@OT����,Lw,K��U4X�f)-�y��  �֘FQ[��3��p���r�_�(q��!rvn�,�^��]̉�쥄��������!�� {w�wb��<���

TE����ѵq�|�>�Q �����:�@��h͜����ך{���H����r���@[�D����.�����L�ѫj�H��ݑ�6��Z�A'<\�O<Ѓ��G,�,}r�5�X@�U��1�>�D��� LƽOgbĝb�ZK�-�?ՏG4XlxVHYEB     400      e0��2�ajQ���mԈ���7󆎝E�]V���
�Oj8&d+~X���6S��#��S6�6a����=)	$8HE5�@���>�!�\w]��0�lN�3�@�=�!U�Y©��ػ�J�����OO#�|�'�;�<�"2Zj�[���_/&j
� �F$��y�όM|#�P!Q������h���O�AF�D$E���cdGx��炢�L���g�r$JXlxVHYEB     400     190��Ů��_��6�{� ��[�t�����#���z�u����-F1..�v�������v3�~0��Ecv��r�1�b��E�Z�BEO&����)K�M����lg��a��� �z4}sef^������8*\�����xHl�>���,=��}�~k�6L\�t'``Ϊ��=�J7i��x>d��7'"��/.� ���cI1ʒ��}�0�܀/k�LtA
--�tG)���g���l���Q^��!���^�IKe���I���l
�/^��교��our�i6��H�����l(!$��6!�@!,�p�R���w�����J��aR�oD\�x���ٜ�Gaٱ�S�'�cU>Seu����~�+�b�>m��h�P�ÿ����XlxVHYEB     400      f0T��1<xa"�¨��OM̫͠�n�My�����B�T����T�gm}�c\�Ro`+�~��s*�@���-�gUi����WW�s��u����H�3����l;��L�����& 9�(2C�(F���7��
GH�b��]�5���qT�%�9�<���!���M�x�F�ώ�F4Q��=��P�QQP��󁢆e�9$�Q��}(�b��Lv� ��M�<SQ=� $�7�rJ�iX=�XlxVHYEB     400     120?�N�>�p&b\���tR$�d}�@�-�JO��-}������zb�e�妸��{�aW��~���K&�?r$�paR�7Xp����]�nGԳ���yUl�S�:~�J뮺>�1cn�ȩ9����JmO���(zy�����
����;�ȕ��2��ZTjjY7�fdH�Ȩ� ��!x��O��ښ
���pf�|�/��_��;�6O"_a�+�a��$Ƃ��>F�R�0szi�������=���ͣP�K'����BI���k:��`XlxVHYEB     400      d0	� ƙ$Z���;;5��I�?�g\l�9�x����_�*�8T(����Q�T�W^':fJ$�+d)"��wr!�*ĳlO�am4K���cO�4�c(Wo��l���v���鶓�0�e���%�����I|�]{����+��x��|���*~2�y��i��7y�o�uw�7�-�q���^��e-P�)��]�\��jG$!��sk�,=�|XlxVHYEB     400     150;�5^�-�s�{|�E5K�j�`�{��&�b$K�t��c�k`K�t��F{�� p�Nd~���L� �������
X��o/�:�h�
���28�gAvd:s��嶷� eP�>�B��!��o�o����Ol�L`��N�����A�rA6�G���ݔ���q��2}-U�2���*��A�0�ȫʬ�$�j%4��A�x
z�Eַ-v�B ��������<���=�h�b�oL�ѝ�^k%���x���. ������D�2?��><��*��Z�n���!�nz���W�ui|7taB�-����<ۭ�_���Ɲ`�~H�-~��mP4	A�$XlxVHYEB     400     180�o����rw��i=e�2[���9��Z��{��o5�zj��IUx�{HJX��ą�v\6~)��&�+�_kwm
�6>Pb��ܧ�/�1�7���+>�kGX�k1&�׿���H�e�%�b��b]qB��~�5/�N��)an �pg���p��d>�S�����I��T�@,.\LѓQ�@����(SU�ܫ-E�(�d�7����ܔ{P��uu��0��ĝ�%�EV?yA����7�U
i��C��+��-_���e����֯ɤ��D�Z�)b���pf�<k�P�-g(T���k��|�u���ڋ���-e�V4��ٶ>�J������T�~�36�O{�N���t���>y�h,��/C�v�e4�a�ERC��pXlxVHYEB     400     120w��"?=H��Ou�b�Q1���/�t����jn��;�����!�VG�t�=��}8��0���^^ܶJm�'y���lf�����
����	�hm������a�;�=�@��N%��_ ;F�>T M��T�ଛ�ܐ���}wv�E��l2�Lջ�qSh�}�b������D�O�C�	��,
�Q�����F�������B���S�";�W*��~-.Ț*:~�?�����Q_J�+����:�|}�(k.���*�P����[�J�ԑ��U��V��XlxVHYEB     400     180��7N���d2�\�%jҨ�F)|������Pp#Dܟ����<��ͫ`*w��i���0�KƨBP�b/&-AQ�e/�k�C��^B�L��ͳ�~Zy��,:W=p���FW0kg���(Ek��k������DC��,AWXIOI[�G���*s���\a�9 ��U������cK�F�E&���>�=:H]փþ{ĩ�r='�
��a@m&�ѝ^���ST�)d/�����c�����Ǿ�0���݆�L�1�J���c���]ߤ鵈 �.â�	F�b�؉t�)P�-���A����Z�KVAO�&V=ؤgJM|hUY��!<�Q�z5Uo[A"�W�����x�|��&g
����1�-.�y��<��F���[��!XlxVHYEB     400     120��'7i��;�t� 	��D�1��b�>���+e��2��'�^��}�l��\^gZ/�d���t�$�,dr�e�?���w|�x��DJŊ�<|�����QԆr������/7�:��E����5|��2P�[ x��5����~2�	M�QS3)� �Fk)�&�߂T���R9�Fi�0���ٞa����(�4��glúo(Z=Y�{_`���kG�K�z@�4-�D�� ��m�1���ȅFP��]ӱ�W��w�+��Ϭ)/[��[��>u��\1ݽ0�]��@XlxVHYEB     400      f0̼�ַ����K8ݯ;PB�/:7M���F�R�
�3Ο�����-�h�ᪧ��y�d�T��B;l��X8�&�u\?��o�6�-�"4(D:}>JȽ,�~)H�����������΃��$�S*v1R��<:�t;�w��L����m����&2�<�����@��L[b������E�9T��E�e�&=��<	hMF|�9�|�W��}�j�b]9O�X��(�H�������XlxVHYEB     400     130D���WV�+�u^��Z,)��fW僆W^+��n�̶��o �/tir�3\�蕾�ْ�e�V�3���+�� �泋<&U���$���{U`��x�x�9������F�3���J�g �:.�ʏ�D�O��m:I��s2E>%g�ޯC�c$I�I��,[f}W4���C�!Fa��b���qR�*���9&��͠���1�Ps_�˟}�-|���]�c6sog�:9����@aU�p�R��E���o!�9r�֘T@Tc�hG�9j���R}���%���F
z� %�n��o8=q�����>��8��)�XlxVHYEB     400     140�*�r���s�r5	� ���Fn������	,(�wh	�6�MU���1v25u�ڂ@G���2�۝|FM*��l�]�JpR�B���S�ħ�hfu�w����F�o��!p�=�E���$��D2i�ѼZ�5�7FU-����ԡ�v�a1X1��X%��T�r���ݦZ��<e��$�B�if������6WKA��)ƞ��C����w����G?'��="_=�!��0<��1*Hᗸ7^��rӖ1��2��1����Ϋz��(X:;����<G@�SY�Ķ[r:��֊��"��HH�]4�ǳq7_�H��XlxVHYEB     400     140t9U�������]���3�=�5O����<}�wYt
r���Y��_�?9�p�M����o�>ͭ�A�������T� �U����W$QƔ<���ۺJ��w�#���|w���'�*PR�'u��$R6G3����$[6��b�9�cb���㼑�j�y��c�`�8ۅ�[�+��VYIJ%�_O%��7�%���nGh���x����ܶ�FET]�<�7Ry1�v8
�v���Z��Z�=�h~FR�S{�����*#ή=�,�Q�K��w����~=:�I���i� VSSu5�!��� |5+A�E�Β��.�"5�TNXlxVHYEB     400      f0y-q��4���1�[Ik�#,z��G������͎A)�r^��6""�=oo؛�=9�x:K)���pf�ʜC%���[�,�����|�󮒛�� ��6wRϙ>�;s�3���\�/�;�ˑ:����䕏��{;ov�Ѝo�*S��R������'�[����h=��y�ƿ��bf/�B=̨�A2"dD69�ڹ�zN�U�y�x?�}&&������/դ4�P���{#@&.|Fb�XlxVHYEB     400     140��F�ow�{2~H*�X|��B&#W<w�)l�L�k��8��Lqik�k>J����.�]fe�;�>��C��Ũ� ��� ӣ���p=ͣ�3y�Ӵf}��G�u�r���`eM�	+���6�
ZF�˞h,l-$cʁV�Z�K�X�9�aNk>�����vV�T���=+ɡ�a2z�2�Z#�݃��1ݛ}��Y���b�Z�@L;+�Ǣ�0%=��n� +td�U|Q�q5�}wE�F����7�+n���� ��:@�U �� �mm�jL'����'���`��yMj߰q�W8񣫔�Z��AȠ$J�Dt��z��:�2XlxVHYEB     400     120�~�,�j�I�G�%(S{e���j�ǹy��+eX:��dC��XE��.��iz���3�^���q���p �<ڽ^}��26z��8�}+v}�ƥe�3(�h7򖺾	�]>Q<Vː�14{�k��Cy����X�=TV#�<?EEq=a7/��р���l<]��9���ڔ)����b���4����o,�"�_\�l����h�}^w�7ʅ��S�N?a y�,g�I!O�a�=N�D�v������
�tg�D�v�X@>9��as�¯ya_F}lXlxVHYEB     400     120�M�6�-��)B�3
���4�:j�3�C��>6Y4p5n��D���);�@��]S�}�/�b�h�m_��Ӑ����M�_��`��<G���Ym�>�ԡ ��4��jB�_j�K���ĸ��[8�g�A3��j��<��<!��˿Y�@�6��˒&"N��٭]��S�, ș�>�WD��ӡ��5��a��+9Z�8�`��^a�Q_:ن|%�)9�b[��e�Z�����ٛ���k��<�oN�ʓhRڍ�U#��ܿ�ï�%�)��j�����x\S�IXlxVHYEB     400     110�ݒ^ռ�U�wZzm���g���?L<��b��R�KK����J2|Q���t�"���-�K9"�@b$&Yx����H�q���t��v*��SBe�Ө��Z������:l&��}��_2o�piNcn�b~lܪ�b?��w����^*�0s3�m(ܣL
�(�^_�#���̿�Eڙ'��?������j?d� bC�8�Y���y2~_Ж �NH�Y� �\��x�6�u�"]!�Ƌ�/�T���y
q��v�|j6;̎tRP�UXlxVHYEB     400     1606c6"v�O���^��~���!�q^ǎ���ִ� �Z�\޻������_M�V��vŻ�n�T�$+�n�\��e����e���e�1��Lح�\���~�/�R�0�Ts�8��G$��}�I��vR�����-���.1	�h<ݭ_(���r�[!��n=ܝ�,!#5�2mUT��r^���(�ȋ���N��mS�%(ix��c^�\�M)�U��;���H6����+��������و�#3�����!�賙��}�=o~�l�̯v*ʪ��k��C��n�W���'��(��t��ifҭp�\�ǟG��=h��C��a�&ZnT�__�F�̤��RPXlxVHYEB     400     130s�:�r�$�R����� ���;��w��)��̡M}�VQ�L~��m�I��u�j����E��Di���ño��U&]��_i���^����_�����l�4`_ ��HΌ�/f`�te��'~�v8�����@qh�F�6�����Ȁ�~t��"��L;C�'���"�%�j<��J�c_��K��}W����S;Y�0i�勃�I�,`����g��r�2�/�,S�,�F�63Qb;�#�]�M��&QX-S�]�L0��a���w�����N��VoS<!H5/8��H�2�s�V��XlxVHYEB     400      c0������� �ѐ�h-�O�ӡ7?BR�=r2�#�M�F�̈́<܃㷝q�jH9*��I�8T�[�
w԰�C�c[�V	_�{�e�G��!�Io_8*��[��vߪ�H�	[L������C�%J���*f��XDO�o�-iJfE�3#��pPT�B�Ɉ�Ƭb}˽6�'�����XlxVHYEB     400     140�S������c����d�EgdD��qD��a+�������Mf4�u��#��g�c� ��s�@������l����EW��HO�&
� V���607	l��Y@��
ₙ��XKIQм�n���Ȃ+-���tջ�3b��>��w�6-��P�)N����,������oI�=�)��=�7e��Ŗ �z��؜S�I8a�%%�f����󉖻L�w�^�j��\(�Q��A�)�.?F�6S�<�F�i��r�T�\�3��fJb������i*Q�'�H]�,_qQlew�q�Hj��6�ߖr��MXlxVHYEB     338     100y���&v�u���8Ep2 ��T�wf�E�Mw����#'����N:���9��|�F��>�)A�v��iv��(`#�[��3C2Z[{��_�f�6�g�L:D�]8��,�Hy�
�&�<�=�ˈ��J�(��M�����R~	�OW���)e��8�x���W��SC:��j	�YzX��*�_n�SPGm�G_1�K81�`���P�9h1!�:/�~%�h��ln��b�'X%�6�j�"Β��58!N�H�с�ui