`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9152)
`protect data_block
7gUddfP/Qi99XY4FsUGa+s5QqnEdID88kqBBQTH8kz4lgRIrdRQ0SuFwEsLfG6NbP0OsEWDJMhlh
DDbE+SuWBQwBfT914JRApKalCDzo03C6mFCeOjqPCIgli43Sj12EtqRTjOIHd7IzmqJlFENZfT11
XrXeCpfi13AZ2U0kKlXwQF7KX4EVKILoim1dOCjKhgp5YrFPcsomAhyRguuoHmCiGbSyFTOQKcZl
OR4E4CTeWj5JPP29YECd3c0sTuq+DCeWwa5oAXYayeg9ElVcUzVN/RmHuSrkllXi3H0qNL8MxwFM
H5Ndv1PyQSqgq/OT/IDNNWeXnM+010w3iQV65ysHNN7KZIJaRvo3UE34soiNZDNR0I8tZtpdERTw
uUV2gRVplLVnvzL2oypvU1I1IXvlZwN9NOFJ7sWuPDR9lZRp1GBH2P1jZMiI2TijWcVJ8fn/sA2y
mqSBZfbTn6KOox7XbhzFEdLzR/ZftjZFWqhlOwbzePv4XugYwBa4wuQLpCZfp2Tq3jte17m8kUfN
ZjCkxL3PS908dcF7lkZkxaD0ta3r0b8PLcfQOTdxsyP/E01gv0V4H+v250BGKHlkOgaAKXHF3Jkn
PEZ4w9eIssKHJBDv553t5pFgoWReEo0EeMzYVme5bXzDuJ77dP8C30cfnyAXHOnoTfB/Lb3tT+So
7jO/EF7ArKNeaFBUJve4HbQBafhzKh/94B8JCEBw4uUWO7RUifUPuzdKwDnUBw6eS6Obk3oKL1Hx
MpGt2nnboWH3OJ7LEQkgFsrMeI1FHZwQrn/NXxKnfVJLDai4ugGKWVCRybTH4vDQOXtZAVHoQK0F
qi5c2wXGWAO0i5sQT+TdnL4uf4KCgvCfCKNASy9vS8U913PblFeJcM9jHhgsaCUJHoaZuLXD/c9r
Eb9oSBFmWNAY57WwXtNd0RbwaexYLjrOPgxdqfrrAkl1Z8cIsweaN5QF/ehvU7K0YmeNzDJNoMyD
Q4xvjJmfJ7+4hiy3WaZjzX5YOpbpiB0JjlejO+TOq1NvQ2aMq7xOjJTEuKskOdSsnpOt76o0qslx
7a6zeMPsSdzZ9/2pvqFe+aExx9bRQGlB7UdUDy4egqe+9Hr062NtFd9snwh4FXpOgNuL3uAayX7a
OXpBmvR7urcOAxPQGXf9oXAyYGtm63ihDPX+RJHqmIBsF/9Ny3F6oetbQ+yg6Ki8zQgfA9Y34Ywb
2NV5cVz3WfV+Egk8VsX3Tjviy53b9otY59tkfy9L6neKgWx4QPx1HYBd5DmCRGbMwrkSA1OddZOx
FsCwY+dmSgoc8Gsa6crYXZvWe7cDV9jljeseeywf4dhRdlmEdlGyldUqiVI3PnRs4LzdC3G7M6Tf
3d7FBBHh6UCqmwk/pBe3WPh/PRZNd3vw00lp5i1ztRmrUrp/6SG+WtGF3cL7yiJzJoFeF1oNsv4X
Td6xLP8xrGFWzX2uD6Tbe6210Sdr7Os6zylxbUH4tZQ/6wwy2aIgOC8YtpWitMDUt4vMePZ+7m1c
welWp3j9Cr44yK25H8exVCFxZn3f9GIDjrS0xA2tn2Ot7GY/PsyGzxqcIVNXzQF00p+q2iOAeThP
9qA+3APjt1SJXSfbCUSSfv1aiIFZU9HMYHStLL+C3p7CqN27Empx9h8h6dERPbDTA41IzZLRNOuZ
3VvRmNYzGl0Xs+F5MImMMfRinn5OA97MxGPNdD+KIxJp8FrTWAaK0aF/q0EppuATex1FEUlW3x53
Hfnnz0TRGfX47o1L7nz1DxC/IqK82vF42HN5OqPROyEX7so+uO0MgAZvQH0IxO3+/FFnk1hrLhIx
aNy8oRcxLSpUSWE8uExmlL6Ra1vqaK1EL2ciwo6gR8/bWmqW79483+M859jsBebNKY1XwldIEPQm
uWxggWwTZtQJy9JBK0ujPdFYa7XH33EP2bzo5gh/PDitrZT6GCeevcwxcOnFU/FScUNb4xMFfg5A
lI/4sTeGcyqdZ/Bd6sJNQqgFEa0kFZ4S/4mc0JR5v/muAMa8C78vkO6ukerMpHDTm/vyNRO9zfHh
OhItdz2NXu3p5PawLgrKwlbhXzj5DDsYH8gndtWCWXm+GhoJG0fnGi+Ta9Hn52/8+A9zSqQAIg2O
lxyIOg29dQVHoL1bKJLO3MGiEKP4nRAa6xCLNv4Wk+ZeSkidkLnbN01WR85e+IdTXTGJEL5QGbjg
uboaNylo/G5BQmdVfGhfOx32NX1Caj9I6HIT9J+idOj0A+mnrV3jSo947YOTtjguXo2CchxQJKOA
/vFRHk3FOd0UMohkok+iqK7RiFk2kEjxPHUtlCpCgnUeIs0zq/6yU+1kHY4pGNh5gR/eTGI5uCgP
A2FEPPMX4Zq3iugv18ROuh8IArS1DNQd9bfBYp8ekIspasSf2fVTeUFq3ksjU8QGczHEMn4tAjco
416tz/Z10gCLdqIHdBWz3NGUIpr0jei9wKwvkPEpHt1kZI4+8xmx/rLaOLau8K1T94G7CT+QKKT7
sLdM32sZxpGG+3ctwSceufRjxNTEKo815ugq41XQEdBifO+OujYvNhlPKknCPUszTffxfdtiYLCB
iRObo4TNtBkQeqNV0JwgPH7mIc98fGpWt8drBivSbzRQ3nV2DL4IjTB1TSAjYAG8bBZoaAEHLbvC
yvmbV2SxwNkfVYzkEQ8mE3Ce1+5SwH3egPtXZWwbKKEA08i8L7H1AEcaW3vEQjwnaoLpXD4NJ17u
PJ9lr7+g60nW6S5tf+7GWlMKcHiyn0gCZTxZ7BgQxsIgUv+6cCnAN3/mN5WvoH+tiwDtT/iT27GU
r+jFHsSchMafmv7Wqpk4iZ2O9P4JEgjIQIwsnNayrEwUTKORKLi2+1vgXPYGgu4dY7JWEyWjsabZ
KQePIE/FxtRzbhfNHSEuVZHwGLkitIAiOqWI9RiHH3+ldC5mdga8djj9SztcZxNGU/IH1VbBPZvA
e/yaUDk/k4QKFV7iDbSLeT9iao2ERoDgAGcCRP6gFbzAoVggQIyT/XSnDIOhfTH7ad3loyzMTKxQ
KcTfO2bhNom703cZOr8Kpd7Yag90UcrOnLhIMiy7ovzedn8l6vbfK7aQSJqHeJUvjacYvbe34jJL
7ICbA9EqMD05mkkNiBwNZyK8vCspBrXgxtDiVngOvD+l7vEifB0zIEP3UFI8SLq0/MsyN9kQEc9V
pqQXwNzjA2PzodAyDzICqaEKyu1nmB/getr6wkqJPtkWO1FG6H+PeaEKTtZQffs4eKp1S8hyrFIB
5obkoq81BFsFRe1r9bRIdZqjyk62ZvAW9JIszR8kMFhn/zFyQij5biTYfbOy0LzlZm7jYkF7Rtlt
Ef7Ysaf4YN0ANwyxGOb0dQszyNifujSIRfrGHw7n/+xar9E9rBib0nM5LPJtJr4akL0pvGpZdxdo
eqvyNT8OQ0Neq9pSQpFLFIbf0jslz94ycxeoBJe53V3Iy3TqZXSVh1K/ZAr432I3y9Wk1WMnqmYj
o3Gt2lUHNFe/WrTkN9JJ6BOvKqaJOsStwyFSfEZcfVCmc3e5mw65+X9hEto62dGu7NaZOl14Uj6y
b81AQ1daxEgE84ndKuv7w+o3p953fv25FpL2O469fHRBssfUi74mn8P0CMRY6+8OYcy40UEU+RmJ
w55QWzDCT4nWy8PyXY3d5VE/UeKnY/mUeAOZHeqeAk29pDDmSVPNUl5TJeVAnCDpJgdfwtpyftu0
i5wHPPpO20QfgYk0m8D+GtXBK9w+3L88mZyKvOD/wGwa9LLCoKtkj6NLweJqJ6lreoM3WFu9K+Ub
iul/ltNtR9lq2nmWvEmqIjb8sDa+1Mu95RYde6bWwSSA45Qa7U6OOZBUbDfFOhAHs7e1GiklPbul
CJA25NURCT+90spgGc/97zSXs50MNNYBa3ig5QSUdnqSqjLfpmfsYLmexf1Ivsu5s5OZELaTghW6
/MbYeEfNhb3Mh2RH/B1PVe4Z8RW1oRifsNCswNh6qSlKPqZkhyuoPTIuKefqBoH45cHJ+o8b+u3X
CYmWvgRYICvlYSyhXMJgzT0AxBB2Oc6B1sqTfThkMwtIo5Ujz23mihPPxL/H19mDLe1lN80N4UAn
qkwuwSrdQQMKlLyPXIi8hUf4/ApS3fs2jgLHOYGOIFbQxpXUrKazEo+UkqEXRPHc1rvicEl0+U7s
xCKa+d9WqYGQQgPm0q0Avw1+AQXIHSy5Ac0TUBFxAfsVTizWObz+03lZxNRbAGAcDn4H9s4utUs8
fXyLK6/KLk2WuuZNL8DQQHYW2lofgJ13U2KXwOIA7HpOY2eCKzPiIaoQUONdXvzTvcNmuN0F98Zf
1kGAjF3azDi8CU/keFWrc0zZQXuKEou0VwbsTaKWuY7XQfjifCUR2GgUD7aJOm3+pOaflNtCu45Q
3U6iLW3rnfYZ/DleFFobDSdznHJIofmThGojpMY0YyZRtBNT/E3YlK2INcm+1aI1vLQGMbv5skSh
1yBPI9lsO8qrV7eY71K+58SPQ2g66XAzDILj0XDVqQ99eCpN2c+5sgZi2r0BDaJ8dNaswY4QODm6
8pAjudFxbHCukM1yNE8tClBNU9sBPfmaqbMvRNxNbP7tWEmBfcpivPiOGyNa2pYq/8TbhMyLQoQ3
S1ZFWHipQ5oNAldFpTcI9SVCzkKpL6xHOmkapHeHsps3wLSBufFWOzJPLe6M0/FHEvkPmZCBbZ+J
N8WXU1dCl3V2hrbGOiOcqQq0QEj0A/gx9JFVaXs0RmXF/WoadqZ66kjmhUwN2ox5ezv+Nacb+q7R
4IbJwANe51mPEdyaEvmxTLpbZFnlHrQciACnjFjkEeAqOnyGtjRTk5VSXItS998AyOFNutHK3XUj
JBhTrPSgCiGl1iyDwz4reNzYMa8goAs07ENiMbNrkaRi5hjh1c6mTkoT1/zZwWxnol6FHuxCMdsZ
b6O/9cOY/HNzXM9q9R06VOWJyTiXB0OKNM0VaMGEOdKJcXqu46Wd4cqNa2bD6iC9CALJHSX42iQ3
HPVLTIp+OrLsbi/pkcIp1l4iz3eeanfPPjhJM48ahhPqQzqm3VAscccwfkl558E2vz0zPkj1b8WE
EflGAyKlwk+bfMd6z9rE8HSk2N9FcrLaefYnocceeGK6Q5GhEFbDb0hO4tIHcLEgHqEJIABGFVMJ
wj27jw2yfYGydB28Gvm9Z7W64p3xT1jsf3G9awxpUs1WenXLawwi8zqjvAXcIQ5tad+N11zfP2Uy
N5s8nEBdBMBkNjKqScTmlv/tQi6dvLNGKwu1equcMDtjDk3Qe9Exno1yTT+cbzkAotyCDDmUdwmi
2IWYgvh0C//Ac2l6M0yBkulmE0Ey59h47mgkann7D1dv2CywJkd7BU4DpQIfvt3whzl5YLC9tW7p
MCiSqgpXDvhT4ctpWsKICiPIEHtEzXcKSe+Jb44DOiinhlgp4AB2/B2BKf7kEEE9m719OxrmRYFf
a6l0/6H8hUUk2Xqi94+TiuxzDaAV3gOGpYkqAZd660On/MBNVz8fZKo0w0CqFOEUqXFwXjXynLw9
UGqbO+Hk769qxGKe28o5w+h+82wxSlla/WSu+YUawpaPv7/SaS3ybfQM7iEgJL3vgqxSQcsQD1Lm
nqb6P9Oh++BlRLKkX0wAaGIBR1V+EYWYo2fq89rqSOjAbBDtH1sOGzCbfKTBbkIQpB/9p0zCQtX0
P+OLBNGTc6vnEUxz7T3uc8nmN0mx2W/3Y3gPBOFamkAGsFbbck/jy4ux+nEu3E46kWmlwsQ257O8
qSfOguuXil6j80IwJNyxVZsDAfG0081BDOICtpgscQpUjGtb+/E36zsOsSzgJkGR7vOv2/kGH6Gj
J/caHVdNptkoJBJr5tMjLYLEsbDGPieQPuZMcgPuhk8nrVmEDpsTVtpZ8ZBwoao/1pa21FIfY0M0
FtzWr/U7Cp1SBdipyNZ1f2+C5Nb4e7W8Zomx5ZP1q6X4Z1wpYaqsJR6qCsfsZ0OZOnsm69mWF/ra
Gy50aanjB8bt2VtELI3hFyaTqXyDpjSee7IYvdXwUUyEGid12eLOsdbZWuLIYgvVEdt82GM7APdj
4lkuxMuASx+ITGwRIHHMChHpV6fPZ9+hbU5YmzDUDoMn6B6b8JwSY9oMTe7qLXBTOOp86wnmVQUe
qGFCfAc4GavO/gpz667RbxJqJlwxdc50d4bu4+s03M8z042tN7oCuSaGidribAyzSqpiWsVWkvGL
DZqFVAMaLb8EbFoEc/KwJXdlQgiAwukEHpJcdpbadfIR7jC6MEEplcQQSVJvzebSkrXrqSa6RVLS
F1ew/XEsBPLw01fGc+nyvjsJ9Hl1PcUy1g4+P4MfIEr816sZ6Kis0fJg7HLKG4BKfmyD/agJw4lo
/mwiTDV/yAotMDJe2JsvsYfT/m7jfDEhzF/sFc/podHVEkATERzisUfNf31WHhVepKDzCyHsrHYo
IRpNdJZuOJAsiP0PccIgvkCofRv9Ve338duUxxa8EOEcx69qfBmqry3tMrX4D1IUuxRKjFOipJf8
KVDSEd25uPNASs3AsFw/TBIidEG5/xyjA7ku+9FL/MT18ggu2X2op/jcj4RtCkbsfeeXu2gEjlye
STtEyLeHlP8Fp5lY5reHKFPKuQVR/m2EDk0M6tD4nnsRd2BX3Ids+0sAXgwhSYlLdPcMLuw7k0F+
M6a2UmOM215SLmUfi3hKVdIIjb8/Xphslkmuw+uPrSHXrBHaRGd8+CEy5x8pKksJBjJuKAAKOzro
PS0MlrrcxQrdYfHbXJKi/zqYAM8hLS/V9UlIoEw70By9SMv+CdZ/PJzoWTxwZErd4VcwDHG8gCxz
HHjnJP3OLg0pEZknMHby4sks2qlph3Z8MSJ/28GtNIC+6IQYKxW1PjYNOrgzA+fDyCBYhaqw++Cu
DHkHkfA7+qlLL0DikCtOwWDvdUtL59rFIzrsYqjL+UHeMyd5ykC47hOVzaDcOdCMluw3Pz0GhxiC
TUQKYnx3uEw+hq4fZHApZ9A7iGXH7gPyFIQYSCFoTOFox4uttYBzeDwJYQAF5V5h21HEc1dBJETl
ZdgmK72N4Cu+zmFV6Sa0tlx58StYDPrXeyHwjozMTvEwFTeMACmC/O6RiMW0Ys0Aq9Fpjut+P2pS
FEE68Anyq+REV9LP1HFImP9aDGxBPZ0pcvZg3nBgSPRZfa7RAl0rfmCRfitf2hnTTuj+wGK2edSG
F/a8WFIVgA3seyo9p6abdtYieo7CM+iIC+o1lfF53BiMnGWnPaKnyagdLxcxqFzvb/SetKARkCUw
jLv7ojDj+ubyDxPwPJnIvIYnvcfp3NuhXY+iV/ja+qI8gEFtTdlbSz2BBOET0Qsd2Nd2/AAlYszt
iYXcbo4SbwHmU2x+j2DZD8cEVHbvv2+2tPLTTQxjBYai4nS6tXb1piIlDQoAl9dXDurLhBKYV4De
hRF2htQkrMZcXYHFpLBgSt0O90d53wWtdg9TnZUeqY2/8uTr2UGXhGI8fV1hsasb8kZcrgxkzoWL
gJw/U3fLEnZKNwAUJX2qb5p8yCiyWLUkMwleWX1rt560F5PDQ3LL01t+NL53nl2RvFZHiZiMUFPR
wwy7OuTarAthNb1/AW6GWTFjN4BFncZgssTj63VPYZygRUAgO1POE6exXx/fyMFzmWhY47tYaFAD
dXo7Ik1bkRNvRwl0/xvNOzMQHS9voi7flABdG7bk7DZaPC8xe+/gRja40ar3w26gQvdT+xPJ7DQb
M5QA3NUsZ6cmLAcGK1szEk3rbdyVOCj9wr57S8E/A+nHdH+OYx6ZOZIXdBSugD+FsHovll6VxJhy
8TSouk0q3JwU6gMURR9P31TK9I0PUFuXBdHwyHrkFJcK0EWo9L3DUfV2T7D+59JrCznTOZHw/9DX
adsJFQrx/ROsxXW1kB5jHUV8WD/oKUOpsMSgXG9xAC9IeR1RD8+/mR8T+F3ldTafXk4pKcwWmKDf
RFRWPtgDP7bjDNLs5VqBwmYU19kEyZDdJXC7NLSZ2X+bKas5A1GkOWtkpG9AvLBIoIRYu8BmWs/1
pjG68QzjRbX1wjjfBWKq6iMgigG2SI1Lmkn3vvY9sXpfkrhJC10pkccm3A3YP9dY95OBDi9Wf3cu
cKR1SitOByg9aVAc53KMGQrMXN8GW+BMxFrrv+b/jrutwExiAGOKOnIVGmQWippnbOHrlCkqPKTH
bxBS+3HMbN7TpTTyyi+3NO1vUh16xxS9uJgn85SZmUzysqnzG5gMAdnFAt5XlyYGqajKU+wPE6CU
GL/1vublGEbbr6Ka2bKST2xeVw4+sJXBPCtbJk/7vpVrlZmhkurTIcRyrH7ssPHY+9VjVysAEINe
M+SEV3lbTTOgKFDiQU+3taZFsYfZrey/FC7TgypCmynGtXtSlFQXp8XqSTwa/E/LNSSP3IiRSZF3
VwNsQnzRUQrpnJYrXEphYr1R81Sq3xpmuau+iJS7mEYFpQRewcarwfrgq/j25Jxsm4/cR32rdvPN
nPVb9eV0vTNgWPz0uYrZa5zNHBaVk2B7YS4YVGxF0KVAhiY4foFFlG6dbaIXbT4lVUYmA0A0LSsX
agmEglGKUsSC9FE3Ckd1KApdJqDcZVkOmlMaybNYVS5uWS6ipmd6kkcSSNVzY69SQ2RX639QTfz4
8+rv1ykobdr3B5kUwMk7boJOdU9ls/BrFRvZJq2oWbFIkUl7c/5oZOKnc8rAkzoC2H8ZvU0ipbSI
hGPKrN3pXZm/6wDRKKKVh83t19dNYMvQeeGxSAjEOmezCAa0kWFtaOx54qmP4JM+Ut8BBu/qvEWo
i9jV38nWo+CSrePY5N9zxyDQOtuMg2WxdSp7OCRbumyw4m70VfhC6sNOGPR9/KmoNs/FDXCAEWJ4
D+GCz1nwlsmRv+bEuwPtgN9reoLqR7csLlHe5y67mn4njDT+9Pyw6w5eUb3F9Oo8OpR0VLOdvxUV
xfjAU1BuMnqGHDRQBBmS7Y7+vmirCJUCDGa1NfSuLqb8tQ5ng8sKsMOUBBwnNlNYytsND+UNfWaq
wUV1lbGEHoausFmrGBW7ikct6RTkvj3LEg+jh6cGwdxLxpF9Jr46Xm9Fm0A7RSFvMQYgmXiHPpTQ
ZGtJ2ls2f1PDna5ua01qPMp7qcosSziNtesrgBCWzA3Y9pAUZ6Xg4GRIbkLJpWBOPirX9Xq1mx9X
NlkgysHesLftJJjvdISiD638ILwqnLatVfLHWjxJq5aF0hb+NUPKWze2b5zVq7eSHDf8mfX33MDk
Gcg/Cubnj1pDWxBxF1FvpmYYBRw4NmSrkmXWTjN1j3XdTCYbcngJ8Ee1DG/3QblIEz3MnBYr55RV
OTVwiu1PZOSChrODCq17lC++bpxqq7FaPX1nQ5hq8JTls5cqceDbohas8F7Zeb2uvxvqPp+FOP11
6V4Q/NwEGc3STrX503Rs4Bnppl3oDUe11XLFdaZZaTcRSGOGoH3KqpFYcIc1PNWEHIB5oGjoERLq
o6p8IMF19xb+NiUS+qmm0rTLlbsGjJibDVBWzxAt7asORveae0XZWRmGX+kq3j/Xq+Ftbq49YEOw
Y82S6KGM96ghMxVQbx7lkoVox1Cp5KzvPxRt1m3pFhbzZnP54dI6k04PDifM3+C4/AVCRBDjzHef
WkghswGWouuzY1VtHr4sqU9T1nHC1J2jMPcyLZ3kwi7bga2WXJxmQONbDlIF+CVID3HVSSJFLviL
aoI59z4ytMBdE3sZJrytksMBYHLri7Dirn3Gll9EBKsC/XGUSwsu9kwNcK/3giXCP4E62giT2bg9
2ycsk/OpD1U/s89D8SgqbeUeBRu3P2mdET+Zs7Bu9k/5B2PMB8vR/b1EITCrcaYkJ5aAY8NTS76a
2SG4ZIYYyqiqpSBV97GZC/Qgd6EmXMu8hwABfUka7cXTzUDDJbFW9kj/NNt7w44rz8NVwUjlum8B
sjwgTUcPgB3twxU7e4mrpOttX2iaoqbSdtD/VqzxV3CJwvv9S4xlgh2lgVAItxznpveluJwHaj43
KPI37bVihg4lxZgvZzTiR1gZ0pVTeyirFji9Sh0hC/uKgEtBFGnqaPVESbYuUVYT9TdgkGoYsHRc
retHFJmL1Xki98h7F0LTGnxZUdWm+NyCfEChxqgYKzsg4O/Eb+8GcvXe3UdduxEtryQ+nVr+Mus4
22zCeirOnoix+5mEvFry7tOXLO6gQlw3orvwQ054kL3C+Z5Fw1lE3wyPRDnDgZWB/9Xkq/sDL+ZJ
v3m7I8K9O9T5BHXNludciQSvQj5VzZ7S6epN8vxwRuhnwnaGpYbmAdvGw0ACUbc3yRgajyS36T/+
K0euwCZcgIBd5/zY+tZf/m8kcLW/qNCV5FU8/j7ugRduB1ErZUFALJekmf1pzZRMRFonCOZTDNmT
//pcjlrKcTzVA44uBZ+zr3vj5SznAF3wUFt90ZoYjVMu/rcjxrSgYaPFGWM1syHbjdsLUSxl4Yju
n/gfSH2Har0htarATwmDz3Jjtgzx5Nac4QToyryWTRqcmyYUoJnCmiSCf7yuQPpAXPtbr6muqiB6
WhyULNVo/aSwCePntNJKUeO5cqFyWnnxhqNEn43JfTgjcpupWGquVo/gncPBkr9LPcSCRgth9jXz
V4souZPwtTHYTPXKGr+wEE3qfBByRdnvZqt1ArquNwx9yChB8qyar3a1MoAAExTYBw+dKsUzla+o
wFrM19NoPlnPmcvtYTTG3jzgoY4dr2cWrDOYNlYaGT+dfUt1cT8J7fEocvSkcAThF6f0vi12SexU
e1ybB17h/j3KZkUTWBBVZT+ATjdVmVzzVp57tFaTAplRsqDbBlxa0ywJ9NtAnlrlxrsiWkbgPXPK
sAPDa14qR/630KqXawa6tQHQIhkspYRh5ejE0Xqa2n0hNnebO1qJqkKsofuuRWXS2tTo44IvUKaO
ntAqBucZN4WD5Il7dIULYQUxaTwcA7d2yrUCK17Hdv4wCKd31BlTsnNlxIWWWWbA1mmo36wmxJ+c
Qso2f/WHJsz91re+sgFb/6ypIXfSy1z//qH+USYXEiSlR8PdnWPCmeJEEyj/qiADd5fbC228VBY1
l8T12e28d/B4xhOper9NpoFHHRuieM9Y3FUPfndthrBONTU9k/PNjlKJ5+WiGj0mRBNwuSAFVjeO
bnFlvLMMY3oz/lCfZ+I9QLpTdEfHcr1voTiRf7Dun6sAtK38Zl5+7wcZsXFem+FPHZ7oM5SMEVHc
gQhMGJZxZJNTCHkiunLFYChRhtY+mD/VbfuLKH2C+8p5s/V8ZTlIsqMg0jegmuUVb2b2oCVd/0Dw
L5kpA2vwqQUAh6NtN520IT61Kpwsw8E8vmXQknEp2GlTGjoSixwfR9CCRMQFdiZdYPpRoK5reG2v
FYt58wKO/KRou8JGI+m5EER4G10Vdz0M56r4rPTQtMKrYJMEFIJH+OKsODtwQeputNEADtvSSoYg
li4c53pQ+AzGz2Xr9z0muBiLo4J8K1TCp02sLjR+G6eNXuLtjSMwV75IdTKyCLiq+j33o1D000ID
DkQNL+HnUuKYr3UlAZlSX0PphcTpKwg/IQnuXR2AhsWSOzpYqzYrHRnsVDnXR7sx+kAtYnPrAq0l
F2tfDUZTqcINSwINhrN7AyQbZWSHr80XCiW+aLMSoMTpdlMjAPpdcj2+hdmvbzAbkAVD0udBzYbg
K6kjC2g4psWqoSJzR3V3i0e3OrlqCKVW9NCsU/MKR3ePXOYTJ6Kjkpc/zjfBMd4b0h+xBgKPtAJF
L4aDrF9eaUtPT2GcNosAL6J6u0nxY+uIcd5R37HN5kBbidviG9CFCQQM9g4tbJEPAoOzECfZ8uWC
Aj5jNl83cTGY99LCFBs8/irnJYgEVb4r3y6Vfq6b6SPr/XGLE4UU9Eevexf/U0ABXkQljYfjk5M6
opmiZIeS07Y99AKh6+OK2ykRzj+YfK1718aEU7Y44yPY/Afo72ZdB6d30ftin6OkJm6P8cWus7OC
5Hl208wPZCgsapNzGFoyTyB5p3gukbc65hNubc5FcKly/tZba+VbTgZnygo2zS08IrueOnXa5Glg
tN+9GDuYZkM38QJL8u7iUjtBrlPwgoAkEVBuEVOrL17ioOxqEjy+NUdqpLsi6I2l8oIcFyaytLZ6
fzpYdEcB9UU1K3vbX8BUhB8scuxT9EmEiy7DvjKTzkY=
`protect end_protected
