`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14912)
`protect data_block
fP0vjVThPFkV/wr6hPmhJhjvK2cg+0y8pB9k3dqz+f7ivPr+FIn6IK1VraibW+cyumzrf14UBBgV
lxTvW5k4Q6W3xcWRCut5lUVvUIUOKlcy1VkZrczcmN/yDuLhptEdKE4wTJVcydnA17lxv4dY7pwf
ydaAFQx6ssTGRejEicOMrisl4amIkesqAm6W6oPMTg7yJghnA/vjNamy/A8wg8wiPNkzacMvUiDc
wFjAiQ7hWP5hGRE8UxZzUM+vbrO/FBWqstVdLQ1XqdksF2CKF/zuOgawSWhHcPG5Iy1uaLpnOhNn
IQRhiMmliqZmBPXSzt6Fepkm8hjFI8Ax0b/edtqzRXxm72hTT94aCcR4snDyOPp6G8P1FA+DKi2W
l9JsRsHUrINiMrG0mJ3CcumEJm6MSrxfX+dtpxDmvJZ9FaACamTcgdC8tvdt236hsfMDbKjTotjI
7kWus5LYdB4TgJXsEywaEfsKrF//NBZui+1qKQatpgvSqyqJRTRqau668oCLqK3a1zO9FYWRZA52
zCbCJV7p9VxEIxBx/yU9JsEaDKUSz9h3bm9vK9xeTQ3H1iizXvoOaFpKnsuAqtzXB8GiuDqVOZIc
5ivQaap+8FLnvinkrD2CYY7Tn4cM6jF7aFe0mvFTtgciZ5jeux1Uu58Y6OKajEkGavA6m7MUxERA
UV6CwHMrjJQo9iRwabsPN2UiffbmMRqvhu8aAHdC+tTfa8NMadsZIYXB8XOAss3mXaP26ar6T/mH
3uaHV9c0Wcj4dPlL4lULnA6wOgZnXkMTomyzGUttz4zs/qQtxx/3+78riiBBuvueatjsbjEDcJY9
H8sMQ9Ah0+M1XMbolZr2m1W7zO9MsoN1IAPXiEnB+On9dyppQs3YJil/G98IOEuPprdI6j7CrFTF
NTUwK5FZS2PE0G/PtJfwOL+2PIRn0fgm1/A+xoGWQt5qkR+1BAXJR/bgIBZUGPCt/Bw7xQISKkmq
zSZXD31/OGgNa9LJUc0b9f6LQET0W8X9wtq3lOOLvaQS3yGeGu+HYusSEJxiJjODxaICPpYXYw7s
tdGiMX2zMGy6ibjFftrktkfyqUMWRa9hgCuP0CNn23eyYjXufdjnd4FKJyZTPhw++M3KaNoS2a0d
MRudASDrF+dtYsZqjaeMNbyI3C8sOI7F1omKqcec76svKGIVhYAhFC6DTZmhbVOU5QBLBBsiy7Me
2QaETAvltqF4QFhI/uPxOVsdZpPKZOIEiIEWAxiMjLPxGhEwz8RH4uHvEmQsF12df9mJmaFV3Rtw
JqByadgYoaQqK8SPGrUZGo7jUk4BL+cKu/DlnqRQavh/DSEVg9WTb9J9GkwigkCvP5RHvGyc2mEm
g509eszuMiQQgLU3hxjkyOz2Vrpzkyq/ZKx6J3+5J/QSMxiNdZv8JylwU6H3OdfJxSubQlh561gJ
nTTyeYu0q7MYSxQjkRBGbaO0jf34bOiJHTpwDhVrnA0fqfglGtcbEoCwFNCH/X+qabaR225uKsZu
jscvblhGVp64cg6ukhiAtTKpj/MpK3EalTzW61P+tMpBg+m6JHONEaOYzov27etD1FnSP5R7stN4
kor6+r/2gkqi16cL0Pwy1S/Yk3eZQtRmbi3jv4qO2O5tloFDjKH0zLVrxhirFb6oi+Ng4klVBbDE
XsYnubKU0lRMzltyJSPx452V3UBCyKomZpxfuc4n4HfcgIGSxDkBccJZpSTy2dL+TRoOBhkxJuN6
UAO2ALFKLwnzaNmiU0pe3LiRep5L2PKM5MOI4+J/yjyOJOhiCDP2LmbINcVmdVck5h8MT2mCSwAg
5Qk9U/2A9ncwdUj50biacp9t1Ko4Rqwr8vNj/1UxiiBgVlHQIwb96+29tQSYRtmHZmEwtYPwDaja
/mFVV/8sXFepWQ4nuxa/u3U2q/kiej7zzou/VdukUZHjQ4QtrOLJB+VUkq/zacuy+3AO4GSQMHdM
jKoXGp6BT+d8cDwvFFMmEDEJIUQ19DDUpvCx/7dNBB3TJiY83tV5pOVDvOqko9FOmrMI2itjWzJS
Bv1/ZvOZH7SGOwkj9/UTWadTnChAMTNezlpgk8bC1eNcUI9Od1KCXwMacCsMOfNktEd+5nFAiurz
SDom4dVmVdP8gQ4lNjYI8xKCkL4BR0moH4meoDuQkKBMj3L8Q4uzyQgeLBlgZ3xSgFEb5Vm5SzvF
0L0/7Wv11tN7fOPFCct88CEQbSDNZI0b2EeLTrqy+EwQCbJjg9LSLOLMaUbozBaVJUMznqdPoQcF
bhKP4E1K2ThuRX899VadgY1IznYYVd8XKTSMqSCD7ye9YMTNZV0nhjoHxDClgoXy1BiSpNwyjLFV
kqZgekh1UfTTTAqKiolXLu/th0hD+Du3StkSQZUdGeEdrCRCMMfnoRTl1eDIW+PW5Yn/U0QY0wkS
UgofvYFdRak4E6pi3f1wTH7D52NS0K1o+ykWsV9BeMcZbkmgysSav6Xu6h9cB9T9mHgN4LNdcXMz
jy0WKtHdDjepQv+Vrgxr9otSPnEqSQ3lhY/v6Wg6IFNxMWEqDuzRvyKZ7NfLh/RBsuJvA10ciZ8m
mQ/0C38XsTcHd+0qWt2qjx/i7+pfz5FSQRXxIVonoa6WW3295FCSYVsOnSyMy+ZfKOjMSNUXl+tf
v4XNc4GKUOPY6hFHIRuu7X64qW61uBl2IkCHYPVtGPcYJzrFMkBffc+JCKet8+rf4RO8l6C+2lQ5
oM8kuKnejZ/J+kBfFIkrHXYI3LuX4OTML5c06f8jjV5wmhr16HofU3vGUqIxTMTB14Y98cbtEBNz
pdhTV5zu0xg7l8qzxwi/N2iCeTCxZ+50jUDPRe9JHXdFpAbsn6Gv0hvu7c4uWnIRmCbYv5QtQxiu
4DeDEHpexiSBuizfYhx5Z/C9OidPsVjMfBBzTgSoKDKv3mimBLoOLKniiNfoFPnW8s5Lm50h5tab
5LJKRwivaBBqK8Re4HoomSHFKCVoZ1uGLKe0KzAY+TdotKBoJPDJK/qToOfmC1OOAe4B3UcZ9E7y
VI2YAK2i3I0uiDhvHXe4rtz5BX1hD7MLBO4IXjLJzyMSdx6pTraLkeoHgPPkK9BfPFjZ/eBtCRej
INBORfbv2vRembT3U3Oj4LpWSHKScttgfpLFy6x8igPFvVy1VN4nBI2Xar9ngfBOdKSdoULL6+Ws
37UZmkI0P+nIiQo4Heh5G9UMDCnNCMm3ADolepQNO10DM0vD7o4Xawa1vl4smvgNX+mXhS6wQHPf
ZjuFXoSjpVWYgCRe0K7n2oSiSYv5z6EQEjhsqSMPADDjGo2s5Gf4dzGRx/Iuq1c7jHsGZe8q0sE/
gFtSqljC7r+GsIhWQU1a2NO43p7h80Wuli3bb03MIURwb9AqKlM9VWUEytH4NLQ7gbFvGeXG5Pgx
9UujMLKCMfCcht6eXgbvyB6UY9GjqoC4jgltgOfQqRuGewDfR3wxJSAM3qy2RZ3brRHmC8P71Vj4
FgRuqiGUKHADgRGZeMlH2z09w47xs9YR8Jz4ddwO8OQKg0BuMhaTAcT3v6hfVFTIAQRG2TqjY6yU
j4oCpbhzKIRjbY+aEoGpx3cG64sSY7evMs+UkR7FGdDVJpRGyxdZRXVlIC4NsQOQJfor9q2GFwJ/
9h9vyXEgJv/gS9XSYSK/QLOb4H8sXlLaeor6YmWuZ+EONplpLAuy3nHAtuOmimSHxBmDWM8stQkT
jIypvj5Ot0TD6geJJSzT+4G6MgazZJq/IvkXUVB8WJkZw5GRD9pnw2XwtrZmMrQEmz5g1DX7hpKA
vmeGGnB/hJ0138ipKLKoZpohVet5OF54e+HaEEMa0JqSICAao6ijwom1AO+dZOkg0LBwwXZlJ4Fg
GJNyu1kfTMmsVZwuF2/3Ec61T9TBgAihiVXN/ohfwSeOr73QSjLmr9mO9FtuAMlGCbfWSsTrK5lF
k9Ra58bh/Qr7VJNNF50wd/kT04g5hCJjJ26N+GQKUHVC0ZRk6gBU+rpwT+RhxJEd3/UvGcKep21H
qRi69DfJz3/Ys6SQ9sDAY8vNHPdEd8AtF8Jm0ED6nJ77ihSUnUxFGAOFNAwD0d9vgzrmkidJTe2q
HpOPCa1yrIJAqP8cdqlGeqA1DaQGx0czS1/5pOZ1NEAqwvoXq56ZIQH76KWOLngaHLR/4v2AeTgU
9SMdR9bHBAbXU5dDHDQ7/m2BZOSjcc/fJBoNcJdqRzB+IJlCFL/jXk4t7mIk67lgKhnFfLV0sLJw
nb1no6Dtkv86y7b6S5bF8G/V2/uYUdxKtQ8F+rOxvph87hbYNERBRWJGQF7OqT7RQjjGCg1UvaLx
LSOaBQo1lCsYSRsJ+gfqzoEmR6DxKY507gBnD/LX+Cl7shi/NtFSCdC6AXMLoJmKYtAJPeBdd33Q
VOh4dhdeI8c7GGv4PXuOgVTejC9JlBcr+89gpslSXcmuYKBeVJcaMVVD9W+GooS8P325sTX1L/Tg
zeTuGHLLaWdQp2LPzo4LiNwoknmFHxOIj3LQkvoV4/NfGrSfKO7YifutDlsfsf/GQFA4GHloCR67
On866++AVPdWMZ8La9xf+Zg0QtmTX6ul59xPTw0Ywu2zuN+Ui773LLicVd7cDGO59yAKFzQtCTHg
nxB4wVsVv12SCUMRkKrtsLA05ZmGxccHe49iupH7jvAs4UZlFUMey11DzDElEDXvsngSLMw7xI16
f9O4BJ1UteFDuGEfsZekIBVGnBFIyenQlVVIF3hYVyAVX+/2TT+31d196dOhBZHTqTP+mWtBIfHi
hHRTqPZ1meQ9VowyaO+xBtnOrbwBfdXpK6M0CRJ0yJiMCw945Squ+27OZhQ2n1wkZhydZNKvcVM8
pk3WxAo5IZaTfxFWjdx/zG9N4F/bCH5hhEnLTcelR/tqs1cgxf9GomSoTv403wY3RIUEUYgpeemJ
MF4Q4DWCoqZszufQDndGmT1V9uMOl7D2cqaFSk0LNt5ASh7oYr8CUHlQMAu10BbxPcVxaVW41fyI
OxZXEvoSRW9+RpEGkRwhlFAfAZJ73Yeo3NaKYjCTD5Pd96lTgfKTgiwGZn8tyU1JhT4smkvzkpAS
rnGc1kdNLQ7NqlM7Qrsc2Bn73xnyPl+/9AyudZM3F4lvDVrb27dji5uubxJhq/1T9g74W2j6oH0/
cSERleZrtWyEVdkdr5JiDqCbIynApmWV+VDjyt5tQnDgZoxNRXeD6FmUeky7vW/FFk+OAaExaG10
cSMYSBJ7VRkpc/FDTU9FnsbneB99xyQLjlQ90WNqhAs+VplAqhLVfEwiL92MQmKIRTgo6mZ9XPNa
lASnVchdP1LrPgSIIVBzGEEbLrZ8XETUVbn6lBuq7sPeZ4/dlNuUqTLP1RmKdK71LnB+8fbQCFhE
1ZeAKlwhd2IiZEXc+SF9oDA05FBAWEQ5LaBZeDx28sDmWEO5iRlYVyYEvaAKBUa3JgJA9aZV4EIo
Cn3Vy8zNLRNr0hFCG/kjvo5b0F7P1tk/HT37Oceyy6KtoRGnLM4mjo0d4R6gcs8A37pvxogmyjIe
GBtF2h0awViYL1jU69VobJZHhZd+hGO4A0fuFhk16QpP6rwt7/ug5oTRwh1l6w8NXFIDuI2t5eBb
uTprQVM/HMIJagzZNp9FJefRu6o2t1sE5VAELORqyfPjZlXm8dS7nx9hOWP2sNvLI6fsXunuYXmB
SJSpIY0ApQdXRO5MQDe0Mv/zO0C2UbK61So7T+hTk4umiQb/T8AxpIzTFp5BiyMezijUvXU4qaTq
jeM81FZI4Fc0kyk7CUoJQn7e9/AytszIIbcrgxJUh7umFZlaP8zXCQmW71eEtk6xiqN8HSd8J7TY
PT/UamqmB2xOmi3m9rxcbRwGgT82WJc73HHztJCjlJzB0Rn3zH7hYwNKzNyUoGiveQH4W92+SDrZ
QNRiwEfNsjpvBydfcO/qSQwhc350sjuysll0C5GRJYK+CA7OzQzCc+U3x53UacDitfZ0hre6ia+Q
8/lDlYve8rx6GUMlP9Zg/LvFklL4e+21sqNjHPMjek5Uoeh5N3cuENTImB70Ehcw2fEoyeXJIvXu
PWeEDrzeIj3rwvfIF7F8lqyTBlqr0bdyZT+upeN5S65gcY4VwG71hJPQ8O5WkrGjKXF2+apzu0Qb
O5Wz3s4YtDahUQSRPoYpGkCLtkD0hr33lgnrCxezP3z6nFZMhlyboh/Fo8gA1r7YWVXqmuLlqRms
V0x+j78ykKzp9HVc6ICAmBPyUbK0BlKuNU4huYOxpss2E/oJLjAK08WjVvy4pI1X6idGvQC7r9nE
NCULvNHF2/BCCzqBYpg60ROSBM/VXG+JN/gYs4673luCmGJ35Tch+WMoe/hNYkLnDgJHcyaS1+rD
9PRzMNqyEk0NvAwePSsYnoESFj//S2FgBtxiQYsCb6C8/Z8Bmdcas0e8Z6Bgbf1yuGqSEBTGOLDU
iA0vCV4m30mnCfA+lcojSa2rabuGZMyz8suCqt/+jWuZebdjKvILsK97Dtw13HjjOMAMX4j1oPBs
Z6Nb7cjvvBShANedMNc5wgme/Vu7dS/0qP3PSvjyEuVwhsZc4xpHYngVltL5GPT5REVtwzF2tS99
xx9bpncOoKcppXmBRN4PyVL8MHU+GY6VQuOmCJ1G+Djd6FhIEHnarrikCfTO0d/n99GKvp7RI8PU
XMxEWldtdpUOtbs+AxWwYQmKoO3UOaSmRP6O9EaHvq9+FnsY8brWNCVpj4qEygKP9ifCGNu6bC9d
gVhTRmo6ZRFDRCqWad1lrt2Fl6Is6I5jN4+mtIENbWVJhK0DbRZJ3+FMNJYovFfarCHlj7Y7I1V/
1VA7nNh/ye/5vQquD3sjKchXQKvfpuz0H7L6N7xdOrqB+dIi1+FR8sA7IxKrsXmDCYXF19ZQD8FN
kwcmY7TDIAxAnXN/Rfd7b7ApRqKFtrCVoNX3/8ztk7PB4wCy2mzua+o/9d5qtBMjD/D3t6bfG18O
f0iAfoG192NqYkj7zK7buoJk0ZRQvP3n3n1VTVDjlAQM1gJjUASor9aHDDO4TOklenislqYJyOjI
1Ni0jWCUjBhHc838T4rpJbmm7yEf1li2BDVfwKdTOEWjB6w3yrXqdDrEDfVdgeLcGvq7KlIgXdiI
dHyB5+1vmVfco0MoK8DjAwZ0jvz8jLLGpoBjucJnnp/Pc2vUyUERlI5LYL6iCgCdi2BwQOMw7DHm
qxHn9ULALXH379w8NbI21+p62mSh3ZYx+YDfPM+8uPCvt+pRdv3JMSc+7XU3BSp/bOO5i1d3jAzs
TG2mc5lpCcYjtDPydyHZQaxb/smwZW3/3rjLSFF7ZUaEvYb/LZ8eWT2orL3bNOfWWLBM2i94uybA
9k1C0Z4IRGAJLYxbA5p97nVIfeDelJ82kps781s23QlWBIrxg16KpXqZxdj7z447xDIWrWyyiFwl
+Wyla6BGy9uYPhBvbjMbXwGZJV8YnQt4ieMx4iUmMbE0M0Js9WSxTMDmyaq9uZLZuShN6CwxH/5W
vTgTH6nejAeyI+uL+db/ANb20IZimFSDG13U53PaM5FqzzDKczc2qe2uHpHx+/hNm0GaHBtfkn4j
lOIvJ2PGOSPYRwH0MUcUbdwpq/tJH3J2UCv/ObAGQjxWj2WU6EK2xb/xyrun+N8E3nc0kbxszI9w
UZx4ZbNw+QL64OvvYp+558TtzsVyl0+6x5w2ZG+gt4QGNtUk07Tv2hWv12rryIvDqkEXMSUMdANq
vPwYx655qjwm9T93gG1nup4EoXeBL7JoGyn7qPSg0B64UwBTY35Ph6MdNTDh/6mnseG3kT9nDGg4
dldHM+sA1dnvU/hd0PROGoVz9Z0MAorRcK6+enxmOM6FBfnYby0rPEzIa9Y41Hz/RPBcbpRbl62n
88xbJP5l32LPH5bnAmAKWuEfxuNVQuabqaHcAsuu2xYjxwoRGq8rQX72j3SwYy6BDwOhLgJyk7st
PPT3ft7jQw+/uMRrecehaev5weRcS+0hc1u10UZ644UoyURU33eoY6rJJ0IUbEpvNEqGR26y+hyh
B1wnNQp7801zuA4w73eGa1J/zA6AXWAgsFlf+nhO0PRUp++wudhz8X9qQhBWuHlwbJe+9F2cMA3U
5YPRC4vO1Ozsm4Py3akpc4m6MeQjwg8NwlVkBhmTeJNJN6lGxq/2in025J4o1legpvo+Fmq3VoEB
8/WD6IXdHNc06UjB2/K4embJVDKDCc6YO5UmA4nybYLhEVYReH+sp3m///lmn/KWra6Mcm5Ja0Sa
b8remJTyfKwKdLnA19NEUeA5dAz8YMn5EsswmqSJMmF1mDrU7dLw8r6SFD3G0UFQAaZQWZXrjPQP
CNTJ+spME76UrkihS0+Bm7zjD6dOVNmK6A0zokH3XDv/68FgXz66fVLj6EpKnBlnZzP8NDCHdp1T
jNWuk6yeb62d9NDVQKV6ucIqD9Mo7l51nX39wyKWgdGUlx8gIXdjkJpD6BJNYXUhyhX0sj8Hv2dZ
VZBdXf26+pLS57vpGD/f9j2sgItyVEixPvDrXfva/KmOY7DDreweruQg84XRezEk4T0URoMF1WUn
O1KN7Bvbu0jOndRBEOjOs6nKOo5L6eCydPxPsFKWlsCcDzc9aO9kUfNXi4eOAyi+C9sXKP8GS1TK
di6vj1JPyne22EqDo8Dvrf6OwN6BqUuNuTtrxL0r2XY8iPJZg9vi1W8waPiOO4QryQhKunfcaVEK
vQUr2UXRnkyHMkyju2d9sr8NZXEoQqWdRJWlndESy6mK0aI7Lrp3WhnjPk2xituQrPfREvtJaGVd
ZpBbsUWCImbO7jkta/1aonTCZxEsNs0FedmqI4V8uwrrGP61NnHp9CLxy8e1jrUKBJObAvIGYJLi
Vb4muCF0ojiF9GgQdb5Ko9y7SMiT29eduGLMsSUKi0ho9fhpCjtiyzcMOiy95T/V/xnQOsObne/W
zZAflRinQJr0h6Fw/4Mu0JbvjgQSaa7G4h0PgQtdldwVcf55afFp6gpYPUazNhq2tGfKllwm6El4
cNlIwjU/6QOgdbXVOftGc9qKCBhITF8/l11fc6uiD5l9C4sw9doU7ft+h9HtdQcmJievtUNfT7js
1hl5lSF/nZ13Q36W5SLkFDh5cmgKSDSXri3UyEbZF44yiL7KWeefnLejnnDMmhPR3zc1hQI01JXj
muUKG5Ja7bB7cX3+YCmEVL4JLVAPQxqCeneCXarlU1M5r1cFJl+XWJ8Y0BX6jo72Z8+3ZwA+FZ2J
M0P4fCgOC0R4OPpjQg1/t5xAZ/faJ6+6uQ3waeKBsVl8Bagz0T6EdkPQGeWjBo7ExchSsoUFH63d
Lo9juweXmrm2l6fKIuR1optkHI92Q1qMeoB/6T2pl/cj8A/m93gNDvmhrP0pzQF/flVmAk3JBlpQ
1Vfael1NeVZ/O1KMKuTryeoVecBMShHgdGlIwObS/hcT3p0IH3On5eqyPtRA54vBAlyKSP/kb78m
o1/cMapBzUyjiw4yn7CvDBiIAUR0DmTziZkpbBuhqF/xCr/eRLsictlKWLj+IrmFxqJifyIeowSQ
++U6cAJ5ThNv7Nu0xNf9NYDQhIs0v737FWoTXy++TfjFcqFJN/F7qRxo+j+Fc57GA4st7JsfiyJz
mfNqY1xitwE4bfl0PR8GvNU7sMp70Sywm/Gs8bxoiLalMzKjWQKJCg1bEH2rWyZOpna8r8idR3bX
oOPszMQuZ9f6Cn7thvUsjzdSz+3HWCeE41Ok6EhW0WuFFffosYyaLSpPphbmbKs1OCibH0sPJqzL
aS8dYRFncLdPqzNYqPcuaET+rxaODBQyWUMuWaa9ktv2pPalb60/9d/G2vsx9yDX3kxyQ/xg1Kit
enbyvktCwELdiGIbCcQ9ls6yC0WBk8CNAXOHeSJVskivxMbD2Nrnu62qXzzCxUsit7YtstkiGzab
Q1juedMa39qB1W78/pSRcBIXqqazFY7lwQA69+j2x1a4Zmybx2dWR4KO0v2BRKHusBgrLYOK0Hdr
l6HPWDaJ7k3M3XAUiYoe9FLt4FTl9yLGPoTtZr2pfcLgkaiPuoNioDQS8CLuF3g3bcElD54CECkK
FccsG0Cq2/QEITNyOKmvS7G/uP+jP6iMQhbMCvElZlGzMyvpWN6NVAw2DFcam8xnXrtOCorhwOfR
76+TysULLwdSeg7l71lkPeHrWFGgzTEOahxNfKvHrs2l9X75qnkarVWAulVk3zHnbrwunNz3rccw
CPmjdf7irgGSE9lgUvS3MUekYMkXcGNXdoosphVVGbd+2sjFG/1vIjvMKceVQHUrpRP9tkd6teSN
Sd4lGS7BfxNJC674Fecm4aaWaRHReGqrkXVO/3XYh4VQXyjENdIDJCo5vdlKV9EwRzogfeBF5ZNl
8sz2HaEzHib9XKbTcLX3cuBhClS6oEx8ECuYlpWkzmxDnN1JIlfEwUob8f0fCir31g1Rcfn7rrh3
AwJu8HMRUq/0K+kIG7ZyWUmZIw2oayHHtQndk+eIX8I4H/I633fw1Mx0KEGDaiIXqWcK5lwyos8N
ebV5i2/IZNdbHAzHIXiIR81ikQygBU8iQeUrT+CMky74QaHh41SCB63cAE2uj1vygF1476cv9Zhf
8c8Po7tY96UgLbjvHuzcXeyxFC96sz3WvZrAUslldGaILk9VPZoTXwIQET8wk2pPV3QbDgmVlTGI
YlyNdHen8C8cKE5h6Ez80J/uvz66b/hddvUzYAyg1lGMe1HJSN/cZPmTSbX7ltFYXEmd7eCoWBPi
IVb1ewhUip8WHjk8DSQC0ZyO6K1zbTzFNRd5CtjzGUdiowAoLfgwv+vq95FbKEa79ePNEDP7xkxE
j5XT0k3Y5pw5VL3LMJVa+9oVkd/xh3pCwYaUUsMZKwConU8pY2e8sHSVWTKRJWvvMbP2xnYM42pW
gIKXPmw8Kx17xLNsoB/JDX62Qh5GilmhC7nPKAfJtc8ZgTfCdcHWjpmqdkrwqKgQhjDXF/0BXd9k
XtpjNpNh912ROhzZppsUh8zQmn4Ml7ZWUqF1NCqYEbASudA4eD/Xq1eCz1vD1N1O5Z8DqFEvugcr
kBU3QO4MRPmxmB1ciBmHSELuGe2HgN/EbbYv8qad3WmsnMOIlX459+krsre6Y3nkSdqTpMyO1Gy4
s/JYej0p20X7J47oC5adPdaw2KxfCg4evgHwNQwE5BrXrwSwz02SNLpKZ2LZKQnrtwldkR3kRKUI
MHO+R+6geOEQa6R0vDeDS4qbTPwYXOk9qVsvB1vUii6jEgYcZSY1K3GoWVNkMUgVax4CBtzrJICY
YPYuvjR+agiFYPJ91g3LPWRkgN2Pk+Y+fcOZpoynn1L8vBxxlIFTp59nTX6fIe4QYcFGoX1pm+2d
Gnpz4WivzyQwWGWgfeUgiGKEkLQooX3K6SIwHEQUdAbhFIsGy2XVkZOQ54zYwjpi7LRNLYx4VG4L
AZ2LY+TpyMluUpFSvMnmCxpVnmNlVRBM8iKsah5CeiyOH/abXJ4vtfCMP6OHBuwXh/1TJt9LCxiT
mLfzd9QW3qRYLA9nOOscO5g8EpzzdR2cE1L6DbVRAj2K5vBBMdfqhDQnMApOnIeJy+Fm5F0fFVXj
avpuX8ywT6er6PUdwNuSNs3pJH13oZ5zLqd3TesiUvaKg2OhrOrJKnmTMeLjYNcizSRyTTcurNep
jkWgitsMHgqwbDjtgdhatNB9MmZm7v54AJYNe/ztGTT23D2VygRh1e8m4eiChuNR7/ESdtkoZgET
vCxTXv1wMwMJgKNZpYoJUR/e3bx3lvFDw025i5fv9+BIL18Tbp31ymvEzL3NBjbX2rw+JnylpAr/
dNRv4pTosen7FRFYwn8wABf+8b7ahBngd7VbjHskFIbq3qBp0NQEEECMmp6AcZJ9VtKQ3iiYOT2W
TKzX1ARS7VcQJbvwT+627ut9RKRE83KlvfAmJnXJ9z4a33M/23Wd5fQUUDZ9NQysw9BBSFaaRsal
XKVS65yC3r0g0Duvwtr4w7PYvCqy9zHzpTv2X86IbZcxjZQNwfcq1dNfVmh9GYDkBKWgmakP2WDD
++Zsjv/YN5+nb9cCVII9KR2ZbPtCDzCm70WsFvo3r3WyaoiERLwlQaKiQYAE4QA81/I5zN4jocqR
XivEX6RWNg7mMZneMk4wupn78As559HrzRcddhrQb6/okvep9L00z1n7TjZFCmCpvedQ/s4OZumG
A6iH2lxjmlBAItS3ys1rwDNtuGiEW1dy5tLOXi7ywFrkGA5KSWbxjtbeuJJ+3+9MFX67+ei961OL
D3nS5rumTUoqnfeTIYe0h7XeEo7JQAg9mRIp2qeh8Ym8bArvEkQK+jOTUxAixp4ZfT0yd7xhKvym
EUTRR72Vf/4wh+6M6VQbas32SvSwUcBQhyi6VrRM3ikiQ8X+8UReEJnytyDssP+5odXxlfdu3TR0
K9QQBIcU5ur74DaRK8Asx69IJ7DnhyndtA0hBBUZcUVBnUlQ5PUGvTsIdTNZYtBZbZVRUI5Ud85F
2iy5MxxO3i9NzYficOpTGtltNpP498XirFB7541v6WCEEJWp29IwXb/diZWFqT7uF1eOk7Iniylo
WaaA2rTYf0OdmH8uckYUuX9r4UmDfMgDJKJ8bKJfLaoXH3O0X1bctZVvkK5HezEky6MU0mdeHTXh
0ogspaVEH5m0movo2Hlpmlz4FrgWr21uDH5kJx7zLqPXmYAnM6UucrQxzAjUT7borSfUN/meg2Lt
X+7D9Qi1iuastLwTjZBeTd9oZvHAR8UFBg4NQv5a1/mhc52d6KjGcYfUzRh5gngyNsSVKpnNjG5o
nCcg3M8MOMrzNTFaaxeYWWtzrQ3JEmIAtbj7gnzvK4ryUcVIodyO/Ee62UkyEOWXhiUZpzBJ6Arp
1+idwc7btiucBlWd/sKPP+iT3xNbnR2CBeq1wxw4Tnv1Ca/I2Nl80q7Wi88P4ETF8BHDWJQGdHKL
JWv0DBta/Bxxl+Qy34gVmpuL28jZS8e1S8edbRF4Axe+cJprPku2UWqaO2M2mhwFjXXn0NLET5aN
3nm3eMYQhMGfxti2sWCdGkQWXhgKpJ3Hmyff3uSq7wN11pE7AmWh4C5PblmpPvqv3GOCIFpQWIQM
0fkYTC5aj2Naddg4s0Vc36HQBS4fodNdovAKKRbJ4iRyE40GXg4m4jEQriF5oT41o0O4wvhT1j1t
tewIoWDYjJ66q0FZACJaY2bL1qGBevtgqCpIg7xLqGNhQiFMbU4JPfqfYQKPD1EsY2tcJ2klqjv1
hXw6xPW5nlhhFriJAtpZ7RY5sR5Q14FqczKULYq95rxJDZG2U0w8Qt4E7R2WlbwB18M4qlX7Bdyc
20UCJEOLH8R1GJcGP7V1n02coamtRzWJ1Q7ve/LOBNp3KCWUUKgdRB2wfRRhIQoG7wVP6LgzQWDx
i3NHug/I2ScGAS0cRWcdIbRg8cbVSUbI9+iMmux2Ks+Hep3QopcpZ8wMxCVtdUKQDV+0vwpLLZSY
TMWjtTMIx2hv0PD6aa4pU1RIEysw9Al30PYQUd45GPEHNedQLonO2L9jJnXK7gBFgxjXsTyDKKC/
3c9i/oxb7wnVNNltq/nH1UgoWmd2DZRvUtpEij7X/UpLEdX6xGznO1bq4y/ivvHfIAo85MCW392p
yRiBV4BozkY1pcOkg0uB+1Xs0H/jBbyZpFFyuOCNKExh6vTwSSHtqFPU+ylSjk7idvsOWmuCTfwO
eR0BoNS8GFKNfjQ93d7WSRkLjFHzggC7nZQTnoO9rVENPEFQerLDAR8TMY6JE0vTa2zum12Ki32+
PRS+978Ayjpkqvd0fpfakQ3vTfqysb+UHut5fL9W7uD1oGCBMKA1GbnTzHJ2jZRSSB9OiJ+VNK3f
mJkKgHE1fEumwP4FpDYgljMFad/Ixg/Q+LZAHjsH5WyVF2tBgmsKiB9Y2Py7CtUmuiA4vY+sNHz6
ON9WQIipgqWl9n3Ploka3acBoXmDsZINKkkhUNKQiUizbK2JVhjonPMSXswO4MAtCAsRgDkdeZnt
0pGGJfX81oxLTBUqiJrFyWrytAa35guBZ94NfC0GBlfUIqZJoKJPL8V8zc6+ya7SP3qkRUc/hBxc
ChsnsAQLeWkvLbub8Lpej3NtSbO0rQ+SfempOUpJKVLTSy83kOipWgNwhNyWeJlfmIAp+Io3g8is
846LyG3HkYwb+Ugt7SEF/aUVpnuKmxIU2YPBxDI5kvy3Sxpaix+Iz+32Qf4fUwmROd1YE0LiXOxq
l4CdztBBRJnJu+ymOwtgYKZCV9vRUlPLV6TaundkhAke7tGsDSVGvm8eQSiTkiQshwhRt/Aq+OLU
QvKRThySfKxx0mn9U36pI0eJJwJsNHLS0dBEy7JYDNtLbIpepQx0TPQX7JW6vAkgodNNVxk+RyeW
Y6ms1GvzQM3nCL0z76YvztRxu3sSGrWby+hkkcQkFwJZUpCyseq/10dpvjMwoIj7btlYaY2C+xk1
jV1DHHkzjlg3VxI1T1oU1Gk0mD3/t/49F7XOVB352oX360PImU56ky/JSvmAUMjutzBInQVOWJas
6fV3Q3OhV+xHAgaY5ZUQxU4FE7POvirBcck16gdLHCfO/G78sz7lfr9Wgikhja+67SriqCLKO302
Hhti44JCEq1APSgisoAica7yRzIwHjj2xQGs3X2TxETv9Ezit64hROdMX+K4KAJ/iCYz7k+OuHQ6
EVzfJXhAFjTbi2vggBywwmeYT/NwgK2VtPJWlV9ZyoUJHFuvDKioZNDqyLoD6z43lv9y6NNAugYF
3agpKDmDwwsKxJ6EGdt0TRAUmLtocqaStrsOXyWI+MGBfmwd6mcxdW6S10jaNI/iRXfqI5W38sVr
hvtlIgOvSUqWbmNdjRQlWDTNFziJ1mCPXOvSpF4erYGATkCSE7v61rfO89YN0cSRMTiWanqnMUps
xWeA7VDh/kzvdPSp0piS0Kjj4HPHqATWPxqm3R5jC3+I1I7vWzRU77HwC7Y/snGCtIWyOgmalIXN
vUySa1CE+O01cLEAnqfL0r89ANfEN4l5gE0z7rNtA1tlFpI8fJPQHn348Pd7n3ixMXlz1mAN+NO0
CzrtuxHuKbKx3/h7SXdouP3yu2JJKkymcunsyircCmVwP2rkYKHONdKYxb6dXkIpW3KRKKlU6wFV
H4aJQkOD3+ufzY1R2T2gGlzi9A3VPKdM/kMBPwASBiPvsEHED8q+B+EOkcig7NOhFOt/ytwbtySV
+JZyDSxy7buK3wkI3EUrxDc7Bp4+CTVsbQ2uKtjE8WgAUUsKH4A+AD3HZf8V/bzbImi7+OVh2OyX
ZxYWrPm3xdmIm36ajKZlx0aFN+1DbUewgZrosDYqOHcyfwIQ8bQHuxSwJ6GOi0x9W6bEqt8l3Iz5
irOFwbRqtkarHaK8vsnG/amDbatKybyOQTM52AmgcqKWOQUe/m6IFcZKqryAOBifwLmkEK+exJuf
5sAjPJzxoK0QFg0oTWqio+xtPdLIa1QJQCBPbnfTTQqMcQ1a1g0DPtfeOhJ/pdtZWiQnXrrS/2C0
4s2F4rjOrXhaYz1UHrub22mtWU87IccsB/uACkNiaXkff5TtfwRymKufSd5bwbbOg5/9xDcriCKM
WMmHg+Gedp4Y6c89NbJxxo39C3vO5k7r7UIvHf4SMOqfGXMO4jla7+HGrWgknEizJoAmzK7Ay27Z
GQEC0juU3bdEzY2UnOb7nppK8aWpLdRHl+k1Ub0xCgb1SbxxqXHf9uf10ZcIvD4+p/s/jmcq8YhJ
D/bIsdu7KYkPuMu7ZRfeBHdn92p2Uwt0Tx7LKsX+nZfpjanVWkiBbKJRrRVCDuExDGNZUr2Pkq+g
FDWQhKJ2PWZMt+XJPjQg5kSjATykLbab4Nsncukayd+wcAt0LpsSOzrmVlhhpAyxm4Kv4Hf4kOdG
JkhfIrN4llRqGrFNPYFU5yL+t+ejsDEoplEL5wgMWO1H9ny3+1XJSjq4PLfFu9BorPCph5r7u2j4
nT2FWljnOim08pLLIDzPQxtCJpCi2vQetn2ZeN9aKOiJ3g4GKAyrXLYr//hxdWgWxM6Ta+qKiG46
TF99V5rFHjVg75mv4SzVNKzPC3hgR+lshsKRXO3TUpT76Lao6qQ0czgukRlhuxHlJ5sRvy4ZcOVs
5hNZdyzzy6Yiq4QX/0EP9t2v2E4I8gtBD8UEicy2dXi4SxBHLAjbTcPuLoaQmwaKPTFE8rxJFwHY
iNZDidzZkpphLXW/5/cG+2BBdnOF4o/xOPOYjZGq8Vo5gaZAnk70ndfVL0I7Yw6AN25XUowD6zRO
DksDkTHOB18JdUdcCcg9vP4jqR3Zt1rLmco3ToFKvr7pb6tgbDtCMf4WuKepwqQsQgqIM3FLt4lZ
zSsW0jHRgXXDY4JYwVO531SPanNSRV9jcmBDINg5+TAA1Ak2PpzmkxHDvyX07PKSIEI0JDkynrwS
LwPt24pV1tDmPvp7FRUHIOgoJE4jcsienkVYdScJbfk+whXzGKvb2twbHx/5xHZw0Ewh0PgaIKs6
JNy6wj58GRNvuusnNEwtm4FEcElD53isJcJZxPAyUOToaHphuxP/SMLxzzHvC/8VzqOK1S/dkTJW
J2RZMY76EzNnrSZoJznMOWZJxXkry8AMIOVrupkx6msoaVU0EKSbIWYtK4e0DxaPw7VBQrsrATXy
0OeQvRXweXw4ymSgMv9h6+1aV06K1spyyrObdJWTKaCsQ58dp63bY8qvxp1iiRj7UEtRnNL8BVzy
scRQdd8d9mHgyS9wGXNj/3WNkz1hVE5vvBpAvYlzOtzMELj3BsuPbAiXIEodrXTAf8GuuPA5EkfQ
V8hYvh+JJR2/7wrl3KTbrWLephNYYP7mQeJ4rjaG6B7hLmQTtcAnpsnwFCAVgGL9u0c5X7H2B5l2
F36CPmseVWFf2W7xfGbiBcaiOp4v83nsOq6b6u3hnhNUNV7YktHMAPG3xzYoZliNPzKIOYueZwsc
SnVQz7SWObdIygAEW1Wlkc9pQqShUBpvpEdUO8grdj3liOWKk+9ESoV3hSiSqy9D9OavQxnAVjJH
xFAN48cLxr3bS93a/SuM6vT2FTihFqms5WVQ5sY0HDVpBehEcCipzKE7wHA15bLCmlJpIMuzoaBZ
l2acxnBGGSyhyw5U4BxnfRXcw922BeQ8PCZf8RKaK1W7vnvPlqyn0Nxp61tKdfj83qAfUw6I52S5
SzjwaEprZNZfzaT6aWwFQ7F0GtlDpsSJmdW4EpQ5KaYsj3Y7fTkNFxGM1UUcIp/KnifU5U1MHH0t
Ewd6vJVxIMNB6waiNzGrruG1tgU8BQp85+yaJvo0Jm3WoiKmT9jJw0vIn5chvU7oNq6dhMAguJHD
/0isW/uCaknHjO3c64VY5KZHW4mfYiHkcs2CWcwG1vgT8/jIa89yIayIUAuEv8hvrX3Vfr2a3lhd
nty03mCoje1JG2BnLluBEDpxqpQpJfhlVzdhxkexENCJxvfdoP5oTiq67JzwslapPZTEw/+pmj8f
9o4R0XKrz9/vGaS93qEc7tSj3ugqbGDqoS925grfaS/Eee7xgRzVuNCCtXJVGw959H4rlVzhoCsY
kyxg6YiEGkXkeaEWJs7/eZRMpwdF0B1+SBzXsq2srC4Tzn8FugS71x0sMG1vCMNU1Y9R3gA5lziQ
2QWIf5RqI2eKpREa2UoTS6N16l0MeO8iFltFHPZl87Z2tKqkLM52Yk6PJoXDRhFgvE/dQqnzpWwj
on4aLvfkqJQ8utMpyhzVLiqZzCXDFZzF67eNoP2NupsSdcNYQO1oMT1/JQ5ECUI/tbK46NgAbnfJ
/UzS5lTSNYgG44xVKYik0XZM3+yEFvTDgmtXqCLj9aXcMU5Cx6WIykRIfrQ08Mic/Oivr5k72Pi3
V4LP+8xpSXp+9eeSUtr8HdjqDtmQJ+XUa8gUIwJVsCCCEnP8/2EwXbTtLRUv8JWZfAoAiQEHmG9G
JZ9mSbiuWB48XEIJW4ViI+tFmstPYtTxheXro4DQDr//SnzZ45AgZdXddMAjXdXfY+HzpwY5VFsb
YJseUoqqDuKIc0gKT1/CMxnDw3jGIjT633gUWyxjeqfuRfdhAdpfGOAYHDOsZ7lcVk1ACACReIEP
NBkDygT0Z+d8RtX/94+E1W2KUi596bDnthttlLN+0N3geeepgoyVGKICjBiMluFEA7QYHpN8RXlt
72e3gPlYTW+hkY8faMlkDchdg8KqQJfFMsAemSFc0PtsjWHa2gYcWxi0t42y73RUN2SXXHXUsfNH
pSRsfhmwFNCe9ut+xFkOTvTDoVl4g/cs+4TE7EaezWcU3fHrJZRaYGzgmVXHjHSAcMR9uOYEU6bs
wx6j1Vp927D6bY+l/SS0vkCAgxQATf4TYTefhSlKpjSXX1UlSuagCQtEa3JyzTw8KWcpKXegBJVO
qrnO6s5iehYIJHz+6wiTk6imNA3b+vduFrzEhD5XWKZLE47yJxIkAfK7ZOBtc6U3TxHfc4aCBVfz
Vlotstlcow96RsMhY01SI74S+xAb7MqedTs4YOBD4xoe8wSpGCdf5vl9Om4KZ0aZNxg3j1VnHg/H
2hvS/ztZ8ZEA6xToOu+9JIFIUi36eDuFDAymSohMQhKKSOFk228njifzkYIWiwhwaFqxQ2IvmG7x
6K7hjatvCQm6U3vLui51bVT290P8sGvRfs0QcInLBsV59QN/SIpRhS2EFYp5UBgO/0mAsnFXY87r
uD78DInPoZJcZcBsuzhK6Q9g/opGv3g2b8jnpDK9mwtDsaZtJesQC/ze9sWTklCA+7kE6RtZ4NAe
qyMyz7vi56o3Zjy8xrHiCcCrTrkh1BWvxcDht167fStxEnHhYqaThnYr35CcpMNpV/Q1H77ZMEpp
2XRewXp0ibpOYbiSLOG+CG0FAP9jZLc8ray/onck8dpQgftTnZQftSkudpJRhLvMnhViHlhjUXvO
yP/A5xmw1ZbSCnbgHGmdLJfdNQCjKgpwy7oUHKqeUoKrUR+nmPRQVme3NhDqwvfml/xP/ZCfHASn
tYJbM832fX5vYYkWIFaNo9OV6nyCVUP8g9bF1STOu/dNYdxwfs3H3uQyMwCWkaOnKK9QD7qiSEOd
j7DR+F+ejdY3KCXNMZVgnZjzGd7LMl5d5dOW25DXh1fLBNBaiuuZTJ/ggAEc5YzJXanP8VUtIwBO
Zt8fP7UvjoAG3ib7V4OT1YxCmYSyutTjxCwB/m7j1jm5YgnXKPlknnE1jBP9oLqx2LCa3rdq/PUO
YtVCdOE6WB3RncSfUgAnOw7EpCGYYzsuVoPkvFs9vz1uWyPlCBwncUU/IpZduXmLcC0Jv/N4WKSJ
Ar/SvNVZ6FY/wWu4opO0uYew947WSlazzwVhkKbJPmGsSA9G2hMAuoYsDLWTXjY4e07Ew9K6MW0P
wDi+YS/ot3wzSS04uohQ50cDy2O0B/I4fa0x9MeSTV1/E1mRDb7JRoIfGCn81QhCmU3c1efAmCy7
axLSwAw0sdtx4kfGoBq6WqtxwFi3NI2qV1qyVM5HgbRozFzTe/Inya1B2oYKHtkgpudHFG44Xx1l
AduJ0z0OXEQBtnk1g5FcXm8XV38ZrowRAV/TR52E0G5s9W3MZaDqOSTcvLeES4GiOuH/F3QaiyLf
AbjXq1/TgaT3zNxgzXCFvaiKtrx+CYjqmAHEEMD/VIGnEqXzBRhKPmucrcx/h5mzsZB62kRod5vK
hYYcimEmgOc+6pilhSDia2WlLKZ4A1KyVv/uqKF05Y+McMhqu9iY8/ImYjEIJHMWaMiBDXwahDF9
Z0YuMMpoJ6s+r1roBwfSxOm2IeD8R0G45/JoIv5aVoWwLBI=
`protect end_protected
