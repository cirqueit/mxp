`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
rVRtrqv2S10wi/QxH/I7ibdWKSa2ESmvtCCH2vSZ/KlV46AQDq7l1PzlaPvPfgxRW4h79ZYCOhyf
X52PFwyEwdrT7EDHM30AQnEtX7xHl/axKasN8idQDWWsTHPeNXrEyV9Kad+4cEFIpYD4DPFs2GkB
tAgAuamQYrjuwYE3VcG13bvHycekZl0f5fAbIMuYmUVEwT/6/zWILwljyzzwqMc0OlCNmZB8G3WT
lZ6QJTCBQ4v0ZJyRFVKwwfPSYjxpwdKjZ5g0Tf4bdzt+eJ/VnlMkm+6Te4+aEFpdjaaVnVhohZye
AzK1J1q0FH5+pwe1DZd9ytCr3KNxDZO8PE8p/1KP18vOR6AnY6WlLjdpO9v2XHlUXnGWuNHaTFHz
RiIgFnfk9xgS/ivyKth9aosG2ALwfUcM6Tp1OtzuQxxsoITcBQBDE2nud3yj17qVWajeH8lvFaA0
Kxsf+99HWyftuRfH5mM9OJKb0WDR8KszIxQv994rm5Ebsnm4N7gknYKiOqLxRu/jSxTrKmjr5PUx
mZRkAyoqikjAwjlSHwqucHzHMrvwPQ7nTpguSq97Fy/KOF1KEkMYjaB5utCyH/vmooOqTjblVrnk
PkbivSCdDGOehtXHAd5/0Md3Eq7f++bVy5X3aVHuVibQmugiKhy+pSj/mcVo/WYQpSsj/3AXURWw
/SBWUnQn4pyue2OR7MA7LTQ2ztcNuZ2SJX0yVb9b9hoKsuJrudVSVnsCOYsPCZi+KE2yENBLEIPq
uDVMN/H49NAZexMg9HgK8hAR7tdUXJD6OBaOBt+Ge/TQOUfgVI+GlLz3J7KXi9yI4fbCDg1oOtqP
ZZET76t0ZaH6YK2hLeRegKMnfHPyrB24YHESjJt46dq/LUkIY1B6Pqj1MoDKwZR+qlev4rbPa2j/
DnLQVGsSsbuST6piwfuKZuVl5warPABrnsrW9q1w8T7TRczdfoArjVMM84OB398XoDjnHS9zIGax
iNLBZdY0r5Cxn/ZnOXFRKjG0qHRqtuKnuMUsQhmLSJ35Nm9C7prEEx+PiT/DNSNbsQHzSmhMcshj
qfecoxWuocotETNkQGo+qQzjjZ48CFcRMroD4BeT/EzXLQ9CJs4D3UGXtt8C3HUH1OLy8XaMF6Yl
o5NaIsQspnxg4rU+S/9+ny9L3trhU+VJRQg3Hsjf3W5/gdh4hEXHbHwjIPKgV+hTLCsUjVNsl+uJ
pIaonRXMqn1pSnkOEhrvLj3ApU5FdqRS3FrGFJVIe7ZYuSLZIAaAwCPNt6p4mVXvYD1/GUO6SsuG
PuNZIfbuX0iY6Rc1250tWLIR6lV0igCr+vRaerAJqoXflhB5cwHba74LvBkRC4S7KlWOK6yb7Wpc
v8Y6SMkzKd60JKEfeeIAJmSzQbHNzt8dvhDw3HCEfVh0sWA3n8aL/dkQCeP8UkHV9JKaPw2KnUgW
rwwo/xsluMe+RFQjWxnRrikIrDKJi6A2b1toQIddcLB6SRL1JdHaftkzqrvZNa9TNqD/GTkO+qlN
/jtHj0MRr6xA20S8hzq+48IEBCz46AHCBec0jOmyNhRLbyto6iEXgsdRNG5k4MM/pGMF9w/sc4yo
+5WtgDTdgoDQGoCg/3bruecj4Z0ni0Oak4ckrv45bdlWk9Yqt3ADhYTCtPEq30xgxIc7rgDWkxjR
aYHrc7CyawmCZ/6jyjk48VdmD4/Z9wt7CrcP8O+wxJsf6DdgF0cnpF9yLjLjHI2ePgVTbYUNHeM/
8iwhYgZruadLltWaecjek/u0XQMLFoD+j2Rw5I9aViIZ957vhSXAVHdtPogstzP2NBIoLdB/RK9E
TqMtll12OIa/JZUc1ZIl1qZNcSfVGeEWMvitA9xkf/YRTUdq1dNG5EgjkqCRbNLTRylYQEsIw+Ll
QZPlGb8ojjhl59Z4OIl3Q3HYKsXzBGWnUw0Z1A3X3/Hazz3OY6P4f0a4mY1+Fw6uRKfg83ZcB2Ta
AFZcUySGkj3nJ4hi4KuUlaQNcYMncFykHVMBnD7PJKKI2zMgrGhoDLFb3djz24h2lKZXAg4cHEaI
21roqyx7yXq0dRHdtMiPAGZD5MFpT2fph80T3aw6zUA4vjjV0iv1hptRQbfQv2RvO8DELMbaXQfd
3M+VMm/ydY/hT+W4u1IFj1vDeCYpAIoboBR5shNod1uQIASqp3hG+sxFH6TvK5uPRMPUc7Ye0gHn
fZTTqLPYCKZqJKYRLi7CPjHNHJgrV7qyuiiWAsjB7GiNe8LH6rCWqPUP2XGlZ2dO+lE7qd6nyuSB
Jzb6qD02UjbwCqKKCGvQyQ9I4YuYRRlT0B8J78YmLTKDAE0T2C3DScW5cXErbeS7PDS8mXqOiJAF
2zeKsG8fTmXGOwBecW/YQsjOuNgZeAFORpyEjmHNXDIiaoCL7RWYfU00y57E0duYd97o/8gK6sxR
sekHTjVT5807B7hC75wpHkFMgxGBjQ2EuUA60/yMiNtYs8OW4ohRravKaq3xfPjtIjZ/TvpJi2/4
YCUA2M5wglSKFj67LRZMEZTRUzUDVTMd0dvNv+HitnKCquWq/9LbEtws2KFk0gZGpNLs57Mt3CUI
s2rvdwoRy2x0qbyMjsOc40OFswU84y6KhXB8HnFndkxXI9KmObv+pDScgEl1T1aESB5pZulc9bn8
XLxyPYYTzGDbpSnLdLkv4S0mBtAikEGkyeHRVBGn2MT/UFLAdtK5oM3470sqmoQ1h+9JcJIT0M7o
0zKlM6B5tGhn0dgYQ002dDHNpgcXmjtVCRKw8UT4k/SREXn89vMJ5/AloCxbkZz3Fq4Vq5dt1aEN
bU/9ABiNrm+8eN4IE3N6xKE1jj+FlKLxPfUymHGIGsfBUOjnu7zu4uGH/eK8CsU13bJvx3obvdgh
R7HGfYL8VYu/f3zMxWK08SyrFFJbXzmMukVBQXIHXnQLWiXcvKNmGH6mjRTruTFsqpTcLBU5PVpf
lqzRZFFRlvJ+bNxX8iyaJpBh6BXoaZrGhw8pXKjCoAtLkrWhB8wM+77LIbFEBjgoz4ZJg2btFTrB
4pfj5b5Q8LbO+wCLv5+ZwIB9XbuwMwy4b9FkWNVN6EaZk8KardB9xh60sLh6NJ6zGF7Zkb2NCmy7
Vspf88ukI98VrwuVTjXRf1U4CfKYO0kuEjPOojKuJoqnQ0ie2xlP9yQzjEvCeQqPfCZxHyvxMaFf
5CP9LqsW99w9Gp8WOKnjr2WUchwe7YoWMcXDdFZu9EAT3kWjchwUNqhM0KxPXK89wTPKkWFuKt43
tMxkwNd+taxVWKPDrqEkS5Jhh8PNsW60FoeVmrIR5oXZH3rzwrWtSLUkzAz4LWn3lbHigLvyDG47
2nnd3vT5/2Ja7QlKeT5/41Mg15odINHqKfIKlfMT4MWah+He4ir/btEVqNOuuYtEDTKrywjYG2T7
n+3atJ/IYjOojsbIdY2cfXbYELTA0SQxOTt6qFREifS50jSB66nG7RpNgHjikYVkV+tGZrCmPeGx
04n49YK0PrPoGrcFls+dd5bWU4amzSpL6qWPPoWjQYBIVJ5RA6wKY2bM834R5YNn2mExdm2tc6iA
8Whmt2E6VotQdOQPd3Jmuhlmb1jh8blw3WU+uS9sMeXmb6cR4U63grIeZaTsdC/zGvNMewf020L/
Ulduw4xhJd9hU/msT3ACn5EFAi5huyITiekawTjCaLK+y7dQ3FcyrTt9KdEocQKKrivH992XBbiW
OkbeAX1fAgjgWVZSwDhnCyeKxpiBTVqdOtkUsi1+UeCdQIdwiXWW76gEp1g0quvphUEOI5Qzss33
wKLEHpGn019b4iL//J0goWoVtxxSEUf+lyeWZCViGHp5gyppgPF5YpweG3cLk62TKXaVMNCtDjy9
TkZ6fjucBr3xODVMgWFBaLPHTiTzZdLmPydJq3DGOqKV1YpH6SfL7AKrDhwa3+jd2J5bvLGdXRAH
MhAPTyX4kOdHPxaulYf6021GUoT/mj4irh/qjiaTSiLaGX4WU90xiPG0wFcU7acrChDyrPQsgb1i
1HbaMxQNgzvGzj1pdU6ROk0DPwHHbEL9Xhaw7EDGOLfo+cHS7wqmOB9s3CiXUARW8o3Dh0OvDw9y
poZbfwiweW1KE6dGALG+oIdCdZxravLP/u31L8gJq4Rg6zqgyKbgnCaf9QS0M4b74M78vnk9dQXC
PJpS7jPOso+DThEuiKerhnCSTF1+1ojRZFN9MVIOOnPiMGtX+AgfVNWu4wdNvDpUZO4nCB0lSHCd
MomrEcK4Q5UYlkbosL3JHOfs7/Oq/hCAIdEnn8OkIwcmOMOJVTjCuwKfNNrfzKOJMDYiGnkuL/hg
U7dVSluSYsv1fCbOreMokVw0W79Ii9e0dwjuwnK3aUwi7CjRTM4gqp+Shdt43y1GLscElTAOTiPz
KDrnsYan/SPbECGptkznBfG7pi4UXHMS2mrnSnGwdg9inw08YSECRFFJm4xt7KzrNzST+RrIRPja
BQOv3Ry1KrqSdrfmHrYesKlZmSKr1YXVo2ZOTmK9YkJ802nqcEXXuc9uTtaMkk/RhW9rrpy4F7GL
el04rjaiIhuvTDpmorkNwQH8A4nKk+29ou8TN4M974oyg2YCUJTdsEVHZmHxDdjHP/D1/osDdI5M
W+nKWp+NxKizL0L47jVeF53vqgSGZxJSF5Ko3SzMaIJ3sUcmbdiawudg+gXM8rX8QFmaxnQBtS+8
gunK7lVE0yRCJmUKOD4Fj9zlRqnD7bOdnLluPXxBKSQrKqay0LDEZwUYSDgVTJaHIxTNkebB/zEK
cZQXedOVscDAW+6Tz/wTv8CDY6NPopXxnwzyHCPnNNmLAOJIEnVbUmQUtRV51TtUnu/qIU5ZHy5q
TEyCw8vPZpJJ7IM2OdQbeTqZRhpidx72O1q8uPRC1yAjIy+v0mdgIRKwEVZbF3f4cDubBb/Cdwe8
gmptpp+FLBnJRksL1HvJH6UiPXl8N2cSsIXMrHFbAL1TPcRN7E0WSBTupq88e+4m/iiGwzVO28jN
Ov+qEktSPlLPhdUkvuLtGoS0/mFzDVGsNGQ4JDv/o8SQ60rrzMlvSd0+5i8Ar42oBa/8f3gbtxrM
8aixE5aao3uBibvmNIi+X2x28BKA
`protect end_protected
