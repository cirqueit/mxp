XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Kɻ�ۍ��,_i�=�PT�bXC���tv�#�R>_ܢ1��/�.��4V���g�0�/�&�<s%�C��BZ��u2����9'E���kt��o�+��Ა��\�h���mW]C	o-~ ��$�!���aD�P����R��ޖ�k��Z�x���{c�5�*��,?�l����r�mM���zAѹN4����b5�ŶgB�A�G�t����pɉ3v�_Eի"�G��@��r��.t���8��N�Үo� "z����@P|.ɞ�	������}��kmb|KMD>Q#v>�s�n�4OG����������C�uFo��C!�g�Cr����W��2�c�����a��}|���/{V�	_~�3{1&w���y����OD���VJ�c)�!��liW�]��a:|]�# �3q�h�7+Q�6������b�D�0��
�j��cd
��)G�HP��lٍ�����L�p���B�����ܬF�72zW�}�_l߱��. [�У&ď��R��>�A+]�nR�,Ta�T��/�J���{���<���
l�.I�Z�Ҥ(���'��\"$	��8��*�|��D�K�}D1L����X_҇�8�M�i����zQX��^��A�=���D��Vl �����d���l[�o�Z���A-bQ�1��^���fL��[�]�7K�J��q����yI�5�q��l�`�������P$-lg�-nt��Z޻òR�c<�^��	�>��Q�Uq0�tڔV"$5XlxVHYEB     400     190+j�ޥ�Z���s\cv�=�GfH����>|�їk>Wϲ~����w�c��!!?�t��e�����^���0�����>z��C���a!��3�p�W���S�[���s�m�4�P���K=���b������"`�\[�����9R
��H��pIj{<Od
�Jq�ڄ(i��x>ʺs��`��i��G��­3�����M�7DP<K`g����Wj�9)����c��Y����,��JR��Q=~1�*�8�&�������Xh8_��6A�3����P�i,�`!7����� ��M5��]{��L����ɶ��*��n�l��Z��mF�gv&X���%�R��襆�U���f�����ʉJj��G�8��L�'���WL��+�x=3Z�"ʤ-��XlxVHYEB     400     150츻�g.����G>})�_C�fa*	yg�~��N4�����P�F��I����"`���6ٸ�:��4"uҊ��N)��(~#�z�v�����őgsS!�����x69[�������
F~^FY�}�m*�l�՘��$��1} "�m��~����Uk�j��lC���!�l����b�勃0A��Z��٭$=���=��٣���7��Z�jGm�����"-�6L"_u���.yƺ$����i�M\  ���=�r�J��t�Y���C4z�p���SA)ֽ��*b��/����e��]Y	Y�z<ȏ^<����\$>%�,�[WM�XlxVHYEB     400     140
Z=�$�!�L��}^.�׆J����Y����m&�f�{ik�ؕ����[X
�rlo_d86�⸆.W����h��2E��ٔ�I��ӣf"�C��v�a�S6w�-ͶA�1.ԧ�_�m @�	s�T�$�YG������J���������&��zu~$�}م�s��'M�E����C�ɾ�l�����n��O����%>RR���>�<�u�L�T��|Ĕ����G����Y'*",cW17vYH�|�3!R�R}��%�W�o��6箟��d]�����d{KMZc����QJB�}o����/}��.�P�K�{�
Qd���XlxVHYEB     400     180��4��f��.2=Y���#�;���-U�?<tl�+���o0+�`k1b�<{�7�j����C���	�:�%��\�ք�[Sp�} �_8�r{/_�c{t�/��8��;xoә�%��s�-�aGv%]%=�^~A�x�����	���|�]�̙ӤDU�����ٝ^׍�|��f)6M���}��Ǐ>��*�~�t��FǙ<C,��$�K�p>{�(�[omt��!�IYd�*�������A��hVl�[��N��-�?5s8�!�Fz{�NO�] �յ!?�nU_d�.���:�:�.HP��|:
�*X�>W����p�R+�d���^�C����b�?��h��]��T�/�a�P�b撚գ��_:�XlxVHYEB     400      f0���Z^O�%�:��*�w�U&(��_�`nK0��;ʠ�w�zL�Ţ�m�c��*��bR[���"qIiɫ�����C�}hB!mx��{�B#%ƴ�^��'����Z̶c�+ﾭ2}t��k���i�i���N�ڟ���"���q���=��\f2�����	��r�r��姚~0������N�N���bh����e��-��?�[6$��7R������l?8̊��XlxVHYEB     400     150ah�N�m��
��`�Sq��5�X\7�p�ܒK;e;�[�Rwi�Π�憎�aG��Z����S+�ҏOL������hW�Y]�w��f��|I��	
�Ƿ�դ���1�B���lKs��X�����_���J`���y�1�Ǳ�\�,�g�_��J\%}�f�R��g���?��ȳߦ��a��m�sc��w����Ō�)p~��+��c��(eF�̃���oE���x�~P��o���D�~sV�Z	 ��)�4��=�z�Iّ����v��R�9�O{��PW͐=i���`j�S}˅��H��v~Qlj���Q+��XlxVHYEB     400     1503b~n-5���������ߨ��~ݞ��;����T�*J����x��U;��~܍7�;"T.���Nya���r�����9]���J�#�q�c~��b���%�*۞ո���0�`Lw�p�Y�YiD��)���'��9G�LF�_���͜G�Y��r�9]����!�yn���o|���5����}J���QqGIg��@eV�0����%U�-��գ�\9޿�t5�إ�g_����In2;;M9��?�1+��R)a���ִ����~,�Lv_�6E�ᅷ90���O��cz�ml����Բ`����?�6��)��]�-m�AXlxVHYEB     400      e0�[ޮ�R�>�_t�����:�2��]�ݎW�3I^�B7C��Q��[��_I�>�W�BF�c��N�Vq�
���^ϡ@��*��_UC$�G�g�q�a�o��uT�v�_� ���JJ4�bk(�¿Z�H�  �M�kC|PJ'��L����/ؖ�q]��q��t����Z
��g��a��Oų����7�k����@^,�	ty����8�J���T�JXlxVHYEB     400     180���|�*���a������W����X@_];�$�0-$-�F:xN�֞c,���]hA�,7q��%bn�+��ƭ>�n��=�^����z\4�a�"p4�,K�n Q҅'�<]r��G(<�X�
Z����EAnnB���L�gkHY�������5y3��X��'�:�Q����Ć����N���z�lbu��}9���$XG4�jN����lqn�[^�^��G����v�g����=�����@$eC���,�d���%<�*�i�Ҍj2q�Z}hBU�o3?����J�G}�b��V��uڛ*A�Ƞ�d�T�C���TQ��cP�i/�ʉ�R�ށK?�ާ$��_P'�J`#���L�La��W�FP���xp�?�XlxVHYEB     2f4     100S�ß����z��5�.~��bdeTx�rR-��.�j����Lӣ�Ɉ��4���>��G�1v� S��ɋ�͛ćİ��7iY�}��[	G�!��굣h�;�� r�`��y�+#����S����p��/ڄ�V�s>�Q��^kGͮS}�{tx?���`��OP��LE�#8p�f��d[��7Lcѷa3�lT�R�Q6h�0G@���?̬�Y��D�K�:�o�NrP�x`��s�NT� /�k<އ�`������