`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25184)
`protect data_block
w2xbk9mleX3F/NJwB0DRg80wY1qnEyM29HkKvAoPWl8lhZovquzIwn2+sAySle2j8m+PYidgeKCJ
WjTb7F1cSNEx19+n7OY/L4GdNXHIVEGBs+eadZQrLPP2sgQgXo9XtJh7mclJZkfR5SyfFw/bGi6D
MfKtasNKWasFwWhuMA94KnMQZjHAX4zLwRJj1kCIZzYjui2mJlHtlFSKKHHSOoQlR+hj9YJWkK+C
ueBH76EA1hiE+fet/eV6AAMl8Tu/0X67mlWdzDS9Di8JmM01IwGnzZifHmLsuyDcHzRnzj/CXeaI
l3nNevEFTZtCtLAE94Li5CMyQrwUNIu3YC6U8zh37iIHjdoc7+3jwd7IJO1gNqVZS2a1w2iyrqyj
oB6xFMcr2jPC2Nd/iX8lNPa/LwNf7K/vXlB263lcJgj5mfCTQBNySD4+QDX1o27SQjIel1c+hMTq
PXKZJwCvCGEgI1kKMPl8UUZ8w1M7cgadiz75ZNAVTkdnH4ZJgkpIk3/kWvQ+ZuJiRzeQSJPRffwG
VaA+JBgLpVB12cnq/TJx3RGJZ39xuBoxLBC/ZjwKqHKSGalNU/SaAmG1YuLX6hVAe0sDDAhcjshZ
Okjthj7ArQaaV6vgONlNXc7grBIdBQZdARfx6jxyy4GYYT0w2o+ewWjOqtWQwIAuO6E+cHoBzita
w+E4OswNSTsZ66crWl9TSBJwkPgIcopEoKJVD5Cnqin/Wl+Qvh/ClY2ZYFpH5aSzzAoVYzTdshJq
WRHapPy1m0yDk3K2RJ2ilrYO6osH3SeqllRb4u/ajPc4wyj50nW9wbBwbxbLmRlIyL+zVT/kiTzX
aym22UZfW3vAmAC5jXX4byMfSQUAgjzRQ+tSJqqpcpf9Uiv7Onipi3+j2CGteDrmVgPMjlp7eUjI
r2JZ0JWl0okG1mzxDB3CsrdxcojDJIUITJYjlGp1IIGI2Hv9X93CANbsP8+Wxt18x+IVwvLjqLCZ
AtP90jMV6M3SJT/NcjxmFJWh3o8y5TaKqqrKdvbuaSUerS7Q+Dy1Q+Ku/1svp+/cnSY5k6dgaYLq
8m1NpaiR3XmwKv9FWTz1VBJfZ42HVxntRT8G0LPHAgYUYCX/TNWUr4F6iSVptDBwZzz5JldpxFz5
fepEbRRYhe9AK+A/R9LfO80hn43LrU4oJAyPgWll81sBwsIMhZZKjgzXideyUIxDNLTinTtUekj2
reit/x8X5D1evfbXzWgEg+dElYZi6ezXZY6NJup1TxMFQa+gMhWuq3GgxPHGGZJIKvnxNdWkUA+9
uWnHZHPdd/NuurJaURN/anIQCh3nBoKdAMjjBh5njAQ8KKZez9OfnxrdVKJuD7CB6eAgkQiHCHVF
y8E6ZxhqsYen6VimgybNgHhLZkl/32GbNCK0pDU4gIxmz/y9yJaK2u7xC4PnBp5a3FixGsIpVJUm
lkvEV7zPH2yOh2st21bVMWWKX5YLbmRx6dC0Ffp4vQoeztO5atXXDxcOiXCkSSdbSsucVPgFTRyz
QOCgJKd8oUir6HONU+tbq5jsXhf0aNV2dYH0CJD7aYFTSVtuqCS+3MOHErx0YcLIXVUF3Are78nf
Spe2ex30zkYJoM6PxBqWe/TGbK4TE5+Y2Lcq5litmmUCTDvLyWdcXrJ4mQjZgf6iYailr60Ws/8/
AHkE4kF0FXTHMQi6tHIa5QdvvFHd9usu0IGTRtsAGQrLGoaNmGs+9N6usI8DbgIc5Uf4NoWjSFcL
QMdywZpuQzJ2kKl/yDV7WyZijKkI2gYc0P+yfbjt6dSQbZNovqlmEvEonQoaPTSKxyxZYLVmyf8W
WgbjTt5EwgCQE6IGEMbCecTsTZDatNn47qDbvEWdZp0qMOfmhXXyb8PYX1uQweXDBLDe9dcSdv8Z
U04ospeQlOcVmLcvsNJ4FHrFHy1lKy8EIxoogN2qI+60Vqi6bofbvQ6lKz4usExQZK5uZIDtkNTA
AwyTtSLjIU60sb0FbNMisammOVUlzsodlimJvU51tm7zmj8W2LaqNhmrcvIgM1sezYERScAxPere
9GP3XIM1FNW+3APe05pkA67ji7+DmMy2Zn6RKD9IyiwO5iIL6VKbpPepltbaqcRN9KpLpuLniDdP
4WAUAJV/QzO9AiuOQ7e+SSBjENfaELlEVhwAnHTi3/ekCnI5G2Sn/RnLbtE0Nft73IkJ76PLm5cB
6ju61AkofPFAOpIJc2BMWQSSA0CGX6JLa5oyoEBiyd1rDC1Ir8LsevxJxxEvc72FKzDwvEb6SIjs
lHiQNC4x2vXPgNyrCuBlsLvija4JNFq016ZwqseSTFcAH41lcBDWKeD5jiypQITp6ohCQame9Sjl
OC8VTwQ7tIl9hrDe1f834EYH+XMj9PjbV4AcWA4b+pO4Vk7EABRE2wpPoXqQ+vn0Qfs8SW3IEu3r
QcLTtZz+8DOLOMFz/TGcbA5rPIhJs/g9dntdS+YkGtqu+iQcqQEUmsgUqAXUUwqgRS62znUoi2vT
l1opUMn/sK/6sAmZZH55i4enHpSXpmfqBi2N5+iEzI6n/wBT33/v44jRs80KzQc250OrniRR4i2p
KuTfURG9cLillFwPQMbE8sXmIc4Dm1TBGdOOjQEAFFT3TAGRPoAd4JuHg/ab4870EtoZmVYMr7uF
7R30uDV1qEJ0oKzFjAmFYOYRN9Tnbpi1vCdnsQqCI0JyVr7dkrQ0B31j6jXSRJ3QV13MN8qzTBjm
Ni+omWW4IgjRBTW7YMyTzKIdL69FAiYQ9mwyhFSzIAxiNMLhVkyGbq+dRSKIF7zU7h6LWi1CQdwL
2JYVSk1aVCqkKDPObIjfV6Pm/O5cmzELLZ04WWZoAnFZwpQ1NWFiNN1JGK8KV/3dgGLgQszmVvVB
tT0jZVpRcb47o95NKAR5/ls3sSpYZo1YPyQPkeO3TDMk1eMaFWb+ZOYAailwqGuyMHjK0ULqrl4t
F7DFr9fEiwJPpMD/VC7it9uL2RNjFrncRn1fGLytakQlyYL2LLXcgfAlIH5dRhdR7mYfg0JcyH7D
p3ukLkZITbwOLr6mL3a5ocPz1VMDcxaDfSnjMUVgQ8RQVlkfe0UqrAYkhzyPGFSZAugUxkXdXdY3
CU0dg+yFsGHhaNTVjObbiHRQIvbtE+dVVZBKhbj3AEvypR6JXh/PiaHpm7a2d+qVvf7cZIC5VkBW
CnnVBcXK+DIATKejMpPHebMeQDWfyG5NFUrH234lgAk8YJ38XR91us3SziRlQt3QCuzAS4zzyZdz
L4eNRUF60i3rQ9ZRKObldVNIDv5loCflbUgArEBoaALNdT8GYgwsOyx9GcF+6HlpM/+PK1GCXWmu
S9L67ubkhk2WD27JE3H84Z+mpRBmd1h12Z7fxuKa+0frbvQiq33XZtSsJGtbFztSris1SLDVS8GO
x7wPiEsHRgSr0wc3v1ZSULmZz1FmYG993cxLdky04yBtrMjOu/L5X3JhcjLYy7Rmw+kcvUAOQ8qR
s+vODHVmrIRfVZ1psRVkiAR1T9DEhUDxF0Bwp5lLS5cdRUWiBeJDMttaABT5omSuNeUpOcbiOJkW
FjQ/7AR5M3f2HuZhm3JbKc8GQeczAS7eVkbkJAuhc3H632vaO3n9v0Ybi6lQCu00UPKQJA3aROk9
z2sepAfi8do77aLQ1QCjG1NDELFv1B6WlibJ/j6QP+rxESotQHl0pR+pYiz6zz0C0Yb3eLawNO+E
tHAm5YfOH8k9x68izPxKg0VvcCxl2jRMnMIPg7i1IJaNo2IT13gNq5gxepHKLuV9SKBmH249Kktc
NxT5anTRK6yFUj4aopBc4OmJ8nWRbnTDPFgyA/zoXRf1wmgkMYWpLPzK0zr6IMc6Dy79FIV3Weym
+GYvQVXU65drp18WQHr29DPL/kDocRb+UXKWdP6PAeiPJONp8BC0si+GCvKSdeT2YnHevKB+2JoA
+qGAiAwE3D37vV3jIWuFk9tn1FxgEHdKoXo8YIOzs8beWKRSHw+qBr8sPkT6/zIXpoe2eUoGLa0F
lPP8cB3AQBthk7pD7IWRAEMX24SESfTwqjK3RskzsnAX2aqsG9KttfZJ0TUjpsAnD8+qp/XmAjqP
YiJiKA7/4NbyaKRwJadb6zaGTMS1YYcK1beYWBppkz2B5qvZTTzOurptS74T0PRl4QPJduq9yPTV
5d8BAMck3ZVYWbmOamOezuIlvTTz09v08zir/nsUaRqGnHGzEsS6V3+rJQ+sLpBGNdv4oBV8G/LQ
alShMhuHA6h/Aj7nQ33L44Hb72BIFBX9kZErswl5uW2//GgTarSoxNVd+YQ7pDgEAm1l3R2HwEf4
U8dQIxQZlUqxXszgvDmRG25FxZvXftnlqnfjMiUHmjW91DBBKEhDCVMhb7bO8G5knTg34cMNaP/H
AfOgGV4KCL+OlUniV2rCGF8xiKfAVi5uq42tjxY9VNR2rLl7g2EfUuC9JP+ZRnOzNFkkhYzm39Qw
kMEbAAVS1YGxZGSkTaZ30foBzqh49kRnMuvFY4uEbwn+4JwdwREx258H0dYC/64veJx7Ttf9qkzQ
l6tdM3tkmXBq3PtVM7gz5O7e+2k33GUHOA+kq5BTw3b4JUa0Kuzk2gQomSIvht8DLkULRr1gN+SO
VqNfgoiwOjTpRgJdf7XFCkBnIH6BOMiNWKDykU+4ngmRqcT9mF/R19OqUuWN3bXAGCZoiYVVd8wG
mGKPtzyvAvoqSmprJgSH0Uxp5LaSMRk+SoxrAxSVOiQkIAFJsYd1vMBO6GgRLIh1UYhZodfXp2Cq
TB8zd2XZuWI9VHhlV/jUyOANFehXgYT3BMbW9vnRD6tWVnKCPy7v8dYUVOdtxtdo4icdtaRBVEW7
0tblgt6EWME/e4uYUoyK27HNzejZAk7nqVenAZiIrFicOQDrTKQqwRCPLrwBME+f6ged5gB4uzXy
g8ryQq1OlngT/iICxdlnFYBEHObontAYjnm8Mt3GM/le08X5r/Cy7xSeg1YQZ9tiZF2Ayk/AFt/C
BFZhYCj8gUxV99dDlImNkN3uphg9mPJNFe0UzPN1nCdueC2u4M0bUXkSd2GENLcEhBkM8LZWgzmj
e/JAIhlx9l1nyNPbzsgNmoyjjmqsbbiFiijUmsel1P8wR89YCwLkOh/4zTM4H2DFT/AAvBVZK1aj
f/fAS2MExOy4Ih2UkwUi9mvoNLUq8IyJRVipUo4bVj1aauJYm2ZBduPXlz2U4F5jdkJYjYv7bMCK
Y4nDBBz6hxURXG0vLpbMnl8D6y30EzfdA7irjfNbldQfVnVBtq8O7R4Hd87Zw1hFD2KNj3qjRLxZ
K/NIcCp94dGzqiFDFYS5qzZ65fDNCGi5j5TtGy97EEllnXs8D6JSgup8+FZOFq25pYMw1CQu+6kY
2gkHUZYUzb/PwcBwvkqPBQTEJti2BKoaMX8Q+4J7uqFkkiiCo42cnFKFwkGLztIYoCEh1c1HenjW
WNMo4XYnsfbJPXteM5c81nq/ZFLa+9uDIQL7DarH75aGa89Qj2Lbqi7GU/r07wAnROJG7HeUYC0r
XD1HTHsRObbGxUB6id4mmkRWIQSzyCTCKWQyReVoYSg4JZqT+oh4T2Nq4XWaz1I5phJLv6hm+sWp
DtuexKNP4RROpeIUoCy1XkbRmyBzgITLulfffPRaeMI8cTabYnPDk6/yHtxCHCKxfhx6wum0D+Kz
Hs1Kuh1jDM2at0Oz5iiJ0CgPoeWfpFB/X/euX3iEJcby/EjBgsRU1yzKNoDeAHir5mSLZ759V9qp
650pLOG9tzhv9+Ykw+TDsi70T7eGJbOxLCpvpmDuV3GBqUi9ZAXMG0HIMidQuhdnkx4gQ31ij6wf
kUlFvJvpCvJQsbXg4ZGR5gTPK6xa4t2qVDiXL7CDvnIFyPTQR6Yobwe2c3+Lh7B/Spgl111tD1cj
j5g7EECRzU/trnuRfNi7JSXLfgXoUCgpB95iKJswn/I4x89dSoSKxv/NAWIh/UwWphuMJiAAdNiB
ujNSM8oyc3koQuRb3+Bwg53krNVUP1gRuZJnc/y2HJ86WjTkKkH+uorNjrQQH3SmixbW1mjCZgKj
vc+Ju1y6n/Be73v/xPTwVT41t3oLLYzyKDlDMpN802Zbou0WyW4F/wb1u3Uv831/bVXQ+J91pt53
oKhKbZ0EpA0uFuVY2VnpFp2L2ZWYNsNcDeVU9hntSkBfnGOScdfOruWgr4Djr1S0eL/GbOvq/R78
kwbz3KG0u5EdXJxlYFhBiZgHic3QBcR0JuVpY4jWRBrdw2pVWE59oJnCbdz6SBPO8K4b60p3hd5J
owtBMqbHMnmJkqxSUAGE15lqDRvlYrxr0+LOYXuPTL9soblT8H3zFcq76tsaeZAORslyJNRneZLC
wXcxAu8/24mF6wy+9ZQ5z3dBREybQ0NCW7FlyJkNN3PFX3p1J/12xcqokVFowuICGEizGZ8tZF11
3hm7bSGTQOvpu+7/0Gk8h6Y/tmxF/RmVewiNaBSB1yDQGZ3sesL3CMTEDd/9HF9JoqUwX/NwZuNS
YW0BlGpTHL40Tp0cRq2cZdSf1vj736or8KPPhCfokHDtGsTRiGBv6gCsjZbBvTY3Yo8CABegVzzW
9LJZVialzLMVDqielJFaV9OZ8kHNxjhLBeHhgdvk+Avk+EMo7VX+8zGF6iBQfbmIYWQMwxCKvvtZ
bd8MynD1PnLK8K3WS+ELf8tAiBUQFVCYD7RboNxIj+g/kUfBUN3A0jvK9pQyb53FYi6janILGT7j
KlYkn07lcJl94273O1JTCLe5x3fymPbO1/VJEj622D2IMlxZZ8CeW+W2/TukiaJn+1r6CgMdIWhb
5CIDj2VpdeM1zLxCxovmhEhh8qRcz4WiXL/FNoNgZwPOwwmxIo3zTSKtR14QgYF48iSycYA9gcfD
o6IwK9LYl5A282zN6nf52Bfzvq4olHlZHn1BbeifAuo/e+/97rCQmPEGNM3hcxL1KKGGVWpy9O+d
3Ab8SVOIwWnFs/uX4cya4Hc1bh+rqIP0UZlyRNxeSKTc77qokLK2WaNvVvn15zFWNYlDHwEkdi5f
GD2qGNnUHtfrxNywmctHoMxz5LH0Bl2vP32Xe0+ZZ1vF0JbFFOgJn/CaPxJdmd/clhG9s+ioaOiA
ZgGoejpi7p0aONNwpRKTgTPvfP8x8fv51y4wWJj9lO/CF894dPH5rMlHIOkj4kk4cY4htmE2/47z
YIvKlD4qy8qWjxgYRYSrp8Q3iCtZAcdKsQ37r2Tl7sVHC24sF8w7K7fzQ8BKW1ugc0ntnOKvwJXT
V9PHNjOtAlVpVV9H1uTHUKsrpLp4AFMCGXJmk/aB86XuJLv8WdcLHSufx5PCf5PsrprITYTevrWt
F0ymLHZXAHLKiln0QJAEbnRfdE7e7cc7b6hCrzcPhlsubT+c+aWA69LygLNfPJwwdfQ1VJNZ265C
q+T1NNuQH4yf6zxZgSvHEtViFVbsESrGth36L+TkNZwhFhTC7oN+QNsaoo7WHzFI1ED1d1mnOZj6
4xMLWp6xt0/yeCMNhSrcmY6AhMTeqXrc43kFzY+2BwkMdgUtUUuFgRTe42mBLf2g5W+nWhrdDZfE
NOCNz1+jGLB3l/U0QimM3mL/E4L9kYhhWRivcRcSSF4eZx1wCj6mWo6WR6ZPaDgMGK2GA3PRVPzY
6X4y0CLzgsx/2M0/qd047PG5YMatUXTyOpUuz3B63UNOLVSimA/5s6PkxKaxHAkMz14r73zhipGY
bk9VPjbIIc6wZceYEGbqeBG1vxwHy173bTH+tYtBXt3NCt+rNC411JkQx9UIF/cssNv/T0Uda1UL
YFbcfoCVjnjo6W6y2TajffBc1HwFYDpT5nsNcutehvd6BPq1nDJbyh30m736TV6F3yw4ZSvPlfEJ
CR7HH7NnYmQBuO6nICSCj8O/rjcI5uqMxI/qQ/ngFnHEf+Bs/kTH1ZiA0ElMwQlf8o3ZdPbQqCzT
1/L2xcIIzt0ELQlZC7MG6NyR7IopQGJh87Bau+2m3uoWpONxlohoT+nK52iG31kVIMvw1O2pGKhT
XD73UVNmjrdtYxqAcUpyTMQy2igQ5nmMu4vYMao1/wsxVwOl3z/djfLMiVHNUzz4uaG7FTkoGn9a
aHpj2rh2sgkqR6lA5RByVGZzK27tcnpbGImOBrBva9ATt0HRCZ2PI4eJg7sJnJX8iNdO8gg6QPvH
iwjQzfFvlXo48yVq6hIPAzdNQgGJj4o5pONzBt1wdwOD2kWU6YmBckBErvaxDNrSCrXF3iEdgljV
eJKhGPuICcWYkn4HdS5xkni62SjUPtQ/InhosXTKZyRtptZmnwzXMEm6QmuNwkVho0rKPI9nbt1/
aP4eXWrOyoljU9tBlUY0r9K6i9gr43KlVJDfECPx56qwGQkY34ts2Ah3+K4E3jXaRUuNa2WO/CUk
ab+RITlc3ZbY0tg7SPCX0+lA8mmwbT2rvQh3/hWBVi3zMqi3hZwhA3GVZj5HRrnKNKIgKxw8ejta
YDfeOSRE+Jh+2eVKnCTd72rS9E41tQljsst4piGYGJLDVpmrtxso8+3D2fUJT9W1M6jrmI9Vp8pU
y2TeVl6JtYpGm+LOR4vXzeV7D2pb04D/8Fan74FhZ27NvyR932Hh4e9lFSr3MCBEE4ZjCrW9mX+Q
VhAZdVmsJDtIgpMnHi01OfCK+VpTWzMT6LCDXCnTGc/kDiKOBG47mHwkrbXoxiqFEXz4KPC4KrCo
LD/xAPENXTjLhJK/ZzSnbt6r3vhUvM3pIfDKXIsHsQPNMesbEJT2eF9Uih202GWwQvHbF/Fj4v2J
O++C91elujDz4lKzQev8w2gLc5GCTIjbyCGsnguLRYpJdzl7tPqHPcFLXRr/j2NfTnQWvM5sHcVX
liaRMulu+l6ZH8hltTPEY+lJnAIvF1UKxjEK3kZFGJ/oZ/I1hdikJLuVQc9vmSwTQm0P4iJU2uH4
1jP4o3H/2m/9tVqXHjCyyQqxdc2++a6epkU3mObv9QT5SxyluXnPMOqHUy95fIrcuA37lkAVk5x8
Cle3le09pA03QHyMDfeFLxqJBCv+yPd1FtxdZG8+z9HT8nFxNoBY5+xAN/6axFNT70cFv8Trdt6l
KZL9DMmeuxAYoV4h5LeLuoGmMPsppSkLUgHtloXus86dkiJhZba0nG5LeFNhLkAF0NMl2Enr9RUB
CDMR6H+pcv1f6b3x18KCMKklF02otP6UdnSWJs8KxM7VhCGDdOeEv2FV4W8/S0HkUsKBdOKAzMKo
mF8J2xLizMbEYSsWHiKeZD8ymEQsaa+yPKpZaITrT/f/GQYNML9rat1WFuTKj3lQC50iR22eB0+O
1rA1y7aXwHfUNXziSjwyf46FENuZuTXZX5yNS0IjlsNjC4wE3eGWSgvozFRXR4nxeJmlg8sGKjtG
WMLbiwN4tz4/PWbJqG6qOpcZzB8aTfW4TbRIlezDw7g8HuytviWqlHVHDzrFsAY28TBs3qxfLAAy
ACon963gPpNQcsw+uZf4Ib3tW5fU1uX8T6Wy1I70mXUR9Kn2qBNs0q6Ph7F7uWZ4xO+8XbdWIPiW
krLCiT58AUsJ5ygxC/a3RJVrKyKc3Fg0odldH3LcuJteNyDtsB+7FVvs3ozSY1YXehuQTr8uYXGt
Wm4Ypr4XFMjwUIPmlqT42BJk/s01jNRHdc6rwFf+Kd/YvwNjjaZ5DVZQ4Ap5E0dkluTrHYSe7uz1
ni+X3LrVe1QaOChM42N+Ehr81ZyR5pPlrMQ5UY0tzAMmhDA4G9FZAicPUiwLlHkl5n63r93tAUkZ
U7/hPtFA7k+fND42CP3R7BlhdZK+GVbrNqk4g4a5LSt1R5TGQzzWzcD1JkBoB/ozVu5FW7mfkDy9
bwQGyz9ZNcYOJXnkJubf9E0DHkI7lXK7FArA+rORLM6yGGcxHcqbejaXMyNgnhEWDgO6ArBOSzg6
4mvTT9OfsiNXRLrHTR2EE63S4T2rYblRe91j3Jlk+foNbZNy2PPtnpJls4/MXhJQL08oZ1V2j8ai
/FJIrAey5BbfFHpkXCWfgWY8T79+fE3Z23nXXo7Ekw/S4rSQ0wsXHN4mkGGE5lzNmJI6IGBfybJK
TXd1fzTUEQpxhgvpaBYW0gWGudiY9Yu2AjDvaCdGPnFLClSO6dNAtQJdUgMnF/WdL055kM8CuSu2
kpErbJoFxmVnsLKWLkp8EUyLaLnCrf8AuHuwDWRf+VQjKk3GE7ak+9uomLd39b3ocvE99tP83lUu
C/J0FTayaguTwoAdGBwEpkP0OPjAZgvWsOUjdP7Ojj2TsQe3Q0+SSdtEDjpWYZRZHg1i+C/x+kWI
ClyM3855Pj6bwjQQlqfvawAq1z8KFIo1wSNQBQm9C32LwVkpoSmyJdllvUPQrChF12ZETf31kFou
iAtor33mRhXVMsAgOeEFX68SHH4I81oP7ZkfLCzxDNTCzEeVe8ty07+McjoW6QNMidsdqt93C6dY
DjkNNBoQFQZ3xrWLhb6armA3MCWwUN0UrBrCi0QOiaTU9ENeitFgYE0yik/wru0rfWdrnPIoCeUu
8idWfdZzS/Ec9oQ011IFY+cbNsw8nztc2KTVwNlgtMzAl75JjDcjgLxodgzFVDQWSXTcMLazqcFt
jmTeiTGZD+j8qqNLL9A7qjbXv7prj5X7jgos4vdikmiVd/mzyoaLewTKb46F4DUYXAfwlS66kxY2
2MLsI6TuxUWeRJV4+dLWTEUKFJJpZBBxDvStfxjyfh7+QxJG3YFpNZw9vMbjbwGNb52cWXRogp4q
SAVRgLwAE0WY8DAzYTLepJXIv8/2AVuUoqZWSrGnDSH+p68mM1GKvlInvxa4RSFeNUPRmPr0dEqM
XCQM0HifbbMivzEke2gGq0keu9lwhrAMbadgakKeOVr8CQ57jOkJ0tmmDspRPTLkbyvsGbRwmoFz
tDr/o0hZx9D+oVx7TywgrQtJDtPmiK+zXAOzqkSYl02nVcMZAp+EkTSnBbkbuHTLShvSmOohdGHQ
Ir1ke/sBY5P+3cm6REWTriAO4wK0Ih0oA23m81qmpl1Io3tRP4skXaPLEtoqXU0FnadLTo5PMrs1
To3hNuxERrS35JiuOON/TJlTEbhqtithA+U/xVBFlt6Fzoffn/oCr9KK6jkmKtWSCNmGJHybMsWi
I9jmQGKrG49YziXfe7JXLAz++AJU/DuzdUBCm8c4rhRQVZw+LdilJKR42Yfv2fhM+VwaQN4zqqI9
NAAq3BFC2wBsehIfgEC1t63nfVAmv2JIB0drZDmbWdbm2gcKqG4a887bZtzAu39U6624SSd2buNI
XQGGVq/FerXCIdT7oKkarPDii2MSdbNqxDO6mAluyjtOYysLkdhXPP+9v0Xb9I050OMR1ZM15+In
5FQSSH4VrcPcC9f1m/1hj/WeJInvNDk93T19UK59Q46rE1KzGSGsnvYubFsnDz5FfmowMuFJFteS
9NPMse3lqX8XXIKqH9DnI/3IRF7o6MXyhkS6G3hSWycN2MA5P2C4ZFhK6gcle68Qtm2vKFcL+Ls/
Altc+Mmnoyx4tfLka1MbVDsqSU0OCqZRCI7jJ9fmqN+Nbv+rI5EDUhPvQpc0JxgBxFSQFxaNFUN8
FSCt7AaZGrS1IYFqn2NnVcYVe7z82hGhwl1sah07687NhOqhdPKO4MH9gG8AMamupkQCEqzXIisN
UkhTKuc3TplJkqD/cYAb2boLLVWCxcSzmvsdmd88l6FJ9HHMSZxtYBh3P6N0Jd84v7DWzGy/PsN5
+43SqrHHy9lWPYp/HLyU4dxZTnBwwrZqGddzOd9TMp2iK90EcL2gU/vHxPwvogwbMeQI9ONndaLq
tBxFIA+3Iv3YEM2bAtvlRwawRfRzJDpRPgqJofFE3oD7fYcwknK4r0SKwg35XtyXedRJGnVXniZM
Zy6ngQ2BLr+qqYDM+fnZzxQ/5b8rL7PiiHc0hpM6XsIEYe0qrnd0L/9AigyLlNyiyKgR1dctESye
wxlu7fRJs2E6mEdwzA6hPqTfs9QnvuybHolWTtT/mvIpJLnRd4tIPGULgrmuQBHvjDkv0CYDgqCw
E35Lhiu+yAlfHeH9YpnNYVmenofNLnf0S4ikbx7AUw+RKVQkx/Ig3+8FkTJlW3pbG9uqpCAX/L3u
OyXkshzsn+c6H8lJLQR1CsaxDfPS9BHRgvb6XG6QoYxNO9dF4E5kTp/5xhvsMCe0ZckVgd1OByNp
yT/vYBaDhS3ScMN+XhUc1SY3rok+Er+gR9r8Pz3mUUpQEylxvwOvDJFMWw6hleGpaSnadr+Q4sVH
j7BY3kX0TEG7tdcZeKyyj92V+gYvm13cOWoUitvM3/e2c60fKzRPcW5J2tXNu8/sQHp4AtGSaPR7
l2bNsU51F2qK14olNN2xlosMFTvUDv+iHHkLfmH714lbpuC+c6oH1IQKVOCS0Ex9RnY+g5N+5y7O
8N5mM8UFLJMefFQAKdHxvqpuGC5Scoakl1gf+LLhOmUmQ76R5lnBJSYAiqcOqkvjioKNgAhrZ+Wa
ebMPFgr3uYhNodFW2U1l8AN6KeMmx/3EHvZ6gD9dL37nRVmr2YTAiyX6IUm3YStluTLN9f9wTDsV
pUouWoFMI9o/GLUjULqYR2shEZ+QbTv5KKD/rnqjHEmD/GaFxHg6WHkUXrJdUiKynmEZO0KbNXYR
FncOJAKS2aHxymR84BbZctyWRhgglGe4ZmZwu46s07+z+r/ANlLfU5sVqAh3fSJHueHrNiRl2MOX
7Vo2SBXajoJUjY9fFCRHuny8fIIjMMk1/24sWKS5Z2nIIUnkJDtXD9AKlUYRGxEKgDEjhDR+JFIf
ng4qNt45kUpwzPLgr/PIFVh1AZTrdHMz9t+BD2wM3TBafa1Cd75RGrlJhplgi8XFI6ezfsLHMQR+
QnX9MmhUTmAgRYfwQl1LugYzPHZnd5A/7TRxF0fIO/iLlZoH68UFX3qMLitAjJ00P5PMtoWWiPrF
ixkMElYp3VxpBPsz0OZh8pALjdRzx5bfYdcSFTBGTl2JgJ9lL+6V678psctNPfkP/a5EReCPmebC
HPay0N+ZF76Gchr0T1sNcZ/0cAZ5uC+sNtIlBEDkRmIh1vtpdu6SbyS+AvC6X00QQZE+yXB/qapd
SkUJ9E8zsRZkaO6IDdYA2kck3EeXlGnvK00C1GzpjFHZWjZpZcjD5ZCSyiOurF3VJLmemMqjqKWr
2ZeIbPCYzmpiZSmPZvu75nQhH63biutpxbFhIsd2vtrM6WxQYzx+xvn5ccYOiWNTI6DVOg9xPrXN
Ki9zvYveSmZTvzc7ORJNeQuHls+Q/QaMirPNxYtpLP1/XfWJyiWAbG1czOEWwHmctzW9gcpoRZbX
1ZlyP1TQfYmspYWM8SelMW1e7vmnZXEwsQUKucuAwck9Xsw/5UwB1ARxrbaQPUiK3cbDVQZCXk7k
RhIDrmNHx1LBoM//vF9ANVVHCBWDj3/SJotSXCAlxiaYyxIveGZrZwTjJiMWUUr8AEjdCJUW7/Xj
7m/ow18dxO/txvM7yer8jmYBCBqgkkO8eCK8qxV7PYdnAX0XgkY69PF6v5+x3Vdf4hovuivv8qvk
cylhLePEHZYBlw2L8GAmmLXWXBUSAXOKyi2NGqtaw/ACT5Jrys8lYLUd+lBiD++Ely2QimSPhHPS
pV0MGidI+BlDGzfRncTJsEa4VTiFgdh4IguiYrxRYPDK0ecA0rq/aVrOyEk/wacb7cihAvCBPMm+
pQ4JPFmxLdpBTYOhkEeTC94u7JV8ZVnZu8HEZLyyO9iDSBh7yqdeYGysHO8LU+c5ZAdyAh0iM+i8
Hp4ROAu8c9OygT0Kv5UYT0Vz5l8+cW+lBczIypIlyKDW1osv4jZNQ5ojzZKVHQV+mqVKmrTTm5my
Gorz3FOv/2RrKaIE7kknigiRhIOTvbSVpc/m8CQYmTDwtsBLApfjvWc3uEVrUAcbv6gvxLaJQ6Ua
YGM9eZbYrDFATl1lymjt/vyiH48wAoR4JSF+ofhYNqU8pQoIb27OMyew0szWzITjxguuN8j+HOVe
0oSa5nUgIKaK97gSqRIyVLBIvDljiQAfkdEa+tZYjCPUt8AUV6ZVD24cTBWz3Kb+7W0YrS+37iz5
DpHDgMXi+fTrfSNc3pssoyTnD5c/Gb+Hx6Qs5e4G3FUETvgLFvw2pDeGd2HVxG3Ph4363mANk5Hk
QWTv1V72MLOIwi08cpVqRZdKryrcF6V8GuaptSprDfpMFOgDp3dtl/8NB/YZIuX4ULnMS/o5A2ZE
Bew3t9H+L8Oa8IafbvfY1Emmgsjoe4CId0Sph6uvJ+D71lw5VIrbpT9ihMGyBojjKRGJqI8Zx2NT
2ztIwPflQ1K2rF8+2Dd9DnSWjZ9ltLBQhiFAtDB5NhGZuW7CONOkCcovWT0R+5fuwToXoDV6/Ipq
lK4MCMT4lNe1UieVVVa8EbNCXoyGyWahBByW9LPyoZebR5q/cRgbAoVsUN5LJvVl8o829kXw/zAO
5jzrGr2Yrmhs/3MvrGen/rtJZx87zz1/C2w20aObRZDYSaqlJsGjYCN43lkdMzkr9kI0cwEqUnS8
iE9TyuhBEWQXGC9fkVP6BhBctJVqyTJULAcz6flxq36EUpU73shRsHWdGWkER5+hrRDfSJ82U8kW
YXkvjs3mI5/LNQ5dSxlOEaZrmaiLZ+ICN4NVrhjLvaqlo9j1GlW7V3y5QjymbUHdrz7oaKAococ3
/mDNpO4BEf5XOjdICp9AAsUDBYCrgcM8qp02pVHo5NEm1f60rHfC2lnoq5R8ZXaB5Ef0CZFtScg6
thq3pa2zd6FSMyQkIVgUwm/yuAdDp6ItJgJZ6SjNuottDtGWYDQSlulZjR+3dmpMsPwvEAjecl+A
GDWQPuFF+ACocr2RkqrP5Ebo6gB+DukYOjbvmAAB1CKHrag/hgKYZcKE9A5OIRHMUz7TcbuhHm77
WjtjVJPvg9EO384TYEpquNbheKi0XlegNWDiOLh0BBMKTaVIk/X6vZS3O42MTpoiih3imWrSL6cr
rtGGKJywgJL4VjmzV64R8VmEyAejl+wsr1jPRrOc8HJ/QAiOrGrUpMka/ETxMURfhUhGZCLikYKN
VzxyPUkMdFbrUM9wN2Igqsz3uTFAxVzJJkX8CtEwDzIsCeabgqeacubITe2fX59ygKKzNMDzUcuw
I1oqUWJgDuRqZZYDEcjj9stVY+LVswUtHCI1llSJ914T/OOklJGy5HaOfDDAejfsl8YcAqespQaU
f/rvWnWFAuThoh0+dULcQTio56MCylUtyAKRpeMSV9GAWcFbZeob16NT/niDWKqY81FHHuE176j7
Qop/B/C+SrBqFF3yJUInkW5rQQgDt/pg6GE4sgz3grZRSnO/l034gEz/yTg7i/N/hs1qGNgxWtZJ
R1BWwhRFCVopZkqJskMIJfkop5SE4ypb9w4iiK63X7iNCJPYPQ4eQQ+XNhxrUt8/YxAPwnmsMVYK
LJOox8+FUjQIn2YFoXuQT7IbrWwezJr7fr+TkTMLNmmJzsjkprpJDUJi2nJE8jghUCV+Me44WLZB
ZkzSVGaF5uwhqBiJwS5O1pfwzbL2sLO7cVClFet28PXxQvkoKu7lixlaoYgT24NLmVyFW4lraj41
5eZFNhj4GdDDWLU0RDeL5wYfSOWtOW0vx6MIO/8pxwkCr8iLnjejHZuhdRdAKCRugwT2PgGIDXwM
EiY00jEaF8KH6yonKqwEtKM/eXqHR+044bfv4nnDsFcwj1N7L4dDKTahsuDf3n6PCH49e2v0RUFO
zgDYUzZ8qH3PBIf2QrzVfADx9oCVduhJyYsfD3pYR1gvX2psFNgz3MkjmC64fFgqKx6CqNp4uAdY
Gnem7vdfDdvayKG/j3Wsh2BuGtLcCK7F12Eh5IjIkLWnQfv1GCRHfLLKCKGk9UyrR0AURSwIPIqC
+IYpUPANLPcmjAxsPNcvCiMyey+1+hVQHqKYFmDpOrleqxpSW4lyhTNTSOERX8qiSoDjVkyHl1/H
K7vWCaPEUnqX4040Uk7BeiAn9aj2Cg9STfS9uXj4VaglO7YmnZXWpaxMQDRpSQLFQHldNlz6gXN1
p/Um1ZC7PlLWEpGMpvO0S4WSSJc9zk5+MA3gQutn4iRFieoYBEHas0l4VewtWyvIltJU9AQP7IzS
vP4udhMNzxIINxDB0TIqd1UJMXTbphWoWx281lTW1evtIzRElATzJ2W483mwsnpPT2pZs2ssJDox
n+oQj9P6lUb06yMq9t8yO0gCDnRPr+K6SgjE8A04EcXlH9NTh7jT2lftO2rDpAMx8eayOwPyr0Nz
lCBea/JMLsMwxTiARs1ygSMgqHXhtM/vlz4qUvbuPsjYcRo1Bdcx85w5IhjFrQBDPQQdKXKy+PiV
acSg4WbkKGb9/OE+HJAVfoAjZcclroQrLEotSAMJ3kll856X7cvsYj2LN4W5Q1Gar5Jt4zv8UOYV
lQoV35adhr7fbIVG+c5OXMxeR6cEBjWWXFynyc0tqYp83qkNTvaPFKJHEBWRk5cKdaDdEVKEzA8e
wqI1hmN3vU16+kwT5lNhF3FAZF5KaJFuu9aEccayM6pJAddsexFWdWHiWWDkaHdYDTCvCa4GNw3x
71Bd+8tc9aooxgJTXekm41NUQiquSJ3K2UVr1Q6EzRvFz/AL/FYjFLPBlpafZ4fsJnP9Uu1MB4Yp
60ELBEIkh3C4RukTi6neXJTQu9JC58ganmAy3oMkX5f5jS5iOxvYzOUuyhq2bA7vRYBYKWeZM1Uf
Ug2H85DLVcbbCktnNnui8NmNxpfmQVYgk059K7zdMR4DmIPmYFYd/9EgU2sQTWlzHV5K+amH+CSj
nEbO9hYSXULW8fn9tmzRVKgAFAtSCu56FS8Cnux2V2PZWCHw79BKoST9VVLlaxeSc2KjDg/xDdJx
hBPErFMWwaO3F6fWaoKUH0a3i03scK3bGyXeVY3IitxCfMzbddaCl48wwafMJwky8aLvCOU1872f
X4T/OSezqBWWIix1sdEgLTvxL/H0VOAZP/R25HEtiBtFJU8lhpnMsVXKzgwfevYbXCntMFQyY0sW
wpOVSc37/tVQXetKKr2nlEokU9M/3X9fMreujgDj/PElc7n6Dim4vnz0mKsybg4UEkCa8o43Kvs7
8iSYx63J+wyA55NjC6ihHWnCKQkDxDkVjOYSMb9uAjLK2XVncCajheeWcGcVcProWS72OcMscYdy
OoArjagwNmWEmNtGLljM/N4CNUR8R0Xpf+/n08jUDHC02BZjXGDKMnEcFj099vtheQKemNav6QGa
gApxLmgumZFpf+nqymsxiMFKzPMg6dRKxMiFNI853Mw90r5772e9Ye65VuIxUJNNsg7RPopQKtCp
QW6/7KLQnpH2zsZXXcQFTE8gPwvH+264qqnLtzazdsrZgH574oaWlhVKGc1BEpbo9g2n69Ryelik
VFkTk1L77QCrEvfHg7l8k3vRrBu5DiEXMmhJLIQXXuLIA6XdkXQbsAUSPhh7MEhNdjhXnuzWf7ho
vPi3KaQTxf8JsrnntUv4AYllyoivBkOFhfJPFQiQtcgh53Srr/njUgYonhdtwaWnXwqKzo7XOa2Y
vBQJ6a7x8gQ9+6o0m3uy4Av8XBqMo4AZlpm9TiqakiMQsOqBmga9Nfz11Xy2AnJoU9P4djntBlCJ
c6sq3h3/6HhtRiHwvfQnRxvqx9vzQc16SAF8Lwbvp0RZwfe6rn52eJoC58MEgHw/KFUszvd/k0Zx
ZYD4wAYkNcNEJVxnN1zWTP93TjK837cFJ6Cr+r9JdEQkYIe6XbO7UhxWfi6vcT5Do39p/YMaNfbG
kWltPnQ8QSHXfV4SUE53X0zlDNjTGFRm5ZisvHJxewQDep3HVcjNsjcU9opVqggFfxA3As39sxwW
hGvHQly6YIGWGMAValUfnMoS992sc0lfTosqZutu3N0S1lseOXFwSwjq/ae+VUq7dUFrUi8wPfUK
fOmKA8f/CVDSWZlzmWN0uJq29Cy7dfboAOfRioaAhVv+DJ8pJ5zedZjmLeD3EHucvGYuMRi0rKsh
5Q2t7rVPTDCUd1EmocztjNXimiklrLzjOWN+2jfE21bnCxmwyX0Jo/lKVRuREd0NQRUBQWOaswZB
mtA5Oalzsci/CdQiaqNtaBj1tSX5Uq1u42UxkC90PXOTMaDbp8um3r6R8RG8IKipWNz3TUHfHqo3
92fIC0YZUP/sxdycRZrMnoLDFlVxo8CHlKJzFiKTu4coZm7WiomZBcjEpj3qJzqniBeMKkM3ZgzY
5Tmhifs8g19ceGVLuEhxnwspodau682aLI7tGcTt+ylPJoTaYTaaSCxBKDJ/N0tKdUlBKxHh718B
vkis3zPorDwQfVeI+Qt/C9+7D4fvastleLE4U1hpx60k4ueUeCQUj38hrjY2c+FfF9XkSUYl9Df3
+diVCxUVlVw2P+XWzKwuEzOweZeuzpvsn5bv7bE6bnS1tg7ls+4GDJawFxzGEvZAYcg4gSMKSj9P
itH5rvEnVQkJAzXtXLFxUwr6ho9LL7Tz8lSu4ea9aTZmek0prKPvHB+yVFcxRNFfzQ2Wc6lD+XsY
kt2OLgjmrAYYyNZp6MKfKmPuRZr7A8A4ZF61hUVXOcMeeMaqRdVhRJheBA1j/BTPL1cHq50hxbb2
pOqYxpdDLP0Oqu/trCDOpqM/VGf7q3ZcX6uu5oIGuyWyf6iBWLTxwF41gDC2XAWEUB4KNvr/zaXd
x7tonNszabbOekdt0Y3FNErTDIimED4isNButsfzJvQDu/G806oWwoj0X4WcfgSiSBNRZd0gdj00
+mwpaWUbJuoiILCNxg78F0PvfcNYckiUzcCHC8C34XxVL90XwgWXjeZETdDknotzHZvrWQlAjkWo
0HidS9HVrwrB+LnSHgaBzyKQ/5Iw4xqCi2WDyhgpd/FOoxptfO8T/zx0YLwpI/g5KDyTFxKgWaXO
X+H3Ms0BInTAMhYgv3hCzDC0xLyfjzssQA7ev2Cb2DWiLDN1T3xQ0cyaHkK/WDrXvXZcPaBQuJee
mqxIkwtQ0iwS3wDJJPzS6bzZxRydvnmA4U8AWjp5aJttye/gtXkgAMx/7EpcXvyZmLW9E8xeKupM
CVDKiohGgCdWL08fIjxa7KBBILbJMvzvh1eLN+ZPtv9BrPx4HVnKalYCGGetCiatoveQD3GYiqtE
aMYPo9EW0glCK2NsiYSiHE9Y4WJGlr5284al+QMfSf+FJYwH/QZt4G7WJfa9AbP6NXx1Lytqsar7
v4rLc2M4motIY9KbHRcW/KmVRUC41zS6R8UTEmYTfNQa7jWnjNJtlSsfPxAlj1dy/5VXrtzbx0e/
VY6cSH7Z2mcXrzOa6jpqLhsB5IqKo2GrQbh/IWSfBfG6gt1eqI7uDZxhoG27cF4qBq9I7ChIBZMP
VrUr/dy5tfxiH0cW/0DbyneEWOCsD+oXUQ6W95snpjcTrYFq8ocnQofvKV863K0NUUT2L+X9bS3T
vvd8moI16YntilAyCdtMz9azVm+ZrxfChurS7ncBWj8/MFEgdIaDrq3omsEwmYzWJVOGSPz+01S7
x72oYDDRlS3L8oYnVScDoSW5ws0IiF1t3E8JnOood7XLj9MNHUooSwCVw1ArUdXN1+PzU8ek4jLj
1E6EUF1Iy5gCAINmQWoOvGHMARRcHEQ1Rc4dlY7+vodgzj680yn6GQ9NN9MCYDE1zP+EZ2zFp3Ld
V/TIQSnD7MB0TX6sR7v5D4QQuwdumV4aq0iV25AMoNYDGwOlhxHbAd7jtrIDtt/96E5LibfyufJf
SZQywRJymvX3YyVnPDtaCJtcU91uy2VlZxwJ99RHzMFiV4GjUKmziJh0jjQ+gRlcPTa5yo2PXq7a
YlvNK+S/GJHcGvY2KP2RYQnGTy+pbT+bpzFKgMMQ5xH/YVM/UxnRvq3J+hGlEF/IX3aoF5PZfzmq
WzpJNuS6UtJlk1Sd+wcFjAVfMByMEKa7gDUzbGAJXfvF8Z4f04KANFrQDN5WcD+IYHrjthate2xv
09N6wZjA59iE32di+Xzc8Rl9CSs1dVq6C1Urft/2nlJv1menQh3E6JUJaq4EthlbZ4FkhlaVomon
M+TBhtFjsgZxp1u5gqLMSQvhuI4DTnv/t4ZA8XQT9WB8FdUNpK1Ye29i7iZkAR3IFHKbWyY9sOe4
nTqtxz0A+KrFs+ZC75Rt3MM5iRxpl110lh3uD03R3LepMXqt7Wufk24VGZ8aacW7s68OykCPfZ7r
9/QTeNMhIECcxyKT4LsGV6TFtcv4FztftMWB9TbgD6jGyS2b91mOzP+Ilzcn2poIZODTbvA30bWY
hkZ9DjL4o1PPCt8t5JjaNwZOmNRZBMBNxofyEU5XxJjMZR0JuetGkI4sm3t4wtNyQtM41+8ZE68T
ZU2+1353BGDKiF45kxTnTGJ5OzpoeXhzCsAWMHGwSUll8N8cCX0723sqrRHs5U2KamrrFKKmL9dV
KCgMk/ZMUt0gwxVsCZNKeXdEviKMJo/Rsn7VfItOUwQaRosPFKFe9kyIt8y/pvrIhGBI+J598Y6C
sdAkVpA7oz7UeUXTe13cQ884s3PGVMptw7RYKlDotqMb4trr/IGEFveHjIB5BNCQbisEZVapTKM2
qg7Dh5gnLL7+3HNXLZdF9Xa16NbRUW8h6ojqYOQ4hzLqWbqxH4aSke7NJIiDNCXt4X7sKkCX7Ib5
BRmaeA18iODyXYM7kqjV8uDz98Vy9awddghNNCSzbWHfgE2deeu3gKWgfOb1q0QDb/Jj8KUhE+8c
LG9RXUnawJN0pMaJbtK8mDcUQ0b3TmoZKlyRpyYNKtRamQ84NGJoGSX8B90dAbIiExFk/dTwE8RM
McHwYE07oye5zeLXAz4W6jCKOFAYWfIMkEFhNM8GowdBAbrXRtelkm5TuU9M5bV9WcUSp1EZp069
yamlkOCo4WwK9fK0RIDkJcWzxW4XcWo4wgWGmvcKZ3ry6IXims1qrDGzcrsp7As8SNNeGscWk8Et
3QyU2siLmS14K4XNyA/ElR48eP2jZI7ulYynzqzhhGCIfi0KvcAO0B+O12xaZHL20OPtVneqW4VZ
6NMW/nloseElj6NdgdJdEeCAEAeZw1nGghsiGe3wj8Daqd1Xg/oULXb9jA4VxUdO6sjy6g2sQJHK
7N2WKTt58fS5GZ9xpr7iHqnkT3FyKa+kqpRbcpUzCxjgldNsLyatlZVsPkZO3bkSDjcR2b5CH14W
S6A6scVISRrOpRmQNmAYtoGGPyCGFvVxiQGaFnVmnN96y2Tfkpu3ymyg4ERDg4h7F+lcBnj9/hAL
2lHsWCezesxe76BJQOf9w/pFcGzCJl2DZ9s6SQDHhgSqq6XI6eDAxTxOeMfwsd3+zEJjYXXoBAmb
HwrsyNq464hs36EQ/XQ1zYtbldk66BQqbcA8RamquQjg9vuaZv//Yca4L7BmZ2ehf7poKvkFoY3Z
t2HgLRw4Jkqhy9h0rkrRfHfsrZxM3Bi9QnE8QDAFWXwBj5yGbbBkdswQMyaeQDCtaEHURNqVW0/Q
vvuIfhM3qWSzGgUqKKFVBS0q6evPfIbXIG8ej5IoBUWfIxEmBNiALTRokIe/19lPCYTJX0UPgkFs
61x5ZcSjTwQy9FkazhUl4bxn+ZTHgyiwZsLhjh/SISTPX5Oqf7XTB0ORye3qUOpFvcWLAT8FBCZc
4Yk7XyyiercJENHphIGhaUYtwUV4UKIOCQeeHfb6m+E6lboaqf6cDBdMnk1qvEKQ7ThHWlTgdleb
cgnPCPOoOy8RS7hVElnqLxTO7Z0kxTm7ET1ZBaOy3PhYw4ovjp1q6holex/JNUQTmSGOQP/czzVF
LiMkfnTiMFmuUwK4OCzS3IhtjbPAhjxHet1u7eMCeTMuRGEDBRbolVup9phRv8+70y84WkfbdF37
++10EdP/Hd0yW7OBjA/SflbNxPGCWtD1sotXG1ZDAJW81YhKrbfogR8UpcAuxbniroHY8D4XrupJ
WbqqPDHYvjmpId+o1LFWPCherro11uA2zQICFlnReW4O4uY7s6NDAc8E7ds8vRH/y2oHV4YIpFnV
pTmNxTWEVSEV1YkeSKkZXD/XWM7yXOGcfzmfodJd4rE16xvD3q2OSKqClGjvHc2wLT3wF8I1V0JJ
s/Np+1WQXg8aoClGkp3BeiOXhErAphl8E2fBeDmNBsWHOyGzqTRNrTPsF8s7y/bm54SRyAsdsJpj
kItEyDMN11RycYgqNrZ1bbj68rEbzWwinufi2pvJpMFTFWUkLXD7I3GbAT4XvtUXEVVPe9FmJPBj
Uo9o4gvHQQJ/w2E7wiTUVvKHl46sA8KXCDPuz+L1HAQCayzvd/9EuEJI+i5HzfqAjbxG5o8Pg8Yb
Ex+xHyfb+w7tQmPtxNYb55EInrK9mA2r8C3IOiBPJ2QAgg3CTf5dbLr7uVzI5E1+vltDUWFRYHfa
HlwIvZdmcOGPh73TOBifQ0tzQTseF/KRTI3gWRaAC/gZkxF9hJATrQzRhVFbd0UAz7rez35RnmfR
jBtCKWlFRmraGGfmaPsbixRRbAr5kg4LPOwBIuI9OmeEqVI9zetO7e0yg2XXTkkzuz7yLIikE8Rr
Vf/UmTb1QbYapKb7xF15uT3FiQHwk41fpiBHFLF/JLDcgoeIE+fK53mApq5dHwetLPv4bN/4Pr+T
SF6Ze+lB/s/zL6LtpsFWe8GRr9Dku2DHidxyYDXtNoHE3N/5I22nzajpyzfBjFXFlyX3xtXXAwIC
ETMQIfJ+4EhtskoAPuuSPqdT7mOpOy+ZqY3wia3f472Z5O9cPtDH4/oJ5pMYJSfrJOfGgMgGuU6m
duzG1p8QJB3Owaq3vNdh+o8FGRfbalRsmWh5a4F1uHmDG6Sos01YVoa77+T9flO6L9pgaBI0R6UL
emE5qIjHfm+TrRJAL7YZmNB4G//plFKiTJNlQYpy+eYYM4NgCo7hh0lPkW5W3c6tLBpTAcl5jRjN
IUoiCihhROQcqBxv88CXu2ElFgj2ZFqnP15w8N0xQpvdSUDwIf7Mq3pxfNsycySR3oGWP91Ducno
o2lXogN2NqsXbGySiwDb6mybcWW5n13T6MV/ymOiEDOicfBmD7erhd3WBHwY0ei/q0UX7XHXxlOc
d/Q+RRew++zWLKFE9185HUMKWspApQTnmq1f0nJQkx7S3hflHWL+ZycFByQbV0JtZVZUSp98VsPA
0oeeuXSVrmASd6jde5dF1aSjDkf0vtmOBEbn7PNNXFhi4xUbpx9tc0O73tgu7tgv42rfE1gT0zU5
gBTYpptcYsoS/CBNUKPlZtK3IQ5Bn/q1QVGGFvRsdf5zPWMZ1+donX4BRsO7Ds3Gabi9PYQNrzrT
JfjmWGZbNpP9nkV81RTVUopsXTFekYz6v+urORorYvWz5WbE4Lbt1ts9aJOLWM0GkwG5V8j4O1yr
+4jrXjXh8DOjAHJZmGls6cK7iVyQdOBzoEU71BgvY9QYPwqCjxml6xwLjzTMX/0KofMzfwnVhLoD
ynvXI0D/iLYJBSrMuKGtvQwfvRZbTB4S974guI0bGGdTgg0fmYH0UNXw8/aT2cKwZtQEo6iGGByJ
ZWswS31Y3HViH9K4uYcz9hl/0IzQZxHCvcCMD2KFED8g2XS4zGpbDumZ08xjCndOOS6zgSWIJ0XS
9iJAUbL/ddCOOie1XByJkucA0h5NGnZb9XLJNCWGlK83tmNh3S0lH0fdsngN1wqnW69VlVXlmJTc
z9h2PlHekBraiIA19eGc7Xwq1GUollUy/qkm1RWWga3p8RafapVVdpJF3MKuTDCmh9sDKg6+uxgx
RHJ9cvmrD9qoHMS868ziGjBZr2k7TRaq/L85fnGk2ZLgzXoqMada4CzwH9wL20ad+0yRssgBeQ+B
dY9AFkv5Qfjt2kB3pllHJbmeYeBOUEIZxJMiUnKrDBRg1OHnubovH2pXrtTYcUKBADJbW0d7qQ7i
A+tSADyIfZf/lwu3GjoNSzGpN51yQd0Uz+2/n2lMg77Vla+ekX4jJDLAYAhZcC2Xcof6Ng388WkS
loGyUBqGabvQ5p8s1kJmmIT0UTkTrcpQLMhj+swp79DFSK9+LPx0xk9SLRGBwKSceY6aiZAFs2wr
dzxbobXKR7C1WA+Xtdl6yhWA8Rxva6wFxeAbtOloUpJEwhRTaxRzviwEvrShcha+874bLBOj2NvH
vHT0P6HabzMITH6sJfiHkr3fEdCFm1WmWpai64LZ2u1t5J4nW0UIrkiG46OqeSnCGxezxfKwqpPl
CgkhrSiaGsLtif+XZoVoQoKw1AAnts5L73LGoextE+CtCxZO4F9jq8vCLtRBWMzmmANx4QXLlVc5
OeeX8NGmUEfR162Odx2VMg90hVUrIOF4q3ys59JAyqVvookH2WK/QcC1iNNJ9CNCskaWAIK26Qcx
VGqAUe1wkduDqaWVNWZYrBlfH8OuLSU3oorSMGsqs1M52Heti1m2+PnPuwTcgnsaTpVxARN4QXya
w3JTxBJrtvM1Z36Ob1sbOhPL2ZqxNd3RAAwi0GvGTQaUaMf6rUM34I5rUTCtueVo5IX2+1O+uBmc
5t5O9Bad70bZEh8bO8IGopXEX1qwnftOB0QsL65mWz0ygqKIEaYpGiFkhI+nUQ8uCvc2UAHlN0ps
e93Xy5gVJMhxjAJUf5Ja+IXxb1u2C1qzwgtqgM2AUbOR0o8vdlcg9o8ZldxZWtR3ysnWNIRz2QCq
QXYfNVEgfUgEM7hCT2F7JhLo1tajn6imtxmAu4q8wQa1zfsQyjJkF62+rojNdWNpn8Mc1a5k/IaR
pEXieq7AzMfB8nvrmcopLpPfAnOBQ8QWrOpx5V5Jar/GZ1ulAv9pSsnm/fWDBUvFVaPuK5v2ytb5
HQ2jUk3DrLaphbYK1FRIFSpr5X3/1G8fmAZCV9R7U+oXUbqaCUwgyel2+PpEOXh6Lo+1akjk83QC
hLmMJZkQn95oJNFP6R+R5wyVwa22LIGHbgCPAx+zQlPWYcsI+MyDuClaXvYUmXF1WHYfLBo6Ce9Q
pw3VNUqS7SscinJfb5dH3gWgdggq644vviNs+MTUJ6Dbn7oh+N/JRWU+xf+cL1o3vZxKvNWpkg9q
zirfIKg0VZiTsyBQ/gK236dWQBvOO4VbDjayy6HLUumd2X055iMI2LSa4L/norQZguzGyrpj/mSj
xWgM2GCsF9GRnYQW7qW7sQ9y/vZEkNKr+km+IK1XZ0AUYq7Co6t34KgGHXu1gCHzWclNtBGcKnb6
5cSyXJbGjiaQzZAPkJulsG5BPewH8neDkWteIRjrT/CzaGN2jQj7pXmE8xiSoJKdWGzXOc3+zEeI
zGQdpppOp7FUR8vAtQM+xicD1DAudkhe2KVW8E/BC3V+p+gB3AR1k1WLYwTnJzswt9bpLv4YfUsD
RlHWzcPbvnaCaF8vVAIKCMIULqxi+3D1MuUzp++rPAwurM1/Do6CF1X2uZOYymxPAjw3cLOZbERT
RwxN+9DHhc3ZSr8DUI+p+6jUBRQfzoXdHsaSydrhF77LGJvMVJ+Uk7QEFRD84J7ZWOK04W3kYi4j
74bbHY5h0Mx54r74wMJi5BTfLO0OBAXk6DKHNEy0l/lHt1ecZ/jZIom8E0J5Z9h//dKsOb+f3q+p
D0h87IrnIJ7UyQu2n10l0YBHZJT0uYkuGVHnnZS1Ysian/v3L+fsMhjWiRwZf0cK9todmltzKlO5
kQEbf02elJQ2q95p1Vm8q4ktHmJ7jDGT/97gQBi8Wm1qNaHecE4hA6mXbpc79SR4PZGKUUT0Htub
WEKiTEHerepBHO6Wj2ha28wx9c+YrVdv4ezR1FhqajG1VkiKX+V/sA8aE+DBLUn9cgR0VmUDfWgx
AvZXtz8C8wIzoz2S6kJbBwHkrui0orTR07agBShR5xpQXb2GQxpj+8TZN4XFhBUh9Cgr3vaN/D3D
CXwkcFaoq9edRY0US/Mkw/CwG75RKgY1pLGcewo4C57LMNc5te/9CyeT1vRJXmuxqIz7SnkogV4M
6LrZ7d22TDdPTMkxAOI2kJBZ5lVObFJQE0U5bvagXik1a5RFvAmjg4EyNBYhaBO1aCD5tyV20wtD
YvWHScuoZms7aiU2iJQE4K0n6CO/2cjl/QENYxK8bjBY5QiQAtqwZ016T+uYAbj0zfT6PP0ClrtN
tgvRuUOjAx5K2MSSx8l3Hin9FLE6Mtd7yIWHx/VJT9YL5vfTMrofz4+9fwptyh0e0m47AC0w6QRw
MQgUTMt1NmUtq05vKP3uiuQnbHxrK/HaDP1RmmpFQeBoPRVMOQ4HKO+Y6GVSvfllSeXPTLJAmgMi
Y4gyCaYnpJ4NngNY99M3xNFl0szEpC2UsYk4nwV8+IckOJTM4aEKajgB2h6CYONpDMDx4mfpNZ0h
Yh/+CJvNs1edCKsuto9pfjusq9oL5i+e3MwH+iA5a+j/IDV91O2KP6V9VTZxBo1nzj/gZrKVYmrd
m6FhPMlh/P081yOPzGgsA7lvePjxISMFCvrSU8avhUvlxDLbGveML2dJIikH+HQMEgETzn18+HEf
3P9n1MB8uGx3ef2chzvfVehAgXXkDXdLmIDliBoKYRASMwWHboL6YK//zwQj1pdrvw/TIA6g70u2
FWe3M07dqMHnXCpbUHc6vcj5EPO5we4gFon+sxZH0skc1M4qjYZ0MoPCWeCKHzaIqDgXuzs4/cnz
DjemUOxpdyYoR20Dour2s52Sw3fI21CSKcJ5ACeOQSlEBSVdxKZblFeasiaEsa0Xh5OLj2kFcGXm
AQfm82KpQgJXwPTRSSrF1EZuiC5OAV2bptDsQQDAi8JWj6ts0gJGiuDXN37rZLM9VwWY8XpYBKUJ
2Zk74MokcCp11hIQGGDbOjFc76T4ZK30J/LhQMhDBM1eJTFDHeAAtEACq4JNPtvpryK0ATEeVGUY
awcVo78TIsJgCXoOrtlgR38J0+cApihFdNgzq3blMQOaX0GE9HDE83XqIdqD1Bd+6Wcy4j0m7q5Z
5F2RfWuvWStEdI8cCiH9ikjqki6dtZ91akHTy4r1L8W+bcQQZo2SuN64+C5asZEMixjhnmipR+Ft
RAIRkq1U3TqlrD2LnLLxLNU8HXzSaGqsjY2TkV6IwS6UM0WCTgVRdX4yPo6Zf4vOVtbCBVrXX6NV
HJIO9BeA9ROXyGC2rFF/oX0KRashU8pYODI5x9XU0dGf3B/FZIMnzbnFcGBTVOu0xC+j72gAXbWP
IXinJ4/mHD4WEczGsnRZ3zpN0WogKBwzjcnKLjcB3zpV9r0T2ndxqZ7rH6bwesw7NtwDNxguDPRe
fB5NAi227WXHcS9O0E7Gkr3c1DTECdM2xQ4sIjQLy9EVEXC90Zjo+4SRQnf2uFEcj2UL0KC2Wjz3
cGlPkyXZ3/kx90eoTq49S9XFH9UmL63fV60cTq9KVe/9/dZtog4cdQYraUIHltRWuhvuQIl3xSnU
xEfPfh8Zs7HBKgPCPvXZILl4yTr06tBAW3yjGfHmL2hvpL0VAV/chkw+r4cwaLvzZRsoZ/vDHpTs
vBeft2L2UsBWNGb1b3U+YK+c8aF+rQ3uAirx1qb0gOvXA0iYbHvfXDXlhhz6/Ae6yVLQjZIyzq14
Sf8rEHo1HhS0HnQ/waj0yXBWNQE+SFMkakqYBL0n3nLHtBlTN3z8u9/5QmpK3gG6QO/Z+cvtK87q
UJvszrJ9e8XwonsBdVkr2FrrCkIDsNdvucsKI0vX4B2QEliVoXXtX1Mshd5LolSHi8lqGs0x02R6
DX62w0aj1qwoTiiH9y3gp3Omp+M1U1dVmAnx6LY/1AQpoxLASzWggH5+jadncxRYhcZhLeF6+Ti7
9EJEIvlvWUXMQucTHQzZiKPBoZ67ZMvvtY+JcHaeMwEpaek+/Ggc+OU95DA56r99AzBJt8fblgdg
B3mnfCPNggZEaquxwpK3ZHbg9DAgBpcEBxkClCo/57P0iwJ+XZO4Nzoc18yEjTzG93C7ohlVvt45
MhNYgvy5dnLz9TgSlJUUeFzIuAANABbxl7INXH+ERB7XnHV52Lsl4ILUJkha8EzWgYvvmmWBnOlz
EdU090Chw/7GPrtDVOecGrW3fxrO12iUrh6hZrm7r8GTUl3G7Vnvgz32pcVS4ZvoSkg5hkKJ+T+Q
npWv0zQcAOeiuFHDj73atx/BWjrVgceLyiDT70sz/HCtvdu+apYJiBlZhFL/RGFEchyJILOQ4bXR
1pQiJdsqJVKxjtwpogFDH5F03CG7YAaElg2Mx9ug3fjjiKyae0dAaQVAXyIvHma7BaAXETkWfOH4
JbRacNNCxTCDVwLFBkvzwa4xTlm9L5x181k7vZ6qkjsxE6Eaye/IY9nVQXMfxDD3govGtbxu7yBy
jDlhOgepDaTtYAM5BtOOk80NqWpTzGHH3It9/DB0lENpBhnu/ieuSNqpXDfG6CYa4o/aCFyeT1O3
wd4GFIyIhjRe8/hbXkFsynZ1JcM47hZ8xA3wkf2+8niy/GQMIJ+6dnpFm1TWadE9CdEGtuz+Khwl
rgQ+1OGqDKRHi45vAQsWO4HUNWWhQfv9EQetke0YglD5R77ezVTCgLOur4+v8zB8UK8C4Vnl9ZoQ
0s6pPp8Y/QGihZPiNJsrEQwQOJ/1g0GAi8JdEGwR965DrTAlVzz2TwVlA/L1G8a82Ag0RRMZ4B94
qg/nFf+0X93F1EGVcA1utNXFuQwyxn8V59gBMCQpPmC9Rx2nkQkTCSUUtB52gHBPp6n8PxEjowXY
31Ma0yC5ps6cSWuPJCMTAtkdPqsdFctID4/UFYBp8WAHOa9IdXXtVa2wGkK59UcD8cOnBZ0pX1tO
Vt1rrXvlzYmF+Vgc1WGihEFW/UltwbL/XBjzvffljNxW3LlJlvfSg0+p5Avlv4o5cTb/DvyTMxIm
llv9hmMONfEVZxY34lpHpY9/mUsrgq+RJ7h/APb/j2vPyRR2Oowt1jx09QmPtqmkGCRLgJvHUDzV
m0QWxyjPLK+mvxNTXOjoetR/fwWHl5hSMSo6AgP80PDIHuE6X2va+tuJgd5koW4nwZuUTRQzIl0n
CdbLC9gK7IXyjMQkyf3NHjmD+jrk92IVfRdQkmFYhKyWUp7QpyC/0W8HbPQLonUyQt4y2sNZm1hP
alBeG9aSNPeQVVIW6pB1K2y/kXm58fqKnKGKnr3TtRECOL678wTdpBBHrTWlUOVeMOhpCNQt78pC
aQ8xvfwkEwLZyI4hmk/TqigA4ez2hasoHa8hEkyBl02ChwMG2rZTVGlKBqa7RmyQP/WciKQZL377
uvOTWhhAgcHEt6ju/lestggN/uEY4++OKC1hPxEbD+IdjVCTIPJMtUV0n4K1Qz7buOm7P9jl19HV
2wqOJJ9Ou4oCfWMIN/rPKIAbulLKabpBaAvH2kVgK90vXZpvomuSnmo9aFEHPbOtw6MeNo2PKJOm
i12gKRpMs1GkDDy0xm5LOoZSp5T5I6rr4UtuCqnnwX2Fn3U4wz9ZOwyQhfqp7gs2G+tiC4r8EAYf
g6DRWuVgVTcNfEjwnrzFvSLxAylGI5gho90nmfheZPhEuLC1j4nrPolicNRJJUMVetW5B8hooZi9
PVgGYMz6t96tkAQFxhBviTLYWYCiKConZPly6BL3acTRKw5/KvEMyD2hIj0+0Qulq7WR59Ry7BsG
kQMLnE+4yTBX4fwaxJPwwG+yF8aWUIb1aJYcBJHcFjayROJN94frE4qVAYe90cpjN40NXmBgw5A+
L5EfQsPhAOY0Cgs4zPaRxSo7ec5dE1j9MxKt2RdjAfL0n/l1SIuLUglpQp6sGylcL+fiHu11VU1W
z83VopJMNQlywrDnrF8+ZA9vi88Ex1u/HcvQs38KXkPgvj6u1ufQDAS5LyJNjl1xyiGBSmsSItgX
KzR+rlLYfpgJZ5Oci41Ozvd9WtYMbNnALBCKpxww8Kph5xPrEh5EiXKfOH/+2ZYZbMNe2ydetCCK
mKMLKAd5/rdWY7tWJnTubh98WD2C2gGUyPpwv1pxYqgwIm/J8BeLQ/LU1txgVbDRjXAGj3buVi2i
lmxO4yLU0kcm+ov70v1tOH04OL0qoHBHwN/Ko8hsGi8H17602iPX0U0YKCxfAbgCV+pboO1/Ylo5
sH+kN1T5Pnbwdc7yDtmKPc9Pl184RLFubvNZTuCxRiQXf+F9NPZ3XCRI5o/tV3KRunRWe9HT7MdI
yTy7P89uIYzAPy91MSYOgamuCtgjWgZDD8dLq1XlHNGg6xcz9GJjM91J3gfPoLLcV3B/HE4rIBOe
ewRRRqd8SdC7l24W1e3t7lCGN25lUpmWIhhcIo75qEhGBhvJoO8qGlZPNgXbE0Q+si4Xa/ckxd1E
Bz5KKUURod5VY/4+qGxZRVxcBsPqqEH98DQhJo4eH11B+waG2TDs0sqKOavHgz9NSaaaGABdX0Vs
7gxUaLTfJK0GZ/3U1/7thj3BGT2JZAf5Oi4qmsNdbBYPUfdSQzzIHNugwDC43sVlLvuuCbbEL+A5
xE/SVt5bhe7IglkxeuOPiq6BYKgHhYlflSf2AP4tJ5YzEZxFk2BG5GEWG1hmmJtniscxdpRmMBr9
EvnoPgDlAJCw/pqvSqkqoDJSLRRApLNstN/qtv4WiuJKY+BrpbTIcK1mXRJzCjJRFQ7ZhD5nONJn
8s/9GgLO3Qwq1kWMfI7Hb9fGgrLvYtWFVLxYYF/6zgX7FxwVWYhee9HyOkRF/PLdPRgpzkqSqrWi
k6P24O8TV439XCN13QXJ2CYYa0zP2g96tlCF3hhTc+O4r+NfLijm7X+Og4obrTWbDyJMwXo/snb4
Fsv6+htS8jNW585t6kVAftQJsOhmnCqS1waPEieKSNgxdfD94H7epgVvEU68DVjbnIYEVjoM2VJn
i6MHkIvLskTeNYHloMf6dZJN1t73mHQxYBRGjA4RoPr84qGukgWg2WVDNGawOjwzATlotRdpb/lY
u/InedNLvN4lodgJEMsVcLF53JrJje0AudKrybmgQY0XVaOEqhsdVVmQDJFgbJf3hRvbn2dRcdz9
e9a2CgZSWcNPx/j+zRXezLLYNlRhrFfs1GH0jFPxnEttJKZctAIKT3ZZmZH4+18yOpN+j/8jgfVO
8ST0AOlWM8g8iBlcWJ2KC14dVXoUC0FkN3u9WFGnlvfz0udfxP0PspWmGkKx3yfoXG/J+22u7ZiS
veFlUv5C70L12ocg9uVSyjEbaIhSO2Dr3WbQO74fafANXdKe58vH4cnFe4XKHUhoge1N0htgJafW
ExiWyq70QuAObgOt4vG5R89tYFrDHY78EnPo8nt/0cYa/wCemi8zB4Ewz414SdR75r6qbfBQgIem
JaRwcfTOMNaTKUrMDuBwl4pKIyV67Efma5C6t0QyPX4zyz2m/BJMXJNmSPzTzNr2nIcS29Gr+/KK
1CMl8qjUSgh8kMvwsb/djSxjnCuN4udQovAb0WsqmbBErth+2CKNLyEpIYqNbcv+cG9W8w+la7kU
i+MH5Z8rqjHN2bHpLaTomDIFlXSx8RQdP2JHB6qHV5nhOhmoL8JnI7H089fsdM4zYDPzFaWgbkKs
0eyPe/3TE7VURUw3P+cuTJfyoMB07E1G6wqczRItWWwd8BgTGDL6lewkFOyGh+3PR3bs1jPGv+yO
p7+2Xd1RHE6SD5Ql2wMzGuI675FeeEaytQ6LbQO8vHj1lReY9Eju9G5rW1qyHNjnSsUo5sV/ViJz
D2SgJIltBNFGGKnpQXeLJ63ulnKkrkWgu4/J/8FlRB6MHGyDp31QWwch2tHBKvGDX2ynAuG2cJQq
m0kxZsCmxuadtiaFf6Fzv1qOUJQ9u5Mmt+JavK3Af+6PjjzovT7K4E6vBMZHWAa5+7mC55mUEWhF
mph1a1wy0PKJDSidutTf+U3+LUXg37Vggb/insAcBrWEB+MIuLVbiCkhFs4X/82MC9trdMc1T2C0
D1Yrz/I1mns85UE/rDm4mHiObexTeqywYEURo68HTz3ArTfl+nknF8G8z3v8pa0kFrkknTbAhOk6
2vCqAJgpaWZtb8zr+ZNcznXgkNpIxJB86thgi6hRxtW+OXstbJpB5MRtwEE9n472+LV2g2RnFcdU
eqfjabdzn4fKr/PH47rL/drlUZTiPmpzcfp2kQ0s2ae03lVFa3x8LRTZWta0jR/MlwvRJHZwKw0m
OSkvPF9ycfkXFBzQDgDD1XPeADjkJTYkynEQV4fvutGdY0+AdzUjBcdXlNkAMuBp8Waq6DH+DNq5
pi9Ezh1jWhM6H+gj7cSZnYAsAreLAsFtA1Wtr0y7g8gxCuS+O2xRTbPE24OEGlf3j58eTqXwtdT3
bjnV95VDCTCHSA4p8EJ49lApIQdw5AywZqIzkU2ecIqNDmxpUibpT4G7BdPEGN5bTFG0/qoFjFU5
6ELb3u3hqu+yo2zORlyTtFugXvrANdR4UJ55+KuKn7r72bwV0Ak5IHO9AbRhxWfngnfn8OZMMMi9
ykm4L+wB0tGVg8/wN9v/u2cfyH3v9b9VRIlyicxmOD9rdktFHy4Jvu+CcGbgT/ipsM0qkW2y26bL
LhzjbQgrJGFshts92n/wGu7y5Z3H/CrFAeWLTt4ANUSFobdFQDMRbR69dEFkiZPf3l5U5HJNpyxy
Qd8c+TKKOo68mtz5eOwXvkUbowt/OtyCWsfeTMo2BBRTrx1kSh0o9ZKYM+1ymlme6OSQXZzYmCIZ
iCLdNtUXzqcciI5leV5jW0G77vOfTEGw0zPDOB6ClceFmALfTAyHnknw8nmomTFVuF5Hz5aI9kXK
jwCazaPv8S6CCvyoXYmm8OTniixmAbiICWDp27HofCz410nBcu+6G+m/6HzEzVgqqwxX6PK/yAVV
t5uqXv8J9ZF1q2dtRQ6tWMKsLvju8zui9REcpR990wqh9qfTJxAWZZIBmyTGgHQ3LckTzKqtLJJF
7hBmFUqEFS8A0rpVlXc0mTLMo4aGb9oAy27Jbkh78AxYIl9YVbk8kIsd1hB5rG3hOu16ea9CKl+i
T7q+UIPbZoPVAx8uj2iuHC6ZKENsswOCnseIFBvsRevYdhl+Jn7QPawCZlq9Vz/R2uSB8Py2+q9n
nvSV3qQHOKYsgMi+6FP7VXWxwb1+p8eACx6oM3W+DIw36Yhmkr4cmWAhf+GMG3Tuw2NGiBy7LEdI
EnhwhqSx4MhjUxamIkNi3dqv5069k2sVIA1Bpyn0kyCGDuf5qwiNmfKGeBOEHA5GpT52uP3giNdu
4Vo36NxKGkwzQUK1Xu6aza2Y68EDacQw2JPsahBg/ZasHh1vQKScYTSNibJGtBOfWnuXvhlwKS/4
cSHzlNmXwJ0+qwfogLYXLR5N4RP2VjxzfzKImzvZNsRKh4iktq6N6SwZ8O0ZEhFJu5C+6KNAr0gn
ntup/2srY9JqHiew2OYzn9oNDZRhcRow90rGtl9bUbbWawzEtZNysxh6vLwoE/CMMg1KZ64zd6fa
ZOZh9oqLrxixuYrUSQzsklytLGHB+P70+uNczeZlQweydBvapchJH8kUd+IQmY8=
`protect end_protected
