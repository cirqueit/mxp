��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��н�q ;܍���t�|g��`O���^i����0m,]�H�k���d��~z`���ۧ@��y�$�[�t�~)8��;�ʠ�d�w�]�J欩e-\b�X�;�.O�2bAi@b`�i9P�?�ʎ<�;��B�_IjB�M3% �ySS"��t���(�ً���v�@b�1���m���Vʙgl�%�sy�77�~�N��Mu�W�>运�>z�l�/�V!��p���?Q�����1����=�7gGu�`��[�Ы"�r�2�r���M�
�c���D���A 0N��wS�wN�M��)bឳ/���-g��o��u\oQ\��95�4q���'��b_խ4��h�Y-��T]$�|��9�Wnpc�'DΈ5?"}�DՇƿ��h%��5a��G�iD�Q��>$��hzP�w)�i�{
]*����!���\8�=��B���w���b�D9�y?�~X)].Z��a��s��MD�fQK���lB<���c�0%-?D@���1<U���Y�H���R,pr�=)@�L��N������U�ml���D�M�[�i�ߞK���Me�;h�fys:H|퍐�O-����r~@KNH�-�]tq��{`�`?2s��=�bK.꠬�HY�ց9�^����Ѿ��+�O3br�� m�R&�Ղ���9�s����ф�?�9 A�K��4L�gƊ��^�@��/�}�Cp�:D�Dk>"�mݞ�43J��Ɉ�<h]�혏A��$�'�#l���*�b
�;� :�#U�B���@��������ͣ�P Q�R_��O��</���J���0%�S��&U)���a��mpE�2�d�j��;W�G強/��3�1�K:��V�/7��Eז�<���Y�.��B� �9���nn�=bY��B�*nWs���|HA�U	q	:�T�&��Z��W�R��I�7j`4'�\寴���!�r��˹��?4�X00ճD�v��245A^�]��{|շt��O!��=�3�82M�\}bw%R�!��"�/�?CSK�%4��̄��m%�]>����|�r��>"&���y��Dw��W��2^�8!��E����Xn���	!�_��Mm�ѳ٥}��}Q;|`�"��n��j�l���RS��Q/�#D'd����UU��DLſ�l�p��*&8E:��u-���K�\�>Y�����m�PD��R���� �\1�:���S]!�aK �2F�Dx�ӆ�JG
(Sn��X���1�؄� �H�Ռ>��|�l���j���B��GJd>���?���C�b}6�V�X>@?�B@32���4y7�g�i7+KCᵕ�̳;���4�]�X�z�����jVme���, ��Iq�߇����߮�r�駣^�!�,:P}�.�i�6���!�V���+û��b��%��U1�V��,����ZsCy)A�#{�Y��ה��;䯯�\�t|h��W�Tf�O����#;�����9g���y"x�H�pjg<$F��w�e�h��@������d�T,�gy��ۼ�H�Er���^�)��i�^D�u����S��^Ԟ$��@X�U�q�Ecơ���Q1y�W� �4L0��̕ߟ��nE�D7��+���r�庀�R�W�Ȋ���}�,P͂�;��g��XKu�݊֔��{��gA���C8=���HP��{�#½�B����	Ok�^�r7��Quؙ�q�U�m�W�?5b�y��t+JEl=�EM4e�B�r��6í�h])J���ϼ�6`|�Zi!��#ȕ#�r��A��A3B=��:��5Ђ\��"�b29pH�;x+;ӭ��߈��؝۸$���9Y<�:&%[{���HϽHS6��P�d��Isu�jjٺ����f�N��>g���R����1E��P�GuԤ�j��*r��[z Ə��2��ͱ����*�%��Y��km�T�Q��c�������q�|�(�AC� ۡ�V!�"A�;)�q(��Å%���]C8�0�e��cO>F��*БG�ł$ U~�`�􏴀T�H9�(.�
��ex��O�nG=�V�_ʉ�3���~�x=F���Wn��J�jw���JȲ�1�������*&�xy=�)������e��W��x���(l1�6Z�3_3�i����v�&\%�L`���1�)/*'�˚t@=�q�N6�����Iiy��cV7�(�LQ�,���-����3$3[�o
���Fk��Sx�ͱwPgb�`�f�j�|O��%sP�I�
B���w�{$��G���k�h��,���bG���!�ˋ����ѡH�u����1���a1�%8�S7��|ts��io�>�)�"��n:�,��WF��li};���Dw��ˉu����w���S�񄿦ȏQ��'/
���6�_��MY���Ȍn�'�V��w�BED|����l7��uܴ΁ۿ%�"�p��� U�� >W�0Dǲ�H?�ñ`R�HvT0w>&�'�.mb���1dkɦGӇ�<҃e�~:�e�@0��n4��;o��������OD5���-N�e]�s�}F^U�6��I��q�g�Yj�o�!#
�!���U3��6�4d�l2ʷ�Q�i���݆����Q	k�g��8��+1�|$����a�Lߤ�L
߅����?�j9-�:��C��-��3���G�����Dj�Ym��hD5��B*A@�������9�˨�0�k�q�\t�q�I��쪑*A����{���PD���xG�z��J]�7_,��ܸP�It���\��ʛY�dkbq0��9�JVHfy��>`!�����:�)�ј:4��pb5�F���fj�:t����m��ຫ�3GTڶeJ����d����w\ΰ'n"fТ0Z��mր5����l@���^��|p�m0����4��g�gM	�k3�C]�ZH{���#��I���[M.$��v3cs�a��y�&y#L!�,Ա��4���󝀀o]��v��,���:(�IԙK2@ψ����B
��q�nOH�0��Z�'��xsj�K�|}`#躕����V~9���C�~�JX��؏X�@dc.�_��]��Ѳ�֏F���F	�E���e���A!�Pos'n5�qW��碌6��WeP�~�_@g"�bR!��5�����M��'7�f���<��VS���1�N�t��f�=�,���"W��R!狥�A48��M���>pA'4���3(=�ﴶ�rY`j]4i��L�������\�z2�.x?<P�JE;u���9�}�n��G�� y�����V�����\�o������3��]?�x怹�)G��GG�����n ���� R�v��|����TM�\��F
 ��[��]#���]�M�rw���6�L�{x��dZ�a\-"�/Q.��b�������h�>,�[�p��8E�\��4t�I3Ut�𲦈��΁-��2�8��:�D�3�N�m��=�#O��7���h�{�M�p�nb0L�V�P��٦����<�	��� x�2���q�#�%�"��[&n��e�zu���8��4J�3��DP���"�C�XF'�f��i�e�q���F�k����w��N��A,�+v6H"7��
l�	�����۸ǃ�'>ْ,��e�����_�� Ԃ�!}3�jЂ���*�s�Щ��o��*~��4�z���>4HSS��y-��n�σ��6H�C��h��g9�scP�{G)����.��o쵠�1X���ּ����0:_|�%AJ�W/J]-8�uQ���>&ଡ଼6Ǟ��0N6���|{D:;���H�c�;�Y��׽��u�S���5d�٠H�����C��&����xM·�w]qu����wZ�(��M��0�9�kqA�$����_��d�`!C#3��M��`��fFԠp5�mґ��Aa�n7�^|�Ѷi��{
�.D��-��H��&:O�	%Vz;��XL�@o�4�p ��^��:��CRC|)�T�hr+m��sE�̃�k1�c��\	��O��@��l��IR3h�
$x���߷�3���bsK9 "��[�� �-_ʻV������dk�q�D�Z�*���<�C���S���0��]���؋�s[�q��͘7XQ^e�4�R�y��f�t��Z�b��� ( �d�&E��LkW��ˎ���.-N|\u-��9U���*8��T��L{�P̺�-��g����F��ZH�B
`l�S��w���ߌJ����P�R��{14��i�D'z�R�訛;K#7�vJ�QQ�d�_֝@���Ȩt�]�<燣�4����i/��}?�f`OvYݙ}�EO\�^�fVD��#�|_~u�`��M#$��3�Ҷ��Ki�0�OB;v�/��}]�-������E�7XI�\�ӥ���� �ze�2�\�|G�9(���9�T������Æ��#n�U	H=�_�
XO���#J�gH&7_?�YEwl��F"ԉ���nK��>��l��Y4����c���/r�7'��+52�K��A�8������V(*x�qL�ޯ��^�=*V�M~-(-q(�����ibn�91�8���ҟҎ+�S��v��X���Q��~*?��Ϻ��T�D�eP��o��w���IDQ�6��X �M��& +��Fjx�0�aX٫:�vu�}BZ��4���j�
Q��g���?m�9���	��:�$�@��r��Ĩ��2��."��>���?�CR��$��6���09S�.���	�_E):W��;g5�l�9^�K�P"{s�����c���,t[S6CT$��.�� ?��$;@D�����[O��������@��f�2E�T����0x�J�^ҧ<��k����G3s��Y9�*
��4��Ӣ3��D�3��B�`}"�$#�A��P"�塟��>�	�h�~�#����%�:^���iA��"UjN�zg9A��$�k����v���S0�}��E���~H���_�A��ޱ��H��ȫ ��~�Y��G��E�C�O���q	���B��N�� ��Qh����c��G?);B���9�$�a�m$d j�g�e�V�=���f[�h�MVOv�t�<үx�n�dU�]�gH�]ן���/;����I)�������dZ��2/����Zࣉ��)+�p���M"�^m0�g�g�,�T������5��<	��i ʃz�8���~�~��{����	�+��؀��#���br�����S8�xb&�|!��xg�g�8Nkd�C�m]��崨�_���>h�c1�Oy/=��)�	��s�F|�s�q4ީo	����3��M����~P���s�`S�h�H�Q<�t��%f'��h3�<��D����/�����c.�/`^v��� ��I%����V籩����ނA mD�?}�[����i0H�ܔN\�_�4!Wq����C�?t���<J���0��׵6�3��(���M$���"hq\ ���:��K���+�9[nZS�_�5u��6���"�k����������K�:�ޕ����Z�I=�6ۓ)��@J3fO/J6�-�_�!tΫAvy�_xR�VX�)
!k&CR_��̑l�����xkJ�R9�#ĵ�t����J��Z&�8��"����i)_i��S@�"6���?rv�UCdD���B�"2�W�@�H���b�S��{���w$�N���f��/����d�EaD��=-�����,����q��|�<�f�za�:Y���9^3�c�u4:���r\w��?z���`E0�;�a~�L���-+����h��~H�z{]GSߍ�L���V��+���p+7 �@Ɋ��CʍU�W�Յ��p�z�K�ݕ�2�f5)U�M��r���O���4��/GGB��BY�Mt_7��t�Հ������<�CLzm=8F���
Sw�]��$���o�xU7��|MF́��_�Wv�e�z��i�e�+����8�}+(�vu��v	�*Ә�>ija� sǱF��I1���C����w{�Lì��O��c] o�Ժ���h��X-\��Um��q��2 �)i�y_z�GrHn�_G�	2J�0H���Lg{��<�����BN��S�O��ְ�l�0����G����ʎS���2`dC��Nn�;Ie0�Z�b2�hWB؉U�ceC]�c��/zC�3�vt�����fg��U���2�GE��j�Y�x���.,�,��6�/�g>�b�TvǺ��D�;�ұ$�x���N;]�v�UQ8[�3=���