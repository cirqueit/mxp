`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
T8WOOFEuKW8NOlGE92KNhhzpdZjzbMEg564Eop+uEjvaOSxppfr/RtGp9Mjw1DYN8scsB4kZMINR
d+DelqJn8vlQnpNMxQ/QK+I9eE7maXbELCq2yeg8ksQPhGVhEY3msVWwA3rHX1pIr1cqx4gb+yVY
7M00OOHrJJ9KT/mXkhKYjWANGljxCPBWiAIGWdKV8TzDr91C0lAs4+ipsrQkN2LmopVF9oK58bBU
ZIdtcF/T/EY8B03NTybbXTb8tVqDhYpXr+/WfCVffszb3mGBmyEvRVe1LrZeXnNXzrapLwbxNo9K
m5i4du2IatGqxbrbedvMAEeyKfC/DDeNpL0h2P2tfOLpZ1Sqcr7rj2G+NaHiUfvXhnvcx0DePiSG
dmcS/JSLB411wYYs/2KBVtjPrhnXV6z4890+Udv0b1CGlGDQR71+y9GYkXray6h+aQmhEMg20Ghx
3yXzG2b/T1QsvWp98JAIPqWXFmf3/6DZ/rz4YUT5OV4KUnpBi/JNeEMFSKFwLmaKLzkXEj+ZRYoF
sopVj32KxCXSuusShgKZTKoLyezOgB3JJOA6HCOXNloU7ZP/WZX80uQQxJXDOTX2sr9+VTdVF5lZ
Wno+EC3MZf1/zfxeDP6wQO6hPlJ7nTLwtisO/v/f+0jIpEHRFRkZMxIHK5e8VKaKZlWZlvKGK9Eu
6cTYXbwsZR+CR4kgycTE5wRlz3CuJ1QaQ4MouZ/tD7J2gc7r+JHGxFjNxU811hSicIACf5yVu0vG
FAaUH39b4RenC6v3AnlpLS67QuT992o1B0q1zCkdydb4kETe3OgW86L63yfHLDKT8edC5X5q1/kQ
kbpYkG7IoykGr8aneSqrz0t21R562GXU7kKagTIY92TcR87w8iSHWiY9SnX823xOHWHS6TnYhmlH
PNqzRbVjagN0zDqvMmc8HgdQkKuc9szKPMx2fs0HoO2z98vfoZvzIe7Y9bSEkHkaGHFIubY+WNip
ygDW4Didklhn/GhVkKttvaTgJk8D740+An/PQUvozXwGp+qOPsC526jM7irhdFAywZJfckvTFdQS
+eQWor5ii65+s4ocj4LUr2IRyeZV8qbq/ib1QZOVbzbOgP1Vy0OvM1/y5qnvR6cwNpNLtvQrHZP5
rC1TL7M6BynsmHDYseTbIYdKRhTuOxSu+KQXe+XJIB2WHXko7DXApVU2XDvpftxlE3sIt9mSKSn7
ERf8f8jyJ7b6UTpCq7RqcmApWxwyUYyRlbdnW/hWdeZjBwK0hIxfVJzfMcuzfjkSoIG0ay7FlcHa
SfOHEc3qOsrbWEhLeJQ/7BhIWB9BKbyCMXJj1HPKtPC42FcE9KhJmmAc/meb/8dOlP103pEEHB8X
8uhsBDyBEnp5Lh2Ax4N+8FNOIICkZhO/+csDtiB30uITufvqMhawGMPebDFmCEu0/zACE4blQBk3
qEaJq0w8B1o193JWTNcFdz3WpCZngoec1e2/GI1OkWSEf2ulGKC5wegI4zme5YsMejaND9eLG/PP
Jo5bVV6H37XKsSw+9otpB/I14cZ5LNEpXllOuvoF29yiK1Mb/L42Aduhi1jkmG4H6vEV/5Btgi/T
kzm6p24dJrcIiaPOuzdqlljqDxgMB++ZutXKehrjwuBZsZyg2ZM40wMioOR6itZfl2bPDTHIHbkn
aqQldTZhwhuaxEEyOxTG1PkxemFmiQJA8EtuSaVPn4xd45ZbxXnvkuYZa9MP9FaK1/h4I3ULXJFa
vxpOJYr+pRyLm29yFc/7mTNJIghdfUPyXXu+U4CUJ506XNR2LdD/1Czl+hZSPz/cGpW+RRU2QXo7
3wFPtKJ8fApBqtouiJ7ImvkjKaOTojoYMiNrLF2zpmhkwFcUHUiik84p5BbIWO5dLP7egyNAfx1B
QkexSCyK5PaW554YIWv5EL2ZPmE7IOa3lKVxrr/V9ZxzFTywYxZPnTKPrtFnbP6J77brRdllWaNm
IEz4Xgbfsad2+aAZ34RKQKI51hG7GWlv/o5Jc9sdjlDKnPEsqcLqhBR0BMR48/ZX6UjJmD8XuuZ0
UBgNNb6Jq0ZBXDyRlVqoY9e4SJ56j2s9DXTTIjlpR2P2i83gvdZfrJoSSLMeDgXJ1fYZOEqOzjdC
+k1kbPmCzWIPo2Z4PNVeP4tvNJhAxLlKyZjn23AzUPypaZ4ZD7ydQ4l1dndVROcK/w8wuklmmYvl
1Kne176aj7pmdc9dtrspC44CneA1DMHBW5uMXQ8NVpBjED2fwE/NlK4FPjTi+j7dS1Z9ILM0LaEa
tZUseVwqi7CvX8UQqeT6Of6YhdheFZejxzsiJ9J21ypmaI6LN2cVzLJ2DCBl5K5EStIheQ1pHnOQ
vbpTm4Ig2AjC5cq6pJO6A2GNweCfiQ0i8Sk9W9vLC9jF/p1pSza/CDiD2vDO+B/xX9TSrIIsBvAi
hhGGBXukvWTSZrFWUKVyAgWZU6ndV14DllO0z6upqw98MT13KK60salOCpAOuCWgTYH0Jlc1abHC
NLGBK+bu0N/HlA5kJuMqUwo5iNbIgG1qOB50kEelWl7B9sznZuTrKXWhM26YjRxQBvoZGc2bq8rP
MfNWr2Myyfvfcn7at9geg0zP9f2xSxrZeWRwIIfB/d9d0PcfEEpPw6ZDSdUo1zBU7qRTP6NVSN7K
TodmRXUJ+Q1y2gJHk2EshpKt512wfyWmNDVhJ0fditLH1eIfWVni2+mYFDj9TROpdJKsV9A/Wlev
NWFNta/JtMXOoRL6SYTOl8B+W/nxh2EIMwllJ69VKnm7CrMpacRELVLmdqROfd6z3+mtbj+6ouNx
VtIo7Ynus2zB8UhDpUOes7rRk7VOCTW7dONBcWI7mKAG+0uDZ2XlneVcMqQXKez+/YxS2yvg7OJL
Y7BQFGEzYZXbsL9GDOsOF9nEHNBvHBRGY7iXWgvHFtOXemWwaUytd1+hwmHAb8XbOMxpuNMP+nnt
aMnNbQSyezcVkzCV4qm6bJXUFbRXPVEUtrZJhHYWOWILGYQ8MhXSJ4U97pO7299QD/s8oZZprFPM
jqP+ZqRoDuDqKFpn4qF2+Ps6c+QbGbEZ2AW/8BcBEoZ51V1C26MaMpp8YBNqGsPFZ7fvOrAPZlsp
YEAUaw543IFzO9kqafX3dNPT2qRPovrCu4sp4cDfr9/l9yv7fNx7kk03ARYJq3zYB8PBEaHgh9YW
oBD+o9rKyxZW4+HQhs46V6u9fJsNsVjiXx6fEL58VfDn4eVv4PcLXsrf0ldiQtnoSjgj69ybim49
p0PUPvLwrHvb7MPcQrkd8di3VzDYB/l4hCE3jFDnIivp2BvdCwQ/xtLQe/g3k0TSooPm8IyDeZgT
efcLf/xIVX/VDWizVVNQKrVI7jS1LOmNuGR9Tz8qXnq3+QIs61M0tB0/+TRtzyBFN+CujCtApLtf
ZcF30WbQDGMQxr5ksWFW76lcGszNyYzxkPoJ+zG/AYvxBS/9PuFTSCI6jKiNjkwz7k+QbnPkp2R0
IkV0KShnYBqBk9UeKGSlnuQFtto8zXlBOJV9CnzMiqSXGv4LoFbdaomHpIqAFmVq3TCMzRsYF1Gt
vj8EkcqM4OYcyDB0R9vxqZZaACtQI7Xtnvd+XlZdlhtl6YOUV/Sy1Zlwt+TIVALeAU+JbQo2NOUQ
x0Z/Q2E3TDGocWWr83ZDIS/tsqAJM+FiadudTAxpGfFVjSwcb+MagDcXnA6CQatJSZ3TGAl5n7SH
1aWMMZhqN/eIKaylfNwabVFATMRjPdf/hEAV4gk0J5QztFIRuDvxaMsP54HiPUYWenroDQ+L60/t
Fzm22KPHMvQ8wn7ryeJiJQYjajJ2ZLpZHg/+kWTEJaB4Eaxr+UXRvE2ZRqhtUgUDuS48In7x/URt
H8VPGRGJH47/S9PK00oGB+9o/RisdvoHp2ifw5PBoy5F87p4Y+W5vObBFvta9Le8zKQOsn3IaR13
6+VYjklcuiXBGkaT07M4+aQ1n1cJstwGxXLpLyeQK7OqPmK5NEUC1x3sckXBKYrYw35G72dzvXx/
NN6kUo/nhGmrKUOLNfbup0fK24uW3rauL8Es4M7V/7Y1BneWSLruPRPqx1d11ksrkDT2k+XibAGZ
g/Qi9GEWJE7pDhsMftvXPmTEc5vE8SsJOpZXtuAQrLwF3MyASYaV95olbaQvEiOHegwnGxDDe2Fg
3tepF78WHV2L1bZX6BmBSGXuvPyu0gxjxfuLAIvh+mFOz/nlEW8wWM2cd7LvzQ9VWTbQCPiteeFc
oCs6d6sIc0fs9YjRa+vssFOzJALbR9LX0s7aFSrf8KrRTsD4X3Ax17dJCsTIZbJFU5Yp3iiT+sBi
tAVMtsbhQE6OIMjIbBcSLRnj2HkOT2KRJX8IeRGZp4tZW0JkD2BHK4PiGnFI7irH5WCncLZxSV0K
1O6ucimhWI/LZXahckWpCVJJyx3eCdqla6IVjz0aBH2yS0kCOcEjkYNsd+ZHBeZlk21TpHrdXpdz
64soSlaAqs3V1LrPLRNPIbhh8qvesi9fcsuCRM5YXaK5QR9/9zBlJphOduLrNYVe49ci5KM6huAs
FcIKSzRDiSbfFBvgbdHsEHyYrcbMCsiVRQRFmVZcjoaW+oZZd4rNjGubaa9hv+YM88Y1VkN2YOOp
1+MaGpdgGDeCSIG0zTyVsiodWjRDz9CgXD6FF6Q1udN/7pUj0757iX+U+BCzRqYM1nSv37zWaJOH
Bh8ep++yHbbyuumVBpH8ERo9gH1zb5b6f4pVlc06YiMJDldgUDwFt1RDAsYw/EpO+VRo+s/JobGd
bMJtsz4DxgHczN7jfw+6yfiSdhCAHc2GMH3gq9S4dk1tNjGoM7k/+EvhquyPbG0Z76jGgWsTh2Nr
daotwBGyDeIjI4DRPdqRFoWGMmNnhH29V9BsXF69mXRQ46qib4h0GnbUuAotqAoMvbsG2LmLoWH5
SskyuY7XZgtdCk592RoqNtK0EJ7bUG2+hxYytRZtv5NJG04dIeyIfFmKg+Fj4nLIlatjpMzNfcrX
CEeRtxMfBt7yX8ggBPLZbQ6dGil3J2dwUKgj8LS0L5A3msUQcwWge+y9/xmWBTt9I4nCLq6Bb9wC
VtEsrC+XOKv7DQyiEsbXzxVJWOlvsW2q0HCDiyDG0hXBswbUTVXrz30mUCniux8T0eWMEoKaJlrx
BamjPyChSKOpSnCYbP4Lc1IZHB9EiuTPivLkMQr0lrWoar8Km+Ekvfl49SLD5jFTkm6FcYdcaxbf
M1MhRZL3dzuG5cIZe3fOybB+44NGy77LIgr0lzgeO55oCs+qffIsaKywm+N83a+8MDuXsQyfBBMv
6GeX2HR8nidbfVoMSIt3NbF2695Qu7a+gru3V/19hwYB1BqBveHvxHrkCmJhIZIu3uT7NnaP0piT
Uyuq8/RFZDynGbJkhLjHiDxlJxMBgiztF0tRfsYomOMI2XLEIJ6M21cdyVhI5GCk7xbcSzosUdpC
EjKFT7UPTm8Ge6/oBpn8SDmqKOSPCyJ+b2Vpbz+Wj5n2bdupYx6c+KkiOGsK1QM1H4tB7OOCUcBn
9i+5DzUQHZyo4AssP6C+yAqxmLbLMO1h8l31ET3jnkDXgjNGQwjfI9BQvxusjjQPGy2jSj8M3co7
ZFL68k6b0T++6AFVsBMjLvAMsMvZIKDN/SDpAQ/sfcC5RAD6DdmmNUGajP0/GnXGhJWuAT3F9A34
Fap5fl9Lwv/RPxMc1gwadXy4r9TNIIGFQ+kJZTtQAbsF2Vsms7LZn3Zo5lDtDLxs0EoDTASCGE8M
sKCpM0ugSsMecrnAZjNDuQz0mK6bcXHtWTHLn1gDI2PZMmZwqGhrUtluMuokDRzNv4llSocUVMrZ
uP4HGaEvy2YgXKJBxf3cZTRmBOLsC4USt1Vb8RRbAUTE3w60zPKh22B1yRMT3/SjO0BfG2KgeQac
3A6cFHhu1I/Lvga4ttB3FUwPBHFJZcPN5YAbmFMGC/KAAko9UDk341XJKaBKw4mqa76xVIyESIxw
P4HZlB9Quo3DWjwq53lh6UphN431UosZV6/8igbRWiclAerki2yQqYIjJcbdgjhlYIQZbnCDWCEo
Oauln4gwx8LhVpy96nkngNJwn9oRuhKfF+WZmlL2z7yCuJVuZTRDnGj4/OuvRF5vYJUd4cfzP6nv
FsGzfMCbcKPZsf28BczzDs1Db7ebbGt2CzoHf0mg8ZD1bTzvOcnA9O8bi37F3KNxvpv3ihGRexrW
2OvA6PHQUPJAKQNV1TQRY7AUp4bSYZ7mMF6EKmlZ3rSD5sG9xnG3OgsQJuuni/F3hVj2UBJsF4Yk
6z3LQzXL61wwmLDT8Jz7LlIDcJQSsEbfnXCZuRmD+qHKi3E5vv31h89BwB+16F8W/bEs31toZ20x
wummwN1cZt0Za/Br5YPttFWGxiamDsUICMPEX3v8mw5FEPl7UHO+V3N6kby885MaiBaEX+93zrPg
g27Hvh5hN2u9Pefm7jH80sDgdqTydQEL5JCxAQ51vbprtEKHQPSObClq8ark8LgSPv7EyvLJbTDn
GLIl8rrkqeq5ZVmGeo4pGpZbrcZBY9HazT6ar/70Lzzb8xrXCBqZa9+oNHCprcL4VO31G7Dd//mp
dd2RtSx8SxIwLY7DioZgMSMRs6WpoINK10c5QCvYp81Dd6QhsYkbvzivFkwnmM5qnKx7dkpQfXrN
UuD4VMwfS6jM4Wmp2ifiz8Szv8SE2Pkl4dbsP7I7zcqbyIbSXVxdE/BdvQruKzHfsQJnEpxTqugy
SyfyFCySG4KfseII+czyhyvLsCadBAdJoRsuiq7IO7Z4fwxVUJ1WcdZFfKIusbfJ6RjQqyQgb+lf
2akSiKNz8JCGfvt4zALS4m8PQoneYKGNyiSg82BSesatD4gYnmvwKFrr1zPSZ8uzvtMze9zfUHTZ
t/57gvWFtNXty785AKkmakaklw79uZXjMzI+LfwtBzLm+Wsy7LTnGWfWp8uzfpzxlPNUVOIAsd94
0rvR1Sc9MqXNQ6BPRSkK+9/6nclOwZ9Mxb+2Hnob29IZnoQ/F5ixEORtCEA7jVPEhbz0rxPphmwZ
cckAGobbLsUHYTbHKIV2l18EBiAHDdhSEs2izXbwBJXtLvd8A6wDbKota41EhOszNbpVV/xLCYQq
yhvEE/fJh1lc7J4FRaRBA3USmsTyHyRuZWQD9iWtAzQFJbhEnV4mVPvurA8McFMQRk/4fP2Uyvye
sxrpfWk2HfBHBhi/hao3XmFEpiARoJDKWb1+hFOp9xBKUBf35vkAKyzqS9gHut3lvMDICdwULkc9
fGeR7nX5zl+rSwzBZTat1M5b4DLj0/oA5JGCJy73Gs2OjTrEG62bgaaHl5rX7zm97E5I+Ikf88QO
UOqhBVzVxeuukuu/nLtilxnb7/f2kApUxwQ0jOcgjZOPmaTeiNooCehklqMayD8B1RA8/FGHCXTp
fBdIuNvtaMvXk28EbLpAeCXOjKzOKdOwo5fMJf/6DaA7INsAxov5dKoqQB74i/7gE626HpYZURLq
DdbfCzfEs/ZNjlaemZ6GhgA8LFIFG0Cw8W5J3b9qt6SOCTXs3E1F0UYW7vVcV3U69gtcIlWTunze
NKdBL5t6LPq2fF2Nn6MIqMnDREKyWh9/Cp2L2UaZDGNDUT7NIsEBzzPE48c2wIFNdZ9gilmB3z4n
IMIxe+FshNe9w0Fkm08usaTnhUqJR+ylWs2Hm0RLHmyROqGnZClb7YMy64l6VjAf0eA6Gm/pSMxq
0cwZ9LIPkKmfy4bBpm1OANTWtKq6T8EHyjhAeGDIxd59TTnx9hataAMhDqrclSMBvbhg6fIoU3Wg
e14mqlJEblNrZmN365L2JrkCuQdjPpsHgJsKN08vR2U5T1jjnjQVMy6B7WRBZgrFXca7G4WJeMz6
XRPAWyWnncuZgI4+85cZ5Hh47BjBko5ThA5aB3Bj0FWxcoNAWjpvkEQY6RLRFQ2wglA9cPwmp61x
wNKgM+vOCTGZe47bExcI+35IIm3/OyZy0+MuJK9GOrBPf+UM1q1LGF6AAeNJ0ThcjBUQnsNuXGQx
L5j3Q1y3uetq0iWL2hGhAel35F2WyMnQol9fgXyHBJaJK5VFedEyzVhbJfhWx46EZXenvUQi51wD
2hOYsOxAjKlviYrl2GDxnE/bwO8Gwu8q3lmY2IzvaKx5wVVMErZ8MNFee0QOcm/46fQSPCzusjH6
oYJYTO+uhBX+m0C56d+ON8CRvNFY9RT/l9644ZoGSztIJnjhc3UjNDbi1f6ErTPbkYeMWtdTBWus
D3aP7O5+Dy/1PSTi52uuZuNqgSyq2I1+iNvkLIgR55JIrqpHh7hBwMLQ+EnjjlKR/bqYzPRkewmu
3wBXphX3XEfiBSnsA2zAL4G5QOaHjKaK/RHHvoyzJhQweA39biYo/r0FeGCUS2HtAUYuqqWlCcpS
Lq/0h5AWzYg4R2yD7QX6K9qdhQ7rJLcAcgAqUU8YRngpiGkqBNw6KD/XXhHJkf8qW0p9u5MVxV8a
khOpX+Tng4O0hgiMfCu29eyGqavMqhnvj/ryQvxdVFPjoBca4YPi+IMw9xH3gsWr/5EC5ms8URBi
AYHQi66VUsyjJqiZRTgp9VGhcmuQhI0PCeBTHZ9Ec2zJt/Ngw/YJesF6cPyTcUUsDrE4qNWBwRkw
jRLUEu7tsfNvwDopIdSH7GBAISBNBtbzsjMgJoM3Cxb1z/ZZWa9CGSr+Ib7muo1F35rBI4HHaiEk
L8fLATktbFBRwD5cLpDbw45/ITX4w7drtrZA9bpAyLWUG3p1/z9rMPYyUz5NFAghNBdmtESKNKsf
X/cYrdIiqqoGiwXlTunjLEhKVRGfoRBa4pFv88vywjJR3i8L+m3GTcVgRUVz2+4KMOyxUrIT9q3B
PPjK+S+jaRKUuyXg1I1FYQ5xZx27/qQvOaQ/x6AtQfchnZKmTHALTfp7el5a8d2jBpEkH5jRKFEA
B2+n+wSNpSwkSevIlbuHx15VSuxqI9xQqgBUlfmUjpU4B78I/gkWHAoAFOzRMgYOOAXcHr7gBGJk
V+2aRHtcvbyls9utsInYugL8rmqrZQECqTIjOeYc/6BeMREoQ2pFS3R1LITgjcADaoY71e69+U8u
Rib5c/p0Uxulye+Rey5X43o0SvXhtAA+oWlVuZCRzZ6+tZjNetjVhOUf6tMmLq3vK6xSxNEDmFqF
XVBuOPH8xvbyvVt7Hxy/YYx86mtxtfo9phK/UDhrd2nV/ckzAR6ZHKavcp7UtDl+++pI11H8yPfD
6EB6J77/w/wkoVG0g8wmcCvGZnOuZA9geo4V6Fizuz00v0U6iobjaCQsFcuC7f6GFI8sMKk8JDak
40a66GHS8F5SeWZF2g040cwSQlOKWBPrPh0xP1fpTHNWOrc4TxWsjgx/CnyCSszYz//SpyCcoliu
20Lh1x9Wt8ui9RXHd1Sj5vv7mVwjnHLskuO5A81AoJdqx+k07CylFiCECdG40+ARWKyQMrjWdCWb
HST0+2z+LRp/R/iAK4UjTsujlHu1aGWgVno5OrwKCdlmgdXtF1UdI55Uf4qXVUhpb/H4BTKiZezg
1GX/fq5Oq5bahuvnjuD3xD96yhcO12j3TZuCagc7u05zdG/UYu1XTgGkpSwQyXY6N9K7jNT0opJ/
rgEit9PG0TUF2vThWwSPtqoh0JK+DP/xubDJjydAyhfh5J7R9FARWktg+nBUtmLKmeoJYR4rFujp
HeAp2I3n4H/gPRwNRdbHrDrC2JHKK1oF+7ZMrNMJ4gorgbPGiInXWmEQx0h/PawNKrAHSn8KKPQd
Q37250/pGSRX0ktbC6UjASAr+RhX9TXI6t7lXwO6L51oE8NP8BR3cjjXflWx/ZhxmHWbSm9Wmhwr
PkqNbRLielUbh5F7MKDmvXzSpCrxDOXseEsb430+5eOqavjYCWfien2/96ZvhP+A9n4flWuk2i6l
AarDMJ60xxhxy8KzzfwHFgFN20/Dw6N3z2We8WjgMaMlPwLXuf0w1o4dg7wj+SsWPh6phFCXr9uv
AaKRq3P35bflSP9n1zKqv2KoFzMQjJCmjNqvVjVbaD4FULqM6AsMxKeIhfH5wjnNiS9KWQohX1sf
lu9gxvs5AVsDlBGQwpBFlEOAubKBsnM3I0/YsGDQcZDLvJ5Z0H2gHqJMEYJEr+hkLBC29plOS/IZ
7VWIHw6PFca7TcFbiLlTgVi0P2D3DO/1ulwPQb6PFr87CoD12kqWu7OQy205KkCZYwQr5ekPwvUa
OqHqvKcY0Tkgdg22F1OkqEYGM+3BQhsGyHsJCRifUYssXS876ppd9TxiDVpr/l+98DxQ1iNcBjiN
qqb1MeJ5sg3b7Tlc7ODZw8MPJ+swvascdLK31q0m5FmfGDXWddxaB9JsnWYukytCAMlu8OpdVuHR
dli4oRK0RBAeyx0RYnU64X7MsgsKA8x5TItU6dKQABZKwUWKvTHJmRsoS475WzbchvtnrzNU27oI
bzHM4AoezIxYLcx2B+UdYgpuipWXaT0WWnWlGNpZ2TwLnljDL6jbz0o+vn0wgRpHUShMy9GFak0J
fs1zPZMpY7QEFxz7XmiWpIjAhCO/BlteTUIDAFg7JJHvP1pVR/uBaJKy6PHULL/Kz0TVkDrZbnCq
pM7hEhR5AU53QUnznZ1xOc768lIAGiqe+PZ1C9cAshMo5PWxIw/zYRdG1t5PWfWZ+ntHE9g75OYu
/u/90oza3kerLjzMhxXdczaMCC4aBU5jHbqRwwQ+mAaOP1707L1ZkmHt/zeGwBhktBBZXLa0cXLm
o8Ai1NvKIjJsOvvDNXC+Y5gLeT1B607ygsj++26by+3lHmIVkQzHgYYdV5f+Lshx5TNLkjnmwZwR
7wYHOgPypI0mlgZlFKxN+M8pZd8FxT7bABcATDLRh6R6OKeLc3doqeuOIbSLon17CL5SoQivgCiz
OsgHyJs5mJO1elGoUjN7Nwv9ZeEdTC+2jp/WOaLnVNnl162IcyrMbFPVSuWptcGwWlRsuMTbsw2S
E0FLAF17U9ybf8v2mnvfCVclm6jIekB1qK+M8er/pD8rfAFVV+2ju5CWmqy1joiY8GHXIJy5vDTs
vdUXlWVJFRC1XdXacC8DKSq8xntTE8hzBRHwKaF+nMJ4mkbbRsD1uJivSnf+WA0M1S6e4rUa3Oh3
pEEmW2LsqJuxrubjttAT7M+eKewz
`protect end_protected
