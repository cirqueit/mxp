XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��n�9-������ܵ{�L<>�q����ʟp��D{5Gk�� 6���hȕ������ёlRF�G*�L�9v���S��t�A��?L� ����]���g���#-��]
F�x%��z�GY���o��H��E&�[�U>���,����Za�J��(S�"�A& ��vl�b�z�e�l��ƍ���ɝl�[�7��gGrf�5���qY4%�t|���W�"� �h�9��.\��t��GL��FD����c4$���i���?-�ߞ`E]�Id���/б�9�dW�ߋ�kc"���W)�&��or�MlI��>&5E���K~�,	��e�>�[���D��uHp�a~��C%:��˚��{X
Vr���W��z'�e��?e�_[6�+�GcC�3�̔�s�ؙ�h��»@)����QH~?��Y���~�~�T�7l�_M	@�����Ϣ�Ao��@���<0�D�{�;X6�澷Kqsà��Y-v#��Fwr"�����j�����>o{��!�9i��������ㄖ�:E�Y��I��{ �s��\�5��F对�j��V���Sd�����e� �
#U;�|z��.���p(�꧕�)
rp�Z���䚘7U���)��P�#�i��ä�W�1F��Jj���*��	�	
��΁'�F���A�7&�c����&B�9T[��ҿ%�).�6����WԳ>4l�Gw6.Nuf*�ӌ�~�ִ�
%�Z3�Dw~���{��횘����-��c�`����ҰAXlxVHYEB     400     210�q5��L�Jݟ{w�`��٫�J
<�J������FO����?��Z"$�]���^�X0���=�QnD���H?:�#���G�]>~����� c基^7���S�g�z�3��;���|�ښ'��yYf]؝e>+BC�v�@^���?Ij���觹>�Hd���u%��I+�P��c?ýT�:��?6�Nj��w�h� n�xV��#�x��G�~n�Ѭ."�bL����)u�P���7�Q��m/��2�������TA+�M=6�J/�A`�K���M�
�v��{�Rf^�i�3^�0�^_����<rV��]������NK���Tů>L�^l�_��GLB��e�3;7~�F\�&��8�}���yZ�;�f��r��<9��OO�Yq=�܅�p��׫p;���r\'&��?�+o��6h�3i���9i�|qbYD
��b{�l{.�;'<1�p0ꀝld�Z+Qͺ*2"L<O�Mp��R$�Ƨ����L��s��Z5Ȅ��_Z�9��FM]99�TA��ly f�(SXlxVHYEB     400     100k!�q�L�*|�: �B��eZ�����D`�k���G�l�1�d��ݨJ�d(��r3�����5JB`��
�������R�����)�1m�Q�\�Ƕm�z=z����̈́���&��\�[S���}��b�B�fH����O�X����r��N1b�l~n
e�N^�=���!���";���k�]3�8���nW�� �=#��淟>2����"I�^l��Z~��T�)�0m�ﷇz^��ͻ���OL;b�XlxVHYEB     400     1f0�i�6/��nQ�mK8�PY@R՚�=7����PH�q��A���rupR(t�^H
�U�3?��i� {O�`�x~�N-��{a2���3<��m��4�C~6����ʢ/����(g[�ڹ������:�s5�I�C��h�K�M��kM�$��&��ir
�3��"���#Ry@7����<c�߮5(<��ɬ����&Wq�dwO�ʚ\6�mll����D�s*	�e�s�>`	��KΞ��GxQ��2���e�eo"���O�����A��H���)-ϥ������@�/�VǙ���[~^D�I����xS��2�¿*`@ 0{%�t���Ư���1�{�WP������Ube�Jy��fRV?�(Ѳ���u��_S�7��������H(6FJ�!��k3�u[W#��C>f���{分��K�v���5m���������;�>ں9�T�0�*�����T��XlxVHYEB     400     230A�戠e
n��z9�;�EE�Bg>T�!iկ
���}>�TШ�h����Z̐�'[�U��R��
:�ٷU�͉��B�oyOF�r�n���!~�Y|[����Y�����2u@���k����9�Ӝ@l��\�h��熤\�ه��x�"�`;��m)�������o�, ��w���;�3��y�����O�IO���7S�r�g`)`�.@�� �QT� �N*+�O��dZ/�rC�j`�k�&��3��t9 «�����q���^��K��N���G�NlZhvh�A����e�S��d�y�勺i��B>'l�����p@���� !�
���� �-��IO
�N�@�Q	r��$+FFp�]�QaSJ�麰��H�uB��w|�������ؖ�*�E��U,��\"��J  YH��9��_Ո<ow<vUXlǤé_Z�y�a6W��M�U��u��PJ�Ʀ�z�����I�(��|]��Z��~`6?~QX�Qb{w��+�5d]�0���s�FH���1Qw�d��#��XlxVHYEB     400     1a0U�0�i#�ٽҡ��%��Tq�ڢ��m�`���/�`��Q��{j#�dXv���F"�^Lx�b���^R�\Yb�6�1T$��%��=�W"�Ž݌��|��Ag�kH5��A�^4����	��s��:Q�����n"�g��t'��!��bf�-���i��Fa�ѥ�^g�`�wದ	��ʛ���S��9���#�b�)ׅ,�d��ˌ�q�����"H2l��c#�
1F2�]f8�۾���=)q {܊su��.n���W�lE�u���Ie�1�]��E`s�mzի�.���$�v�����&���$(�21�f	qT�Σ���  � ���f�c�^z����PeY���D_?��r.&�܉�Ȱ\hϝd�ⓝ�����CF�J�t����XlxVHYEB     400     1a0�l�y���g�M�#H1]mf�xgɳ�ϸ���^�,7�-�1#�t�����`It(C$�F�%�o'�n0!��
'��_�wIS��|���&ԲǌUDP���E�h�kT��]�h��X�Hبcٙ
Vv��ɬ����vy���@�=v�4V²��1K��#Ų%��VS�˯�C�2,ʮ�ds���@P87��M���1,	�#��R0�o��d�է�Y����K^<��ya��w�����ߚ>=�)���k=i���dLp�������BL�~K@�(�*��t'L~L�G�؆��Ⴜ��b1#�L8N��ֹ(�	n~}�K?�dX�ءjE����(w-�;P7��uyu��YF�T��!��"IRh��::�,4���4R�=��]��,v��k���J��XlxVHYEB     400     1d0�_K��g��t�J��
�?'>B��kw�柖����]�+7���*��D��1\F;�}��Cc����\��"�Z#nT+���^���"R�!��2\���UZ� R&������0�C�ҵڰ�U�������FQ���Eo������������/�^���-&�}�{ޭ�M3d-Ó��滔���eH�D�cj&x�&m=��+{�&]e$�~��!Kv#C�agn��0ޫ�s���Ew�"C5�W~��d,�!}��j��m�˿�w8�ҋ�y)�p��if�
�cz�䈞�3�;��W�0QU��P�i,��RCո�/P��AChB��M���z�|ݫ���ig��* �	��9+�
_���ʇi�&�8?�/6|	h��0� ��)��m� �+nS�7h��i���r�mx\�'��AG���zֺt}G>�.�K�1��C��XlxVHYEB     400     170�u�o��)�nM�P�raw����c�6�e�	35�ſ�I�	g����!i�H��Pǆ���f���� �6jҞ��ǲz{�o� 
�T�

ɹ%R;��=�Na�w��Fltd�"��N�3�}F[�v�ǯ�JK��{�g�Ͱ��,[Yu����Hq�1�=*��2u_�`���/���^sy��X���>��V�\��	Jɇ}!]:!f���e���\��~D�c�Җ�^K� y�7���<�&���KJe�L��\0,J���_a����f
O�7�O(�#�3�=�#9�3$
BL=-�Sc08�n9>�{,���:�~=�%�C�n�Gw�m�T	��ڟ�:cf�ii+�4.��XlxVHYEB     400     1c0x�}���ŉ����3�]/1|�o^�%���$3ؼ��K1:%6y�}����3�3�4�Z��5	�Ŝ��5e�1o�M�#7>����c���z$�}�8��~6��Z)#�?��h���q�ۋ� ����p�h'ޚ:��R���CI�w���u/z��u�� odh�!�~X7�o��a�ښp��_��>���&�Ƚ�e�h)��0�k����F���i��	�)��Κ2�)l���(5�����(�!�O��Q+Ǔ>���﷽�Z��
��4�+��q��K͵����������I�9�o%��G�<�؛�%n�V���;]�?V}��Jh����l�7�!2Y��ٟ���HCe�8y��o�gT���Ѵ��
�ABk`Mv-ЦP�ZB&ܾ�9�B��X~�&5P��4�Pf�E�ӡ��)O����-�x`���h��XlxVHYEB     400     1a0uU�-�j�,�D�%�]Y3������d��>MX�a�����9�M!9_�d������Et\�[.����9�������>�G�h��=Aė�������ҋ%�N��:s�ܑ�l�_e�Z���	(���t�'�aV���	u���y�}�R���78/�<O���	��+j��C��市���Y�]��ge���}�W0�����*�6<���>"]��]�Կ4����iڴ�&�Ќ-��#@h,,!ޠ^��A_��W����Q�9%��b>�p��/b8���Ѵ{�GW�3ב� ���B����?lY��Z���B�D1���_��afW;̀�[Y;
(*B��%'���ۍ���� �_��3kYI��ԟ����x�����K��z�����e�H[~��vfXlxVHYEB     400     140"<�tkh�٨Y�Gd�!JO�����V����Kbzz����uqs�1 �����khZJ�'͘"o��&4�PY��xBґ��$��&�ʃ5}"����H��9MyM/�5�r���W���D�?Jٮ^[��!b���qY��x��@?�1�ȱ�2x���t��A�ڂ�$9�F�K]�e��>(�p�0�&�� ��}���&���4�pO���<������8�X�?=6�򁾡GGP��bA���fe����9��C�B��~�b��ț�d��[O���lo�����EK�_��n����Y^�t�=���PXlxVHYEB     38a     180�>�ɒZ�pn u�	[7d�h��}Hh�}�:"Qˆ�g'3N)^�c�C�}�[c�	�K�m;�:��?��?�n��t	,�����~����y���eK9�(�Eo�+>��$�'S���KF�ȝ�UhY�-�p� �n�.�Tĭ����RlْZ��3Mn�r��ib�l�=��&�"X��JV�ڲ���&�?�ة����JZ���(oqV� ��{Š��zn�D�z�l�pI�)��z�~w]���m���O|�K0�<�D��`��T6jp��ρ�νLL,|)l��_�1��N#�)��m{��Vۉr�����%ə3�g����B���ӣ�N]����>*Բi��BƯ'4~����J����i���J�9u,�@n