`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
VewG8w/qcB4bNUdO70zkTvNhk2CnMLMErUjPgRMmb/Jot7X9NSWH01sKtChqLWsFqppO8BVHzzv/
PvU7Dw54UmfD+hmPrpmkhJbKze4Ab0ol+w4oQktatp8O6VCdVEN6txcTVDcHahAsQ93nP+tFvnxg
gNxR1e53iVLyEDybJdpwSue2aqkP+gwNwFeVgH9vwC+GWrcXoiaU/G9PLSPT9qBKPm5BGsXJ+gxa
+KD5r2DMikXHoUxLkjdxRkHXszcP7X2LT922P3b/iWBAUnGsuZib7TBmcrGsGiKWv2VUNb5E7n00
E8xAC3hCQloGbTk5rE9QF7merfWe9C0HhjPu/OQH/j9lAubkNH0u4NejXocGp113YEB19lsDlPGo
hT+GiR5QyNndCxhp+d+KrqfgEk1TPls8QRbgLijB3L7mm3g7kDIDdoAA0ct3u9BFYF5lr5KZSeYh
JYZwNZnV89s6hYuNIhVPdfcn8hKk0Drd4J5CITRVdHoxLRSN6tk2e6ZJRZALVWrbfH1CYGyZhQlN
onOqCySXZKcTIRGGsatP9+W9GjejsXQp35H3s797CuB1VlaNshO55Cli1TabMfeF/Ph5WRPi7cFF
gdJFi7fYKn15wm7ekSP7rZwnyJxMszr3tLUazuwZ6WRAbOmu6AKnlFfa0Cuv3Y+evDPEAiLKgS3l
LBjo8yh1feDgS2FPj6ErhPCCbSZit2BRRlCwyr9uTcFXJ6b7qkEfBaNad4TkOfazJQjMj2h592uv
Rep7a/HRbLV9D2zGBRtkYIhDZjsOS5wnviIrhOfWibwSDe0P7Hr+dKXllnJ2aEzRk5FZWQHBG7g2
IZBUL/t+I3TJyRsKOpaeCdHUJS21k7XfC3LIBp3PqDMjddq5DSWXIbcgELgmndVZmrZ1Vtv5iOip
wj+4c9dGKpP5xT1l4nxzC9Kw6qTKo9Glwtabkedq05VkR+rXlPgqZZ9DIBgcMNLjAnMj1D/gsocT
M/BEj016qmTK1764NJsjS5T3wd6VBs1p9rwZH+AbLUl8U7877eCMjdENs2BQ5N5CW7P1ka8oB2KN
TE4azOPacIlEZcqEb0gdQ1SSEFuHcbpPrgu7HZFQAoAMP6TBUPsbSGyYEBXFVhor5UaY8hSdCS2E
i8y9S7mbVIShZoFwrKVaBH3Ql24pCZ6IRywB0benCsjvJcXNcj1rT3cnwN886RZr5C1afFQCdL8M
96Nhi1qFiZNEgB3GZS7raqNhCdsWxfUH8400dtaFitAwjrzqxi/gnOjURH1K/7YEr5UrVfsWvcEa
mVFmOzcR5Rwhb/fAWjay4UoV2JBlJsS6YW3sIOIL56LEzrURkhAZQyp2RJn03BsCRePPlYOBo5Ee
6FpCstAO5e7gTZnYZkpyCKTnwwjxhMUwGghf0NTos1hYPvF0AYVG4eU9ZEgTMcUBsTS5bjWeT756
d81w+rjAtOtbu2KZKYNHYEVTYo98FpKDxF8eqdXb2Q0FSEesYoyw54k2r5imdDpXyXpWQZmUufhI
IfSUG83RSCjk7jseaMBXG5oS8o4T08o4xDu6wNir+678KQcWWQTENhvTL1q+/g33oF3M+UQaikdZ
FFc8531oUeKKYb1UR0Woap547cvcFDTWs6fSgNGhV30MJ4cEGt34yooasaamLtsQbndGcrQnQtRe
9+pvjC0h5MC70AimfWzHnz5TX/dEr1YyVb8+MGZe/LQjy0BJUkyhDeQSt8nfB9q6T/B1IpytYbk/
U5Mu0avAgtzH4ylt4ZuU5nfnNATOhwjE8NAGAhNRltMKaeGQSYHpN45Xew8g04tV5uhK7n6dRW1r
oz3I2ShDz+oIkIU+3+al2yx79McGJiXnUYaKl4vLkbRoEIWhEEQHH1fKLIVpKg4JvxvTdRynZiba
aUTJlhLz3EbaE/DfUUUz4yfunth8Gk0LHDzGAgNNVPcV0/zOIKDRtOiQFsxR21TaICwUNOfbMm5x
zYRLfZVBSnryHEe6oDzDWnjCqntovqESAVBRdASFF+4IN7MBB7ZAJtJwoOulxLmW9B6ub09DG0TT
0WTvwqxdT96mJO2Mz9nh0SMURLV06phCTzUCNDQz/nO+UTfob4CSXAdx3nk4Cjz3nfIi3d2T56/c
ypShb8962fKr5j9SLV5ZJNW81uSUkIi0wmr51B9aO79WJuC/1rkigsUgRwAK4+rYoiQq2pcHdMaE
npiNI/kDRaKzn9gQUfu6qGBa4PAzYdwmAB9DMbrYYxPEuhpuGJy3bRNOsaTPu6Xs+jQc6N55U3vM
4PRkyhe9MFFo/8lpCsesiEp6IAz0ni7/gap4e9fqfHS5k5NFMH7GB2VU7zsArbmyNAtwpVtNSMMD
H6qo797A4xTvbCD+mXjcnfZQwMHVJKBEvznM4s3x07hlim/f1VzOqLU43pbKX24pAxk4wATZxqWX
s201XMPZ7L9jusp0gzSZ0W10SVVYkHY0sWxk4/5I/bjBQQq+dSPjaUXHk2jkwXsvg+1zrzeSqS5f
FQKjQQDTQktnWeT0T4QIcAPndChpRUZeIi67gIW9y190i17+kxu0fUpxJNq+D0DDf6/6x83IuMIX
o+r08BwcKFsoawZJFHEKJ9PaWNnzTUiKBhzvYxu9twAeoAgdxzt1yyYJXVXKDVVDx+0mTbKRG6BI
cj1ZRXDaFKjwDqa8W4x5owbvNCRkA5kd8SrzI0PuSQNN4znQ0S/+xTiDnFVSwGdsMItZMD3UA/VW
ILjdJsrJvczSwRAut60KHC5oRHEY7Ccy2ecNzX0PuZldhmntuMV0Pd1cd2TixrM12SOHWH3K7hra
tFYuevWuBj8rrTJYRoYw+WzV1Io8cAGjaAkR5cXkm2G8dcomqO8WAu2u9fqaKrUep8VWSWRD+Cvn
x3KsAFmfkIugSWsZDU2VuhmVGunzgQvztjST+LEVkk9mBY3KHPv1zXooy5u7C50i/nuiuh4edeEe
LJf97qUcjKN/NSGFq98EbKO9N3oiFbnLLKKQCJ8Kg37qLX9o4pLsXYplTSfcwan+oAFqprkNTDBW
5SaFjA7lQnqxh9C+HqWFSwcmBPWaku+V9ZjSeqcqAL/3USRHBYhSJ3WbO+A2/GsKaUOLFKrg+N52
yRerPhUa1m/LRy01byN1V9qMMbFhd9IVDaf0mqwIsy0jp9QPAcXDkSL0vFg+TrJeJ08Xw8NKxTzU
RcxMqGcmf/19Ld9xMjmcElsGaBANXrPItroQQ2HK2mWsrTNo2d2H3Mf8ZY1azsp+4j+owJDt0UOa
t8VvPyhjgbIJo9aS3NnU+3/PhH7PN3IQsS4YJGkFvFokOqUWdMlgi5gc1MMuuW9nOJXW6LJbMi0/
qpG8MI9M5+IapfoVPdXxHrxWF+P85ppQscUlPOYwJ3kvVEBUSwmd75kSUDBEfF74PmK4J+rH2Oiv
N6Ah8bLsCWHo/gEh43gpwb8zPeZJCNMT5toGa28LBfH5rzD2/CM0uMWj6CKDwaH4R2YVXFyk0f09
hw9GtgHxgvICWRo3D2c9s4HfFE1tW9k0zKVocvOZeHwRUb8mS5OzoQ6HKyJEUvT89iXxqzh3pH2+
cTVCgBgw1y+XLsCCNi/OypF8dV8ycwpIn9SnoJ5cJQ32i3SS6em6MAGqxp2VxoF1KN3LoMbDVHNw
WjxF94d3gfG/9suvB07CYddT8nWt03hDDUwVqv0hKy8SguOVivulEz945ZwETCHrRXoC1eyTpXx4
Ix2BfSdR2u3UVF/HtxZqWoG0A7TKN0zIYan6hzBET4KnKmbb0JWtwvY9oL2OFDWBVmeuxfpp6eQW
Ob+zugbxy5fg2IBxX6cVHHOMwM471rFD8iVVJl++9LjGmqsVx6YpbT1IX8leJ3vyHnoyHlNveJWI
mW9UEwtZCw7aT9NyFfzQw6isukNTlMqmx5QrfRJFbEWXwEP2hiPd7ckHLOf1HtYY5zPCV6NPTjpx
wtB9ELRqYJqjQxQFSQKktbhGtU5mjshcBbhtPv6brtjMwpq5b8x09VpBJWdZWRgCunxKp7dpzS9g
4tC9FdReIxxFduBndmB1Cac0aLT8XaGRwSwnlDDtAlbct/YqhdFIT2FD+jU3Lrt6ZPCsBi+HygqS
1CNkw7zIG8s71LRg+Da3nIZb6hC6Ypu8yD4MaS1V3v/W4fmFjV+8OgqNzZWjPafT/QXkkoU1rqSw
hYKgJPGWeDK81gB3WY6NG+C6WsuoPXBmDG2x0SVGUkzVrof9pBOsft1URmHvq67oT5yapM+Z9reI
xvmIO221svBT4XECQYVFjPChfeLnfr8+DOmvwxPYp5Al5ogr60Bby3VoP1ctnOnpnw5Kh5ZhRz9V
+Glab3KKW/3fmFSQ567sTSLuzS/t82IFQqOeV9fQZlw0yNJSuluU5BwD0F8ecHkC1AKTh5GOhkKu
kHu8sus0PjMIp6FbwHQ3IL0kq161gORKhgtYztsPhfQQYfNb1lfhJiozUKMBDrLDxmQTCFKo8x+y
uBeWdFgGBkd25ECzUevt0I5xjemEugPFw1ypL/JvIztp6fCI9dSiQBN3CMGaxO/XlpRiK5AR2998
xcdJbHd5SFI1emJVwu1MNCVrAVirvZd2kN22CdaaZqcH6wkzaboYUiOO+ucfxKgWHxnDxSLxJ8GL
4EzZ+2DUCyB2ZqitqEwXzAnvXJu2r9TBuI0NbtKvrPgzuyrikUxs0RfvhawdtAzpmzFbiWZBR6V0
Rq46tnoL0rw3FYsb6Rhp3zCCDE6Sdjyu4LyluQsSu/HahHhAvtAHzq5fXCVCZJsAKgCVhcoYgzKN
lCtJZWl9osbM5WMbSiaT6dBkY2YoVjG648EvpESzofmlPthJzy/H1sf7iBaL/hKP2knkw7V8SkWP
daqaaOzyqgHDGc9z2eZzfgnzFX0XtxoPrpSMnBH/7nqUcu5I4IJC89nJ9GRcIQ6cHvjir8QbeP+E
Xlb7FZ1/p+E4awjp5xWF2//2EDp5gQtUCNLC8NVbjkZx5hFOW3RAl1a4alpcrv0JqyZx3XFk5wjX
DQSt9DCkeA5aS8qiWY9m/aXRu8srnIXgm6I7eAAKLnQ65lSEro460zfh0pAstOQdmCSqfciziuvh
IlWoHHQgXOWSuw49WRbmVw4zpUCmvKIwdKO65skopKh7TgsDxK3jdC6hzirG4PBjooAHQ1XC6vzh
qGlqfeyecFr1fAHAfY2GljmNdpw8RG4p1ZSyBBAigL/mqPHp7IY7MCZQu67HWukquhr/VJKBpo9t
aDlZZH8YBS9kZREpZIWAdhT6WNLdsBIlczn4XlkXuI9VXQwzsrIiBZLFLm4EpyM5DVyhSp8hpg1f
C3vIjSDwm7hhTpvy1id9dk7CSg3NPyRe2zca1t7whetEJp27aBJEF9rS9IKLBujhOCHEz+3l8p4Y
M9n2gVC1UKtIbKTJP8W1wYOkQQ1MxsnzOCpO89X6ayczDEyC2mYutcWXrDL1HcXJXOPIyebJxd7P
nwbQA+RbWjfqfFkmo96sRXU1RWFrZdlMGhBIhbplhMTd3BsRprSPbTf67rQfJNFkWo8o7xtLrhYq
zS8CdVPtjrcqEtKitq7lcW2BPN3vTXgUloC33YUh1NeRQNF4fUSTuw2AUBaubWLOBg2d0h5aGq4q
6iF0/GuvNIsnXfixvhLDOp33PKDrhJdp/azhNaKnmOGoFe7vhkZ8vfoS3kKyVJzZkiqCOhv1EBIm
eNRFVH3SwG2aSqJHM+4yB/hWfREKjKOyoZ7BsOpd1gVbbadXFamPoVxSI8WPdn58Xg6V8pQgFnIs
w9MHE+dP07L1uZs7YvtzW3P3yHMfTD65erjD8s5h0jP9JKfbS+5nFmsT0svztSeLR3BMeiMaJCCJ
zaQNpm9C1cuiB1UgWILXe9UGWZe2wFscKfpE2lcg+M6S516ItEHx8GjAiqp1GeG6tx9cH80JEpA7
mb17kDXI2YH0in6nkZBocFg9hgdxPpRE6U69m68QG6AZEXkklB2ZQgRgKx3JpGHe6y70S/Ie/a4A
w6+mgpfCaN9gWgxCYpe2+4gkVk3c5zV6d+t9kecss24dcvOJETzQNAYsBcH6qp+pEw9M3SX+YoZ1
w/y8kqbYRy6wYk/u65BRm5BJA5STHTlCglDyoWtwdrXrXZpyFpo7wcmxrJQWyYEqH9I4NAVsH2vg
NfcFe4256qqev0dIZmPC2AymUK4xG0abn9ol/i0AtBjQbufBpwYjRpLgQccAgpvluUxHtQj/rRBK
1KVhNfz1QvjFywKCxYcuNJQf34m6MKihZ21D1Zp5Dq59qx2/8W8rqZs1Kt5SMSOxapTFAh44jX6g
J5KXnLF3MxP7pp4OnJKuj16HtXP3iVdOuIZyxIh79xu7QMi0Ua1kQ1NnDrk6x9x2dNr9VvJsgV+G
Xvp+jRZceKVnmhdrAmMjhQzipoCr+aPj2/znZDN5a+eGvRLrLHxWi+ks3wnGsDuP5kn9v4WTAj1A
QBli/BoYrCQQmEEGp40L8qo7KiIcooWE5+Ub60klYZtPorEWkQvl+KTPIQ8FdDloBFots/fGq0TV
2fqzg7fHGrUBlIv//r40um4vJWnXcTm6y6eNMe2G/KWil4NnsWNDFbFXdujc0kKOVPGb+0A6AZHD
+66Q+qTXjU3ivTu1g3P531dHElsBrjjxtzqcJT6aJ5Ol0f7xMe2jV47q9cKBZ1ssyCJ2C0Uundgs
JmHXpmhMAdtr8mv2FdmUijLBX/cM25YLnv7aQ+8bG48+YsDkoj2uiR8pi7ty1jcArv6VXI9Wsw1r
yghSsnQy7LsTdrDy15NcgK3BD1Ync45RIrrv9xxiE6QqZ47djHEN1HCNhFh86fAcSTBp5txV1Gdu
VrhMxJRwE8/3DEcITjYtfZjvmN6SdYRcUgHgEWJvEBCNmo3hQpViN/lrSihYm1PQlZiRFOGGsiEJ
6ABaSd7EuTUckbHCwBwYsIcDPj7PCjkW1q/5ennA6KAkup1hurCPL5WmBNCbXHrmIDc5BFkqi60m
l64P/2uWkVGq7HLsTvOqDVknr0WRLWvIWQphPeRCtl6zpiGGAVwQx0b4HQ7urL7sp30rkrLH0DMH
/4wfDv20ERnTqqhSUwUO5PaL0iYObFi06H1Kzk6cRCMhGenM+vcT5VAdKg5zpiH5cgTm9sZMiA58
Jaz1hz4zmxNulrVLTMvcsqJq2+GZ5IJhiKv+cH+4pASeVR76S1PskdExuAJAZdtdEkVU2QHXoHC1
2I5Vd5Jc5cd6SIy3Wtb+1LPMl3gwhzBJIp7sUzhM1j39r8bBo5RuuZ+ocgl+pHAuXIKJWUmi69BB
YEKLUquZaJTe6ZOV1D3cfjlRVGjE6s0StosYd2G27xcVH+2mXonICXW+kpkjXqYESQKarFLTzIF4
4DOSCDVOu9bbT31/NCGmJ47oZgV/7GdEc+pOETl1O+Kaq3kFOid/v9T1Ea8yosPUGhpCcgpn0xVq
/sbrEEuKr3ablErl2/KgY19tZsuvW6NuVdZs0+7ZRUKCBnI8wFabeaFEeFb//qg+BAzBKg1B00tS
PyvIlf2aZCQm87nvd3Q1DrnBJ/PDI2Cv8dYhl48VuNj6y/2hxup1PbZ09mDOadlJyudL+5kG9sRw
DQqtnPMsG+DEF0tZMrWhK9RmoUwHuWjvvr0PAO5nScfvg8iW+08MKXes9LTcpSt8/DNqVh7xFuBJ
gm2+//6zN8PDPxb1uV90mpL2vEowus4VEkJb0AHLsB+i/N0dCjMbn9AQYZn/bGc9gTwaFeE/Z8XH
8v7tVS90sjZ6Fpzkl7LWdFgKdEllESVtlUFEq1hXQlVJj3Otuud9QsavBRo2RKb6FKyoVMq/ZFE0
w56aAwLW/dOYYjPUIsWK/85UoyzMSp+kLdx37EInNg4CQRD90p3DBZwFM/swhKXLfLUFLOUXCohU
rD7YuQCR/7xiACJZvn4ivfcMrZPLjdDERDemv6YAOw3tv3A2I0dHQOLrh7ZCKPSlZNf49Cyik3mq
cm+EED6wJO3Bgup+v/htLMvTBHd34X3liKUIzHkUlnUGvNgNHeNzeWg4Uhlrmqz4ljfmsNK8WyUZ
GggaMRUgGO306apgZSeqZBrVPh+Lqafs8yDtm8fgmTuXHlva2CxZB/mbDIL6ZiFjI2l2J0AXffJi
kC3LsgNTsp/tpS1BU0CR3vbxJyvda3A6FafHqX/G+buXTTjkrpAAGSDlurmgRlKubCOq27H0v5IW
G/R4zCUwowRsa47k2DGkCqazn4i2rZ1mEetlGyHciY1jkYeGWHXSbzNkzwsmdClwq5BTnmqDuMGD
1o/DqMPfg4LbBui5Rsrm7Sp1W6Ky6ku9zpekbeVcNxN1IBUwgPy9DMFCm/mkihoO8UnFu6zYi3jJ
pCPrwZkPTkNMceZPspN/Qfobz5lLptZDzlxupO/sei09LOvDKNoiTSBdqMMBHr5fW3xQrcKSWlL9
+Iaeyb64x9Ak1SROF7UkPWfPOKsBw2HTAjn3oqmSxWiVE5kvFZr12IB8D2hglFAJp2Udz8zcR/HF
ZgicJ0DPVlpWfWt4bT6R703XpY3baqYWxXVJTCCGLpxoiBbZoYULXsY0q8yD+xFNIiKe4D1Ovnxi
TRy0/rwPEEchDpyWd0MSwEBu1L++xERlbv0aDApHK281XrPOOpW2Ft2BWluX+FHxW4DmABE+vMJZ
PTA0DHZ9FtWuVci4x2GgUAcr5qbfEt0HLa0efiQQuYwG8y3qKPKGzTyo9kQDPaOPMbLMXlj9qOKt
12p5ytmtZF/jTEKA3KMs/pdJgD3UYc/MipKdl4HDoLbA/40y5n5zSG/3+OoTWEy+YyufJntoErQm
MTNLcAIug+bDHP3+iICLHm3HCrtBQQbla6CnmuBXa6raSFwXRFydRfS62mI3cc6yYYZ/1hEbgG5Q
BshcZvQDPa8PpyNwWhleQqTZ3xwxKpcweYTOWIJdxm5VbYlFaiNeI9ZfoX2CwHuTL5IgBxRs/Z9P
Anh7tWy6J9+PZ4QXG9/d0/WyCtq7ARZP6PgsDRASAAUDHrTDT8qdC+WjdHleKMYHZlBgk9rArch0
6Lxjo0PBf0iXZqa+8JQOPIwW4fX4RZ4d/wSk50IVuTKpC8IQWiKncJ2nJYv2JYxX6Q50/sl4IdCc
f9jbtotQHIVQpm5Es7sb8UsIZCM5e+oOHLOFzYeOiHgL0EAb/T1UYU4Sbz0BmLWoiLfrYszdaMn+
DutyjDFAYJFEVDr9RhLExqmsog9ipq0cqAsChigd+ScRmXbRSYxklVQgELhX+mk4zdyknAnc7jLX
u8HWutIon9g9ahmA21qWUE04p2z2rROlUQe42o9g9h4WcEh9p6rDmy4It9Mn9lbDbNbWBODMf7Zg
YnfhLEsrZatEo9IwjS2uAv0M3pb+r4mSmWTLmcL1NMsy66IEJBnbFHEGlhPBfgl1PUKR5LIeAxlU
m9g4C0F8JCwQgTXQX+kzgAFE6/t25zrIA4WaPSeVBUh+Gavt0DAQ898XGzU7aTk9gJdNhl5FQW5w
eCKD71bOw9pUr9DdjhCrqzID0sAySu2OfZZOLaMMfE4QhV/Xt4qoHyI4x9cegUcg7iQLLmkrOJLd
Rw9dhvi/pnAHc8tWJmk4o+h0V3z4m+Kmtkp+UZPKURJO3Qa7fZysBcxyv2xifWfHEKV35eAvg35b
PVtpNgRsuRQLnxlQ9CzG3vEPaVFMGg5FisphmksAi/+PEA8lV7oWIyi5UnSNP3JBKF9PI6BP7EZv
5Z4LQ8fsiHA1Xpxo+3MRoN3w2x4uNOhFlIry8KDpPay9xMnQbhINxGQlI6md6Stzam3zAjQPahO0
+962oSklahLbAiaTjkkblAE4Bjdb1/aw/6KXUb8Fi5zmXmljMCQntZ7sKgPWkzcEGWrXSo4hVHVf
SqceTF9cFLjq8SSFGG5fFlliACE/BLffUMaNA/U+cUTMV0YlS+W6cLCap9TBCoKZ4RHknfiGyWsn
vw6onEQLynPlyPHBjDRRC80Tt795qiDOnYBlkP0K+NyksPAtvPONFFbSJ9VFNFG5eibHJ4eKRaTC
cduf+oT8Z3IALChab2QCfbAT3n3pMfXEx5quFBvFFCSKaDdxu+dAdMYCAXsfa+h3LecONpHo+Rvq
8TW597QLHq2xCyL4XpILgznH8xG0qf3YpVvp56YEmSUpz2A2Xf15wYPRg3hNMj3Jx/owGdApZiG8
gqXvmSyLyW69xt82cwCw8ExBD8isFfp/KFj00zo1zdFdslJhIbCmhdpeBJZOpzOFfQ4fu+yUZm9D
EDYYmoj3As5lXYaFbhmoZcnJf/+OOCHpLgHXAuZByp9aBIPNENlntVtc00uq5j5RCzG7wYl1WaUu
FRygwl33CULobzLiqN9gZ0wfN7uyupO3bPmeOZmSlfJrB/TtGzByJaTV98DwCm9LviDNf8aQoLbZ
m7pO7tocBA/cmg15XMP7/Y6gB2pBvnliwPYbe7gi7On9H1L1ipCykNpDJmaW0BnR5KlCYMG5VABr
q/MpU5No7hXGENfv4eRjeuiksyVmoEjua0PlUI6oCDq0rh0txN4hgKIDeQeLQUv2gSbR7rpK9gOy
y9A/qHuNBeACi8eCUASZFr2vAeqo6R09seWviMwQ8iu2L5B41vlDUISZbMXh+7i6beg69RNjL8C1
4J+h4GhnJ9CU2hOsYRPuJYrxiViTdoxAYuS6LXd2l86bnS8s8Ef7SlQ2O2Zk+Q7YKFyELy/nFEq7
QY+K1UztaeDN27Pfgz0pLMs0R+noIJRH4mpfTPP5RltRXS7A1fcVg3rzVg0IBBn8kL44jyW+Snjo
x60nxgmQHwEdT0S9SkSsl9IMzXEYp/bhRP9EzeI1+nt0fBWh7p/KdUzUa5gzS6G8OMOX2BTYXno/
OY8NeHtLXPynGo5FQL+3lRyCNNZ+Tnei5ZEdsZd1ph7L+bz4jyeuawqfjp+Qgj5VXRq7gEF/zL0t
RMgfCkGgoNRXaJyPpoOTBRYR4Sgln7ARS29oBtFMJDifbO4Gq4WqDXrBd+Oam1rfTEsEl/OrDGdT
SjahEmfjJKgIaGxxzELKZLypgi+LD850xEogtysF1x+JZowWDg5FbWylO3wKxsnO1n0cyCjOyWaT
Q0vSsUi122jwtj/7Yy1/7jo/FpAGratsohBWoGKnck5y/9Bvvpv0X5ilMDKoLASDMEXyxIBsWwvJ
m2dsqihZpFI30v1S/zksBn+efm9Ms/ewa13mqPQtKfRwArGfI22tuKimL1SKrmeP4H2F6+y5j9P2
n4iwz+GXzY5crL3wTyNyd+buYg2H7J16npCyYoJGsureTn0Qi0R6FPk6YlX4SnkocySYoT/NCXQL
2mjy8LUvnVk9/um0LK3quBES9ILtYHzFMLGS9k5sfbEhsv0awzGwkdu2fvnQKEyNIV5QMEE6hOrK
rKDi7C5dn8AztYVeKY4gu+MeKBVktEld21jENHVOjROn2HrXTMCIejy7k3TxKuWf02nK0/LGBOUh
hx6To2d1J8TU26edZi+ateFiil5LyeIRGpdIkKJB1KhvCSIq2qs5R31oLMDz35932ZJ9zqkQeXFR
hYELYPvgg+W3AxVGQu4bqRhIO155bwihSkw880KX2dYAX+Mc1Wx6x/XrBCuJk18suL06rj8MjxIL
Uu5saHyuM5hrh9N5W+P3kE7dBt6ULQfzDNu4U38vbmiE5qs4MXKipu6gIVJlRNFiN4tG+UWZIE/D
PNRFHBCVmhp/+TiuYeB1CbzB6O0q8M/wQHrp1nW5yZPuivSyNAAzqpOuVWolg+cqJasJoixrItzL
deaUufhchDYlktUxueRhDo4dz60lpEhG/wzEI7jcixNk3vIt7FnQbNyV5ySYNYTl3qs4rqlmShv6
t6khwIW2a0W34Q2QqXt35icIH0MjVheIlovmJKwQqQalQN2Fqe5unC/xsNbklWNKHvVPdpGROIlk
U5bXav3V2B6vlikYHIbGcVYpDOxHtJC6MIAgxCYdAv0E5H7WiX1P7X1SsVxcHAaDKEIns59aok9Y
yTgZDWkacpaSQ7G/Fq/tNmC46hX/u52PQwslHBW2gEbCq5h5YwWvNPuVYu4b76KME2qOyDKioNZr
qTqTxd1CnrYEFnYVxxoROPvGZb+JfcS6+yg/T8YlebXYXjBRfGDTx7C0peVJo32jAvU1LByRnnSq
o3uIJ+wVTwZO9EvRdIvYhaJwx+qIaGPVYzfkRtAjbAb/Ngta4WRAh8WWVfTmiUbuRPr5Bob3fhvt
HNC+JzoMx3YFTTI1KGIhvQbehKsWe4nUYlgxzJhtLTDfBHsMjLypng0VZmfG0geZMpwC5S00abwt
mWasmDVPKu4GY6Ot7jm+CUlh9KUIGBKtOcn9zc6RcESGAtM6UNAOl4NjZVQH/EmZ45lpX+9XEktB
Ah/BXIYDDbyfUxemFHKsV25AS+Ygjv8bFN55/Gsums+zLeRHMtop14QVPmptyy6ic+U+RgPOOAqY
KrttSuRyo0SWnoj5vTMSFYBIE3AoaWe4aYol99AD84XOu/ibRYjp1Ja7aztBfepZKDO1uxQ4qfFG
s7TgC/ORgMS+YMw3qea+RgYmdWOj/vPyi2bENqnH3hLmdIQ0i4W8aV3gBa7M/SWYUxUd7vrd8amZ
ANvd3wMg5VeGSZEu5vlodmmlSfRdMgddvjqai30jtJiWPfP6Y8xbJPRdAf70i+3EX5P/kwhSIYGi
8JucnYBk0yWSrEB8Y+SmjjKkmXXnTFUWazknTMuznzRAQuzG/1QolxSKbnC3OzMzaiMyTVLlA3PI
pNFuq0lN/lUeqkKTZ0rNMmXjYT82wYeU9MfinQFvmRictRu/KPK+JEnnGm7CQdttCpbViMO8Nq7u
k/sNq1KLE2utT0i2i1kBzpWqbK4KKVpFMteUpyXg/cl6xog+4Jbwk/BtHL32/qJUAHYs/8seMVGc
HhzoMgNiBKOuEQ3XVvio9twpm0EtQ1krY4qlXbktbBOhFb1d1jZgIdANFFuWP3JkZA0nRSeoMmiT
f0QN7ECaaAwRuWqV2Z4wxorCNNxa5teJUaRT9D6noD9IAkqZTK54ODFuaaHsnhaJ9aAJweb+a0es
+uCxMa0a6nrD1GXH5JY80SiAja4iS3l2V4+GuwgOBWvwMx06ZNu+A0vb4EAgIyHJwK7vg6oTlqUa
2aoPv5s7qsCpTxNy1KMIYCLgT7VrAbznnW4ZkJJU+Mo4RkUxrvndlvmB/5fdMD+kZrvK7gJ9y2aB
zM2LDzg5++78XhbBHLFCPeiZzt0TV1sre/bjrOivIlfcMeJn2lRye5StBHdrqOXI9Y8HAH5tDeUN
eM7z6YArFbGewvHQy9bnDyh1txMlqurK/9xWAU0PSz3exFCDvRVbvC7QH+mPzsqCqdWH39xj4nN2
LHd9RfwzzEPHxdu9SU3+hT2mRBCcfRRXH35qROsZIV+kE3Eh6VDW5AAJ0joS9+RYmkPtd0H+f3ml
TgHYZ936WCgZqViYgj/RL621rpLSW5t5NkT96lh9ZhalBMY5o99PU5q6D8mXAhty5MfxoI0Y5Qwe
B6R04w5hjKu2cyQEsw0HrcEwyK+ZDZo9taABXQchsDghGdn1V67JeQKUT8cZTUzHjQ+FWe/gvVHp
iKfWEafUUOAP+YycZuAG5B1GHw8V3jvSqevmo+/vrRu5DS6daCigwpeJCSoqYAFs6zTNkuxIW7bX
txZ3mqSx7HGqczJXT3RvDsPpzoutnN0TnNaESomQ/1pBcCZl2KsKHEm3CZUFY1/CuDCOX8ODQxAH
PYyxiy9Nijg08J/zo+cLM2T9Q6lWMIvq+/AY94pVouFoL2fb3XxHiBv9WCkbioeyfW5VFpdjoRCw
5KZZKjj6UxD49PuZiu2jL4hO/8D+T6Eg0vRXECp4a0ChlMpfePVo38E5tiQQsuUGAWVZOSwy2sQ7
e9aguFqyZoJOF7u6S0+/PbB1T7SDo9sJQSMFyD7BCXoESSZmBrcrRLcj7f5D84HNMgNi2xuTtaUt
IqBw4TN77ml8V7JeKWL459P/5JXvj6PDVLNlz/N6RinOZvaL3Gsheyq703VHG5nFJRzKZ57Rd9cn
gMsBceDmRkLI2i53J8c7qQ2iHL2hN32T13mvguP50QcC7oXZml0RmCEeePtYiX/xrEJW7ODQogSt
Cc0fOK8o+JW78IzNKQNZlanIq8NGxc+SXsanDfYEDz/FvY1hNrQ=
`protect end_protected
