XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������b�^�wm��3|R��kv����U��_�
H����
���&��[:��;��Ǒ ��Ļ__����^d�f�ؘ%����(id�  �c% �|8�$�x����>��Kӽ����N��^>�vt'��VgZJ�X9� ����5=^�<�KM���� ��,4��T���W��w��Maʌ�!�	>�5�N�5�^,������RTC��f؎���:�@ln�W%QlaO���(i�Xw�SFG���a�B6c?����qƱ],��_9�@J�x�$k�&��(�ŧ�rKYs�B��ݽ�〳JT(rT���Oc�K��{NU�^bU��R��2���2
�G�afr�!�G���Η��t�^�s�p���K��ά���&�+������/��I+�H�׹Og��hjv��DC�C'M�I����bU��|{��MQEƝ��V�WZ'C�_�9�^e#z���!���X��8]��,%��˸�Fl:<^C2�Rk��,p�?�-A�k�nO��~3�G�Į���R�Q"S��M�T�$,�x�Mw3�+����}z����u�B3H��ld�W���hb��:�� Zf'(�[Q���b4�z���\��!K֯�. ,Vc(ȁ��6 �;Z*G�^;�FP�d���A� i�.'4�B_�F�������#]��	](׃�s� ��_ �fz޿��u���I�(�J>�CA|H��_O�+nR?�Yԏ���������4%~0�J�� 4@�iXlxVHYEB     400     190y��g�����b��_5/��=��m�c��t��=�{���!�}[U�2��#ej�m���Vb�l��G��'7ku7�m-v�
5f+04bQl��M���@���+���4�-#���R
<�V6��I���(p�Pl�3k��$;��N{z�6�������Kkm�5򢻤p9-W��m�C�Ef!�����E�U����ӼO�REe�6�vb�x�Z���_-P/&+%�ڱhu\��·�By��7������#0l�Gu�2�--*��k ��R�o����Y�R�Ú�G�$��G�f$*X�bL�����[���l�z6/�SB�P��}J��c�X,� ���If���g�Mx����wiI<Vw��`(��Au,2�,����>)� W�fz�a�XlxVHYEB     400     150����ޫ$��,� S�R��Q��5�2�),��uj�
T���֘M�Jbu5C��*I�Pt�WR2��-�SIy)e�ˊ�vc����L(�<}���R.��-&�(����3c�,����b/9pт����T�ܥ�/��}�d�ν��]j4d2+(v��6��:z��eF"�M��rq��g�dx��k����~z�2�\ț--�+�m#�~�%U>����u� ��P�Ћ��|��st}��5��	�J-�ut�-����.b�oq=�. �^/=��Jy U�i)n�9y$G]���qJ��\����w���0IqL=ӊ���` �r�:q�>�XlxVHYEB     400     140����V7�fm�?Y	��^��P����x�џc��@�!����;�AgS�����-��%�;U.3�ՔO� ٴ�x_ک�s`�u���~�м�1�ֵ�@['��c+���T�M�O��a*����s�{?%���կ��ZP[�)���m���gVf,v7��c���6�eD^�����sY��̻��v�$z����f��~Dgɏv V��&�}�������t[�3~`�s��i0�<���P����?������"���Z4��o4wH��Qu@3���+�/���4�4��gO����Z˜Ov��g�>;7i�XlxVHYEB     400     180���ۭmww�^�Mx�ȁ�J8�cZ�� JՈ�&����W�Z�D�$�C�c�2w�	x��@ª��s$F	AR00�'4��Q� </���{�_��iu^t�N��ef[ѷ��t~C��y�Tľ�6��ǋ�Iu���ma�h!;��h��>���r�˕ټ(�Ɂ��/��Ҍd��~I������S�W��,6�XUo���&��L�@ ���,�ls��zG4
�B��Vw�WKAy�r��"&�W���5�\|+�k��6Ҥ��%~�X`_;��̷�����P����p��n���F�)A�:�,��n.� �<�ǳ���A�)�,��S��F��FwW�fm��8H��O믣X�8j#"H�2n�%�{XlxVHYEB     400      f0*UJ��)�0��a��I���9�	-|ή�2l�b�(������T}#G\����~.��0��)��4�{�z��Ɓ��;������g7q:.��Q���?]f�M��LDX���Z��&�[�5���>��~�ug��BcHv�\?�q7N,@��s�]X�0�߸?��3>=E
��Lp����|�u^�����k:��������Я��g���niB1�x�B+��U�H'XlxVHYEB     400     150��F�����U~Й�Lm���Y��w$�x|�l�7ǜl��d$\W�XfB��w1.0H�G[8_��$f�֒~�5n6��	��M�.����H�ĵW�B&l�^]�xАo�ʤ�f�YD�Z�* ��U�'�<��[�g��u��x8k��3�U#�b���=d�3�uU����S�9Ս,B�$�n,�J�������e�78jg?�rx���Y���I�U�Ӊ�z��.�׃1�bN��%���xؖ����^�a�1Yv�n�W޵��H�GG�dѯ�.q��g��p:�Ѓ�CAf�-KVVyY����Z_�#A�V�����I���xR?�1n�RXlxVHYEB     400     150��j~�L�7 ��ي�nO�X�$a�`;�qs��}l�0�P6��)p�P0���ڦܜx����Pd��Ʃ��/�s����oe.��!%G���?<H[8�	1@ ���f���?��_�e�&���1����g������F�PUZ��D k
�r1��=_���Ո�������*���E�@���	EB�,��eQ��lP���,Gtt7]��������vty�*�V��^�yZh�s��d�࣭�ĈN�$2�X���Y�T!f�l�R�L��>ᗗ�D^X�P�h�Ez�jHr��xpd�[�*�#�Ȏo�Q^r��MU��)�_huXlxVHYEB     400      e0���=��c��[G��M�l:(%)�5L��:e-VC��Fh ���hxE��9�ȭ���'?����ߧC��nD��P�d*�z@��Zq!V7�;� ����є�t�psܪ�H=����}���C�yq�3��Q%�G4п�Qe�:���V�wP��"��5�o�����S�:�A� �l��	=f�4lҫ2q�,z��'k"5G����toW�����GLhXlxVHYEB     400     180!���S�"��G���Ԋ�]�� rG���jcwS����cYc��;��O$��&!�t/~��d~�cDIJ�mꗍ�c��m|ˌƶ��:����;On�v�&~�&�����w�hS;��/Sky�ٰN�hwD�{_IWu�Ja�������A���!G4��p`�|EdYPU%�׵RdEU��h$6l����6�_�T&��y�o���ѐ��5RTMR��u��{�{u;A�V�d�,|Ȓp�c�ն���J:G�x�sB�!L��AO��-*��C�ɖ���K��d�wB(�Ux�B��~��&²�H�u�&��Wn__w�>��ʎ��"׉��A���=H�]q�:���f��<[v�_�Q,�(���Z�(��XlxVHYEB     2f4     100���1)i�>X��"ֱWWi'�,��[���V�1E�;���W Kh{ޥU6���2�{�w��8~Z>������>0DH�M��>1�����iUO��zq|ȴnȠ�R'�J��0lS����s�Ϝ�TIpA�����'�|�$8ZU�v(cw֋P�4X��%����51��f�ab������]U��&n�cT����I��;�h|�_�Aԝ��!�؍!>	��p�):9�����&��O�}_