`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12016)
`protect data_block
Si2oLrwrefNkmyexfp8ac58phKV5bJqawCyb3BMAoBV+rem8u6h5SIg1m2xKPGpDe/iB8cAgcGJT
wSaONxvxr/nmBb2fFOdpQdPAb0cfaJspP1DR0ZPtMkq6B52suQopUMyJ/mETLcXv57q7mpb4sXbW
luYE4VpCaED6D52uXjjYMBmPpzJyo+PkVJuFrkaG+lXeyrrKTDWxC55VG9WsFmAoOQ3R2nNMp02K
3lzvSrvzAlEdEMmu+f3k6oGtpVEM78hFK34PLVf2b4Z7YZFlTvQBVUGFGiY25qtG1VQ2eeN9L0mK
HQ1MKxXk0JeFjEKfmx1R4ijDdNyo2Yww115NfCzLHmIYLJPrUnsUo4B2+0SyT+D3uRWvzZWfyfiC
O9Cxyc19SGAcn4udqxGOLO83agP9agyffY7stmcnPdW3+1i1iMgRjqnQYfjBsOiu2EDklutHudWD
PTvpyN3hr2080cuQ0sHuoQN6fKpsX0GXE4k5ry+eLEQ9WH5Ky9pvaYU1Y2tQW4yVjdL/4tr6+i+/
cQZ0aD8WYNf+75cdgUyYk7dYVcASO/AhYJGnw604fVTfQ7J80LvnPPWhhOWI4XlZIhmYPRq0Kloa
r7Kc/9ihRRxOlEt6ehEUAx1m8uGG04jP0AEjndxS4eVw6nVQMDD5Wz4WyKsM31NW5BSoeXywH3zY
2rbpLf1n5xcbVHyd38ezy/jQbXvX/ZbFO714W6akkdFC2NOjtDAIE28DErw4TE8a/sH8gGAjE0ru
aMK0nGFwls749/vp1F5egz3CETEf15c/+FUWJ9xFxbr6Y9a/6wCLk0EwtlEQHqY2HPx+Rh0hnPL8
4LY75/VwO8LMW1VBTYrjDvhvpWCjSHBh+Vtnd6WrTCQT7GZFHg1tp9ldMt0hvxZnGibzYvVs7sT2
gKzFQykhi7MGR2JkcZOG7CM/MvvNWcE54JTMdmysVVzifwKUYD88DhYERm2v4O/SueLqzM2G859c
nfnPScpYoDorw3gkXFLZyNWMyvk/ApyyFPiXUEbT5ieyfeYbozhrW8+agYTBRWPn9Mtov70rSH8i
GQ6/zKbf5OH3Sy+YUtka5N+y3ZcHtLSJ49A/j9rdDbiXZvHlpaN1cDZX0FuYI5c8LILRNHVarg0c
Rp7ghNWX0yj0F4989pT1sMBTpc5tOC/FO7DkEhjd0StK3K5TGks5y0yJdzfxs5ys+CVy0sohPGaM
H5z+yBXt8LCpJ5UFdAG5KFlXHLsdOHl10Sq7qZ/DGzUsa1yB4RuZJLZavlmf3bWOojEr+HVynbgT
wpWtt0efawVTcGJoElirYdT8jSWRto5aAT5xpV4TUV94yEQp3tNk7NLnjfWEQFlPy6RS7o0uzTyV
59Cv2YMoUegETLI1MjteIl2oTs7BjYcSgCnA9flwh4f9JTwKt5ivDpPK9N68GeD0fZxBEQ5SLCPi
ipBvWmiszZfgn5CdodDMQBwyU4hj0q1NvFxxCtsNpl6cFmpPgjIhMlNEz8RSyjmaBpDUDCDDalie
A5xGp6M7b1K4eaO4owUuDZ5s9RGoi58D8nxErNeh6c6uS9AWPukGPBpjysDKccjzcizHUyRw1J92
jTR+kBKZ8r/f5R5rMUZgC8KpialUK+ICIuECba98Z/1z4zkCdWTKMUO3ZCmfeuc44MC2jNmrvnK3
1AUTQJHyldQfBPNzWOR6W+XloGYjQqCdexi7h5hRBrUQX6OnXmdgCY2b58CVyHiinPRnpcPKrl1J
RItrOQWmC8MZnCmG5rqaf/WxFWhP/9MSTP07vKD97bU81pq1yEd3GrY+ni1sJBys1vTmy3RQJtMO
BhyZCNcrD76MQHaN8cXnbMXd6h3BqWYFuWP9WnDtaHD/OgMveeQkdbiZ6fcN8AG9KdNcI3dXlutn
U7WDGTtK7/lcyosMC22Endgl3ZExIrZ6i+05eMk4Iull1gPg7iEmHPTD+WKo9mMDBisTmOb2TIwy
tU+tLdhthMWwDhXDXit+Xg8ppYKheHFLRhLsR0fdQ9YfV3Ent53rbPVHkIdvws3ka7T/VY1klr4E
gPfTUGCKCRSrqBVMh4USa/Vw8KEs9NHMWlV40Eg24wWftC+S6ln46b2HWlZuzCxtjum/M2o5Zrxu
zq0DrRvGTnuidQuXQXZRqU6rhvZlvMkcJIEmMhdextHuAmvdJyqHrxRAsWif36dTnmHjFh2bn65T
xsR0n3xVY3xsdgVZPCYlIChjcLR43Q/o+4Oyp1IaZoLrGeiCCry1UlcHU6R4UtQ8H4ztoDXP53BJ
eBourzb+tn2V+yyfFVZAgkddEGigsgN5Tn6jUmR4DbtNZhmGghWiFCmhFHUhaSYKugjX8VO4Tl+N
xf/3BVDFskrCR9emg5e6FQuY9LU52HgHcGV67lGmeGA2ERn37piHUAj00DFR+PoKKXiwcryQDpAX
0Ka+E9H4sm5FW1D6b27G/oZTWkU7kmGylPEyFIB41YKjjTTpSWufuCORaDsGV/bqIOnWAcN1E9CQ
Wf8ZIjyBOusQrNc+0VCc/g+t2M2KIkPuo+cl4a8dqDWO74z0S0RB/Ez12cQAehWK9imgRBdhTy5X
yStsGt+rtAf8/LP6IMVbpGtMeA6MgdHWTqMJxNmROW128ywuDMX6QAJxm5jVE3IXRzyeQLcBZ67I
igtsQooqXjgKIxUyTAtjAAnZKZOFYmnkj64Dxghqh8LiXPDu6lp2PQ6+7jEvwE6To+yiFeJLcbSC
qCjiZcPB9uWDPnANmzWU5bMfll9Pg9kijYN15gT91BfdcB/EL1fkWIoUwMhWTyfzVgDaE/aQTqle
IfvxchpksIZsEKCHb41oeIws0bDg2L6ti0xlon2FODwFeBvLSMiPV7vyCk98QcMeYKekRbAlRlLr
IbHAGUIDKpab79Jfza3FnYPFXk32d4pD/G4ua72uAZXxFUzSVJ0Cvtc+VIHuVvIxFpFK+6s69ox3
Sn5xrbeSBzYzMzqIjlueI6XmQdbXuLzz/l1+3l4+VcUvvAlj81zB3vR+aLZAIL4L8DyAf/EEwgIb
z1ToEZ9QcJcM8TrDtVJc4zp9XKA/lRGy6zmDMdPZKwyqmPtG+Rk7gPruuI+6cQIIhu/hVZjCni1k
/myps1hS5j3cbYGT1l+mBsx/Sc9NyHYWUkZHwefQw1Sn8+ubwfifRy/UTYYCcPj2QLmWfjrh4Y2V
rXuowp3LsArx6YGHq0X14SbTiMBP3axuWZJPUlW3cOhgV0g04IgmbWNGAjhy/TKpXgS5kmeHoNy4
BE/Aurf9fqjXCp3sopFrN88bM3aHR/LS91u/H/MRaa5TH08mmGcQ0edBH7uC7jYHHSvkFO0NtAy0
fvGgxy6PeUp7fZBPRDdj1HpWHx3o8fSNBj4lQWJXPny3bB73t18Ho+Rlo6tR/pmfypVkn9fw4BNH
pNS6dr9RT2EPvt+JxqIF9RU40oIWeCB8HZjSnhJOr9VvOEyNkwaB/NPAeIHHOg2TEwAPKQ4RtlSk
uk96o8EMG8HJQ7N6v5zJoqbCGQgWLzMjLjAttj2NiIxB4GJkITaADYg5ka2rZHiXSjvmnp0jz1HS
qjWKDa9ClptX/inOlrJBtlIFKKmW1X09DHR+crqXSMNcO+xkQIYYDyjJeXsv9ShwuQqvDYjTK2dZ
d8o6oygAZi+FjscdKIXIZ9P4BZRr2ojFsoCvOZIXV2/gncRGSIHReXIvweMURxS9K1KtcMKVWKvP
tPWiIoEdXnbw/pCj25rLVeK4xigdYi4b+SMIwMLJVYyrRL0d04bQ6W1HXBsoBcHT5NFv21QXmisX
cB57rtfJKNsrtPeVOpfM217CcGusovmB/BaKIeMvwdRlJReI1RZpcBJvscNIFY0qBYf5yutfI733
8mou3cIwaWD8EZs0y9hoHAY0obNrS/QtcfnR4QBB/7fPqLXjdjGzPrDYV1aAGS/CBd4xxcXX3dvo
9Kt74Nm/U6hfrEcp2ahj2lpN6B++v34Uw7mn94JlVxJIue126F6JEZ4B0A+Vg1BeDfuxip+X8Pbz
AwhOPkUIZDh6GViAbZFp5HLLS2/gvdg6qNhPGLbQ5xKpfeFeY3az9EjJieacx+uy2Tt070x4Wror
bEpxyyUmvPZQKrSSSiABlkX2WxdfNx6wrgTPtRSOyJOU2X6QvRs/HDrM9Q9um6XE4Oi4PEx5TFvy
ctRvcU7JqUfbJ4D5GoDfbvvyu3WYcnwYoJ+6YNfHy9T47fY7v3qCTlsNU9kyOecpB7eRrsI25HHL
Ghmx25KtEmm4rKnQbTXCS2UgRPrmyW1fQMCXDMu0Bn/Os6UIk5kcJKDZ8xZKXG9oj4+VpldIeeEL
BeT1AhbgHPWT7dG5bSTeB9NXOxydZzwiatGBMrjcVSxgHvGxdaMrUnFXGVLEgE1Iv/lPH/JPP7tx
D17x/yhJO1ZNj4gbSaQq/o168zG9q9mYDo0riNDW2MTKes4dzvpmABsH2m1AeyAD9jBYUlyjxA7d
jZZ6+iwCVjtIK91F4dulo8OaMkbtIwaXhfVFWFA7lp9Fk3N5wmIpOshn6zcPE4B1UyKAHLwS6ggQ
nBP06LIE8A9vKoRJjuVAtA2YXPyt5QOJ7OMeUyelzZ4itcywqFYxYKeaxckmQXH+3+R31XbTkgPX
xOmA1WRMlBS/4wnTEuaUayDcHMfi39T6p/MrBXT+wqkkbtZv2DxaZ4GujVJi9DTV+JsnGt5uin8d
ICbEI4Qg/2ulS2L9JdsXI81lYo1yUP8j/12Ft8pJh6NMvFkBhVoIHyfUxJqSN6ud7EjEyiWJMYvk
gY0er2LPQDZBBrclnnn/rfyEb09lSGhq4WxTQVHIP7ZacECrMZhO+PXZ4vuXERZzzut1TUKa1YYf
6tmHNeLDnxqYHHXRy/wPLxXM58Ht4AyGMtr/bVon/GRrBCf/NYIvahP7n07LA48GsMJB8zg4gftL
SobkMQJgaavem1Sps/ztoKkQ2Hf7qTtORqLFU1wm46IutrwDu1jEhgq944U2cqtj/uoeIBFciSJz
SvBT2KgpvN3z1scbljMqrXrE+7VDeAl2LPNzhZ7h7zb+D4qdu5B39YYgP0fE57cvrTJNH23x03fD
MwMYDi+zZW4Z2gqYd4eXa0w+NIXOggvPSfKpV7k5MNKTfhagU0lAtHtLVKHocLyjOo8h2jGZxhYg
6Vq3u6rZRN/wE2aXBVT+fxlqFYDDFWzkGH6r3x4IMhdnDk4L9fPj8fbNXHyLiZwglsZzLXOGpppp
zSiIx1i4HFnPG/qHdl2zlejn509Zoky78gljegdY/0vWwfWWO9tsl5qZrvhcGkSor8Ns4RJpLkNO
DWcu/U9N5n8DvAuuLBzwyzVI/E08sI9StU03+xp7v5ctXr9jP+ir3I6o65Kd4Roaraur3qEueilt
n3gJSuuTLBdgAlwy6i7XIhlXbYae432koXbNtJT2ZbbmWP9+07a2WQQiDB2466jTOVmO2F81m9IK
k52rNzqLXUidk3Tthe59SIs8GjC0BtjJ04fELuD1QJtQiwCXpIwTRuw4IhjfBLMdtJIOHI5fdCWE
b+HsrDhHHENH/57X9kw7fCNtJPPizGl6hk9hm+DLHo5kyao4i4eSfhBSEcr/CZOprwlgPbkzO2c+
Hm7Pa+BTYKcpMi8Okduinap0bHGDxc+g0EuIIh/D1qm3YDqMKq8s4Cd/fKb/m2L6cO2hSSriYDzs
erB7uYOMTtwlm2vpmnGbeB39eF4Xb13SZlI0SYG39VSg6KVRCEitG8KcKLGcpEXzatBm1P//3pj9
y2RG2jeWA/1PPWmxUeM9GYoqW8z2pItcOBC0s6G9Jj/FTRdwfBqwNEUVYUccBZT92dPLmYnwJ4DX
ONIiwBXDwnEIp4TwZsq7yCzIjsrZjy8jtiKQJ0JbGWITKWDwjik94Injm22AmMstVCNvub7+ZFnG
+PSFdFC75rSZ44kd5PPfETXHrZKQDTcGQe41vqrTvfbbFSwvOgsVBJ4Q+pfma6+U+qthw1Ijlua2
j/kC1i6JJ99BVe3VX1UsHHv8AeGytTY9DqwZWrXc3Mg/JXUvsXcjzqcvlensp8HBog4BWkEO5HBt
xw4lCyzy16ZZBWBedEogQftXxdFZwfYbgv6Pn6ge1OGLl3GjnLs931BmNlb+2ol70YcrxmMvK9yR
dRb6shHQtQ1F37RVdUO1ZLR4Lw5deLVz1kxq35Eoiv+KXQKALPgvIpfEPTBRKAiJGA7UvnWRNLXe
FEMq/85qW3k4/4J8sXEuJJ0T86Sclm9ffUwiteICrBwAz49LVdDhfM9AjW7eF4SjT/mwoiXiMR/i
AxrQw5OAn+pJKHWV8okcx5cwpOf5yGjKouaSpt6QkOqnt3EkREfl5aFDc3rEZTKXq8gFFq9WlaFX
V3KGA0jOU6cncfriLixPPU86GxWkMZKSbcDv0AxL86mNA5Hy+qrzM1Yi3Z7Ff8j8fx61WIBvzXTv
SMmGJBYrVtUu/akb0VC/PLaTnGZIB7I1hLegzSV3njlvFBX9zDrKH+/ooaPEEnFMmonUN6Tw/rq7
9oyhy1+uonQJ7j6uxrLPlwngmidWCYXVgRmwIasXEqyX4pWnjMFV1HlQbzIY0ISQxpCxy8epNWcz
tWKa9WPJKzeSr1WtxlaJK4YoJs+OxFG4yiLdW6JsGkNJfC/XjHPvrB2gW69XykCeY+caf+1RzoT8
QxrYIpu7/GFgxuJBJCkdf0UuPIlXjvn4PahEJUbi4/108n/37J7R/WFOyBLO2d0YXBaXqjWwvaLD
VuUoKBUxbL0poGHq3bxMA3l5IIfibeV6vdH9LMt9GDMtIyHgxupHfkIgM8SWH4VzOaE1UgHTFEBC
mJcCKpA/OucIlVs+clltUDMakbSY9wy+U0NbWAvGJNuWjZJU1p26TNILRC7OY+1+mdRHAnX54RtS
iBQsO+YgqXTR0gG61Qc6O1a6gLi7qLSGw8o1mCe5zHoBYb66N7PfIkdrRDlRoqtremYvP/hcn212
Cp/9gwl+U3twy4bOk+O9oNcF1IlkD5vKrmanfXH/ueAdLt6sfjRzdWvxmCl7CEwRWc9bA3vBVzk+
scF7/Y5ktuNTJTTXAOt4tk8REfMslJfExdOa2HhuODf3f8lqW2mjeRtA5ZVgN9XHjNJ9B4qgyX+8
X3Ls3pJpMJopFIpRgEp/leIIk2rHVzO5weE9wU7BI3/dqJtVdbdbydXPevJ+brrzhux+vuaSICwz
2S4Pu6HyH12BYAX/yVQ70Ga1jSN1XLUVIQPMq3silGAHs0oVZIHmReeRJqhSfNZyLUBY0kFlOWDj
6kP6W//nnw/L28FhMy7TxiWZWhdLywJtVs25mQX9R29wbeHVl/MyYs79BOsrVL9oUN2a5SW+lu5a
M35ympZrVv4mZVArjkFDdlsCnCDllitSkd4HDnUlKp0ohAYQkrq1Vj5UlY9Bi0am0OH4x4MuxqlS
ZFHrDJpshJJm2uBYStxBKicPOzlh7r8P0dpiaTc2gaQE82hPClR4LQsm527CkqYTRZjCwA9sE9Qa
KP4jb9vl+5tEU87NjtUTV/CnJKQ47pWd2OHYg9WYH2OEWslaoumpNgkHtrphurC8mzD+7R48eBD9
xEerSxxd/1xeCENXi4AQoJU4dBzny/euPDa6Wk/xlSeBYJILTK5VBl5qzuBncv4SZ7IM6qHFtXOw
9U1h7tDzMrUxHotONv8+QTkusPDzYGSpTiqueIw1bRsSQfyRS/6DBbfq1FUtD9lU2618idDkMhZP
U+sg9qLlatH5P5sxlStUQd4KuIJIcKhm4RxGnyW56+0PADqp3lRg/c1pn1ZcJ4echJWVDcoGjCK7
Ldnvb+m4FLh5em5kHtaFJLyJftGEI32RXnhVY4Dy4n2BRoWYCiOs948aoKXMO+p02H+xw3pj0e3S
Vv4PLUN9BTM6uU3duxn6ahiSlcybxi43aoaAdOZoHBzE569exIBGgoamGYO/29PlD/+hBPU+CDCB
p2lq1kcqB/9ttBBrfcrX1cmAmZpoXY/6jp47cFwyeD8QZTFcxvmMXhYrjKcPGOF+genhKqIWUwJX
tl23cmg7JXxTkE/ZnSP63CA2eJonMB2q/cSlswwWHM2beVKn88x34NIYUaS2XmvYQnXe6vjFo1tU
7LOwHcvGfbRGMZDl6p13x9vbOWaAOsl7Fet47lsXhfrciw+b4R7/j8gIG9n0auv5qvyvsBkt9QFk
RDuUOZp/rYlmNYcWOzj5TIQywdiTYUc6CRs6IMmoV4nHhFBhuH04pOEbhd1N+HDvFJ7vvu7ct1vO
BDQVcD4YXYF7BZ/I4SK7J6ptf+DK1FzVeKNz8PKlpbv/MVjKPpCiO2MKpeO+NGVopRyZjRgUl0xE
JIWb8HdScxKMz3kzTWHzo0Q97s6xNVY+eMB34QihQunPLLG/MoQuGzLyJfsu6h0CWtvcwI7oyU++
g8n5WHq8B7KhZgTxWbty04x5d7dblnvtjJjchkoeoLTko0ilHnjZswmixJOtYCN1EdJq/TRn8D0u
1n9VdKLVA3kBRBA2zN5BjGfP+yjT+gfqSwXjtBCfzPmqXm+yPArMWAQL1tb+K742rFqmhacmyqE+
O1qI6TPqHwvS/2DMv3RBlWyaLC7XvMrLprBLwlMg/cV/6HhY60vrpM1XkCh4Tu8dE3fNnMUXS7OM
tKau2tiEAaW4DKOqL3gmPlMuPUxROAjmioDG6TtsibbyQfC2aATXoFNUKJ4hoPVTMYGmHSgOl4cI
G5nIg0xSrHnurOU3NZgxlnnLBJcHGjaqDNAqFnVFHqMdukUTuz6BDok8X7gA9ZlJK/u7xVMyZohb
Tn0ytChwl3XLuPPIY/FBbL2A+vfgZS5XddA/innGanmwaFhjAQvkDVJ/fEWeFrJ2PZmyOvle1TeJ
Y9op2NXDOsNkS07aavJSDhruHZ/lMvjinqDhp3U247tFoIwZB2GqKOSMW1CuPsjGtNQ6PQWkaF/5
bbm1CRxdux0rsZSZmIgNh8753gI3Si5LuNu/MXFzoyC89IitmkZK4IGrxGLZMq9JSgnSeUzMrho5
CBMe9PmMFZmpzKhH81F6Pf7oZGt05AawIgE7qrPlnQb5RtS8eZivLq2ytW05Oi4Mi9bHTsGNojT5
2v/03zkXmjjZOB2J4crupLnYzUFg1rSCZuKikqu39UMKDyir+E7VZeBl7v+EsqrWIk1saodZNnmR
Hy0muT8lR1xvjQs+qCs7tpi0FavVrOhmsaYVX9dypoMe91AJtB1rfIYq1LgsOkMLNt/oFdI2IGPm
IDVOIZlZkkd//6zRS1SnDzPiEk2XQQKnXYjEPoYZJeqhhHoCngYHOhCIMOnoSCHL78tbBKL10igH
Y6gHZpLeu8dl87cLg4aMjYAmkB+4AzCsBJv2LXnfEkny9y59P610Cd0IsknLXKM6+4lmOGhlQpD9
qc4KkhSQ2FvFaoKprfHLsuMD4/0QS1JKwy8amvBb9zPvnzNneXSKIgB/yi3OQa9QDfnjQbgUfyW+
DZNKW6sx2QrxobIsrumcQazOnRmjJaR/Vgc7YIiXvqjscZNNRCkhyRa5K1WRkrqd1RmhLOIY7hrY
7SNAMguLzMiAQtn/UfFvmrWBF8Zl9oE5pprCV/bKQYGe1j2mdcn3MlGBQVsaBZyh5ENL5Y9P/0Bi
/1rj8W13RBUaQiQb2sNdsOlzhR2gbBV4nvOJo8KLNHvEAWwwR/ZMjCimMXxut+ZFyAiPmzMN/qeH
UcgXRBQJ2WBEALOAIqfEi0oihwHF6VOPjgAWiLNzJrz3egqXmJ+BoArNY/lw9rwmBxAEg514aHZl
hlilDOL/ErOOJYolwjGe/NWTp0s2HnB7yKa5baTM5CdtrTqBGDtYrxQ5ABoJmpr5CUmun36ceAUw
gSuRuh7VzgIgdh5fumQq+WiKPml295kfxpqbKHM62hvnvRf4NYxhmA4uRaOGt3ES5Muk40bxAWK6
FJ6GO7/O6qNt2Ijge6x+YPqsBMd3pHRDz4f1pmXDzKH8Abm0TEpgYkZyWIzcr55s0l8fMgYKxWTL
UD+m4pUzIH+8NSOVWenNGbAtzhNtvj4orvPstdacPiBezsZyURrroNqTGIUeLFakekulcLxQiDaM
Rtyj8Pwhuamq3Ij7nCC5CB6IP9XesTKUxRk2iNEXnuXN9Esk4QuP/xdFdIzgWBYp6a+uhUjYCb1Z
/Nx6qlxcn2qrFccFCzxVMlqFLpUjAbS72dKpUnxQfBLVnw1haQEIkCawoUqtlrdzNTRby5tzNFh9
ADcHr91/4sUYFy+NL6gliFet48cCRdEyD3iQHKBJd9kvwzuWh9rx9ODRdK/nCH49/Jv1QGVVqLWv
W94eTdCxmDUaJ9smVOatY9xQWtLJ92Bd83XU+8WigkXe1Kcn70qQpD2yz3NBv6kQbSDM/uox3Ys5
gljz/iRSR3lITZY/3B6SnSCSc1O8cGKD51kVM67Jrxjo/KYjLF6JYvQ8TZH8ZkkSlaBM+7npNaNP
Z4z1UwYcpZe5b4iE46shb+TXU+u8BGJ4R5T3PjTd1N6k8cD26KhVeQXCgCrb2oy76+gyu+RuB87K
40azrJCE/xQUVkoJqQijSNtS4vyna2VbSTpa3GesWtEk1k1cEXjy7xmYWR8wGQS8YcXYoejUInSw
SJp4amxZuVqLhEDCBZ5A2px6/4bpLNfXr+u71I9VCxiJcOwjy6bDe9D99IDPIQ61DuDcgg5qLlct
XqgP5IxGHRNbxHt1CFX+4Z72C4qBsFJnHLXzIfy5b0YARTdZ0YTAnHSRxwDre+Ri4oYtAZ/fzIEu
XKmp1seu489PILXY+iSJzalnLOKOE8nDdbDlldbmg3Dubj+qbU75VNO/jmmOWTd9UezbGX2Y9XST
mm1wEN957rXxN5B0CMzAeA0sYg0uGeT2PyrXmXRxf8/sjD32ox669USNs5nB5wq2g9sb0euPnnqW
bOBMHK216zaBzT4oafiBswle11HRkl1L7YBly663f/EOq2mIzeep4JmIUc5QCmAJK0F+Syo+/32h
8xP2JPC6QGV0zYpRt3UNowvefUkRbaRDbVIuuFFKoydxhcP0ErXvGO2/pV+wTx1yZAmLqkP4geb9
9kSZPOr9egWKsQybPfQ4xAXfEop6KuXNMCjhbieH7NlfG7/1B2xITDRaM8gKA/kuVV41pBvfQ8PL
2stNc7/P0TP1a+tcN41oOpyjxG56g3hHomCcCULZoQae9HgUsiVxfnz9AzpahKg+bLuHkLX5MIBS
4aB5aYvGu/mjg+amn32GWfkoOD33ycLnsjnQLzGKVroTbgpkrbiXmUrUkJxn6nNnpvFqR+7KvP0A
8gXyxaiuYpwUm/TZACxJBzx1j0aWNdwaVjwYR52PwT1/GPSxREWj1g3ar0ynOkjNb8HEHjk5cluB
Pt9SAUPg7kMSulrTKLUpqCyooFmWBG43kv8P8fNH0IwF3BooVoPjW07bY+f6jQcKkajFpc0vwkKf
O87NLMP97xXXvv3KnrueoVmMg3S6q6ktrvgKXazNojMWGXcVUcIsIVzqXMYl+n8avwASAfYp/c+l
WkHcR8bVPInjfOBL330gDwdtNIWm+xvLqC4nJrJWB9TF3lmEnGJmaET5xD8uw35gfEckk9yQAoxd
dRZPxIYRVoaO+I2fYYDnzg5Nsk48rS7LfPj62JnM1QETno9AuNrS+/8itVDkn+q/JXZm1oJmyyXX
0Xd/iBd1TJ/dAAQGcSvyKKg0mU5mjymZT26vgCrS4bLOUV3+ToolNMiV4V6kf/94qVM7jMPpEKU5
Vb4QjUrx1C6MR5FaAS4djmpv5FPxvT1N5udeWINsdi6omBF6wwd94jmGh06EMrIqiUL50oYMw2bU
KsMN9ShSJPGY73LnqlIzkZSc6P1yHFzPeNBpdi3c22p2zL1Sj1mrJSFX63b7d6GgzBijhIGU4rrV
2SOX7KKTdDPUQYPE2xvq0WvIzD7oUVEGZLrjgXSvxCY5kV0xmYhCM6N19qKhIgsG+oZGaXRJAwxh
v0QfHkR6ipLhOGSSwh1h7/y9MyIml2PkOd3obq9ZavUgGhHe9a6FFcuvExs0QSSfxsxEdxCgz4Ui
b2BLs8vO2tQZKucYs8niKBGg/u1YuqUGk3ry8H4s+LYx3Q7JPZ9KFMHlGv7oECU9fJxEi/gIgZER
00nKWJnth+RJ+73tN0Jd8zvahc2/RXxndHOOppb3/yhABgveeGdd2LJAE6iaDsNTODarhfBUE3lt
Y1XiDvbNxIu7y+bOJbytnLrFJZOzzs3CTWwEWKnb8CVX/1xYTDD6hoWotalLtTTBfId0lEfSiIQy
R6BREGdz34uIpadoDBZHZDJKb79KVeZcomCvWOf2OhJ0hFqrHzWkad9Fj1jBhbpvRs+AKLtz6L9i
CE6vRSoj8Ve/KN8yQM6d5XnhOnM/xmQd+udkbylrTxkzVI0FAP4lJ4G0H8E9QyCLfBa1qWKuDu71
AZxZd4Axq4h2GbLUfzgoPbJlN9Ggy7MlvU8ypoH7PpYnyljShBKXyBweK62ibkGc8dJFqX8av94Y
zAA2M9NXH4Znzyz1WwkGsBSG/y4zUn0ulI5Sar9nTnSA6LmM3sHk9ad28bC6Wg0dN+7ugLFtnqS6
WXA+8YFw9wfrmQ+198x8eqBohdDqE3Wvyonf3PI23EYDk6/MjMFB6AV0zAIJAWNjTVhXQ3ihiRNK
cdsE6kcgV2Wixd4IG4bbQfXdWtdkavNgjiIIxc4UxlCy66b4wrvRJ8NHHYS7pdS/zXvr7nvpe7wy
Og3uN/bgMLY8uBquAOmdGE5VuXYozlcHPBCGyZQ0kpEvnwbL46RCA3x5JCjS+sfjcym95+aVvT6G
QGdAMpVAWJo+vrHbchWKj9ppI1SI9cLzle9mcS75ZgJ1veVTtEYjzON4nzzKEhmV1QofHHN2Two8
oa0XlHvi61/RbP2IVlLilHh9VD2teEXwE0mn9SgOMnASYHpKYxm/bfbNUlElfwbb/YwWfgdQKqo/
1hgyFzqPPTwCxhWZ1xn+jI/8L/jcOQo//uqMTaPa61orR8ymPBVY+DgckYjjyLJYE/V/xioBFjIF
3FkHi5iGJFbuNBMr57WtUIAPnxU+IgKzISyAFeUsrZR8HrecY8wF4T+xCNrlh++DQ23gW6SVGezO
4txKe0s5+d50Y7ErYAb4lCBkyvP3m/QOqN2VKKvkuOaAEOgSJ3UhLNbRMUPkQCqoq7JUfwJ4AthK
LXZff5BKvnXRWmc/pOOublBWNivqLr1RgpvGiCep1dvHWXqzlrv8G8LKGyhMvdvUkFCqcB7F0nke
IsnB2qLhvdMTuVnMmnxUad/CLX597ABnrfJuk6Pi+RP6sUt0mOMpRd7JxVD6fnQ2YF4X/yektv7X
KkbGUvyCyfG6JKHQeYFCwmvOTXtn1iXnAQOFgJucvWnTWcUb85RucThyDX4CgND2msSUPbvKjn+B
Xo147N9p5qZgJIGR9jcVs2DoTsA1Dg8Vag33nE6fErdl6b2IRAfsPM/YUMzrriMugES5RX9XA6ld
TMH3Ey6NkW7XrJwQ0hEa4QC1iHfZN4rgv6ZEqyfpLvgyuHPJEMo650Sb5sY1BmOjVAw7FACkDSJ0
jNgcVCy/2ZYAlufdWO/vdw8i1jAWr49h1WEnA7Ft/pDUCArVFIYBytbJs2b9A4onZrGpXGmykdfQ
kJ1LLqo7bfk9TeEYA37ucplAiNu1c6CAOPL7dinSsycRQsZchm5ps0tW6gNLJjIMV+35+CLq6BsA
f0nggjrDyb2vOemNE34S/9WhCvksCW77Lo6q8zksWGk63rT/Rp0kJoRkK0r84kaf/Nrxyy+sP9/D
DkpI4zSeLSZK8elvCDJUHfargXfiUQFY4W4xoN8sFy6z4I85pHfDML0JBzdwSP2JGafEUxrE/619
W38YdK1ANan0LW3XpTL4mY2y3pa102aOJL1nHO4EJt+KfLMilyBfG1Xa+ozWtiw4EHoYjOp6BJUy
n4chaQRD3kuTJK0bigr4llZuMCb9SHV8m56HTGuSAd3uZEAEfLfsbqqf7sXZ40vK3THr4henubuW
Wenrt0TpgejGzumVY7NXNExFOeHehFMsJTYNC+eHLbjgKSgKyQ/0C46PVisuVHNJPgBN2WVu9lB5
CZqB2xf9sUsh72MZJwO8wg+3nmDcx/0l8azfR4w6xOq1NtxXu27jtZAQ9hIOENMO0nyJSWg3Fbcn
y+5nKFTG2gHdWOgT22njcf7iaVucd5I6oovDduG7GR6JmZIqU5m4r6CXwf5K4RQ0E72STdj/FalA
ccuuZkrxr5i3S01kRKzg9f5oBFMrxA6vGd+J1jP0RBvlbo52leGa4IAvcVcsNiL/DAOYr8YVVrkS
58ede4RfAa5BWs51rV6ZSafrjn+ly4HpFEAh/PwvIhjoJOzMIEzcj0+qN/8zPtD5RBq6k/ST3/Xf
LQ/Q/zZSLRe8jCF2JtWoI5Bt8QDtdG05rJEQ9/eGnybGN5ln3idt++Zi3ZjnXMU+S5Fvngrpl3UE
chT6m8+gCvcaR+OfZadKvmzFQZJFQbV1ulCrTJQXPASBB8/G6OknlhF20k82YY2TcrQyfCcnMbys
hBzhlT3uq4j1Oj/GRseSv9PK9RGjKP+eDZlrh4InlGG01BVdjalll+K5u1ivVfZtOL7p26Rr+PJG
HNsGReqYWzwn6SMWqkh+XX9c7LvwGrRjo7rn/chlNZ/nAUrvdbYpe8w4M8N2YmNGLZ5G73OsUrvc
xnYL/cu6v8XDMM4z0ir+fTQQ4ouF7puM3tkLrOuOfrOrN0BJMRht78Fobjg1D6If6B4ecFuUkv+d
d361AEOklk4NxFOWeaP68fj3y9Pa63Tvu+RIR3beah/3Pd5FYXecKjHDWsflOS1EN5JG1vLjX2Qj
ACPfpsGJJYpYILwDprM3nAaBryFX9MyxjO+iNzjfs0a47I5oUeZdQwfV3Mw7PuDVvNSNZNzvswvD
AKs2kyvRbC2CDcnDCanx+jVYi0PNX+/wCtIbdaOAS3zdSk0bRYPnNKq6xeVjaIx/6QuPfk2+Htvx
G68CxORNXmnVr48g1cm9DvuC3OjJXBp/NCbO/9LnYOnIVGTbDJbi0kOiwSvE2rkAu9xUXKZP5Ftl
o6vq2ZmUZ+yjXIiNtgl1vbCsOQghMXjFHbK+TSk7BNEUTJms4w4bripK7i1mEKgMNOlZjdr0v3VR
Ak04fniuDisi0Iar0FdWDOIQQLTATvYdNWPOOA+1ctcPpQtQKGvFipNiX56I2OCX6ix+EjuzpxPv
Z9NVAgqWmHwlZGs2LPHmuGdowOQTawANbYmvAYcxsEuYDygrqY4oKLUk+gD1yhB+JCOpGzjsMuXN
DNjMLV4cwHIHiuoo9AC+Qkd20pMT4tNgbSb5wVx4EI9OgFDZ1V9+N8sW2GSqkkAeDBMAa8UiWEx/
5afCAC1msqQzx+XJL14mW34SCK6dxmWc9KCjoGBEw/WxUqzlfrTPBg0iiRMBsDDRAE4EZ93O0fi2
t1mWllJQXa6KAPbFCLA7/fT/LQ0kmGekAQXwZs9Dz4yPaM5J59qXwH2+HWHB9la5v8c6HZPO+P+D
QbkXn8PnwusBlofhkMZEEDUZWqOCK5IK9Z18YcPC2lW6Uwcpz9p0CvdXo/tGSHQERPez/6QdsCWg
0NYQynMleKepA2ovLtKBZXU+lETluNOQ75LR5cRoq5a40tP8R1P58fO88Htb8jH1OYJ+mk8DYb0S
eLDtEABy7uGPi5AytUe2Mrr+9VNgsfHPcDB8mpbOjAO5tqF2Qc2mrWmCfkMk2fstpdwrsE1UTUuc
i/inNsiaJNagvCPHP27mcAWYuYGjzJeJCJ9jTiX0IgFZqau5Fzwy02e8qV43laLJYGmqaS/O7GvZ
xNYUPasbF6+4IOMdAaL+NdEw2d2GSptPL4bi1JuuAMep5RocJoFeU/1FqZCXZAWCps1J5MxTRkeE
IBv8OGMNuFptvPm2yS1MzkBTc9GvmlQpoqJ/2lZEi8uQFkmcZ4S5BQUaVQioKQ==
`protect end_protected
