XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!%�4Swm�,���?�G��@�7��L�\W��ɺ����]�Ϣn�w���4�'m婏��qRW�����uI�����������a�8HF�:������ݯ��+�X�W������
�,<B�5�0�;�!�
�łUށ��=���2��F:G�g��X������Ÿ݄&0%O�O&\���gvLwo����z�Gj�ʗ~��<�O�	|g1 ��:�Xq4#v�:��A��tW{��ł�v�U.;!���ɴ��}u*��3�?b��[D|;������Smq�$Sm��k���x�W���5M� ��=*�`0��T�"�*�Q���(�������|��j�f����ˢ�Y}DU޺������d�g��N�ۀ"��E�ٶE����KE ��+i}�s��Igz��J^���$9ߗ:�cz[+� J�dK����Ӝ�X-�
<{�?-�����;��S�AD}t�A����\/i m�C�	����\��;ʘO�,����:{�."(:CW��<��w��4[�c���D�S���F�0���G��Lk���dV�!�� yo���|Sc�#ڶ��#��4���t�@*�=���6���L5�W:? �W���]���B�k��%Y)�۩��+�g�a|���na:^���>:�(�F|{,�]��Ę�(v��඗MA]Խ������gVq���y0c>et|#��@�-7X�Đ�Uȸ��h���7Ԯ���8G��g�ޯ!R�Oo��ͣ�lXlxVHYEB     400     190��\%�B��ڶ"`���2��h��«�5Ua�٤�Q	a��XY}��r��j�U�� ��mS����M!A=-_��l>��q�v��{ZH<cc���&�f�j�/t�܈M����My����������y��x� x,��d'�8��TO�!�Ct]D<�3�!.�C��cub&w����{���g|���	G(�:��Jc3��ʚ�^v,@n7*Mc 'O���)\�"�td�#z Y�_m�n�J��·z%w�9mv���u�t$�u����?Pj�B0�<߳	_�y�s��X�]8��.�:i*���sh�[��Q<]�n���v�\�0�<X�D���R������"U4��Ӧ�KՐp�;7�Jr�$L��k�$�3�����3%r�:���)Ӿ�XlxVHYEB     400     140�-��H� �� Yn'���5J�E5Zzۋ_e��x�7��Hc��]4rB����Q��.��(�=P6pY�v�cs�h�B\����'����]!�������Rv�(;��i'������?lV�}5�T-ڮ�� ����&N�:�r%�x ��BU"5z�;+\n�ĝ���v_�y}���e��]��K�p���"�?E�	�Q��~+�
D�r!:��˲̙���.��/�:�a�10��*�����[�詝��Jx��>Hdm<�0���Gaٚ![# VW��ܺ)��?:�o�b��,lL���$�v�XlxVHYEB     400     170���ŉ.��B{5���C��=���s����i�*4�	�O��tT�hp��
���G���M){�F���)�_�"�d�Rcc:����E�ȗ���ʬ���SV=Y�� ���*50\v��0��!��z��(٭��*]��5���`������hU~�W���i�s8.��ў�e�N�i�A4��v��ޥ�[�eᵛ��'e�֏l�pkc_�L2+g��ݷ�������A�`/Q�od�0o��O��v/�i���0�Ⳟ�n���>qJcW(�t��҅X$���k~.z�1��e���Y�/?vaH:N��Be�ݣ�
���������"�#UgY�I�����|�d!��T�T�XlxVHYEB     400     130�cǈ��E�Z�0�Ș<(���ĕS��g����	����Z복~΄Ա���E	=[o����W<; ���/y�<�|�����o�����Z	Ľ�W��Z��y���#jl??�dUR*+ȪT��vsӑ��葉��H��$(f�����fI��y	ѧ�%��Тk5;-�� � �385�V�}���z�܏}�ed���M�v�Kf�^u���TP6�E���g�+6����9"���ϔo%�z}�|kwq�z����V�<�:��5��s���x��JXZT��tG L�ݯ+	~����'#��XlxVHYEB     400      d0ɟi�9�Q�}�@o�U�d!Yz��X�b��j� ���w���iiRz��P` Z�Rm��R��G/�Y�D�cԝCC�kƤ��U簼l�Ym٫���AW{�ӟ�m ��؃tr�>v��_=.��)�ʗN
���C^1��M�nܲ�d*d�#��>�S�A�����f�n4��[��� �VF}��cz��f{$V���v�b��J�G'��XlxVHYEB     400     130e�'1��d?��o�T��Q��U��RlĬ�b���:#� ��S�C�r�2 �6�;QH�d�.��i�fN��3�F�DK��Վq�g�-�
�T�V.�`uo[ň�/8C4�FS�>Ag��	�<��{�tYH���g��6Jv^.�&Ԑ�6l��6ށ��i�&6���l�c):���f�? wzw�n�9����!1I	�|�.�����.���)�Ua>��E7Ǽ��D�-�o�1!�9f����za��$�������-L����X$t��[��(�+#Br��*��Q1*�gE���AXlxVHYEB     400      e0d���K����4��]�,ՂvY~i(S���V����o�)�桒��T7W���In�4o���-��߅B	�x"��B�r���*��	�|�͹��,i��[����Uě�>��zV@&���A�۴�-�N���K�N��xaM�s��F�Ʉ<5���*r�Z�Û֯�_�t��W����������}�r�(��N(�Wt'"^�F24_�L�T�Y����XlxVHYEB     400     140��g�X�J�l�T�c��ŕ���N��t�'`ݓ��X[��j�j�d@�"�#3~�ϯ�<g(�� m{D�)�Z`�����Is�+��V��I��������"�Dt���x@�@BM�����&�^Ԍ�!��qW��d�T��_�taֿ�O&s�T_;������&�!{Sv�1�?�B� �f�	R��Z3�̑��s�oU��~�}��X<��O�)45��8���ac�CDNi'4vEź;R�%łǪtF�}:p���I���ç��?W�<)- %�+?���^������c+PͶ7��8��⫤K4j�������=��DR�XlxVHYEB     400     180����{$XD�(`�0x{�,��Jȇ�M��Ir�����R(�T��Y
+�oh�b6^�������69�Z3hG�5����)�M�az�R��g��e���D��d���_;U���$e�\�81C�_�4O_r�w�hT/�c����N���U�&��?CF<�(�8��Z5A{�B����#��RIЁI���my�mCqԢ��۟	�d�9�����X��T��M]ש��bI�
��I�u�j��2�LC(��`�kfK���R����Sj*���7�����p�� �n�%���$g\*܏ϻ�ю���c���I�%�|�l^t�yn��r��� ��S�d^�{�Rf���*����(�?�W�l�G��:RXlxVHYEB     400     150[��۳¬Ɍ.��uR������]����_IH�9s�3�����L�Y�$�}Â���E�/p�-�wڟ�Ӻ#�z~� ��@	S)L��O�e
�����'0��1t��~'���X�Ċ�-�r�K.��4���Z���-�x��\����^��y�jy�Y��=�md����2+a��w��n=�է�'v�veы�&�,lI=�$,�c�ꨖy�>��n�ﾒ�4)ܧ&�T@��!��D�
���e�kHʡ����y^�%��x�{���}�I8���e��,*�������/�މie4�-Z�<f��Y�TFk^�������;'XlxVHYEB     400     160g� ��j��w.Ԃ�������׵�����H�Ǯp��1����]�Y����Ij�i0	��Eb�����}���9��W���`5�` ��zȳDJ�Q!�D$3埂�rq�H�[��ww��b��"B�� �Sc�FP��{�͔gRp�-��sN�=��C6����|����2='ꡳ4NSV$�P�C�i���M1�"�n�����懹]ա{��h��g�\)Jy?"��U!�b��~��=+Y�� ��M����B���)�B�mqh��� WE��؝Oo3�1d�����F�^`T�j$���;}.��n�r�_���N:t{�B�8�[f�њ~d��TF2LK�XlxVHYEB     400     130��W�&{E�>�,�|����D�̟~r* �Au�M�bGH��\�u�X���1
�=%��O�XF��~�D��V�x�������B��,�gr�K\�X?c����]�|���pV�Ymd}�>�ɮ���l�@�s��f_�2�N��Y,<&�����7�R�\��^��ڣ���	���l�^5�����{��B@_�i��ϪK�(yVhӢ U|����<�4��^����.@O�}1�i�(�%z-|}􆍖1��\��W����p�6��k(����C&2(|W�S�VƐV�'�e�R�w�SDXlxVHYEB     400     140b76{�r���3�.��F.m.�>g^��u��:� x�n�S4��Ո4v�^��2�y�D/�K�(��5�8�~�;��B�*)���#.&_/.h5EJ������O�H4Ax�@[��O�YĹT���
me��=�c}+�z
qMJ�(P���d����dE_k��c�5�uJ�~H�V"�@8�QRvwq��V�jeG�c&T!�΀9=�mJ�&�֋���^U���f�Bǐ��!�]c��#X�J��;��'��^	��_t��"'�n�L[D���y"I�Z�J9�$�@%.�s!�k�$w��,>���	Hݣu��CY�XlxVHYEB     400     1a055S|(��`�iY�'+��9D.�d1�H�Pc�������/3�Z<:_���;@J���(�~o��Z`�� Jjiŭy)P��0պ���r��4���qN߈I�����1�+�E�/�0�9�`$(��Д���c�p��_Qw����y^��xp�g(��N����4���/��
K[eOt��A`KΩ���dD�I�\�����\5�`�(d�_��(ƣ�8XcL�ñ�K��J�4�U+]8�}�Ac��Ǖ���x���rH�������Ș�hw��.��9^��)��~�u��~��ҜAc������Ӥ��go�@;%����2� B�75�!����4�^4�8Cjm�2�P��	T"���95)�Nz�n�a���?r���u�|ӟ.�z��6�}Wv���Z�wXlxVHYEB     400     120�Mt��e�ϗ�B.�HU�V$լ����uX�P?�o~f�q�K��-��D��c��T�E�P��LFozg��tO��.H;n�K�׈����X��Q�4au���@6�+˱pB��A�Y�Gy'��e�Q8��Q��[�ŏ��A3���z5˝z�:�ޤ�~��/3��й�g���u k����p0�֪c�U2��ѻ��:��'�Z/��6��
�.�cl�#�+�>�Xā�AԪ����r��ZR���p�}.t��[n߳2#O��c��zU&J�`�B�|�\���XlxVHYEB     400     180'ʤ}G�.�ae�L'$��T��{�%yU��a���$r�ɜ��ue�%�T�h�'���2��=���مI�����+6K����6�L-I���HEg�\Zض�4O~3kr��֪e��R��[vx���)T����}T&�r�y}�H:�5ܹ�-D�s�$��t�Y��-x�fs���ܯMVED6f�|>F�+Ĵ�h��͘8�Հ�~�;��AZ��M�ܭ*�Q�B��r��r���04|�w��hH��o3f����8�}L423���9>���2{�X�Ǫhբ���p���:7V��-m�	��%�@u��"���Y��#QӑEm߷I���8��[��WQ�+���&�!���pZ)�_kn1_%���u���X�@�g���XlxVHYEB     400     160X$�s*�<��/�����[$��4���}'��g��?�+��������e�{GC*�dä����֠g�t曉b�sy"�����R��0m2����h����ߦ�"R��g&�٧�)�`�Q�yI�!`c��)C�BO���OU��d�+�eo @�5��k��R:yA!���r!a�"�W<	��Ԛh�-���g�C��\�4�v+p�Vc�nT��"�gO⓳��|���\�C�f_�N[��$�61�'/�-�F�l��9½�d��hΔ��T��c�R�tARc��[It>B���R��h����7�ɲCKK/�ެۥȃ�c� �
���ःr��/[�ɺ9�J�XlxVHYEB     400     1b0)+��Ku~Mv����9ܰ
,��z��4f�~������x�~T�t�GBݺ�E�QF������L?�#�g����p�V}�J4
T�����o���K�4��(�H=���A�T�]�;&8�m,sPٟt%����F��S�M~_ȩ8�4(���Oz{l�GPyXO�����~�+� ��6&&Bf�dP@�E����{���� Ⱈ#�n���#�U�B7�j��!�4Ƿ*�"���3�-c*s�A�.���Ȏs�~����N�/���Q�8G�z�#sۼ]�/�����fQY����� ���A8�+�}���*�i��Tvں�~&�RVp�/�Ó��b��f}�=`�|y���!�"��x�
rRE�39�]�oýV��%T� ��<���J-������y�@\º��G�U��XlxVHYEB     400     160|��x�e��IU�U�f�i����U�N�d�sŧ��sf	Y��ό���% �e�+3�䨜j������ ʿ��j�ѕ�Ow��$�L[�B�Z�vJY	å�۵�Y�wl�9�����sj��ve$1C�s�<���m���mz���K�����]��z?=s�[�D�J�6��L0*? zp��:'��R�cG�_~�����"�S���N�T���AF��(��WR�*- ��:w�.Α��l�hV��-������Xo�%t��ֶ�!@uS�Q��8a�!���#rG-��d5���4�\��u$����z�|���$�@Rͫ����ӗiFY��y��XlxVHYEB     400     130Xq��ןS����>�R�-E�.>i�4{�k�͏'�%�y��!��юzP�R� �xUl��1b�K�HҨ^R�[�o��'�]Soy���-��%g>A[W�E�D-3
�%�i�sp�i��2�� "�p������!n�	J
Xұ�RunDK��i�����9��A������>LX0�P\Se�u'��'��XTV0ܲ|��� ���Ջ^@H�,H#/��L�$B���!�p/z�@��W6���:l�!�������<���0.7>�}՗C�9)� k�=�A�O���=ڒ ��"�EKV�XlxVHYEB     400     14020��̞W�_�'����}a/�'��El:����a��!�j��Vʘ�{�w��BB����q#2�?���
�'ݦ��<�>�J�������79_<�B@{=~�	=}Z�j���C2�y��1�[�tL��'��ɬP(���xP�X���tpִ�y4 ~~���wD�<co�Sg�����?ܑDhh/c�3Ӝ렟  QS�JO��H���*}<6�l,U�u�o�`o.%5�T$nLv��LB�9cd�Q)\t�&`�`��a)=�y�<�$�1�6*� ���������R)���{)V�XlxVHYEB     400     130��{�g\��8�a:ށ(S'�܇�ψ٧����Ha:���@�8�d�ܻ�n���;��X�;1�A��|˳?N�CFĝ	_WD`�HYO�x�X���0%b&3��y�1��l:�g�JL��F��4��\|�xNP�~�u��M�����J"<&��s����K,�WR��"�Y�!?+���/���(:����J�MJH2�Ə���	4�t��`*s�hX۰l�sMR�.�<�v|�9qDmW� BR~504ҶWN:u�/�y��C�D�r�r폦+��m>������������XlxVHYEB     400     140��g��Tr�Ǟ���������S>
��I�&�p��V��',1x0��'i���Eݥ��Tͥ�%��čp)DeX:}�^;���G�����@��uZ�L�a��z]��уRV�M�E�/�w�b��o��.�Ă�ge�r�Ij��Q���	��0�Ay�*X�׹Xm��,���-y�O�'U7�;��LM&;���B>���aK",`M�(��N+�s��V�/m`:Ƈۋ9(Τk���1�q�b=��K����T�L�m\:�� Ӵ�k[Y>�|dw�x-�9�dɼV���l��_����qC�ϝX���`����&XlxVHYEB     400      d0����-~v�}3�-霿׼��y�Ζ*R-U���>[�Ŕk����6l8ea��k��Q�����Ŏ3{h&��-�7���)$��UR�"��# �Gv�d���,��rDԌ�L[vMC s3z�=��rX����KX������4w<V�B�9�����"��{z'!��T㗀ճT��x����3���C�_.w��D'.�� r��u�B!p~XlxVHYEB     247      b0u�Ǉ��^Y�	5�]��N�0Z��p��X�Mx���#�(ေ�yb�M�r�"�Z��yAs�º���n�)�Ǩ�G��u�j�6�G��c��f��&Y9���Hl�,遥p�T��%#��*_ĽCx?���B�K.HPE�F��&Q3�0��ч���1�}����t^1iS?�mr�Y�k