XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W����X���+&�����cx�� ��,����F�U�	��7@rF�m�i`W�Q��V�/(���`���[��������i���%]eS �2Vh���a���!�F\��yA6�k�lh��ll�����
}��z����D�����)��b㔍���B���3�v�%�N2��h������7l�l����efP��]`N��t��=D����<S*�]r����I��r�3�P�Z�ٵb �����f���s1W��Qq�nd�ez�/���̯�_]q�8|	�!V
�%\Xl�v�a��f��r[1f��#�Z{�c��?j`-�\$6�o̃�i?��ɕ���Nϖ�r����:4�-Î���((�mV^zۥ��:�=1���p��|�P2�ύq+�t�L>�#�-�0:��T'��餳5#7V��K�{�3�'�]��@�+h<��NV<!��6�>����ZoT� p~7_�	Q��`�H��7qi�YzU�Н�����2��b����9ڔቧ�{�@zq�����m�6aW5�X���L��"@NȐM�x�V�L��d�/hOx6͐M������O�|�B����kӷ�P a��;�'�A?�n���r+�\0E?�#g`��$��u�@��E���}I�u�-o@�c�^i���� �(�uʣs��D�E���I�l��N���+#��x*�H����!�����W!�BQ5ka��0-��+R�T��m�3<�뙽`30�a��XlxVHYEB     400     190̄���lY��"YJ���3��bRQ�֝;��k��	H\"��7�ݧ��S&�p��@�s#���b�o�5TBB���9"{U����-�N��X]�(	��<\����=�b��1�>b�T��R;ILƞ�D]<S�@"����~N>.~�yغ��;�$6Y�T������;�Ц���{���F����#���	���R����L��adjJ����G�5�tO5n�osCs�b��t'ܞC}��4����&�a�J��~7������D�v]�;���P'�Bq4��߆$;\Oۧዤ!ޙe���Z�ʨ��܊�2*�ehL�~����9na)�|.��$�,p�Fd�m�vՙ�����b�(�ɞ<U�I9 �r��i�nn��\��C4��I�fXlxVHYEB     400     140�!i�:y[2f�*֪/��<��[���j툃�!�"��fbä�� ���BBK�٧�,U>�z!uK9.��L�
�J����xØ0c��,��Xj4e�! �`w
����<�B�ݫ���ā�vr�b�P��ɉ9�.ޚ���mB�_�%q�yu��!�v��Y)ꏣh��OJ�0��\w%^t�3ڌ���CK2��>����)s��L�Lh_X��<ڀ� :�]	�M�g{]�K��;���dp��]��p��M��x�Pϴ`���y�[�H�=\�ۦt���_���c���n �UL����Ers�XlxVHYEB     400     170������Zx�O,Y�Tv�Y�n�D���}��g��l����N�C(�Yh+f�b�Z4MQ;�|iH�a�
Y3U�Bt\7acʭ���c�*�>�j�.���[��-؎_R�E�vIl�%iGOIt��1�rZ ��������&��mM�C����Ӳ���ǌ�*�H�!���P�>x�ql����鐶��6}����4�}�NYP�7��tG�=�|oT�,�A�|O�`�j���n�w�eBm�LF�BF��������9 Xc�����-���ґ�2��6��ug�cG��N|`��m��	�`�!a�>l$�>��S�j�*G���/��:q<���f���EӾ��7N@��sXlxVHYEB     400     130�H�n��������\}��,�q$�~�F�zV�8��Ea'��c뺮gvYv���{<�!nt;�3^�:cʾ	@MeV�U��ؘ������	�>P��� =�c3�ګ�Ι�Qn*z1+��w��7� ̀b�i��ĞW}�w��V`~�k�w������&��ؿ�m�?��?y*�mK�ϐ�=-JY?^LA�q���1���������o(�{��'��(%���p@���aSK�Y6��n�`-	�m=3����N��9T�
��6n7{*�@`�Gfl��
��4p��U@A����L��-��!XlxVHYEB     400      d0k�4� �Z�j��mEn�X'�����%�H�#ف���Qk�v@�K9����vK�Hr�(�
�<\']���h���/^��^��%w�/�>�	��^��c!a��ʁe-iU��0��v���SHŋ'��x��8-�X�5F��呆Id5Ȭ��*���Ѽ��,����-YQh|}��85{wƞ�1����3�O�*����L[�G5~5�wXlxVHYEB     400     130%�B�~n��9��]����7*�6`Fx����Ǌ�$�g���=���-�n^Ҡ��3Д!w�f��z<H�pt���g]�1� �	�2U����
l�?���u�։)H�R�AQ���q�^�	�zg��G����$8Ʒ�7y-���Ԧ�Ԏ(��;t����\�yI�x�V�D�qj-B|���:�T������ZS��ڂ��h���4TO%E�+�B!n,����_��=Rփv��m��N�[h�=�g(
�#승���1��A�����:>�^���w�m�u�b}���r^a8* s<�XlxVHYEB     400      e0<�!��aJ����Ձ��2��Q�T�3~۲kH�T�t]���:�Hk�ְxa����f��sm<�{<C�C���L�����(|��~��%)dc-r�'�%�K?�o$A<�P�(�[{om{�{�����ӿ�U��y����y�'W�8�H ������������3���Œ��A��uՄ�O��#VM�MJ�=vJ�-� �C�J�u]��XlxVHYEB     400     140�U��6���s�>oѪaV>��պB�)�+h[W�6kO�{vC
ǭ|�f�k/�N�!���[����ȡ'�KL�UA� �?�`=#��-V���,�WզL��4��q����`������	�X�Ѹ7��L	6��U�-*�`���1U���0��X����7��2�u4���P��<d���)�9kUv0��H�M�>��V"���;<����TIf����jԠ�=б	����>�=�=� T�zI@��yB���p�.#��cT��y�ζ�r�C	�<6�Ma�]T�kF����XlxVHYEB     400     180�8� )ө礮�p�Ci��9ӌݒO�Wau4�x9p������*����8�����|ܮ�P���CoV�������E$�R�,�����řqA�C�K?����5q����� 餯�\�Xg{$@4�{��8�7/��S��,zS+�s���Yi�o��g��@�����-�m�i�09[�S� Nt�jy����x=7��xNLNZ"���CS�B���^o\ˀ�*뒒u{:�E<�<,1/�^�n<R]E6�:wO8Ҝ'�YAD��	��"�̮��կw�5!��)���;�&��-Y��O���kE@�� R��x��L�uG��1����$����X����Ey�X�Ϥ�z�}.�l�UH�wj�+XlxVHYEB     400     150ax�K�(��.�MeK��c��!���� �ᗍ0"��I"ల/L�9�����K�<<_;�8��P�{3/�`X�qo[S:����º��3$�;|���=�#>���;����}2��@4f<�u�Q_��4�x{A*DiX�'�?���U7UQz2.�i��85��R���>� ���D��	��	cE�]|^f����+�
:^�Ə�N��e>��,���#+l�'$���i��8�h��nU�2�H�U��̮��96���C*J��9l����^E��\\�(�/�2]�2�n�9P��6�k��>w?wp3�5D�ۂ�7���Ėh�$F23
&XlxVHYEB     400     160>�^B�1��O\��
p㜚{=A퀮�#ש�JRJoG�<Uݜ� 3��Txf���%#�qo_�D+k���>��g�~�m��#ؽU�h�N���1`��Wv@��2���	<�Z�@e�P!Ԣx����q�G�+������@�ԋ����\T=}Vr�������	����~�GpD7��q��}O3-.:�RKWj0��.W��ѥ�-��_?�n�;����2���V��=e=����逦�qJr��T+�_�����t`�+�t�:��d���ə_���+�����wu}8�n�M���.XJV��@��c��s��B��z��J�T�r>�)�YXlxVHYEB     400     130���0@������v5-�&T�ܩ3��fb��(|j[���cG�[��}&P�۞80 ���3�-rv�q�;;\����ѧ�D]0���8�Ų-�z�OFy�g[���4>:�U����;�&�Ԟ�rЧ��V?�O)�C2w�]n�V96��K�p94�x[�Vٕ�7��[��$h����Y���Q ?^�����kpj{�) 
��v��]�ִ�e`�
;PX��fEtk�A{��~����f0��v`8��Rv�Y<�A,и�l�	!���7�f^Fmi�dV��H�y"9K���XlxVHYEB     400     140<�؟��-����'�C|�Fʣ�	>�wF��3(�ܜ����N�*y�U����hrس�x䩶;���6��u7��t���ṋԦ׽Te�����.��bU�j��CY>N� �6�7
�k�%Yٶ5z�����- �����K/�P��P_����Y+&���V�[��&X�&/�uyh���ɧ�=�Hw4��l��'3�E�)�����3�i�(��q�@�1�2Z3�X����<5(wL'$��t�.Ԅ�v��L����Q�8�,�������u?�Q�՟���=e�ׁ�1��5��C��) ��������n�	�XlxVHYEB     400     1a0��d��[���F�F��r�D���qJ�/�	�Hy�W(v�lmi����f���}\��.|
,����M�"kZ�]��&[��D'D��T`f0���3M�^�K[A3�b�Ǆ��.;& �B!Qvgϩ�ՐÃ7*8�j�9�<��uΓMUyw�j���(�\Y]�^w�9�C˷����$a81��)��=�F�ſO1� "W0�H�#JSW�c�e�c��4����c��|��zWc�S�+�i޵c��t���t9����?��,�5a9�pm��p�S�]9ωpst T�yd|J��U�m4UHm%W�wE�%M���G��`�~f,�yk\�9֓VG��o�������'U�%2�
��0�%�Ȝ�oz,:g?f���7�[6�x�@yT��"��¤!'��QT��c��݂�2LH�\�EXlxVHYEB     400     120��p��=�M��+k��7!�lB�cJ�M�A+�%�����4*�oI�Lʍ=��_�H���&Z�������|6�@'���[��؀�'}i��e[|�/W!F�?Ы)�"�����*q�;w +���#����S�<�!�M��=�����W��U��sU��:�E=��Y�67��4Q�)A��X����4~�qjI)}Sh�"mU1-��Fl?WqRqu.YC�+`Ԯܩ�P&4�L,Ed�B_�/b[I�i�Q�X�ι�ZZ����%��+6&�c�R��3n�5��5yRx?XlxVHYEB     400     180K9�|,��߮l�����?��4��k�z����:�����i�Yb���0\`X<I�ZM̢!#��]�m�@�5D�7����'��܀��G'FH�e]��� 2w�2)�]b�����x��j�s���C�M�SLm�<�{��l���d�����>hf[�)h�iZxS��]-<�����6��|
�?��ѳkkΰ�Av�w�ᓴ4���,Ͻ�
}�)��P��6�|�j���N��"}�>bL)S+�}Q��{�oW�� �.��"��SУ
�)�et�ܽb�j���>^۸W&�a��ȓ���]p \��ޚ�Ɬ�ހ��{�܀QD�)�D�H=���7o'ë�rn��� �la� d�N5�Y�Nc��q/n�XlxVHYEB     400     160�{�[S���DĹ^�x6�z<��{��=�l�Ʀ(�i���h��U�/��L=���XW��E��|.qz��� ����<�A�F���Zф����4]�s�0�����3��:_\�s�#X���v�b`��͢�1C\��#�o���4�e��u�b��,#����xc��Ȓ�	Z��M�Qp_�Ht.5�������wjeh(?s+-Ax�
B��Oȅ��ъa��,�?��u��g\�cW��G�L08�):& �HK���ެ����ju����ߑ��η��RV�b�6q�	g�RL��y�f~�J�( ץb�X"WZc�4�&��叞t>�EU�S��v~,%�0{�:Ձ��XlxVHYEB     400     1b0Fa�w�h�|��v��A�G;;nj�))�W��w���Q����qS�$ז���7MeU�4���*��2z�/C|"Ͷ��t����r]6�4{f�j�ZUNDr?1���yz�l���`�h�f:��Rn��:蓐K��C��n�k���h��^��^
�4Q9��y�Q�˃�5��X��4��S#tKq�W�4`��B�����UJ9��G��8��}wcoXqj�Z߈�c�
(}�.��AApn���	����sN{��v�h��ʏJ<z��k�˄`|"h�5�M��l�dΤ�l�|?V�,�2��ֿ)!Q��}����=����oc�]�c�+/R@�drKa��(�tV�� �f ��9�LZ�M��%�ؘ�tw�x|"���W?E`@��C)��k�>��r�p6�'e����;S�"м�zU�I�2XlxVHYEB     400     160޾����7j\o� Q�%�V�9��Cq��<�w�3�.��`�C��zv�t������t�'��h 4�n߼���6C�H�;ޏ��Iq������h�4r�����7=��Cj�z�G.Iu�I�p��R�U?�A2�P��h�k��]G4����hu��d�DU���!`{#�1�P�^��d��bq��ms2#`t��y���Qz�1t �LL�D��̞,ԼC�Ӣ.H|�*t��<��K�Vfj��B��4�AM�T�C��$�j�V�!eK/�����{��ޅ�u���iA��9�|7ͻ��h������͸�����;��/��Є�XlxVHYEB     400     130D����^�_�S}����9q`�\��p��i6�$Q���|�9���/a�8�Mѷ�=���=�ь��J��Cyr/2��`�)Wv����޽C����BY��o}��� �sDMM�l�I�U� H��0��e�-ӄ�>z��7�z�NT�p2ס�d�i�J������o���>�PL�I��,�˝�����J���Uj��rш�� )�0���L�>�}��G�^l�x2(t��!b`�Ԝ6��{h��#zK��@�&��2D��}L��*>bc8!�+�g���%R��XlxVHYEB     400     140�w\6�AI��p�����Ȑ�������,����}. �l_�YN˥��$Ǫ1� �0%:�?�x�T���D��p͘JJA{���}`� �t���'7Qo���`K	�[�3'���r�/�2σa6/)�#�f��=�p�߆�O.���C�����F�a���Ӣ.Q\��oqb5���Mxse�8*�O�ޱ��yI\��˽�b��V) \`��``8���bM��`�����Ū+���'I<�C�]��!8��H"$�kh.�	���<2���̾_W�SnϿ;���eF��3�A�W�i�_�ö��gVXlxVHYEB     400     130\:�����"5�������C���ǽqE���p s���2�|Y�pW�0r�l&�U?lb%�z�YY���kE���Nl���is��.RzN3Th�;��`��E�{�;�����v�P�2F�o���e �b4�p�����@`"Ŷ�%�ڎ�R%w�N��S횑ȷ'?5{��`:�v'a��#n��s���C��u�/wBx�b��m,��׼L���0�� �)H f��UƊ�_�zA�׶��eѹ�EDh$��/ռ��O�`�_O��,�+������X��8B��K��pM~��XlxVHYEB     400     140�ˈ��7��SUoF0�I}�d��l��Q-���_���Y�O�,�3�� ��78�d��$Uϙ�P�Lf��a���gV29�<׬.	�P<�u��~�F�s9��&�>�fw=(�O�wN}M�iWX�-e�~��.����Л�}�����M[.�C��C�{���09�����:�C�N��Gn!���F�SWb�d�g�3Cz[X��')��ٝLUJ�Z: +{�e��F��p���Y�{1mej@�d�������3P�{�l�|h��O�VyHbuȗ��%P1�]F��4f���V���Ok�\�H�r��a�����XlxVHYEB     400      d0y{���I�؈&���r z�h�k�����0�A��V�
�^�my�Q�h[�#a��3��j?�4�2��q�)�kͨR�F�H��������7�]�j�Ir�eE�\RT�e�,�WA.�Ck�0�ĦW��K$�[x4*k�����Sb������
�#�ҍ,gUw����)�8�� ��C�VV�BT5!`���,�n@%�Kn��XlxVHYEB     247      b0�)UeڠA_I��o +/�t� �"�+�Dq܊��V8L)�s��_�J6G�4�I>�a*���ǯu�0{���h��Z��#7�ʲ�
.�!�Ac��:��枏�P^�"�Wo�}�|�;�:D@��eBn�YσCi�M�#7������� �#;�%�Q��\(܁U���q�o�