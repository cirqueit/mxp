`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
SJ3ZZLhl8ee8Q6ZdhBGYEOzLuI7gYh/BTZMK8gQmjSOrFXyPxL8iJTIgXF1wkByF/SOedUbM4lET
3zcG39b9L7KVfpdoGFpMMlBWE6R0vVKe//fyxGiVj29bWgrpWT/pPK6lhTzgQ1MyPruQWr2AJ24+
qRld6NYmrnUyTMb0i3YSuCMsXtvfqn6Rx54jJfSV4jNlycZZZOJuqFwGWuM7iPba7FYVG18OGA4j
dkvpoZUaJGyH2hdVgdl7dUwhLzz8OJ2q7BVYd9IxMvxKqo0/sEk7940IOew51yoAFPbF0rvj63DK
8Ae6rMM+IwXQq2t2/O4nWmGeXcFcrS2sb+lVEYy6SsC/g4AxNnaXFaX4a10iTRWl2S07YxRS4G7Y
IwSmI5StNpC8du0feFTbJwUfvmULs5742p913YvGjuNnhx62ttLObCvTurR+l56v8fLQxqvmmnrt
79EchjF1PR73WxHlQ3YsKCPWoV/XYm00csm/+BxTEQdGj5EABg6pn7byc/cy/sP0vKbwscfcYgQC
wHUKzPTf0sXZ6Vvu+U9d6dwrPb/wKP1gHb7yFNE0xqPMjMkb/9DdILv9+bmT14W08mhPts6JLOoO
5XFID4Ueyx+vylDiX7gbuqqcBwMnrOc53XFAR4ZEJbigaJpj4ILduTxy7GERwNk1QYoIwNQ586Fi
iKrkzsElSnvwvynlWxS1Gv9bGama+J2pGMCI4STvLrqdDRLRZclIO7HKyg48w13KJPpUVOQqWeDE
MbrcELtszSabifq+fFs8R3OfY/N0VhhedltEoDJtCGf7ah7QfkYLUt0oF67obBtgMTqikxc3Nbmx
5IEteKwW1yfyu6IowdmzB3SgscMZGsRoyb65i6KKcggR3q7nZaKuvT4NeLMatFycrj92GKRZc7CL
C5yDOf2xWDz1II2KH9cbQPhHytkP8xsyPRjUsCh/9a4fEkF3QW6UQyw/i4doPmUgEnpuSbrMUCaC
nRIV8CdoYQXssSw7VWrkwov30tNjvdAqXK/DLqVts8zXTDHFaXDdkCbLgQH+MzPWDnQIOHg+Kd5e
lmqkb0zVkOPoNn9AGR3dXnfIst+d9kASgue6Ae2kbd0LL4/IhfXkNTKGPfW3w7a0SP3/OWokn2jd
KP6PH9/wznvKvXGz/kVi1gsxz5uXo0wbBaEWYPW1eXnewKZqPod6tivPeSwifzul4xsPEOiQJlTT
UIOoNj61V4HJL12VgvaJ5u7dYzOuq1Q1gg9Bkpy5TEsBpXyp4TNzdh5zUAuknPwJoR7pDqEEY250
eiLX3Bx/oMdxcsxAkiIbrn04QNZzZMue+VhOcMlYgMPJaw+vsYMssRS/XRgU1c1xfuOcEOQDXqP8
YmPmlWkysbmzUDqfpqa9Fgg0pywAekH8Qyh2/IbetAWwzt4ktWcY3EzMOnoZoSiGY0atQypNq04/
K2S3oGEUopGmlSoOngckHGM6I6p5kmoG6y2NyZgz1oO1lnxNi3lpO/MpHCnbZFG2XEGS6J1+Gdmu
n1yF8UyRt9+rOqISlYYwpSan6aEnafPzWdG12Gy57H9ck0/XNfbm6KtxlTw6zZdyPQb6M5SoJaoL
23U0mEWrUwbtQlyFOLsQ3I5BOoFB5ovP0HBn9RGuwl23XWQh4SlRksIp6yZ07xDn+8sVjX5f8ENx
nUJTHudSgoHzSghBLcpKxClYsM5652C2NpE7J8wVIjo6ofqKAqFRYBbomOF9Pg1Fbahis6vj88pM
wfrgnuGg+7mTUk3XgfUUlmMmPAoPMt2AmUScq/qvj8YzyTXu7xQ0tvZXlw/5uHDhKcYfdZD+a87w
sQ0lkrvStnohfAAwZ1PglReg2sMwRtHAVXN9y5LO+uo3umA9x7wQoeE2wl2EnRvGzEwhOL2TFabz
/aZdQfmisGvcatjD9zyyikgVaiQhunYU7Nt0EXJwU9zVafhh8xEuZEiTqyyRyLchLYts4wqEb8YE
ZKhuMl6KEWbp5cb0n64BCKhW8Z8x66SVqfIi7kPpze7yC78uaRgJDcEHrwTUo9McdjK6Pv8uL1IX
a+e62FeasoiabWPK/P+pR1IF5+H0tGP4Tb0AEhPebS8nPkAhbtAO9fqHJH9aH1xmEih6hwun8QKi
9km0C4j4o0klS+3hVI/LJAwMCFOcYuzBgVsGFngg9MU0/C0+AjkdQItzZvpqLHj/muxA2yJOSqnS
2cBb7pzlsi5YgpB2VB7V4KCmJ7UwYCqOp3t27ArN+OE3NlPMpLJcNDkxDxqtDEWG+GDTdRSLckSs
76jg58nLOETpQwyLTuF0ea9sSCVonhoAhsMASXWTiMwEX42iNI+7lo3ADM4/5LqJ8cXCnscnruiM
6iZOKB/TcuGlw8u4V/bfQafP2rY3WrxHFUdQdf8JVq/dzfjfD1AQSQvFmKTo3cUT6NeqXLw76jeu
U0OEID6CTtIB99SxX1ieSPspwHzwGGaAHKo65dogi5vMuTnnuIFUOeLgtwZBmPlz4dmD5BEYw8X/
LTLB92UGnh29K193NUGFXnWawxkUAE03AKmiNHtJLvJ19/t4QwPo6MwqyF7nA3lY/DzUYJtuYgWG
UxfIljrcfoO9R/I4GmG1o2FSPkdCTVHtiALI7dR0e8z9bgLFZTVDhsai7EKx4cx5qgfiDh1bEtz2
X+wx5Rm8EHcNYiw6Gu7xIZJoCYMipa++173fMDDgzNjf8GUljC5tf7/ujbaSLVlPlBK35VvGXNER
npsUAPs+0vklNz7lQvEMY82Bscd4OzBLXGI41W3TPQofxcELlKDWWMJDwDEhwGHihjwiHf7bHOzo
Odli4KQZ/qBIaTYMVnYc34kl1kjbOXOKlb60Le31lQ+bTVCnqOshXMTUUvzBYcc7vA8nswfZ5urN
300vJlG6J+vU/a1A+FW8VCecDair1GtTFp9WXx7ofeuoYdqzhzqy3XMTD/OQVtWtZhbbYttQUbO3
L8Jsp+eATy0iX/SHUZM+mzahg32Kkd2qb98GWW/i8dqUn+pIfPLSyGTcXVpSB475rQcmqpba81ga
9AjAkeNWn8dG0B1J/QSyJreE0FRd29CrCCtl9GPfOJTaWBo8L9Sp0RoP5EgR+1xziKS23VfKolBJ
LN9Wf3e8YiVDMpKrxQ4wnRcSAoy2YjM0kS1w+KPsm9RFhH2d1EQOXlx92ZbOTKGl/7qVDJtNMXeB
Kn+iR+8S/D0w62vc6UxtVEbNX3qjK5camCnRPC4sNjGQvTlA4qQTnd22lbsrfIgOKRVBg1LcMQHJ
5c3f5LFuxgEXhAlhHjX5aOwvCIETgwnV/5aKpNQyITknWOl8wSj3K602GWsD7IDwKEAJuldbdFRr
dm7CjazQ6pLSUXt0K7mW7SnCi3Aqbbck7rKCGusaXfoaFcUoaJ3Iu7rCnvTsH/1ADFIeruGAnGvi
Vo0UhutnDajCe1mayc3Y75RdpoUfZ3EqTtWqmwzElybVCXQ11Epv6ZYB12GoZEpbGZL/nb5Quusp
LC+TqP1A4h/cBOVpmchVeBjmaAmJ7aa3u3fo97LlnFIiZjdps8mJadVGAOSkCrER/F/G1buUIwWT
t9grdk4Np/9AEbGzCCSNp3+tuFzasdHqZljBXn0umP2UFU2aAf8WvkLehxa6S8FwyUtiX9jcSPSV
ciD1ItvUrUaPSGKaj+FKpbBuywPspulCsLLEK+yXXkT1x/28upRv7q3LgGEH4MucaECEksQsA0mO
R2+UFDyR46icCsyddfphR+YRv9uq+I4NUqVXKy3RlE11hB0xQ9ots4mOBb7q7mzXwEDzuZha01y6
pWytPxX/2xbDtQlNvxx1nznQvAUK7UZRvte+0QMd7/npQcKBlczHRhukxbtFWyjdiP9yEMU8U+fg
t4nhrSd436n8nLEJVh87EahHw5jRmf61HmKrGcS6vGcM/KPMqCT6f4KuTKnEHSvH7/oIUtQLm5qY
mFAbgP5x1CsKNxDeHvybK+aNl7JApSdNLmwqToX0GQzr/guTUkb40tUgX3EDFGUJX/RIc6VVJxl/
/vwSDYR8vTRLdlaZ5n5f4nrhTDu8wCfmaNhPl69CpMfKsd9QB9HwgXLC51Ldx8W/nR4zENpFm0jo
RgsN+osLG3Uxa6H/+pRlsFMHC3Fb2N3FbmOnuBnfGus099TgnXMLzwp0U43imFbQhnYTNyRjbmCN
Ek7NjhTNbdzJ7vQ+TDPUEeiYPnBEJcCjGjY+Tw4aaHcQDNDO2pg34Ee5td5LLV+G8J8QbIVBMM9k
qjCFs0XjqJ8OuZIgakrRglHekEDziUihLopssdrlHn9xI1dNxGjJvIdTO8On09N9dTD9nJ+X5O+w
j0h5wpT6E6OYhaKT4t4fZtO3EOfLRmoVH0gdEqEXqFZtMKJby+PQJCO8uBt5qa3TlRg5eKaVFulb
nBZ8q2hOF25VqAqFqTo/ETCySlKqD3VxvuuY8YqfW64yMgeVPROF1lI9PuU8/CWv5GiG95Sp+T+5
vzAcz3aZP8S5NXa1ZrhE/VpNE1njkD1X/tUfv1kGEOC08T4DwHOGIhAb0FFnARNwgo9SnD2qJ8St
qLWp17AWhAKSyIL2Lk3lj2fpflRNsiDUCHQKkpomU4bNh4SgZVz+HsiPfOhx6ixae5krANLJkNF8
uy7TqShhhMgY7tGXRi9yWywSsjGUWYQbpxNjAm4N7gTXBKB106JCJcyf8KI5WbzXzJN6IWSBaQ3k
RyCExWT/DShMPrQSzHUgba99EZ9HQCCZWzYsc9GhM+Zc9lLpVIlsuAz5gUIF2oBrfA3xegWAMEJL
/wQKPPMc67dSHz2ThfRlm1b4NYIEKIivegmgl7mTFV7ruJVfIGNwol4FB8W0TjxuTga5tzy8i9dW
BCViV6+k/U7v5z/2hvEYcQ==
`protect end_protected
