`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11136)
`protect data_block
qwi4uiVUI/eKGZm6VAZEOhJyycr2r4RMjpQF0cHBXRMSwSx+a8bXIwYS8g26BrHWkM2MxreMjz0I
Zqt8vTc06bjmJLM6fdW8mHFvMqJGj7ag8f65i4ixgAtCQ+NnTXF9ILdNB7AqQ5QsivrZHDITPOJx
4s3Rn/MZUZRnSUHa3hSnAQ9JVkk7ibDlYWXDgvmpMpFPwZggEVJoaI5vLIcLkHkoceGt7Cbs6lNa
pQXosLB0pwqakjAJV+uVGQy4GazTmysvenBCvOHC8QryDWikSM0UyIhOhYFXhekk1U85Lf08fVJl
6tScxjtAUQnrfXOybrMSEmUiofrVt2+DtmHaKIZHKwGh2I3/7LbEHrJK+nW/hEZb9ChRWheeIPS4
IB85u1Kf9J63J2BMJqS2daOMnus0+SyjWSemcKONsZKpQvS3aRbFejdmLcR0hkF0Fs81i717GPY1
meImXwvegpbAGyvDU6tS00OOOFXSpdyLwea9Sdcl90hiQ1LDDSQWKGlgbSHrN3YsOb1u9MxyMRpD
scJakO9LFowI3ESGyaJFFMAqWF++6TkBVzhQupi/MjSYoEoSTgtMCA+GUXTpuEHn5PQArLxiNoKX
h5njjM0wAEROtTv+R8aK2TfpoLGYdZzisEwjqxSxcsOyVLZ+XM/JH/vFsxRqaoW0jDmX+VO8TBJ+
h5tfgq9AFZEwazHf4OzPO9wFnogI4unTsClnTz2+JjDA0hqpwwYTZ5HnCVPwMBNfLAy1gMpCTGzz
pyi1x08AnMAvs1UFIUTuSKX2cU6U6LJs7Wr7tZ6R8E9h0pP9drE9jnasWVtFwAXReU/mgaVvHSuZ
bxpfRSIIfXepAVSqvylmP4LWb6CWCZ2Z3/wZydNBDD4/hE5bDMF0QccBY2qWzisKIX59FygmA2HD
3QIEDh/k6qvUXvuokplpVKFMuwceFY5jYITxVkDcm/eJ7a0x11hJ+E26lJYdGNvc+jh1szSv29uG
fI3KFDIorwPQqLkxsQ3q1HLg7jvaN5wAg7gUH0oiqnvyxqotdfW+6NMA98stj/knAAzMPhaF705l
a+R+3Dcu8f56HbTirL3nz+v/A1tZp7dSA1AkhUo0bnA5JLRLqo455TdOKK7eIy2AJFxWBmz/ajRG
twD3j8UCb4tTX0gEf1tKOJ7zt/UKXAd5ovUMxfhBAH+4qgshpE0T7PtRzQ0tW7ULn4cFGiy1Cuz8
l00Dy9MExo+IAN8oX2wiABS2F0ijx8RJ3WmPfSj8HtszMPiwYuojrGazwSDqjUt0mrvejEGN7xOl
ok3vSgZxzUdsVk+Ly8eGuqrZAlc8/JsMW4odCjsJPLKlL7Rr916JDAvOO3PNPF81xvhGXjlriDVw
4OjZztnUhCWPySe/gGvkX2TEOVnI117vcMg3R3qVi37gz6Rtl11pwrOc9jg7Igwp6fDL2aAXi4lC
d/sTwgKzGJOkD+0xC0ovitwPSL9quVZsFy0lSIPuWmPNig1JNLaQfVMZttW2+i5EzO2mldZMIX3A
8kIBGL9EY+IvP7oAomuQUJc+OO4XcahfMHPB++2a2oUaq0hdSfmz80MmWIhLOSWhSwMeWUPGLkad
zhuSjQ/BVJ6cNKnm9+lz/ZFwBKCB4esamTHLekRxhZAByyHrnNMrtW4TOAwAmH3dCbHoIHE//144
03vxTffkrXaqJEnlPJpgLM+CBGJ9v1esnUfEJfgs7ZikpFgeWLeWhzeRTtuQx4MT6Z2qPX8xpSgG
AaOZqiO8QzKfdRwToMvZe5+xTsAa8rO9MD1zI+427Dh2bKleS9ekRbUCELYOb760MNIO+Oy7tOIv
D/LPKLJ3VK/4G6eh27RyQPoPTINM52QZJU5bSv6+COkoH3aVA93RFbJ/7wCXjJWhElcJkPhxPZsc
k2eKmLuNspu6x5J8QrB534Taivq/ULFGik7hBPsFI2ZHkKJyuW/EDKMmoUAZsBpbeftsPzEkkZmM
DzEHTic7O7w07YVZsTAnkkAWroEhJWnGHlbbG9gzWTtnH6Mlegh+yVx9huuTWpYE6A/jbUYhIb1b
cnu168ILVSuJ6/Ya69oloTb6KQR3clzgpK0DDO9wY/Kg4mDCh+dWpiJ/934iirnOb4kRwIZ9K8Xx
QEa0w6Mauu/S9Y3VgcyOhz3HaGrqYbpyPi+CiiBRMGwK1tDZJn4CmYwst2PO6S32/j/MdBezVE6T
WbK1f+ZQpI/NoKSdKEyOmivg95HWmqeCYccn4aCEKJ9YUT4+FtNVLBLhluTdSBopdSHQ/DztpCzk
dL/2gphfdZJHgtG41c/AkByWQ94XBYZDszf7S/25yMIg6XekzyfPfWzerhLcXROFfsR0DFsF+6JX
Z3Wq0YmrM5TdUTEirgVB8oi80NzWmVXdG+lpvNKKDzrPFL3lmkR2nu6H7vlbBRZsDTu+F/XkM0NT
xkMeOzsvBjHKBEEpH8n4xkv/nlwUG5HchzEaity1uZMymBrW6p9sQbENKPwbkwD4Z97g1RQdlidW
FaLZeSXZNMAbJzd/ulS+2r9g3C6ybZSgxpTjQoAU29IxBuJD5BGe+aEnwLuyLQO3cz45BFlukkip
vs+/PNAnRey/0UqJXqrQFRiY73NoW4PIFnMbn50Qxg/MEeCS7oBX7ItN+OzQKGzFo+jnua1XELzK
7dMqF2eJ4LBafbFe8Wf2FwzTcUZm2iJZ7WVZWmC4xd8rHMvSHVmoyQEH9gJMQm+1w7vTQglQdNfl
0t39DbGNDNpqvqsIZzKftea/pfn8RU1lAhl4300RbpMu2fkEMKx37IN/UmJiFgCuEupYq1iA6JW2
dFAopmNIMkRC5TRKe4nfM/UoLlAWzlM2d7OchOXDTS1k4CRSK5LSoCLQr6/HTMSBGlucDZr+toQ4
OPneW59xSE9MG9Sr/3SgQum2mjWkBhtwZfQXiyOXZr5kRDUm0CoY4mEHGzQtkWF7SNw4jbxv1SlD
03Qk5EObKEoW4tlTwy9vWCWzVnpidLmxxD4muTNj1DyQu5DUdrRz3VRvAjnkOj8UKr5sLhYxlXkK
gFugP19I8Hsrkyd4P2WGANMRYEMXNULn4DRfgMz70zRqciApF+87aSTkzLOfgbO39CkUuhgSVwhB
ssDUcqiCwCN3URa5IpCr3zJOfgCFVPXUZHkicd+R/u4hKK73lIGLxzcre6bxdXZeXssYrLCfNBmW
Io5BuCjKHBU3j4iR5EwuFEi5Z3rfprh9mtiv//4NYoWMrNZrHWw4nSzAHooB7WBJi9sxG/ezkX6a
jb12qeB8QaT4NKk7gKVJpafjyexPgco6HF+ejqiSBUf6RRznDTjI0ZTuGYaNI3c7bNR4xpROelQr
+5jQduLKMRMn8iV9mcKpQER43eGSNyfvWn5JfZF93Oq0kt9QdNfPyDEgVwHl2dqMPCED2YhOtPN7
wt+3EtVVUV8HgMp1JSyYR3CclSw9JTx+8XnVm755nCaePVOaQqlHHjTVfpLoGHt9jV8rs3qLpDtm
Yvz+xmJybP34Wtq3mUjjI9cZouAaLWBpLUY5vyGcAbyAHa9aZMfhKMnhSvaQP/X5ZzapxTrkcJUx
J2YTMnO/oSbweR1H9j12J62J1y2kVW0vUqJQ/RV5Cg8lesnH/4Rxta3ynQhlJXrDOekbfXT5Jaj9
YcjeMuVwXfTlxxB5Ua+tln40FdnzL9lvbUW+MmLvmatfv8k6+CVxFJXOo9+xPxMFjr0MziJ2dysZ
fBTp20RnXvn5ph6Z0Pl6cPueozOMdCLamZtiooWOLBGs2/60xcNG9iijS/73X7XEF3dpfdttc+L0
fq6f6KElmTURlvqvw9QSNLrpi5YNjvC+8HhTLYX+vDuisHqRN8jwgwdSiEITjXz677SZc+WD837t
YxDPgVriznYstHJU5QgFQFtnpxgJjWB0CWBS1au7JCn8glg3J6IRut8mpvQeKou+cyUOANbzPhub
4lUnVdl+OV3nMOJ54SbaHUVRqFenVSu2Gy3HFbwdnPu2vwCMNmPyD+1TZg/kkvwoWZb9WpxInQTN
SfTr+JVPZZv8HuNquBCDOxnyGjZgApXu3tklZUktPxVaiwyPcitBNAO5loPQVC+q1OIv3D6cRPBi
f7boP/Tm7rsGYWD9AX7R6c2V1IAcggsk7NyJj+35drCqQXdebAoMntwFYk3thHahbqdk1hcMg6bQ
vbqiJ0x6aT9617bDWmknBxIe2qX6bEtOEE78qM9XNjf4y1IDp/v1Q7c5Z67M9z8lt93P7lOOevfe
xhxmsOeEO7izxZichvj8LCi/N6Qy9Amk3832qgRkyKYNBdw271Dkmq8ntma6SsZ7+NyttQJbiGwJ
VC8NSrsGpfrFbfu7fdwFj5ZN8gaTJWH8TJT6Zd3uCitPUoRUTkkPTDLrxwA+4XBdWUvsvE58p5CW
HTF6f/bHdzLpqihafSTvZp3gS1oCrZRClCAVDHpY/HwqA4xdnsywq07R87Fsw9mLvCzI4T6fjdi0
0DSyceJHsTeCBa2YbcE9l9qjBMfrQ1Vj8ehJQsNyU2BAh5EO/8ltZKYDs3lo43Wnh54VWtBhrRwG
TnffaK/zBdkWRB5y9F/DrR9WVsNRdP9/42YDmLP+SEtKTWSNqI8NPMphnhNce3nRg3k0qvcCmgnN
aU96/HWjSObjmV4u45sO4GZoMWI8+hlTogAi+VcQ+qzYmT9zvzKGciM3XGFTzbvlZCZ9V5plJsBe
R8DHs+xu+TTyLptdpqOx1oLHZtkSUnqpds/55oyYBLQnAnUUcWXrwduu0++5ohFcBWk83uA+xP/i
t+Ap/9BwG20t0KoJR7Tkkue08lA0R/1o1fMPN07luA1MGhFs+YB8U9gmJoHHc0ycukmAjZk1sl1c
zdA4Sz+0UaWfx+l1UnVRb1Z7dFojHy0WStwBhjSY22xM8FfE7fiqKJp6kbOER0V1WO4MaQ0UtIPf
sdAgVdgZnyHxNfn/wd8jw55YvL5TyzQHuczu1fEthzJP2xW/Iuf5fX6Py3oBCxQ+qwvjrn9NdmJ8
SiAb7/GbEXW5GfSFh7CSoSaGVenRIUv6iUOwn9cpHaP4PFavkoCCcPwsp/zuUSm6NNF8XjXPlSRc
I8QOgkvC/ypBKkPizP9mYunzBTLE9vNvmf9Fcv14N0O2L0oaqROlad0Yc+JtC2E3TZ6gBvbn0rXd
ZM1+1RYstvli3nPxPbPlpfBA8R2Ndb6AKHjkRAM4NLRrCL+Wv0dpceBz/477g+1MHQv5bEfUS6P8
vSrBN9WIpffx2PxjrjZe3fNPTDrdM7/PpSHUnuNQgxO8aoojz/GX6Zbvtss5YT51iUA+Xg94PPo+
KpMzR+M7rdZ5H46UoF5Fwlug/vdpS9yM1YmFyHU2OrgvGcXYnRNI7b5H9vjXdsF9f5bZDQ4EFlIB
tu+guQypGXKvtwqjsJfOh/l7UVrfSD7uAiB4w9g/Bj4skVA3FjSTekEeJS4uDh4pJGiNHLqsgQPq
6wQAcAkC69rOCm3+eTtSNU1vXZAuEHLMA6W9sMsvNnyRG0tmNUCJ/fUlN2UfE7RUMv6pz0i4jbuS
FebKbGIAQS67psoYNHU2kD9z5506iMz0EjqYjTsCBgb8otqvsIaoiCAG3qWGXM5yBx7/1P2lc9jk
5HKKRO7k8+oiAGpxYSq0gB5DG4SKkxNrmfSU0/WvbFgEG9CWjxKf+h0yY7oOyTRtVL7T0BGVT+ZK
58P0WDzLn3I6ag8GyrigWUPwgShBCpSc0aCSlK29dG4PmbV1qcmRvI6n+FBKEo1jZAJUnU53Klxj
h5sWOKhUaff8qeNc4q/qh86xSDPTiKJ/bU456v60PLNEt/wgq3/Bq19C5PV40hStMiPv3XUm2gv2
6gO+nQ6MpPRo4wWsWs82pvFrWe3kuG7i9xBuT99/VRpql7dnHfmjDEMTcbSXXEhUeN8gEbv5ALMU
uSIZWXnlr75kmEgKkDWE8eIsJfZtkdlmYGF9rI5HRdQTf4oi+TpW1DsgJmyLQwncOm7OWfqgGsqY
GZOJKARQ8heyVC93YV+7HAAiwyqoAgqYmCfOdWS4vscGEvvf1NJGSbyD/oooa4FZ4GkXeRdqvxV4
mFBJJ0knFuzzHVW0VpgU57E01tbBuSiabbKIiJfBwWBk3ggxMTYRLbDFgfIXXVKBF85CXh5mZs/p
Gm0rjLvwC5+vKu+hXfC2X/es8q+mrev2x7ySRkymqWSPcg+Jk0F9gTFB9WLjgyZ7nH6rkw/h2LbP
AbiUiyrTsJFo4mC41MfK8NW42I54uix3Klg4M3o1xgrzOb3GaUC0mFBgw0XlEO7ni68Ww95SafYI
Ax+OZ1xRZjVz8zZLNbbMX65kQjskHTWI7DqF3VegXUNu6FPkfCY4RoMcFQqb34rpHCjiRmhZceWI
oQnyyfpBZMx9o+pXg5i7K9wGxZsG7gAQgI2+tvVvfVxvPxey0leIFwJtTAaWMArurmObjLrIT76u
zG4NlSvKwrjlIw2SMnKCMGz4ueMGdu5Lx2R07o8gnkwzIVwvdPIBrYbUvhdkDcybIxd6Un6xXyPL
yQ7UFQXij/sXQLG0999GWjVcNZwqMRFoa8O4K6KK93P5qNO61bonH3qumH8clJhzMF2QadvbE+HD
OyoKgVA1Oczk8LlSGg5QscWSIO0LGnncug2L7mGJ53x17WPLT2XKlnBg/4t6BVKOnCnB4b6y+sWV
MvwO9AQTIJOoic5rhU+nDeMGPH0ROjOcrRaTA5hU1SegUdAIBV7rYTx75xWRMSp2gaXeS0nN7u3R
KBer8nACWZSiD1TQL1VogQ2Os2guG3ep/bImmizVykmwihcLm0EH2zQkDPDCVim1afpJhlBLmcWQ
jujkhjxwe/JP/t+OoIb3uKzTOQRL+W5Z9UGs7pqMZyMAolO5yAeTlVXss8HLuuabQGt7ZnkQ4daa
ZYbUFCMBVX0I3SiEsH0orUtmFL8E7MlDmHGf6DbbOvIB1V6FNbIYPC8ol16X6S5Alo+LsECT9CxJ
pD3ULLjMQRr/1TkypVB+/i+v+pyvkyi9Ag0D4B0aRxC78dZx+0X0IO7jJrOrAKTG4arqZkpozpkB
Yr8Cf28UyBQB0HZn+Hl1zNv+bIGoalTFKFZwB4GiHTHJX8G5x+7gghwcDs4kfIpZmEV0NQbkmMTk
NB+5jfT5FVgq0AyFEpBZ5P6Mb8Ww2Bw2oANz7iZVoG+U/bdJCu41oNnPwKwSqQo/UptbQRr7c7QX
EmjdJ0FM1K4ME+OGWuPCalDX3Ybyyi7Gx1TNymKygALUwvFHZS20Kc+a8BVXfr0MONqq0fiObxZc
EOcAMRW0+K3Ht24iW7p8TWSOAY7lgSGB1syXI6H1keDRwSgkqWi7h57QFI5CL9S/YX4jPiG4sBPF
CoW0/SGQS8dTn+H5JO1kMvGHRHdWjgPaOJ7jqldmajblvRR6TeSzWWAVxX2ElrV9yGUhyALKnxjN
Xbbpx7QC6iEh9FTtzKDiq0VQEEsrh+7FxDmU3sqidGY3XZqLrywO4xhsc4ygdbQak9CZ7JfcjxUc
Bn8L+6S/cxC7H5IqQSxWJCkWCS7Rs7T08P6vGklSMTAv635ZIU3Q/kYarEKw+F2b1BqawzKzqnrP
6bBWRmtyC4BvI2a0y8JyqMTwWfXDuzsnVtB0/yr4/c9WVRWNqgzRFP4juPyTk22g9sklb3V4JFaK
a4lgAbrSNsTB1PuwMbLVsbk24zVKoiOyEypA+b0lmzC4NntIjfN7tWh71EWA5LtsXkN1eUBwO+FU
Jtk0j3p0vTTIIjDMj9pELxFg8hL2cHOtzdiy0W1UjsYxmdSPVHI+4Xq1uQDL05Ybph3Hl2TC12zb
NhO0W0GFRNLBlcPOdDcmNpBapC6rC0LxZUZh1Eeckdtml3tYrT4T/Cc75nny2+3bTbcFucqQi+bE
1RUFCOwfsZ9rO7yUKxuwSf9TvqgUoTyh3Qvs+KMTaVsep5qOp+3WwIfCJNd0PuS18STvKYddpHx8
bVXvJOb77ljakrh6DwIQ8JZVTJ4RbPh10+izH+kdrcJAl5OAThierCkW+uoGqboHt1Ct4X0poF1S
AcUugD9hsX3pSDlPftCZ3NZAyYJy/J/68nEh2lTHo4ZAo9AocUb+7WLm12nhaveHF6Nrc0iF+u9k
CDjjPD1l1T1qC01RRoDHLp+QgD7DtiqlEk03Jq6Lv66Z6jwhuR06JaNi+dvsNdMOyVfJIgq2DH13
tqJkeMSegGIccBnY3OX17fK5XpHIYIk+7v/DTISE21ui+z2CM7yEyNg2SxwNYM1yO0CQ0FE/hHvQ
c8oQ+XPDA7JDPNhpkBs4PmWGvbPvG5pAObjdY4/3zgN9pa4TFI5cyqGY9RD8YopFYuUkrm7IHlCg
wPUYCMNOl7cHrRIZyKx2xr7hBobSQk534JhzxI+KR6EEa50CO17O3jji5LEUnhKZJnXhstPAumyK
uxFDXep8I5ZN8uS+0gHRVFcygkPmseImmg1HYdB03qEMzrwgAHNUBkaBEmJVB2X/jHG3wCgfPuIQ
9M13HQBkn7G+tsXm0eu8Ilb6DUdBDRr/krij4bRMrhiFv8O20u6Zrc15xYSkp5pz3KUXSUwpkUro
plGaGeZq6ATaLyah681DcWAsrPRo5plFg5pfgHzlVkWjU0VwIWP7ji8yMqOaTO7N1VNY1xkxMgR4
C0wry8PTTg/ZYhonE+O6T567BErmkBFm3nib8chDd20OTy+fM0SPA2XjZQ+/mhjIEBSYi0GRx+Ba
OYmK65XxjqlQxY8Rhlyo69RwqUZ61bLKQjHlqUv+9W15Xv4Zb37gBDW6ugBuKdl8jrZd344FXdEd
xRjFfuuxAglSEZT2Q6az9oirza/4Vey51rcs/RJJyeqIiZ8fOZtpMHVULBZb7o2lzHyvI0sZARNY
uA+8osXuS9sSYMBjkIJ2Vrp3GHokOgqIB2apiAVajshvmR7Jfpz7JvnbpcqRVM42yVBH5yGR7Rqz
poeuM0lU5RgZ4HSdia5TkTMHYdSANmI7061NJ/vqtLXUEV4/o8rcZfRllqT6hSCiA7oCpmBhL+ol
shoX1P0oAVqKBVrdapvSmBebRTgtA/Fubm+euSOz0vHkQSbbi/ggc01KuxXNSeGRdTfReqYImd3k
qCoz8JIatD7Uat1dUO0WBSaAZyRVIcGvKB59/AN4iQM9LIwSMc+YAgCV7ZzaAkIcLJVaUz/vuYpp
HX/D67SxfxJjW9+WPjGA/1LFlLJi1W7ih61R2/euwjQ8LLP3Z3UmPGKEtYaOauxSDXRE/UBM2LdG
sNj0LIebaveT1uJCZ4/EgwfGXjCQwpRaSqmkKNHSKGowCS1e0gRb4Ge8EkvPAsmma/6mo1Ab0mEI
hd4UE8piaQZOB0D3LMcd1cv+5HaLkM6G59l9zoKS/9WopsWJDOUTx2k9DiXlA0vh/VeEnafwk5+l
jd7D9m4ctNnlRS6ji7W2zKMn4IlHvBYil2WbJVQ6jOy2ZoRSjWwkKGAXEfLTu21gL9GU2A3pvotB
+O8z2nXfe2oVnEjEhGteUI7mURRn+thxmzbRZVjhrB43JIgYB+dpcQsv3KnwUA2aPpvh9sGJELx9
BOLLVRQ4O4VnBY19ilNy6xeU8Fpvuh3598UuVyyK6am/sy72GXF0TmX8HtxsL3+gR3zymlpsuX1c
8zhgtE8Gy75RYm8d29anlrB0J+UqfmkLRH3EflBCNR3DqPj87nLGVLd9bCd65zF19h4mcuKkFscD
BeqcUPOFjuCQOAQxvlwOzTSKOcaNLvye6fNknD6vkDsXw8Syy86OdcfGJfd1jM+zbzQ4J3gM7tz4
OZqGT5GG2R+S2Cu3PoLnKQ90pwHSKI+/cjicU8q1Fh4b4PrQvq4RvD4NC8otPAaYfmfaBKgIBk47
l8Asi99XfBYj9AsKLSui+he9Uqp0IHXAWejAmUYSUNdCeEZv+srrIK+lZLRjIa1Nx79/1V6mFNoL
qz1GLBvFRa+OLSbik3cGCEC94IbBXIf6MZijWJmTvjPsQsdo9vkrNtR22UHBFUT28ImI8oj4n2Rk
XVfk0IVPUv7mln6tYQpuVLDoaGwo2m8vZAmqL1ppeY+I0Qd1adxkmjhDJ+AQ8u7f4EnxKob+nHIx
OOcafzPpOJeAqUVg2eGxKGB5iyK7bhxr5slezkNwksU5ZxDCZ743azXiAy3VBU63/78otcDUsYNZ
+TVJ69mx8D+MpKrWjHF9egumHDdYmzkR4SsfOTDSHz+yXN1lz5Sa89O0OPeHTpMcnjVgmBnP88wa
bOKRwePsGjnVKrxPoQq840Ph9mnZfyAR6Qw5/y4rFcSJ4uMAXLVf+Eocxckp+8UieeArnCrKbKzJ
xm7Az+nHv0rXY7BYFs5eMrHsh3l714BZGiEB/FR6RuUPJoDMCAUtw6gmQmvogWtrEeUBw2QewP3R
QCLt3Drzc03pNQtBJgvca/OLKuvxGIyG5LBpXAkbyj9A1Yki7XPmjhr28XiXbt+ffVyAYWcyExaC
2FneDMLKpUu93Wo5d9dpTuPI74liXic2bEZXTQ9YXDdPyjEYcrYALEQZf7FCzfiQwShaTXP2Iust
30zIclT+BZ31FcsWftp3z2Y8WRwonWZftGsu0ok1V+rQ8fsABuBbsgxO4KDANIP2NTgkWYkDhJnI
JNaFG+6FWjNPPcmGpHCOYtD6BMeHR9UKTdNDCkQIbUoP6oIdSzVwEy0DEDnF+o+JU+gdXoLf12dB
pmcqJs30t7LVhuVNEdKK4e4v4lTzWsjIGOdIvoSXP+gR1FFRCBb++1pPTNycf25q8Wuz9q/vyyjV
kF+qWSNy5BCYeGfeekrLFNqlZ4/LpkMsQsRroxGTuaw5YxcM0SZgSTHQ7JLZptw0Mdzvvqee7ee9
n/JVz18QO451z0/wE9Cqf2iV32Rd3WAiO186Hv7amaCu0i10yoJoQvzfQAkOdJJW/fmb3909TqUM
ei5P/avApgmOYkqI3j6IN29IwzanqAaZjcrJV33Wcv2pwL68eanPiuj2MXPJYEdWi43ESoMqg0tf
n2c109Wbsmod8L4E6rW8tWJUnxlp1MVgl4z1amrSlI9nwGsYUYylwFzypYio4MEKNSNSjhXu56+S
ZSoXxRHcNNpVXKxfb987ava8L7Gd3/se4KxlRvYKQCTFe9bJC6bzGU4QPvFVNJsF3dJNsFv90YMC
K08G+KHBOtAlS2aZu+lrQRM56ZvWLQ7n0mZpwXdyTb3bCbJYLmscnKBW9D33vB7IipNy2WxSX4jJ
DlDkLlNSm13bVHyWKcSn+leviR8xqknVzxiwY0w33Qa74Puj9dZ38G2pbK3UarpvqRIjtYzgHcm7
EnTBQCUg8HMEEwZi3dKeJXpJrsSgT5OERAKzZ0RNsVv4y/OsVQ/dWivMVOvu+8HIqDUbIHiIVvaS
0zCc4SS8S5AzmTM42AMaY6ydpsEOTcIjOI5nQxXF6Kt1B8mbcdr8HNMIwyEXLpqbMnFaRfOVQ1Y+
4oMGOekqPkWhPPzLvpyJsayWldE7VPd8gFqJi1dSdwbkfZol5YxLu8Y0AeXQS0zSwAvbxeJiG2st
2vcOoIa1p4ji6txxtmrdyLTajDf/b5hdMIKoKUH+9wYJ9HV31uvr1+4TfFDB3+YmA1rLndY0M7G5
6AW9oCHOzLyknY3cfZofKzRnnH4L021xlqLl9VS6WmuHMTUY+OauGjgCmxjJpuqeBULZRZyT7JfG
x3zFgBHJzh8dufR/9K4xm7Zc/fkrCbqPHsCR2chsQPD5ZlaJOqRDZ/Aehuz2C6E/TKW5HoBbaLC0
tVwf31yrL2e5VWjys9bI3VRtXY4G8rwnYd6hEfnQHnCkXLEaFy03bQd9zGu8D2/g2JaIK8PUuoRj
U8w9fbxjVSPDfMWA/UR4RqP1cNoLkXcow5AEHI8gIeTVybV4EGyLke8N7fxXehWOKAd8/gGal+qj
HRCqpJBs/VZ28/CykYtr+jFEwTxTGqQXzK0O3CWFwKtQ5N+X5k8SDvLmdsURAieWSlDmBm6mmcjG
oYgEwL3KdgCj/Id5rJ7Xz64YvLP6c5jIBoMtCY2x3VxgAVoTUnuhJwC/Iuav+oYf746qspHT7QPD
KRvpErojeOxQZc85JSt2m566jqXwVA4604OiWCrL71MgTPgppALBnyCOZsx64n+KtTAmW7F3LwYd
aNxzq2rkzO+/KXd5BLu+pljCDqQuxrTcmiZ8qE1QvvRK57Px92k8nJSuXW4t3tmjk9WFA0idgHzX
7EZNfShzRX95LhmVawVvtS6YDk9TK5s/HSpgw/+Eb/x5Mbej3UwuqnDuW12wFmoX/mP3PyROcHZ2
4Sm/uGwyutryF9QDNcMdmK3lsOvPI3kbR63dzdtdPB1wFpEYGhXnFYZiS1S2XMjWWD/UpUcf6fuS
4Nz6w7LQ1u5yKfCtOj/dxwaeGna7S7ZBM78J+CtdQJk6DNdhsSG5TUhMTlsbF8571NTulkjgS2Qm
LKQEOfxnoWaVSzxd05r0rFO9BlWHsi+osnR7neY/snp5hiZR+U6vSJowzpS0dj7KWf4xd6P82+6d
b8WvpqbsHDkoYT6r09PsYhOxM/YVK/+kmewNQcmP0A2aOTaZX1WdfiPLQXsFTvpXO+/DQoW5UtZs
Ap3FQTVBjN+9Xd7Ev1sdV3oS5isPDcyCAZiG/vEuwwv8C1nL9tPgpnGPso/mQha/3ZbOUGCk8Syy
Tw6PhLNQirEMV+2GLcs37se3qa7NQz6m5KM47YMqNRzHNtcRbzX5ZztswUAbVMI2TTdZ9sc9MceU
Evrj7jZECqXl1gOdQdfGPbpmVQQ3elNVlLFUlkhocnYLGbcP4peil9Vqtyxbz03ydbHkqkmJuMCs
+aB6q1divcymgVgIlCcWCcU1t35ak9abvfwxT2yNjLxXKqcNaM8UfGW2hYnFJEC+mI7lT5bFc5/f
1axa/IGhkk+k67QOw8/PsFWF+pyA8N4eRn+sWxV+imBjb3U3jvF+CfvKLD2vNPSTDr4a5VLQyyup
ozy6/V+ItAX94eOP2jY2gcMzKzkNTA13l7iuDFhv/aP7ZfVES5X2Fc23Vq2S4QT+GKVcMJShm4mh
xj0NAa9w600SI8J7v30eu+PFl7QbwjAwICTmRTR308H+osucSY8nYPlHWReEIhIt32hV9vAQkDnr
G0DtDsNNXZrEw2V0X1T4WdZ6wzfl/F1YULTvapxnwfTmPO7W9lgw0gwrKltE/ooRzkrLPqueGoi0
maGmIZn/dORltkpSVLKblNXj4VA1KqcAYaMgwrJCDbFTInzMeX/lEeWtEMGj8aBGiA9T0oJUrZDc
JClxTzx37HcfS+h8AhzVurS+gjgnGySwKWN5ngIa+TMQ5FfeixztJAfZuCSKdZtvfroMgwR9qna7
dxiMgdqrSvTd9+wNFIHwMGlTCJGO4s9chOw15vp8277JASTITOYDQ/QSh8OrtBs5YYfCO5yjxpwd
SEXyp1CeO9C+QuBTctNio0bvooGRRFL4GCm0tRtWEGv3itWM1c1NI5TlCMU3E8ibIDnw9m0LR10s
nUgYJ18fZbtfC8DzOWh/ZP/PEi4Go0cknHCNPD/b0giJTSe6IqRb+zKMwb+E/bfEA+jh67mnic3g
0u1jQAO5gikHYqMlr1zqKr3ACFEkaV7MfoD2oMHc4FlOubsBfEAiVVv9Y+c1I2xBRMXnlXznoWvd
lO5/FC+pj3QDvHcsSS7IM62sIpHYwra5cbpYgCeWtCKESX6gJ4y+fr1FDcCVX0sEI/ssa1XXWcGP
7Vc1+Zqjr43aAqwgGqOAndSHTA8qUEthHPMPiqO3Ykf76/kClSWY0SGi+Gg1/nJUzGqcJLZdHyxY
dI9zOFeYyeJ9tyfl4dP76wLx1Ba0zQJ8dWeeiU8bYPwJIfbD7i7I0osg/HXAFH2nvkapdyKIqa+4
5hsxvv+ZiB8G5Ned9IjSVOvX65RAhlob4Y+Mq2wD9h1OwXcq1mdAQbTaJ2tN+5XxqgbfWGdBLY4y
uXvpfEEZRxB0EsC86E0rDlFBMpv5YPh8X15AyR+tMr+2rIhXq4FW7qAyqdcUL43l1PVbJDX/cFUi
/TV/OxYp8CxwpTXOmAEqNApVXZEx3vId8SRSsykC/MfOWpBk9rMw6ZNOIgo/JPJsDagy57RMVhNe
Y2GgNE+j1Maazvq6MDto0c2asBz5UhwOcf/Sb02lI865IyfOxN3LPbkMs2NOyE4SRcwnH47UOgG8
FLDECs28tBEvZRNeomKOF2/bNjlnKgtir9vCEjQSHC8D809mz3suePMjKJ79muB8Vl8Rf/apaWDF
2CYdyIaCYoe5MN6EF1EbEL4xuHECZsQOzJDeulg+9bGLluA/rwWFYbQLuaIGNEH6gjtm3ttOK+41
zfp3+hkFMuHDj6/hCXdb2l3ObZWP+XzNfXSJCVURaNISU+/0nhq6oWVhTlpsrtPIafFIA50NsVhP
j98huRiX8Eo9BY0yNKRwwkdRoueYFDeQhh0qOyeIMbUtgveQ0KMpHi67MuMbvxbaHpmaiHdsTtID
FrCzsuSh3W+SK7g3iXQ9REls/EggicnPbxgjr+izFLgQAq6OypUOvTjbb7SrW8RA+PWu09M61/K1
wUpCGaVNhDQjpalqGN2s58wRVuzGBZKgw9F+L1G4ZNekIgGEGt4Q0eCA9QnDK0WLe8iIKVJ5O+DT
etiOFw2cDFAIIPXZMdjeN6WEmVXd6QSrN5nWQpkvpedB+ZMoG8RMTL/ko+HSW0Z35ewRcri2+EWB
566YmFAM9Z0GXRWDqSCwhhhf0gwmjPDwmeJe3kEQYoCoYGnca9ox3TB04LALdOlwNlCTuWWbXKQ3
FTj3NxiSDB0V8ZmApBauyBUhEyhA
`protect end_protected
