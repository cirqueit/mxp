`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53104)
`protect data_block
0HpBwuY8CzlHdr0USFIcMKfx06ni+Tu8I7Qduk9qAA/haavNq4EMYdXwRFe+g3CFgU56Q6MqwTRQ
z/1XSnETbT9txiK79uMczEnoCdmQBLmgz0J/vEbbJwITwT06lc6D+7vV08GLeszTof6HrEZb9PLh
IqQ37W3i0OPqsEJxmNxOXYH90O/MsaIku+XF6Mit3hIlNioqHdLyyZ33VEMhdQ+FlCB01kdXbX8h
z0zjFmHovqRJvEIjRD5/G1Lv34rAZo2ZaDh8EGbDJoGigjCFBuhI2MzUhzMoSFP9kCIKx9RzjYgM
lvO2xUa3XHH905Pl2Qr3QM+TpsB1uv5k1Bc5g5/ZhXSNCGQ/3U9HpThjV/xj0zrQ5hsiIxU9hkL9
dbSuYjyEW+sZKXCQTVqBPMgkh1k5ULalPyhVZ6bvcM52vsGZAuUWHs0V0Ok6Ulp8D+50LAK21tJt
SiwzkWCiA5S860t6wI7enFgf/nCHFgXuFz7sJyTjokxjhlm481Yu+iwhztgCmPmfhvIO8kSdpqHX
ZuIKbj93TLixb47XMDusbr8UnA3pamQHflgvuWeKDzeRVOUwDZomoPheDXFrgjNEFeS/jNtO8omd
8Q7ZD7v4jSOY/E3nL+L7wTP9XEibhAEMzyp3Nnvx8b9zRNyQqQ0hYVEfy13em6gT8GhHuDOsevPN
HapGnobDkZjUspo/xZnc5AWPHe9MBPx3PnCA6uWHanF+b5u7d9DF7C7nbMctfoLnJ3ecbHI8Aru1
JqvFYkhpjQ97w7fIn7Dr30sMO4RJ/xCzQsleLEjQL2NgF+UELvR0AhL6e/VCIkmegzROVpTI4hI9
ukqUB4697a+tU4LKHO3BA5evY1h2NA3Cjdjb2JehVsGp7cke4Dj9NR+nzDoTVob53XxJHbeccZ7Z
hG9C4hky7MHABeejxW9ikbSTZF9M/3CVfA9ukSxem9BdTczJYWkB2PwLvk7Wcyx0BvbDCpvaHz/0
u35jUIETEibBNHMm3gZ3mQWMK3MXn00I8NzPn7iXTd6Nayd4FOJ2KQfeZQ6X+j+ousRRkUDOvrzx
dOzlb3/53ikruNx/uMB6455TyV47xo239uIzQfhivWb7Obph1c5bg4FC0ljKMuIZGqfyvN1+UdLt
mzbcGUAMJLckE+uT+318tZrphYMfO2j2mZVRAWNfZDCT09iX00BoOw0K0zqcBEyDWD/mGZL08zuu
sh5/bC8s/Ni3D/2nggNjapVhFCdhWlHoNNVbJS8O499PKbm6ktmj6dZhP60dlu0JK/dr2RrqZ+YI
YJw3eT7dbjMHxyP6ISXDf3KMLXvgZk+fT1H08ytja83pqjgOEZO8I+VMKyIBZMGMBD0mgGQidH1l
lwGC2e6NKZ9o+soo9SE1M1LgiZGYXdh0wReu5L4b7nH1JhDaUy9VKU12HpMo0tiVJHGlM/kCD8UK
wgFDuBCEC3PCwlRKN0HVQvtH0zBwBA3jqj86auixBj9+IWE79yT0fwerlpcS5dRUn8HNaLFCSaGi
3hZcRN+erugj+Jo/0BBWSOF4QcN4IBfLZbI5GksqhkP4YWbQ1GgbZ9eF3CmgpiUHFXVFDSy7BHuG
3kPD7fdsJDV+7dgGFaeliwqa8ejC11fHvllE0X9EpQ1hj6XjcJlXGiVotCKGSNDSM6dwfgvq0oPL
6YUQpEd8fYDuluvrB0Pga8wRG8nMotXo6CTH1b0YPmLHx6XSlCwftAP8PjhovAsVksnvdq9tUghd
IAnUOvy0dDTbKqoEFOLsHNu3XFhdDicOsbZmt6YSvKmbbu3vXnvKu3550oBZCy2BmzGPSW1AAQK/
gu+yQncheqBFFXxgqSAxwWnpdxSwMpwqVo1SCswhGkpjj8KgC4CjpgcB/3UW/YO4TpMn/30WydLq
A1RB8jliF/ucBbWpTim94ftBRz4rzZejMs+g07MLPFR0tbc1vmioGjsll/TW35Cw6EWydz1S3xv6
50EFQMKq5J7psX/MRj7WhaElzb35PO3dk5LbmVnnYLGDmdVWQn5MqCf5W9h1Bs+9Y+NrDXn41FhD
neuY+Xrcd8TFBc9EhdV2gS6ONb1zsDFeH4LOxI8dsZYyZqkisI539UK5piO3bg+q1GAnhF8DBWh2
vPiFxtG4fkqSYE4CwrYn6egROqdqShfaqguT7SqbI1EFJDnN3fH1nPRSwuIJRW8NCEs7jwi1jY5D
ZG2ehMQYH/CyWSKnKokksMn2uNP3sWPHD7rkEcB8W8yYoJEvAexThHcOXquP22R0rxY7afaJ1ldA
esBphEE3l0A71yDmzubqshSei0SUDN01EUJStI3ggoNBWQBb01onVEfCZKru/Ip1VsSK3rc3ZF3w
kxlUrkQpKwFN5ep3rDLXzZGuDCzosn/FvhZxffl+9zbxCSt4toRZxWQ9Cf5T0ynrIwknqrHBov7l
dzQ5j7iLrVvebU/m3GpPSRI5Osh9aBtqb5RXK50tJKL0siZjl+kyMbuJWQtwjfLjf2Sq4IpaFyT2
rVoKeSzwTn4PUjGAfyY1YJEBRan4UhZrXChB/WWvWIPptEUypyZUPfmaV833CPnczBtXvtZQfV7E
CctzP/WCLqQTMkArYG/dYv7GQG6e2/WLlN/uUiP2YJWX61oq9LilnFqPMiczgBPEBbTrv886Slz+
8HI16b/vgOIdvDA+00sfTffPfmjqJ1gXY0qplDHm4kJYQAeCm7WS6eJADeFh3sPcCUN14uk+/fFS
Vt+FL7szd/myJSwxSJI1dsHa/9NIITHEOTHahg6RDPkqgeG+WoyEtT3Pbr3pWdA0hF3Dzaf/BbT4
ACREvRtkKgnTdVqF+tnm4WpPCLEvRekuE5eqEFvTxR8RmP6OnsvqHlQt04ng511DJeYkEOmXDKLN
CQfC3t1oIvFWw67hr1qcKA11xoWA/2sCnFkcDx6dcdBv9mrk/tn9GcVUQ+uVexzYzKvMgCnVqKUq
CDlo/qe6vJ60PDtG3S0W29cDGApv1jxuufd7nFmb0gePdbJ7PP8tOQeIKCZayGmXRWXUnMQgNeXa
Jx038G/PlGA+BqUdbhlbjPLGkrzYG77HyhlHxHJQld49+1LIYSpc1YzIu6Nj0Cq5dEWktmtA8kQ1
kzK8jiHUiP9IEc1oAqQymqlddA/B6nT3r6k7HVwZAbAE0iOuSpdJJCGPW5rhtGvtbL8VnCCbDAN5
tbqYmV6u29dscFM35sjg44zMWseU3PQFyWGAEGLaU/hP5RygqkziDSdJzlLgEdMF2FmrWE9bSu1l
pEgdc0wntA4505JiKHalIjwYhHsztVpKC0PLfi9a1L4dhe5G0FzriR5qqyFcvQKKGt7Rc8YnrggB
c6RTnP+t3todnmNlL/x7GSmFEm4rNNzXiRSACg1T79FuYKsGvmW5Ya5BYrBkHsXYMmY1Vnp6r1BB
5IX7pMrUGH6xL7DN6Te9Zha5wsKngkBBWiDxiGrxMQQG1cfUGNnW5f7w8qPngEFU4/xq2xj7LL2C
p6S6YI5QKeZDa07vQ/U9FFZQTEkLwvJ7jNzCDgxjm/XfULPB7HoFSC2ymRLL9T87vr3vYH6dT5om
48G+hBXo7pgElznD3/uHpmrkGnQ/vobsUx7ikcpIo0zlrKw6F+K2ywlMkRNVhOVD3EP/e67cbM8i
4qaePwka+CUfLbRNwoATmre6OX34d00PijT8YaSsFDTk08WVm8Uvwq/XRA7sEXTt+auZ5Szumf4y
on5KPt5QvXgh6Kn1HkOlDtM4QF0iFsmKsFak2Qlg2bP9Bqe8qYiU2gLq1fwqGjbKPVbFlpr1bVTl
NGTW6eEtSbxMVCN4kj9f8ah2Y5gpw1chZGIR47e2ndmwO2x+g4DFdo633+EgJ5a8EPqY2UiqZe0a
a2cm7XXtJFJlLIIMuc28h4hkdIJwIhwozg5qZIx1ZfuPNi8ZS1UIbGx0O84INCcfuor5zETOK8Mo
NdjG8+YD+sDXFYqzInmR2kmZaPCGsRU0Z6wT3UBfqoaIh5LHEaP+83657FpyEbFkgV9FpZYgary9
Wk1ocI3EkyLGzYPJ9Ono8lppcn02MCs6m01ZxY8RKNxEix3ay43hdV7n0OZp4E4skK2rrgEKaNZY
8USWT+tM++4fE123ezeKAjfGmYJhSiyuCzLAXdx5jub/eiRDA84kjE1fa+qvDkALS3NxLGgWnApD
VixDPK2Adl63tXTBwDwCDF91eNGQZkbYgCZJAto3qD6m0jos7XzUbQSoHFmHZGNYi3qI9BcxvYNb
xJ1ZNBPFjb4vRtor2Glz8nn57L8qbMYgWCyKOJjhNt74YN5Kw/cTF9ZgGckoE8ooWfMrbOnE8Q6n
aKbcjRXKMaXKOKhEEhuSBFXIVH/VvJfnHuioD5wekjxcLilUKrmxhdowtY/HJTqctgmZUpfV6diw
ABInl97nks53N/Oi5vIKwSjLQaH1mPhZCeutxgh5xPzlfva1enfIgxqqctYAuA01Wv792pEtKu3L
7GYPPEuLPj5hH7ZJda68GkFytdyoWzzRZplqOwG0wsORn3GahGH9IuvzgOpsZ6fi1CQfHhaPoSnP
FbDs9TaTYBqPVL+tW+uKweUeHJ6WKrcxTljBQVPr9VhBlfX6VV2PRRaGUvn2CJ6ax7zJ1ca8IUtW
YO/JnLAKgEUqb4Wy/NVC3fdDXB5ByBXbOGmTAfcVWgzqxgG7dGCnBdOTlrZxIcQ1s4PkzxiQtcfq
vkwNqa3sV5U1413yuYyYgiimLkj0oE7k+ZrjBjqHg9ZAjoAsQ5El35gZQkTTK5EcRC2PxrJSExRU
I+bKir98shjA8EG6lQW7b5BL6G9P0kXtbCIf6IgAIV9vB6FyYeSuLBYE7S1y65OXRzBRqHSbF1Tg
A5I4mGvuvA6xatCQyNWkJ8yegGDRUkMCHAF5kWuP5ocWn9fiBSOSVeG5seDzRWPHVct93akw9FlV
PPfyy7Ll3+p5j21c2LVua9rfmrokPEoWyv56zzww26M5EiCF9Pz8HX/Wk8eXB9oQ98o8AmBpISsm
eZV/OEtT0cRjvoylOYgmk0NSJMw6UoxODNBEiCyNB3X3PkBz+0MnsKTKMmZXk8KPAh4Jq+sF6NVi
1vYxvRtYizZYYis9fpgqkx5mmycuqAvojwJX4n9R1igiwFnTlJjN5g6ctm5l7r5FS2X0GXeOegYl
4GLvgmtK61mWfRYMS/CnDekZ6nEBedQB3Quix+k5EjBcrRuA25nrIuOPZH3ImikNgAWb620VI7Ar
IEuU74MNLXSRsVKn8goTOO71sjjcZ4eqtTWOuWpd8Qj8Zd6rUA97u0nkfJqbcnzQsQkiPxUH41Xu
iFuoS4ZbVbRATZ9/gOGYJDxQATa8ctuW1MSXySV58Agrg45Uiy7wMqnG6PDZEFRuvQ+Ig4+RqnxG
AbqB/kmWnSw0E3iy573iVm3/npXMEPS1+E62b1TAU1IAE6jsYnbmTAWs6BrDG4833eT9Itsd5eH1
2zenFmZ7dXdTroGVQKXbtxoOm2H04ums4iSvk0o0tjIv0QUnO95o+QVw47+JkjHX8QGg1k8KZV+X
RzvU1l0Rue3qfSt44kM05xCSqygzDpBujxvRQmiwE6oe4OXCDygJH5oPjGR/Ct6ypoU2kaHHlRmS
0sdDBTlipLpUM8z2y/oZwI+Mz0voBT2Wp+RTYGuMTO5kQaV/Fy0W/3Z2ivs0gT9wH8W9OSaKkdsL
LJjgBcUL5wlpSGdaO9dRagxvRoMCXUoSHpXDhPjMv0QXX11CeTjmXa884myR9yKcQG8IfnmhCnXf
8MGiN5HBuL4s3PSWVwODkBT5nVbvAfcN3yRaDcGHNqLDBc8Gwy8WH8ZZ/3g+ZEUbgXfa0QszGlA1
sJoUDzEn6aK7rPHta8Sgk/+DGhkRu9XmlL9M9v/4XzWzIes5hBtqdjsHNkCeuOuyYQwZdD1B+UT/
Q0z8Ai6TUv4P1oRsvsk6/jNJU6lGDhBKliupNcuWi/Je4QIEhkpw3KzeI6G5UuFk3E/ztHAkB8dn
MLy3amayTrePPTt9pxw2BRkbRywZGXDLHv9IaaqLbpea1EiNCqKbMR2D8nT8ZyVs966gVvpStKnw
rSFxFgCuq5k2pVmsSZLqlqOcG1mJla4JvwFeOUwexUKDJOtRLYWiAdfBXlnHs141RG1cGsDJgya0
V7oB6f6+qpg/OfqHDBjxpspD36slfyXwpSJO7m51/wbFG8o2nzs5Ju0/RtLVdhq2mkBwQr0lr4hV
OKH0s6pQzQTZgLjGqkiPr+w3eMFQ+TUiuiVpt9xa25x1lqUkcCBYF+nQ1JXen+C4XzI9cSCXrHzn
6gQBtJaBVkbc1v/BpzPKwd6d7xWlbQu2fqxFgGYySJwMAgGfpQrtvzxXlpuk83Ny0MxLBEmugFbA
vA7+4/dGVu7JSrXZaOwLj+4D2YgPWrD/Qek3zS6077afJVZ3oSUXTR6dvoVAw6bQpWaMrXCrRsZR
sNMYnMufhBNHMecaW8mZdm8hclHweEJZlAubvQi4C1oqhXIZTdEktvORlovk2l6CCQ+7XNj0Dhgt
QMFRqPxNGzjGpt9s98pKoT6lwc5bAIp9gFdpMwLW6I6CX0KbKAQL/Z9BlZOM69oYSwbCqgqaxbhA
3Xhxau9CYZQfHLwWXiHngsXKp7ta1A/hcuKoeLvXAdWR8l8xW/lYOYVo+vA2iFFt+m6HheuCJyf+
jeYDR8/QO6uZo5E8c8pvULnl3puq19IXaCHGOj8sPbYOQmxwA53wfYT6Q1MNV7J1H6BiyW8d/QRF
BfSGMuILkHBFRE/IXSgYgwpILhLXDtPBy7WkDIGHA9WTVGrIr1+ltWLgnNyyeSz4kB3Cj5ZY4tMf
rOWNfe8AMMMPmVHZE8W7uaEgEGbqIucjQ6CFqlqFSwZQydO+R3MUYeiqWRL6cmPT9CCeHwfnHDlZ
TM97k0m7DpQMvx19+2A0gAF69umx0KJVGPkjh5O5qNUh9FFINrUoSPnaC+M7ahNFdAglpXuxUZBl
KUlNjrHF9nW2+It8aZkWz1C1kxmy7BZ7SeZ8fjAANL+HE1dfEtRRZwLKYQWFD0EeQEyAWrF36W79
rAjf0SBz/zJumI1Bwgty61zfwvhc3vaAVFJZjDCDyE2hMLSeQIGwHbVPk6bso5u2WteqZ8NliUgR
MShM1ck7J72ZYqC8/h3Noq40c8HvtO6BBrmsG7w1ji7lMl7q6CwiFrOrFaACyK5/nEmN1suiYzcv
M2GdU7V3whPSSx6o0SOvbRR1jZVDwMSY7XHc8iVq9mIKSlD+mIWq1EvpdLOnlGxT3gZSIm3Xg1eH
ezz/xfUxv+o80ZcPQw2/XH1n9tJmAy0oNoPTZOHr/P80u4gGGvXIQvF0Ke5mzfoNrzmk/BFuR255
WCvGq3XEmZpPV/YM9Y0XRqpQwmkW9B3HIsiIYxhtl2Nti6phgnk9+NYFhmdcoIrNuRxerVc7k3Hb
zypHMNKr8qiesGcEfIUqU+EKt290x73YC5zlAw16oHz+vDehGNx0bmiGqpRqKAGeUfvObELYQ7ro
5ENyxO5WQ2+o3kTDZGMbn1N5KjCyEAY/th0gFFHTfaaqfuxd0vlV5IGtBkkQBBCyJrQg3wuBL7at
rmEERndBuH7WyfLHaJyh5etrcgKANLYRRauxY3O+QY5F6lv5d9fR6GxEuaeJUmXypkWGRorGznh3
qdEGB711VC764+Bx6LrLV1wkXAOqWCCsEP87dvnihyJWrpzwrLtRwQ56OPGg1RHnaqIQJwfWqgxE
iBuHGc5SSp8l0c/aM0XQq5xFTgWpLBkpARF34HQ5VnFyw8ZIELY6uiNmGbjasbji7qCZy87CSdD+
2+fC31dCmAAAH4xVli/iVXnliqrgB1A3dwwsX4cVnWMIWD7wxy8lI6U7U3bQEx6CrDzJhlXkyQ5w
rYJx3rfiVbpLn8FKrm77rVeCr3xxVL+imQa+hVSO/R8A1mKaUIrBm04YZXjO/6TV6Qgkoxc6rD+p
cZtntH6jTMXv6MhyJ89Ev51GzV9inXMoWVu/hW+Rs0fJc+kHGoQUTAdg29iYiXrLpzqWkqkEfdaE
7UT3oEUFT2kHL73PzGtofT0KAzA1D8/rEOJV//hHY06IiJ+KAkBx3sQrGfckKzXSFqycm8bc7Ky4
Sg/IioylAEh+z8Qr1sDt8ak+eIBijwm0YICYvqgxoW9sXLC3TFE+j1uyatfJkq53kxjoCzPwHSdb
w7Y6Sk2hG4rczy11WCYt74s4WpZ06JEbWkLSoF8yXovty3X34gDCoWtINV91+Kc+feyhuSt52VNA
HnZPlblE43fifTYrWYxLUiZDaKqXoGuE91ku6DubuJ4Vpm3dsPDvaKkKgb1/19pQsGTN5m2tL0YW
74zpQ99jG4lXvqtlhlkR2xhs4e3On7OetifZs8D/LXPflBKUafvh8wcUzVdgfCMyoIv06NEEcxfl
abx8EhWAS0PqHS78HdyzkFL1nw2vfaXgjxjXfe+JuFtBs90SEahC21IzZvWzZcfm4EKG+cVRHJ1F
5OBk1GyxMkWbh53zpS1d6DHHwHCsYqy+AM6mKfqfS0kmRqrkHbWnSRccbT6ti2eH3iRmuZfcxQbu
5JEbdjX/mYnk+shPDKxEwk8hQMNMsY2ih4qEtru5FvkQIGi4N+o/+wPyPfac0B8gt1LLejZbK9F6
fdLh1VGtV+xNsfb/WwpM7+4KgPZBd97jKUd9zu3VdhCWyTwQnsQcWJQjBr5G+WgmYk291n7fQtEG
YMTOXbl3Tt5gkH45+jpOHgaGPkVtypYn1IO3FhGEoGPJIP0zuJI1BqtHMH/8tPLrFEo9tr9nfWpo
LVIcybOrgNtAWOzETEdqN5m0S/dxfrWR+HfB7imfEEi2zM0hBfF7HuD300UFG9zFroX2d3Ntg6ul
pedJiVJV2pfWzyXZpH9Go5xgh1XCOdsxzvmnjs3nAsY9iqXPi7EqM622MGl6rELWPy94mJO1xPCr
I3GIg31dTWa5iqT1Wk+Ue3D+pYc91L0nkfBMyeaIRWZJFX+JWQSGcr++a75QkwOHScWgrfKwegnB
8FtEjJxVjx7h+RQdJ9hXzNstMQiHV4gLyKC9kCi5NoNkE42iJl1JjS6YFyJcQK/c1Hns0tjnLV1N
9Mc28oHQkmfHIueInE1mT5uiSb8U+LDWGAd8ko/+RvsoOhKhX/nQ1hzPVByOX/hK7tawM2nS0o7K
SzdbWvxAy3OOKZ8vovvnMfGmm5IDdD99EEGX6Pd8Q8xYwFvfASbNsav4pTrUC6zrncxLwy4EDiaV
5O7ufXImn2MayQoYS5lMhlvc3arMz+lg7CElJXG/xxE/d1QPxYHrC5j9W1mYI53IRVTVsTvqF79k
H1E6MsRxYqXr0DI45T5V6RfLaDdl+hmUj7Y1JGOYvl1nFMNrakaPtPb3R9xrVPBZP4snL7JqrZtw
/9YAbzXXh2NMuHqBeUb7EVq681/U3EWFXNLJe9BACvpnb7rHUsRIcDGVYG4zkaIf+LsXD5ZGeOoQ
JfwPDq7g6XCSXcJO+Ogl0/qtl3C9FunNWbPKJFn29S3Pcc72lsnbA/RgekW8i8cc5ukl4COKX58Z
W+SOo/msB5Gj+J37K5iVzVJZVFqiZLlmSMpTwdkf9j65imWupACHYiwOyjstPQH6psu/gJ6YDfYr
Y4EhmhNUpacAhJRigOrpexfmAXQPjLrXpkYfagy9/2PT+IFnSZxsu0U42bto9FU3tTUkTZTwUai7
cNAbd9tY9Eakq0GlQkJB2Ce/M7+FkNrsj1IuTX2GIzWwIAu5+ugAvKwWpsBvx06wQCXHAL8gcIio
rq/2lNgcE2ajvgK4SUYBwSUAR49VxKpe0pVmPd3+/q38x2XxZVboon50XT1pz/lOD7L9WxknwPIO
YwcJglr9f6c1vrNtEoTHkU5Dj5SKVDUVeu2ugw7df2XNItpEzhN0691LNB3mLzQxE2Del0yElRpw
pV3Ds2PpkYpgHolUWXqKmTqHINDi8ol3iWUzqEtYTBmeAjuoCNq3fCoPhndRu7keZNk4Q2GUWDbs
CYwEzbYw1peISpPBZ0qc8J5nOOm19kyEMvF0ewXYDBoCp5ras/He9V/wI+1axXrrixWPmB1TCian
dH6MNuHGEEZ50VylzrWv/uQ5XUJsydNkN++GbAnZlZ3iyn5p3YBlWM/dQrZrCG2Ltf03NJDTNtt3
mVXgsT3Ia4uRZS2RO24PVSQOmZRDV2w1DXHqNbWf/qw0MxeaDoGdbOa1R/Y3bf7G8cy5SbNUqFdA
Y8fiz2fNK/oG5IUgJPvvAxDbjnVgHumDS/tk9Jc+79O/L3YxiJk18Gpl8dssasyxHrD99UplIzHo
8rx9xXMKTJqNgNQg0cM8APXjcQdT0xbuL0P1qq9eW75veqG8FuiTrXx7lHVmmrjYDGDrSh+FyQeP
u3dx/yXLuXsS2beHZzOSKaDrNYIwiRlPrLWeR1UAw8AmXHAgwpthysWhD1e6JCQKreKfYEoJDr+a
rFIf2fEYjax0IkyoCbzqrbu0VZhKA/qVPLJlRwVMWQppUhSQi/IrElO4h8mbp7JGCm6ksFHeZ2uq
tYr/62wYhmA6R3+2ra6gJ65XyI7r0crSv/9UBbotsPL/o6+nww3w/X0VB/nzunuqMA2eFc3Loy7i
K8DuhZh6Yo4giRh9yCt5FXY8CkXa6CudX25A+mrynrKM9BAmEb1LsDAhRPq0ylZdU4oS/Yb313wJ
UhPU8nFqCYRf2FNvvPkfI6yz5mmSSV1iNUL+yXIHIZqrjs2Qrz9ABIOUkIjawuz3DahP+cVhjvPK
hT3goYajGWQJDwLAIDy+gSPWPacl+rHaDXEeSzxxIfp1v3Wk2W/4SQ4DgPsE0CF/cynDDvp50KjN
6yb2rgsRwHvELcfh8ZbPZ47P7jXNe+isMopu/zc5SoK1Nep23CwcVxe9gh+fwWPjFlmXugZh6Mg0
6kxvy7OOIt0IS8Z33+ZKHB3o9Oc7i43E5nZlBH1xlkeMtaVp63Yzkb8Ii18gEPY4c3HjCD1qgn4p
LSbZhaUwl8lR6/Yms+ypIbZvZXZdB5Py95g/5OJxgW/iBRTpCoSdZC1dBX/rm+kZGMe0UWbgqygg
T8t2D1PGO+OgIZ+MUcj4NGgS49NHc1rPsRjTTOOyW+Qm4kh9R2GAchOB1aE09LV8Yxl/ZS1H+P/V
DqI31bEro81yciqTqMmyAuPMnHYVM9jUOwMVwLs1DVQUHv9Gno9YtrhCmAb/ogfh7Y7uKsqFsbo6
vdgjc/9m9O+J7y/nG11Dfba88UUrMibsS1aHGIzyoVtJwhtTm0Fi50nF8o+fPzcwbutxfN2bGXnn
MWRHSAGl/q469gdaJALuxzH/txtlI4rxFsgZpxTWZeTk+dItNpKPXjMQJPlkbCemv75dsJ6Pv+uT
O/mnBvl2wzlJWNHC723G9QOXnMu9REyj26PcwJaMVZAHAkDXir430Xd7eaJsj1lFH0LOCZjZaJe3
QPn+l9Vo8Q+huMklkxTzjHG76B1zlHByLX7qpHgDxYT6Cf47/M+ig2eyfs0zAy+rD92zXpO5OJJP
5GkbDnh/FMN0Uj3uItx01J35nyyyM+Kcl1cv2CKfEKh6wanDeWpVBUKkx7p5BSOIszAaTeWsoq6g
4EbqKNWPD0GGrr7SypOkq+udUummbo/yH8nTtf1E7EqM+jQB2gdwyuwFSSApSv3/3EhFUGOSGMWJ
hpsCLbew7QihoX1z286T9t4YOWRWJ/vKObG23AOHQ3RSOYtZmQ6Jq9wffPwiAihS7Yv7/ix2iBGu
/GQI5xT8WoMZcJ3LIET+E5pJGYxwrpzKKAxR9Tuq0GENNMqm0Af3qzVojTzmjl9VJQSz+QetgoIh
fZNxopy0Wa0HITf0ypvf2MPYgSsbx44DPKqfVgoXfDdmPii1e5Xjz+Yy6kvOtHg9auzomRpeny+N
oamReqzknHkDcZ3+E0Qen/Z7M8/ChDIh8tF1C2FHdBBs/ii5uVlItjUkpdpsSbBkrv7B5WJTkF5L
k/t1q/zq5K7e/K1Pl8/j/DAUji7m8TxA7LvpyTAbGuE+isYt2gIDUGvE5uXynWuurA8fkX3XpJv7
zdeSDJ8KtNL0M5j7Md5NlcGClPhWPILFQBmz9qeBfdAyCS+B4LtjEf79wycSJoZG4SfqwjqijiRF
JC7gOb0PpHzHX0EVxkgzSf9Mz1yNzNkHmnlZLeVB8ZSpQ4U9hle0ZtFUWrxed01usuaTrohwrw2N
BOKwyUw9n0QBYP6phnXNqMUm2eNJYIo26oya7I3YE9MuEkCeB9sa9isdMlWPKVoB6aRcR/rkmj6W
b1VvBgFxyjuGB70M4QnmXjuKxjSKjNVZP9LktiJahODGuyNfXPN6T6QA6I90Qv+CTn7dGyOp2MPe
nWoblvW2mPwWsBrr7I8CUAM1fV2tMDmE4oyl9ZKUlD0a2jitxo3ZadZZTbrCj77oh6a1vjXVGLkI
E3pSN08o5s9FgQtcc6lzS1Yc3gcyp1RpnvA3VL0RHjvArY66pnl4Lmhn7cFBDf5c3bUjHo77oiLy
d+8gdGnfpmXHFSmOx/FXhSOidwcJkFmPuT5+vpzx+zr98O4wV8+bJ6Y0Mjuj38lfmfeE/Poc1EBI
6meAFFsf7I595EGZgM9ZKq8TLbn79Are7HWaMLPpZqM9RfnFVNXPCkQVWQ4u3+teXUjroiO8H5Ly
2WLi75njsjz+xR20NKioBupgImDhzgfutEwoknRpNW4OWPA5oP8SOQ3+kSlxAJqYQVONul97Kygt
V7L8K5tFyLpMo1IJCIS6/LCb3hieTtirfQ/Dl0TNKL1hC0r0r9f4ID1D9+/lMOVoWlip9EjZBaoS
L3I8ptY3RADW8riEuKpzEduIQuMqXSRqb5uZ4uL4/9wXE+L6sNo10ADSR+BtSUHhljV6WYbN4GMg
at8WggHTadiOQO3eowAUJlvcRyCaNoVgd01s/zX7yfav1tURLzHNVoslz0j3wowmkv08c/fb35Mm
kB/mId0brMECe+WML9C/gB7CxKThjedq/HukmMJmDGaWAFpdCVMec70gZ54SHMU9YaWdICkQv3eQ
gl9NCB7zlXf64GhZsf8O20VQ1BUvV79pkGlUzC4E6D4tdnyYiHD9UxL+hHIACYlO/kojBgpMkCSh
uvw9AQ8OthhTYF/0a20lBC+GY3NZP9lYHR0xMokXI4cf7M0PJ4HxlGJRnAaT/ezoqOz7IZB0I9Eh
xav8m+HNlo8ZaMZBdgrdVwzEcEAHpZQ0sEBsDfHwd2RMSLqxmeRaYFaOonALsj2WV7458bkivktF
fJGB3jPoEpo5W1oc1+r1qce+lEw/4GL5mRWCbQ0HYy12v7oQZ+Y2CTZqo2rfSr3yVb8s0y114IyD
zQo6lbQhBpnFHsSiMraJRhMHDIlktG7Sr4hvlKEAGAuBsNwi4XCVYW5xQeC/md4iBBsK71jiPqGQ
4iTVEhX4EdoTqe41txQv0OSdnjc5gEU2YC6hSSyBIgvR53OpijeXBpFTADDSvnSRhPx9vTTyhWk4
oVxy+ME4pbPrQtda0blwzXt0WWSvFWS35HR+Rxm49MFZNH8hNWzBzy7Mw5bYVBsbXdE4oqsjmf5e
p4EQVNzbUjL3vm4EFvdUr42mTgkbW9na0qfqX4ja5I6W/sBCEdOhq50JZVQCatbYaLdLD5rRQBxR
Q5aejf8VsGBoqfqRVw5kFgPfSlZRwKg/YUgrYmebYXnnff15DCuBeNbqiMTlsPayZb4F1sEWQA3X
miw9ojNF0I6dEJuFhThBNmgHGG0ZLKq1bGFu/cHEoCaZiPkCbIElVh2MFAqcyhdWaIrbV7/DWm8f
zZHeTK+U4m+bNRH5EGHv3HxR1tAiK4s+IsvQ0JM6Oztrl8VOplhRTjDHJS6jitj23eng0uaagfy6
nBqrTSzVn5h8+CBlazmQqS41clT4uzsiVYQ7gjhUbjmR8xqkKRSneeF5DGNWMS4ZOTX8YCwcTlfM
3ypR1Q9dr/oa1lCQfp0UpAK4Ms4sDIPwtPawnHHMKdwI+1PgkQRg4Qro6oUdwhuZbXpS+0HLYl2G
piLBQKdb3Hcd7F2+xjWStFF7SgPut29rY3eqHWBEBalx6KDomTA7HU0S3P6x89fcr5uS+l8HYOfs
68/XG0+kibWGerogHifUV+4RiKSTE8vq7khaUn4wXfv778shJKIgEQ6EX8B2OLMwj8oYonKL4niO
auRjZtNZGYIkacGhkLgAqJvqZWwXw2qF/T1onsnQUP4MVeR194dqMeIG6OgAEp0JufMYQ7CKsm+S
Tw9cpLbg2cISR+gVJiS90N3VuhcvvC1eWIRbgSbNQ2LmKUT7B7kX3bGwg6rVEIQmWeXeoz7FPbS7
pbzVY5gEwZlPF4CkMJQdg2yUXSgxe8HB7rSKWenpcoiisBwNV0af1QbqsDHxm6PzXLRvGYpjSXDL
TbTeXTBSY1effIC1kkqIt36CARqd6XZ7ODDmFSBDT9tEsWTPVmGMTE5yTtD1zy8Q+ItEA8mXluTk
TbL9exyjD3xiaDR1duz3SMOxzlCqYKlwWqqeOmp/uoWMFdDPl9yUZyzji0JqtGiSiyU69fMzYU1C
+kVqU6rbJhQMXRqOMrLC6BTm0GrVtFDpaYGAYK143sab9V+i58GW5aABxToO93EwrgGy2YQmFJdk
L4kGoHIp6NC/7Vy4KvodpREZH7SwUHRXHP7S5iu+XW6mqFqiFpSCITWHqbDBbSehgPmPCfnz41Xq
bWTRnGAcROPKESpZUjPkDIaeJGvcz5wU6bm2nEC+L6qfn3timmHcxTv1uDM6MHx7NmWFyaWiwDzV
jk+LD+bnhQpLZu0MkPEmFu8jwo9WqG2TXoNKyhJ+6+V+/mBai1aL4tjsdw912QvC7l7sJzykNRqj
Vg0JpVko0LUf1dy35vMCJgu4EpI4oZWmarAjptgYJ8t+kNNAj0ShtWLpIjV4pMVvSAQ6VbjNM598
yOvIJnAwDkfM6XXMWANWSRbG8PclzvfE8zbV/FwaTezoyEpUNFXCk5UNnRp2zzI3m0nHsnzjnDlL
llVFBL32liLDnzz7Wqd9YyvsluYs/bqkNjIc8dvTJjUUmao9/qAcxILMbyVb2oL0tH659DoTHNxj
o54U+NXEiSw9CXuAUW7QDpe481JCjsDkOaj5OU62sHEvPN5Dol9vVlWDNUT8Kj63gHP+rurrwKcA
yTwIsVdc2sr4EqakTaPYS2b59kYCTsMsncKALS1FzBD4PCkDUpVqjDWDDv/5XfdaZRODHl7ofkEr
uVwVjddQppPltFqLq28GRX3NfVgP26LdxX7djHH2a3/vMLy/vqsgHy15tdVeQeOF5LOyKbrDBXwa
pqxQEWS+ugBTY42RPvbOotReM8V4YDKS00A/KdXHtWhTlFQed249KngF/wrRei1XAovSnR6Vpklq
L2P+XHtnkNjmNNEHvSlWul/QFLdarOdsPEga0VAJYfM2oeQzo/YNFcfutSGC7cSesWnZI0AJWNes
kmKJEs/lsavehZSVAg8ZCWAkgdCvfga8AwLta7ZDOhavavKTD4CGSk2EjxjifX25RJgpCiTOLQLc
1so8cEJwwIBNbm+eY8Yq6lELQCARGb9wB7pnjmyCxLD9rcFHOXcfStQyIu1nC6BYxgD6CrDyZ3or
kpscSvro1tLRQzqjznUEpIQy+55yK03/INWU8j+Iu76oRDk19/9CNiLzX86bvuLxPMwTr+5jlBYu
S8Mmg9Gi8N+dttw2Ws0SF7HWA0zpNKGFCJUDNs8VTXtMF5ikNuJ9e5tr0wuBAK7cP3K30NY6bXjJ
SyUu/KrWnT9dtLcZxqgeZgB46cTGyYkFWKN0w9m7xg0gKySKywDR1b4Xb1lQgqNoxJ7M7W/yBmGS
JZ0MKJ0E8YvRfMmyrgPnFSK4mxLFrloKsPGlv3imtUUlaD4URm9N2CFxbBeGf9fe04CNyDIVW9dZ
qTPFtN8+WgPCHOIU4Noxr9cnnNZ40xIK9lRjqRR3odw2lySHJIfyaQG92FFoybrjfD6uQ8TyZUME
b+Q2I49vMywCf9vFjISYsAZLneQd12+zGtlu7vKSSx+wNsGoBrVUB8BQqvq6Y2dQIZEBp3ef30/o
GPOXhvIQxGs1N5f5TjTN5HDdTumX7vMxJzoLFQ9/1Z/J/8U8t/gfA9ocPfhgHAepBtiGuE4ASe+/
sAQYUba1/7fMNh22is+W8JH2CroWNDaRseBLT64kyjMISnLC7rWfr6PrpdtPhJvORVKT14GPrebn
aKXprn1RlstKSIw8soVf87AuYjHmLku/a0DRnV+0Q5MBtctE6F3RbG+0337pxHJ9ljjE3gugzAYB
w6LTULapyK+3BPV3g/NlUNW+eVe3yCxvmNEcpMq+5R2TJjqKasJ1cfuEXWIvmYwRuabGHbIJz7NF
bKGg93uOEbZOJGtK2DXBX1AUbftBHLuwlS4umLmM1cFhyFPOG53rWeTf8dosZnlAd0r5Te8wwgSp
3gdYofG4U+pVtHTKwJkQHt+3YOwpt7WoGtanAOlmdSa2db0H0hJM8WcnVn/hoNe1oFoEm0Tr9nwf
fdFQ+AAiPueFQ3OFjLvRQgaXplSh1NqgWlYeXx4qyJvIpqAP9iH4NssrugFaEqx9p0pJ8hZ0ot8E
3x9tYS3/ORzJFhYzr8Dev7JQ//nLR31R2EiP8Ogin8BIMGbv3kyeHKyYpn+MBrspal/KQprao1Fl
IH37vBeOIEHp9/U2h1OVwW7xwgDele1XcSvZ2J5WOjLs7gEVLJmMLtj/08La2HW7J6lE9x5Bsm1A
E6qiMPSoRQklEaig7D6rXM1sZira/bkJYu6/tfqfvAWXb2h8wvbSRYM1IE/sn3f1cogDK5oiGoaD
C2smtQ1SqP1tEeJK0ouowWBII7R1FgRHCq9DsEzvCdlPIzgt1a/1YdBgpCDV07TqBrclIQi1GyIx
XNjyo0xTIWjDhbCCvMrOQPn/Nfk5ATA7Eir++9gu+0Zm+A43HieVxUk+LfTCRRlMKjts9zLCd706
WJif1WEzA5lve5U9fwVhAc41EMVcpIFc8E4V8xn/fgQo6GkNRXn8aakQUyb18c3Oxf8vASlCvxUo
QMvo3VFpSuWS2+Z0eF1eGJOYCa2yGdEdGno9HyQSQ/gqtW7n+MPfUX0zjWk4Wr3atWWyNfD1m166
F8M4/f43SLD6X5HHyQGkxDi+5aTik/AzegDMIPWSbvy9YD3Owup0bpSKM1k8gX5jWS6dFZhBvQzA
PoZD94ZAIcIv3Q8j7kz0KMAgXDsYKBbyOzO++8ggCUCbVYljV4yL/ffMicXJCYXcZEAZxXo5hu0t
MkwCFPBMYug5Sch4ULyPOiUxz55GtJEfkGzl1A5ZP3MLHO37MovwSaXu0WnqTcunqSvydkk0h0D3
q/pPF+jA0UwpptJAD0WIJNbYd9cUuER2eceyVb8ZYXud84KoBWJjJVAgXJLTfzoFS/nqSxlbYe7I
3NM6Utx7rwR/bU1dm4M+wKkN/WAYT5B6VBcNBwpIsz5PlaqqPv+fhTm10JAf4/m1YcOD1dfIZ6XE
D/1DN2O0Z6JfbnBhvCIalDPtSqqSgpIBtzWuzsXDMhNOhV1BwnL0fztOt8GhMoJMfB8+NuDng2bq
i/Vr/mLdA9NQuXNa5oQPHIbaLdJbD4S4s063FdRBhPAW/webedc93qqngEKVDmMNbmsDRmSi0VnH
BjQTm2aKScj3UkERvIVKfUDv6n9TINgzD7Wp9RSV+s6W77NmZxBpQ8LwPao99qGyYvxeinmGc1or
hCw9/5aq3xXDyfbp2FOzGfZPEGHOAKVRLU6SQXO3vNuMH3OwgzlS53/XGngUmsX2m2UTNDr29cTE
jbaev4tyK4k705x7zDQM/xv7sqVbgE2Zoh+ycipYd09aBm9KQC9ZqmR7umkLmyjEFJIKXTjdSwQ5
NRBkYPNgkKPERtSmQOR/PuIjtCdmgYGbSmJMKvImJeH4nUN3VNO9DYUy/utYLRzqa0iiadQoSxvD
Fw1MYf7S4mjTazRneHDI61xl+katyDHUoARiVGH+0i+HAFEmcKXJ954VWCcZUdaORgc2F+4sbz/w
+hQUPgBWAWQpY/EVXAGi30181GbonI3jpgls2TU2W9rfM8xuiUqZ7mruFQhqXRsp1AHe0099NVmw
jcd3ie2Mi45wdzg5MYZLH3TfmCo92sA2+XnO6drGX6ZLt97MTTdSbebjely+O9QKU4WsNCKJzYY5
wEEGV7MnYjnJdQyXJlJXSrUffzPiWBYhRgVaw77rIdChfdSFQVycp59zQAS3DHcukFIdPmfLBsxL
AEpzE5ImClNxk1aoaAY22edbikmO8Ssr+j3tupGXUuahOpkN+nkIUAIlyRk9WwBDQZBs4pWzw87g
MNQwk7avp8M39/YuUrtst910OrPjktACdLCoQlBZVNL0sKpL8qb3C+UUgVMW1Zlf1tbXv0KZxd1X
EV+NLvZUdtqxbmVNgQwbtYlmBKxMc5jQ8Xz0gWvfTFrPl+GbhhZU1uBQyOTumi+zh3llazdahuBN
jamN+Gw3esr+h/654evXx317XZafXQkxH3JD4P8Cr69khyFtwEt87JyAzwpvT01Ay1ph50IRRB1Z
EFaeuB1G78A17GLALKC9iUy+Z4QjuNFVQ1s9ZH1D4hSPDIdkdNcueG0w7HHqmVURYzr50kGw7ohD
SL58xA9rj9N8f1oPXvC8hxXWctlrG6HQOom/o5GqRvcyvw0UFwG6jLHVz4HK++8qOxdEwz8iUO/u
2lgEMno3nCUB3j/IzQxyegfG8Vs8RoAlmFt7ALl6qgJ65X+2904MyBNR7T7XcGs1Dd8yW+h/2XaZ
ySsXqiVvwYGN8YocLUfJkCAn+0Gb33K1zxImNlx95DCakurqHeGwc6UFXNYT2iBFz9v/VWBG6dnV
HJ+LboZ10wfm+qmeM3VqXJs7cMCABVf7KBMAKrp4Go0vVSXiEJG3S9hi5BUmnNmb0pssNkQhz4oj
yGOWis5HoCRO7SO/e172+RjP+qpX3xV24BiZhqHI6o4okMb1kK/N4JAc+Q/FamABxFp+Xz9u8xeb
JbBHpBjyKSEftiNI1goovwdGcTaCcDLeb6Bi2W90tPT8eC3nQm+XfAI1FZ4JT1NJbQKzU+AkfVPz
ZwohP06cJU2W4ZuAQHcxVqajHRt1OocXaREXTFydMim7SUfb6nk3xiSlKLcCYMVLnM05V4QuCo2u
S+P0rV/LX0Ijc3gJ9J2f74WEf9i//xi4/Sm0ibmQL3ZzOpqoztxwHvuIc4vbrgrh8lC6x55PVuga
YrR80hUMLdLqTy9C0G5oflKgZodUqj2O359LQesES4TBYJl117LKTpJqAhfj9U/Vn5BNgzLCIk+C
AXP8JReHGmr7cjEmWzh/F6YYlGYpGxJjpPqi5G7FtAEUvUcpE3+61jvdjY2/8LXP8u4o7dItjIfI
udLQGm+GvKpMLybMTK9DxVAOmwSVXhSV/hzVNSt7RBGRDzAUcdgWCT4twQZdN1WZCOYbAOvCBlk8
EGuF8IBXVzueLE+O1yOq16oZ1VTBhGB76bAgvpjoTw7Dv4g3RXfseVUiYYHd1dt68BAVU4xVXmw5
AsHzCzSOOkQ7PdDka/vpbQPgyKDGzx0GqBGVERTyXPBjCILDebhN9xbg8krLa1gNAxDiYCLdHWOv
ZLdvSloVN15+nXEU+qVCfz0LoR9jiwQfk8b/fnQispsUUwXLIaCeo3tq5Y86ls6Kg7XIiddZrCkz
omAzRd702PjQ/5JO1hvRp3dA+ZgAImA38E0CsIbLJvi1VSrZhdaPM9lMUvCVEqDECkhLkhUPzViH
pTKBA/YQwKWc0+dDIkO1vBop6UGLsz8osxrGj5mUsdh6XYeRz1PoYEltZnq7+uEfSXCB8VibPg/q
lEyUHSxhQXd9Ykc370ppNTuGTNFKKTJ9wwSDwO0TqtBT02Q/n/S9/OTOzyLWyJsBlo/6VkbXG7Nx
6UYHgoOe9f+DvT/XtinsEe6lVlF5NIGCG26jeMcB1tK1F0FBg/4mdnyQaMZgGJNkPJJUYrshQuQu
HaoNGhDGwbhVIGWYAqjGlLmg3WpQrRf0Mir7sonIkDk+ut81I1hSfJQ9USKp7WtCG4JBBHM5mKKy
lzrnyM9NTe1wY3mHlBZ/OBjoZdMr+ftwL80CuMgBVey38i7poQ2C3JRC74BE8C+NKSy9XIS9Rni5
FVP1TWaxgPM+b3FrGLZRcY76pZJTQItVIE6bEh/fx63b6GTtDiMw83BaVEB8hiIio+MDzv3QXG1g
00Ie3vih3qkmFZ4wgrlQgoR+PRfg0nxEY/HuMzr3XCHnm680JKYZQREjzhyMJjQgVJqmAVE6YQXN
PUOuJtOEjii8aPabHrCO93/v12G1tb3Qn1G+OxU52Gz5X6cPft5gHgLpeIOze1YyI3+iOIH4ej2W
joBurFkYtpJJXNME5ZMA3c1hZVanRtcP7GlRqtJpw7VeP4PnpQZFZ9hrjdPPoxzgD3k+bzNOlBfv
BQbcxyY5Wg6MrmHOKQMQSrAVVK1KAYGOKVExkQzqN5gPKMythUqshXim59dncnZegdwTEzjN4WWH
gAYBCEd6HNWxN+WgasOo9CTVlDD6f4sn+dSJxYrgMwSa+cf/M8S0ClrE1P02txObfD8sH6PoL70f
1bID8va33GQ2t76CQqf+dzGpMrqhhuuCrGHASDnXQI/5lNzvxl9s3kupW8DMshhncCdDUE1L56Fa
q5viNsopI55jabxTkI3rPTMSGEQ26BHbdci/o6lDbjDGsiSFAUtdRrgVtWqezmtZewWRSf4GVg72
w75HvrJoi1RmdXiW6Zd0Uqh/8mPnkK1Gl8rRJ/lH+dIzvmMhm8i4IinnkBjcnYlBAk6Twz6UWsid
rkkIaDfyW2MsWgMs96fH3mEHN67vwLT4S5D4SIFD8/df5LPC6e7OZrfogvrMckANGHy+te/l5DN0
/D+WNEmv178lwOr4FmJVht24J/vNrQhz8Sjh2Tv6+9IdOVurlLq1Jx+awGEzAw2m2PRm/UEsM2PG
hX4iawe1Phi0Ag7VF9HSKwlPlX+K3b9QQQHMRp/4BLRF/9Vyi0S/WJA44JQokrXPBPIx361tZUnf
CxIj5un2vltgD8/FA0dk4fgoj0RxUJnmc1Fy7NKPWJMiZTakR9R8qW/zf9SOZ8lVV6zWgrbVUVml
I0A82rOpN4hp7T8oKLd2icMxDHKhHgfoENTxLHwcVBYamEP0WZilkvaz1IQAvgzFWsEAvlqnCRPI
f2/AfOCmzcHF9/Tdzd9K2SvmIuay2jCWMTBxpTr4M3vx+oXPnrNWeELM1xFjqIpt+dCYx3mR9KmS
T2sL8f57WcJI+8k36GTB111dlQyZr2U1rAkM0Taj1rGUMSpYwk3wco2aKBXZEFqWDlEsdyueWNsS
sZqSy1F/N0P4GjLmjBaHJGGSR+RzbuiXpEKC1gqL787IIutbRdrpKAa8hiyHcKZJapDD3dyTpV/Q
EBSMbSQjzWoMv2YrV+4DracDHPj3HAVtPNdfOM3RRO2qctmDzitRwvapprCf6gn56OmEz/wZif7u
SKTVw2tIb9TFOZ2e94Owsu5y8gDLJvz71HrGgVeMujkt5S7AqmX7Odcgix0PirIGZnM3YJMkJMAP
3D9K9ihpCEPqF9RBvJuoc6AojPx9K8Z912Srr9PvGnHVDUQlHoQjABi7+eQOveiJvK0j4LhqG7Ap
X1P65jNx6zyJbC2sL/q87U8/Sy8FmuOMlWx9TAE392ZfkAjgItqyfuF9VXJXuqRx1oOCqj7hy4R6
hTKrQBnh0jaIqEiWQHPDl2Dgib78MsY0Dvo2Sw7EGYvupp9sRq0LjAZ/juqAjdFxAOpC7eADzj1F
xDMrN+MrI51bG+vFLtX6FEVzzY9ZyYmA/8zENEbMQK63RU/TW9wQAm1LcWVLmVxlCUie/4sBVchP
RSzfiUQ3/ztS5w4zSfVgPNf1LoC1qRsN2+AMYKVllpk2GGjYfkRkYTW+CxtAHq3wjW/CjoADbBWQ
AyUIlhh3fvlMUQf7WAGsLZojy6F4NM5DXWZu7ymNcPI+rg/mEI+7eviVPT1Z6Q3MAxJCtMIK6ycf
7eCrDv2RmALB2Pb3BbREy/lZNzkSr0ly6DgdrVap6D/N7rQzemEKvOg2skf/Yrkdw7dabi33zkIz
v3cHO6nbcmAarFuuQEzgAvCm0wVlLv4eUSMocfveFAXLmaH1gGSf6jDrjrs8aBldnTOi+ZGfGgTR
81wpUVA0IfLjF73KSiQGkZoPw/6FVHo8nuPKXuoR6b5ip3fif9711xm9V9oEp1lG2GwHuleHpnZE
pbPzZ6lLh04TkbSOmrzpDHQRqJfb1oDGpIw3E0b9NSzd+M+MHocpq43HPuxpNndZYM23pF38TJQD
r8Vo49bxuWeDOmLjRzZUHhpG4BUSuZXpSnd54OB2F3oRCXPvPbOzpNgu3GcsANB27/K1YgTdGs+W
8asoHhPyRBXcWKQRxlAHMRgBMyXn2dxKvzZO/2ZpB/UGKmWMcgbn0ZfK6NsrK9A6/b8N1iOAHw37
9vh5GtMerK2adz09+3O1xl42k3LzF6hPhOr2vvx4YyalNEOMHRArUYWEjCGB+Q5ZIN51ubSNULH4
zYd02NOR6QWPCB2hha8U++kb1+SkI3tqed4w/psWCroWX5fPu+5EUN4pek22+OlcwXCInvS/G284
AhdKZZJFPkuHq4lvX+pKyH7UTCvvGDnWAZTW+07otq0APRJYYp8HSN76WP9Yw0wNFFHH40nkCme8
8N9WUkfWWbqFJEXJDXtsL2Kz/WEqnTyfMDRNgW9MXnxMEGe6JHGLeZfNlz8uBlUWjnCHxRktEeQ7
8ifMZ/B0cQwtzfO5OjNtQwr51pQYg/q+BOj8cH09q027++yXeYHSyRl6jFKacb0LudsPV6Ty5M+P
imlMy2YzQ7VJbu7I/Me6bCGtd80iYKASURLRLYzjDPvkz6ZwBXzRDH85AoptqYcd30HbfJ38mhL7
/CkEuCoGAh4eEESpXxyHGkILU7oFfq1TJBIu8ceu5ct2C9BQ4nYwGZEKHw+jshN4Z4DrEFfrGxmN
bpDOS4Iaa+GBIvh+DLbYkU88HSorcBvMXptOo4HJ2G/vApa9REkujPBlzt7y/W01UjemSgGanjgd
krxBA4HGnkxCbr5n+0x8NdZ3GZSXQUcKkPezuiRspkju71r5H7mHnsgCXl9+vlcYEtTyYFdJ9GZ1
wsqFHmosJSyJIbqeBTGTzgH80Ko83NJMjpTPk0V9RH/rFauaffeamk2ug5c58UG8P0eSZ7kpl4Sf
eRGq/2dS/Oq4fOAhach67fKkOJwAL0wZEAn3J4t3splt6cnn9ivvrWxkPS7m4K8zIRJq0Y1men31
YilqdhiUSHnFy834fgt118Aehxl8mzrKbKv2M+KVyYDXyI38fabNhveS5xrOZvjL33Sd3o/wFBoc
+lZPT92yjuwZnfnylL3Kd4rfiSOkonLCGpaTf9vB/z1pUPEUp9AuwO4+Xw4dSoww62Ljvnvuk1tw
Z89v2ISaNwXgyRf6gUnVysN/tUljKwTTBLjhSh/CChTYuEOhj6Rh2GwRc5l7MFjYc3hckHcxTB5o
aPq5zFzzroO4shh0yMNKklMf4V5nMioW5zNsGXwZnWRPxfS5jsDtXawr8mTIcS2HluRqJsARk+wp
EGNwS+8NzSkiH/IM5DDEFWrK6GfVQS6N2t+CLmta6Lv2z/203W7AxhhWnfhXHIhQ3EmsTRCvSt6+
c68qr/uMibVtihPXTuBLgnj41CnwKkzk8wOPCB0MFsC4/B+u3O9+wdLBoBgnJGRMp1Qz92/JvP3h
6qgRmbFWd4w8CFzegA9tlEjDsl9t/QkZUdK+kQMKb23eq0YFSDEBQcn38PIgxWy6jad5xuGKyBNn
HMKvJGgrDx+Vxw4Lxhm1lV5GnxpLNk2Tvx6EshVOO9hWWJI3OL0K0uIAhywKn8c+r454TWM13c9Y
igTBQZ3ODfS37THSW5Czmh7q8Gr6yGsOGRil1mzjSjZa1kjGUok6E+n3dky7j8D3FZoQdlqsURQz
Ke3R6flqGhsXwDa7gLLAzb50G/WMyVi5XJLomYGjD395TT7oMm3SSylUcAsSG2N7Eyhknc3hZPJ+
316DW+B25s48g+risQJsD5r4cyGXZXWPmWaliywAEtNurFp2pULK+yiX/sSAl0Zs4ZdSFlYBQ863
MZmlwwJlLtlS6r0XOvAHAaQj+aK+fIf4a7IMhOP0oVE1uZ1DD/K0xQEiuQlzLeqGB7ZR65JVpIuV
5fcY7pD31C5tapu2sNYqAWFhfH6jQRAKuQ+iZbpxBERBbIHgU0jDnqoCfMzcWMxn5mj9HOIKAtBG
XTvLpDhoSGsroTK3MhHtd/0BcQbcmD/0Jl4zX0169q0D2WoOi/F7XI6V34a4efakSod3rTk7b1RT
9jTmwdiFPNQa8LexnlZQb6podEJGZF9B1yUzFvtM2N5XRYGDFfnnGwWGEO/miXtFMnCGJToHTI6S
CcvQzmIf4IOVEpIz0yNTMK5GCFBOu9lQt8oPCQ930It00BUOCVUKC4cNwvuhiKh51jwHQJpcV90k
+FkKNjSdUeNBMIPddzb5bvpnTKqM/qhgDTgN+946OnNOqnOgRVCK6QOmea303EXkB257Z6RdR9ZB
KU8TWemhOEqULK3oFoPypQ5jfVoc7NsMuF9w3ccaomtJSEU0gZaRRfZb6azlOQu4dsVTz5VInMxb
JwxtlG70j4DaBIpy5vFqI5DXn5BE0hDP1oerKBr/wG9fP61DMwc4YwkXDLLqsdaF/ubd1WfWh8zg
G5ApSIKABLz2jnJlXTMB2pS5fH7nDcsrg2ybUJhpmPSlItr7wgiP6zoCGTzEtCfSjGj8N73IwDMW
G2YwIYC+kX/pNNZmQkRk4pwX8VFcilXtgD+KVB9s0ydaMWduMJxajYfhv+B2vXFj4qq/7AhwU4A9
q8U8W83R35t3UdyabfowYiLuc3C8k6ko8xz+msU9k/9mCRvlnUya5A5lvF2bKb52p0VzT3W8r4BK
GiY+Q7xb+r8B60beWUMwViUJbYSJG5kuTFtOCltqAKvy0+XpZDrMbbQy2hw8n3rLSSvWK17Hw2/X
NiEl7N+wP1ktsZ52QDEbNV8mOCfIKFu3YYYlb5AkiyHKlSJgGK5h7/iA25thHY8zt58bRvbursSG
YecAN4Yvil49Kj+QU5yhGmiShk91n7q9N5iJKGYqQB0cFZFkcxhHR5IbmPlzke1xnwicLGuUyU8+
g8/0Cdu5CPDuglFhpTGv1bXl8q3BHv6niwlIqZP/LukDdEi3pF6SlywREK9j5cJg+puUX0luskLS
iKudwSBp9eGckfwY9U21ybJXniHyYkuNt2XagccvP81kUOvrxFvnb0W1I+E1s4Q0AdA/cfRHjvW8
ZqJ+Qg42chn3A3zOsVeg8esxzWNIRyj38ukgkWl7XZWFH1GTgLytxehxvDZ1EBnw8IenpLX/Toew
FyvKh6y+f09toemvTzYDoShcvAB+Y2O3Pqic3xeGJxW8at9ESJRqk8yarFx4obM5t37J3yAjLrr9
I/jdIKhu9GQNtNwQlrURpm10FZAyFKmaWgrB+pis04l4v2abtMWRtbzqZnEFByXldxk5aF3LvdV8
g0nMX+/nmBUZI2nJmPwdEJ+RwVWWZs6+pc3dYZfISCN94DX88or9Lg25+/UPjDkg1Br/CLOqMCZX
/fAGEftkCdSXrtpiwtC+lQDjP5bcKHdRK6Bu1IV3mADr5OJfvDd7k27qs6YWYUFaxp/dU8fEdK/V
52DaprT8m+gkUE8uTtN+Vr/q2qA5w4ssB9v8cfy93Edgh9Zk58QdQnOllcZio1Z1VizUzK0TZDCe
iKVfEt6Jf5FPSK+s4NvPVD1p6Vhip3up4R9YGT1Qaslr+tThyXix0tacDDm2jfh2Rl2QuWugD6tx
1eRRaNww9Mf9b/bJ7f5Uw4JBxvScHpqZPJZD7ojZHUEUZFiFco0uFwSnIAo5WGzAkBKMEGeP9XKv
B2E0tzss4jI626luYaBxVISgDr9X/q3Dps0e1uivqB1maUAaWqKzqWEF4IZnBFCO/gcwI8K73su7
3L4GjlThqandu+uBmwH+/I3O/PndvC++HSUiG9Tz4xSDlM/ZEwgH3+bpS2YVcKSRNo/c+2j9FCR/
xLvu22hZWuzsTZbeJnDxC5P/lUHhe8mixBaLftF5/zwtsJ52Kxpt6jy1coZhWXbiViphePCx+sKz
9ABaiJbjXb2CNNgkq960YuVO8WYUfph29UqHQYmvjpaJHzFE1Dy3NXPJmBhtCSTl4nFwoDst/4n6
9YJ2GSo+zG/+JNF5CnrGKPbIk6LaVzSv0UApZn/2/4xtMIQASyp+DVC/HAzQitH7LlZkuYopIJVO
K+ixxAaTHU1WhFAnooh43Nc3N/rBCW9rJMBwEgDWgb9mGcjKXVmXNF95mCxSUZwE0aAhm1jAoyx4
hzvqH3MzWRCUo9XDbpuqGD0eFY9f+IZ8ygepGs5jb7j/c+MK/3nQnOU5tAJ1BCYs6Y6t16akfCaX
C/8cK4EsAm16OI3+J1VM3984tprUNfdV5cOHAZ2yAkftt/FFVC09Z0vjb0ZPxKrzo4zArqwrZsLt
GbYjuWqyi5qq60hAgXzeQ2ZK81IWNs/jphjMBWbJiOmsf3a2mbf0Rjraova5Rv/s2pICKq0z2pBO
PXicMOLfnZPP/AMi9LdH3H8O8s0PIxLLH3nxM/t3PcPClU4fj4qGYfpX0cAcm9lx/c/raYrehIO+
83zN3uJ+tARc6zF8r2nWbx5i2Lw1i2KZ7gT+qoo+zLyMA9E9u5+xcBEuwopgp94b2rcMaLOoD34r
H5ercW9SR06qPZPIE8KQTgah45LE6ADGuD9Z6aV6E641RGK5sPJ+WAhpJdzKNt60bqt0IbHlyjzJ
xgn1W0TDNrfy5iWmIi1tZ32EbK+lhVsQYc9R8D5rHWwFLPcmACmmF+7D9S0JPOIb5e7BMdqbJ3Zz
BsnYjSIrdU+9qZbcOigt8LCWhrpYJ1gE/Yuqm5sJrSTQIf/MY3wVMpiC2u2LhCRsm/UWpuSjaJOH
YsmimDxhHE71BMkDSpgtDwlBXfT4AyEXnd66+kKp5zabTX3yoeqLvXpIyncJE1dKT9bv3kSoYPsH
GjvDVn9qmqlpB2tU8ltEf9tqFAWIQKlNSz01fytbkPlqT4VbD1SNSpK0STpsw/QOgUoEsEloW9xZ
89BRN6Kl6AGPBoyWn2NETb+8WpuEsbkmEn72VMnfypfMp0J1Us+JyO7golGnrA3MHvhS8icT+iue
C/2nEWAy22x8dQIxZ/tFGEIFocbqFg8pymqApdZuRX1UE2HMvxQhjd65wqiXQp7orwSlAUlVGUFS
eaDo/fRX94Dlvns6t5SXQRH2lGnHT2uQcwO7rRVkGPbjda//omBkEgnB1jojbIa9JT+aEPs/1tYX
jfq6ohdW1Fi5bY+XEkvOwyezFer4vy4BjkHTClXAx8iBx30cD2cmlJW/kYqXp23q0FoqKnkHoBr0
gZcn1gh43zwAt3FjZ8GpqTtbnYh+1kDe+3xaYiGe7tWdwDyJe1yEuwgaFqc7w02zfkGJgC0GUz3Y
tsT9+sBGpsfthtPAr+FSjHr8Wja2v1V4lF9j7z6V5JC7JwTHG0W+abFu2sNtkBjsdL5aMKqgoyKA
VJ/KoHpOoUrYra2Sw6JU8uWSbfhBZnv+PAZLqHWM0+cUMhPOMBnTMXa0jIhyFMUinis4ffd2buYT
hAoD/XxCrIpbM16HDLg7L983dEC2CbxOyvpldnF7+GtZOLpWycQ/BpeAJdIBpzao1PYh8xv0uufG
MlLmD8GRUIAJViQFkuGryJo2nTzFreGdj78fdjQHkaCueMgbw6mR2aD4zgPbMGcZ5rQg5Yw3S/KG
My0FXPKCOjKSuXH2+TfAnRZzzHU6hj5M+0nrrsHIUqpNpiKAW7Og2bxZSwV1MkWBHeCpJSMZvRnU
Y8Z7X7gPK2XELWNNCuKzl+ouj7OcTMqfxGBiM3gMMw6xNj3TdPc9ClyJ0iZHvIynHO/K0lG/0Xpv
zJ+ttEgSGxRALcWpMZl63X++uz02pxEWUPJ4Tl6lHTLKa1//m+8a1kFrx9haE9JB9cb+aJAi0eny
3aqOGPXZGSXHR9ADuEkLRdXyjUMHDa6H4M9KZoiKuvZrMGzhZFNR6mghXWQbYpQU+Rh/RD7fx6de
DxVqYW3rkEX4kVzTjy+A/XbEyasXkC+Y/P+2byp4m0yunCKaJV1A0SUA1RAYPg1OggHeWty/iLaY
hQk9awnbYv2hXAGC9nmvzUgEpfsZV9yWgw6dtELGRMvSgvGhpANncEacmxVYuT3vqymCApPKDf9u
JIFfry35KPSTZWTNFVdJ855ZDMLYO3g0gCsxu5xDi+W92mcbqeem9/zOqiNiaZN8yorPpplJN44N
8XnVVJNlbubcvhNGyNthBpxTlqbmNDJBhnlYNI1cgMsIq1OxiTxM6OT4f5WKFzc44ZaPvO/fpUMA
PCp/cw5y2la8paT131DjnbBe+th6i7u4hdaWuWJCj/CWo7y/TKPhwmJDebtBZbCcAwGGZP0uH6nY
cdgXXx/WCFUpyV3hl2J+DILsSLoDEdmBybFYQsmlfd65pbqqB2JQkQipMeAYEtZZV6iP4Hm/iFoM
aeNAnBueMbpMKJwWz/3bh5K6vM60Vz2Ym4rBzY2RnjFY3qgCL2EDhWg0huGLimWmXkUJ5CYU9YBW
JxIDpHSXQV8AY/QrMCFYkgLxyXRQkCfPKIOqeCLksBOdNgSqPxAP21Lvk40vPvhQ29PhhF/bKjKD
ysKiNDiHEyG+0MiNnF8QBO6z29QtSCowTB8+vbjXPJUzj6nutXbdV13RHULD1XYxnDyRkq/MtmYh
rcMlrAiPKahrM1XlWpO7Rbfg4E+xXiFZpApWsaprzGUVdYoTYDvu+/Frwa1VQ+lfUKnegZS0PQbB
XlY2iaV9iid59FXlNXYJSzontrH4btMJwLeuAgqhrzO467sg1lKuJFThEHfHad8a4v5FWFUD3Rff
blMs8DItjAFAny3cdNDPP7Nkfz5XBF31mFJDbkOhNPKk5PMVDT5bu69b4MSymMM/Yg8zpT8v15S5
LjQVh+62fKVW4ztd2MdmLu78bz8uJU9ZfiZmsHO2Aqt1Qf5XYAdGsgBpcucOsUXxvZr0qE7cTMLe
983lk6L193yvzxnbNgSaGDH7Id1H4wn5T9fJzA1XAeYi0xtzQBaGMAYnIkEqf0rUmKre2k1MamAl
0Hty8PxFyzOUGfuYK6N6flBxUuCjpNiHV1wOtSQ8tzYVgPOCewV6o6zHEFU+rupovVSmoFkQBIqE
peI7Mbmy6PsauGgRgJgmJYXobGBFBdZ9F8hDbWsUEW7OeZzGn8VhojzBL2F8uyE5dZKuMrIqtSH+
ewKXKQxeH+S5xWPmtx17gAApxkDEi6NrMYwIPOISExvGqRCOQZxsEUJhZMoqz3reDBYf0LOO5MpR
0PWbXPKk4RmDHuKBFVUIQ8OO81JQiCRm6oHHE4TS/PNSdMTIeN6AAUBNiXyFRs64n+bcLflPH7+1
WV6mzPjkI/5q5MMioyVruGgBq1QdKqnEIFiP01JBehFUX20EA9FmzVDBgbzXX/Wbqf56qV1hwYpT
bviYwWqYg61OQTeZm8NhQmANYkwyfkrmHFkLIKoyF07IKuzjW+8w1ze8N56Ea5iKx9t+zVidA2lR
x0/PsoA3ZCHcXOSflEJ+nhbF6YeY9YCIkyVzvNJHdqdxvripyKJMlJcckPd90abgID6LZRLvxY3q
fOdBW3anFpn/LIYmHvfXedb+B0q6Q/X31+vCRu/f2PVtkoBgqkv8bONH1P9vdPZtNXuSzrvtAiGZ
v+DJ+vsi3GvWsvcf0WWnMPSrU1EGTIXKh5JVW2PrqTnDzCrTQCVBNCIbbSjQWMixRj6S/MkP0PAF
/BQCoos38xPLSHZW8dhPecD4NerlFmnmHWL8jMY7iD0jotWohxqjKDehFOk5nIRaCHThqAeX85pA
NbFj78ayjtZipP3XhsLW2CkvM5vHSxhOtbDFlOqDi/aq1IAHkww0SjZ8Ls7iVj3LVuF6xoTwA330
0NRWAqFiGxxEKicLrogMHEEaEWP2ui0XN6Nr0yNra+7738B+c4NjdeBoRNNI1PHdgeoLQgQV6S2l
QWcJ5U+0+7O5L/Bi9bUkMM28a5bYG56LckA9Xv7hmoBPgmSGQ1MK0hHjKiFwoIsDEquwVCPx6IDR
CYn82H7+K/tfmedMff7UnRKP0oGUUl22H3H93RSz3/qTfSVsNkNUgpmjlgjsatXnKimJKyOiqs3X
ft/B88zNZqxSqmHRZRvDP8Z0DIYcLHDeHpTtSV5if/d1GBsaXCEXC1k+CQUiNl8SwkHZqHlILZoO
QUGsjOQwlVZn+UZsxp1VWqDDHUKrkeoMHYfORkyD+O0oQbK/USQvKbTGIVU27f4jp9wfjeAyKQOG
MmFyQXWu4DN7sFhKseE1eQgaS+9UK915LMMwoU6v4lXD9bH5dFBG349nTQHd2VNgeqSvETVjwuND
Ypo861tmN8/xA9SpUq56+lckqLQocmmsF2TMExKxxp1MjhBVKBa5IE9qSG5O14OG5LKXlHzVBO7o
r42oL4qGfhwN98umNhu52+/fPvMITuRORRTUfnd+izTtZXKQCZ8U22UALccrhxZ/T+59KXbwVy+i
31RHJDTVoEUtnAfxoCScjgBfullBg6B1yiolucMCFRjMD/tuB/Poia6idGgKcOrnjPRr8z37pOhL
zyrACr8kNyr7hthllt4KpA63WcKL503pg/D9qHCfKhJDuz9F7exoavpVUPcwdYYvdBkFssfp62di
np7xj6wGREMF8XBvh2MpPlx/fZKuxJDio2+6+D8Ad2tCjajJB47dbZoOy1Ugx/NRFWPTfwSpbA40
kjgV5QGW4V1tNT9VV1d0nkhiXTbNMVD6iVhI05aT5FG2+j30ncvv32eP7oDkLzuJQtPz9cc19Xk7
3zbDe9ps5gd4LG9MFmtejT0uFVUJPuCgmMpDNKsfVP2kSRka/gtHm+2Dg+NFguKZGr6/ech2LZP5
dU2RBPaplxsnDhq3o/FWhmNfnNpHF1QlSSdFLSQn0T/grOzc6mTwF+czgsJDykyT/9fDD9DZJn52
84UuJJbbuM+FFVTr0a5Wc+4j/ItOpbQneEYCSn0cM35+yYKujOkFW9cpdV5UqotqNTO4YpYnlkMB
EPysPHREtCw7mDZgteXYcjtsKgfX2Ze8KJEsdAKpHK3FC/LUzdSS310t6hFrCzO2Ug2FDxOnvae7
u8K/OLaId4KCg16DXlAsuRIpy0Fl5U/ak/mCI7KnTwDc0RZyvra7PfBTwwB6t+p02PdiABINZx69
jQlgfGxqjyeVLKAqieMRFqUVuyIkV5F2q6xOshR3ADbJYozZ2IzzA8Q0zn/rqqmbVIrvFEdxR6S1
i6z4Z3pZLNTViNeuxU/sLG/DB9V1n28rWYUPlHKDJahZ/8LvEqMggw9V2hbamqk5n9QbrWugmP9e
7O9meGdf0vmZsko/CT4szm2Y9XZrjoGF6dHNK1iH8WV5Ks3WOhVE/+2uYHJqtKj4rLsT6sJhDSqY
jvS7yKSdDh+utAdyJmRUVCKqrW5d99kuz9Z6TKZxUPTEcTSjOnnIC2Is4YI2MXuz03QTHlyrUGE7
SzjmV92z08Gd3PAFdc78m6pdEOT4C7HsGnnTm09HCfWG2fCIyG+qv0Iz5jRiKtdah+4NTQ4sP3x3
GEK/h+vofOnz31bhdp2JSaoHBYB1j15aJwf13wjjdMZNRc7oppkyaggYijeA1s/TjoIaWyZ3hRll
NSBy8CWvNMJEOA7o+uMrhpt09of4tjy5/WwQ4YPlWpZrE8lwPYWHNwuAbo+OjlpZDfuiqPPcxoDs
jVfM/XqQORDOY4XKoRoJ/ZJskd6bXP3IPf7NJD4MgJKwApk3UVOEyvDLU6yY70/iRi0CkKoNGtKj
IvPEudxgsyXfKslShPGDPvzzo5vyX35YJW7WSXCqcwndoMUwC/fxvtbr7ulpqFFGq74GNFVYsup0
E/9F6V1aD26v090JCiPoCJiwEtniHSD7esuwhgX8V4ifEXgZpigmV8e+bl7nkjj/PHTKQ5UgTWKK
gagVMk+Cpne2UKKhXiNCqzM3y7In65SA+NQVcIMDZ9UUIMEqPNYuGcGK4reVoPozn2D6swPzQMSM
ERxif9jWdu00Byl8+DVqFk3wTZmkuAv2dkoc6BzHH4ZIs/jG+zhKJw0tNPGKCaITH9A19qnmf5bW
6GYKSteWTi2HeV+6G6ahMEovSSV9pFoewW9gYtfSqPz9s7qVVSfc1WkIKFx2drcUyqhdjppaDKhF
LcnxJDeYoTCwmgDT1mL2/o518vyt1YGNNHQ7H1sD3WyIVbuq5ltO37M6JPMXYB/N2ORRZz/uf9BI
Axbr5q3FYJOhuy/cRxsPcE+iKUO9W3Hx2cf5zYwmV1JjYWmGlabD81Y6YDm2OWfYK4FlcLLUKS8J
DlOkYaw9s9eMO8gmSKJOOqYzaxcjzgDf5K9yRGNz2S9etG+4iflqKYajXsWBOda1MBHFYfbkxe4u
1ct7DrTOGPbOcxmGD2XJJ4V0YRKIJm6py4Z9JjtSn3H4rkJcHLIjesNkDA11kQptHP5xy60J6hRW
YSK4bon6l458FhygITWkc238/A85beRhhO6qGP3t4kOKkdamYDrrVqYxeTdfuTFYGRGFOOL2sIU6
qk9OvjWY2AoqW6ze+apy0MInBFX6V5+Oao84/u9XsiOXudQBjMUivNDl/wZv76F7U/n1pKXrPZwS
4SHIsYqwUtPv9PkMRvV8k0Kb4NNZw81Hs25qro+DdEoImi+JXwpSdEsyUSQPz2QeelgjHt6zuCWw
7c7nF4FEjNjYLOdrS6ASZ+B4rVWrvVe6ZDV18LJVWXwlpbDjYnjWy65GFC7YFOuWXzx1ni/Z4Azj
IvX7hc3mpZxBhI1X3di/GoNVjkRQf3xIzJ76DB42mNZU2JmFHaitmIStGGusNELViiPXj3fIGd+0
auxO34aMaIwblsJc9Jir82eq9hHdHC89OZgxN7xB556zPA752j9dKSi3xZ/9PLmNi2tOvJ88cvde
QROdkNBxOFroCi1xz1c1O3OWAktSrjdzWtwMcEmPrefqgRpKE9fEqWMJQm8/aBHgHziIGt+fXoiK
xG2QPvD4Hy72Gv4NrOn2ert11qj59OF/r7CNxFleyWlFjiCD3m8xZ7ib7/7X8y97igj/d8XkRpnF
ITRIHIzHNUhJugHQzptq92zGpnSdWcvEx4J0pYEScEiAvKEHBqXtw002FRwmbnZEyZTuHt2/T0xX
ewniy4xWS5vKLQVwUkZGaS32OxvF42nnb31JDX9uDcStr5tpzFgBR1w2MSgITRMg/gM4S8jVZ1aT
ExRGN8wMq7QyFg/vQF8vWflv7lDmQ+n17bAfmH/b5YQAZWzVJYV8Yw28+U1XRQtrY19ffgCeD04r
CbMuuf96JsK7f0v6KjExlkKgjWChsC8YsPFXQJ0bsyNiYzQH5Tig9XkVrSprEl57pFmSWnHf56bZ
ijOOxTuvBI0+gbZz5kpg0sCCTswpbnuQVFneLaNoMtZVLrl+8DIXvvYizqAseSBc7LD3joFOdLKl
WbIO2IR2XwU7X7VAapIhCHCGASBjDgKA29Cq14TMhQG3oa/e7OyHj2vuGOuDS0JqtyCKniP/Dt/t
BwfwACF6uXFceSI+6P8ysryDuVpWIY6rQ7SVnlW6HDLEueNdOzQ/RI3B3MqkHJu0/sb3a/ZCzOC9
SMklQ9sZ3NKUby7jLFZkXr3k8lMfzjq3+6tqaS1J11huWjoqt8v1+hukhGV8qaRYYa5k9PbrYWg5
I/qRAtZ8wCFMUAgZuvI3n+qoZ+vwUyH2jdlyRbghAk74Mg+JulV6lv+8MlpDQTHDlmm+WGXhtJZj
1HQVWhsDioVPuTHSi912gjtSSVPZDX2e8l8aINnf8fVDHGJopHyYJeXuz7ceSPXeSivZpJaGU3t/
ZPxEopK1Jj2qPWN03Yy0zzXczZz0GHxSTx4hkC9IGOyTAqj+XBCIMzGWLWKLduZ+vzRJwOYS/zax
mQWXUiBdZpAJYqwGaWprrYZ/tpNFl/g2ELWqeLWvJLfgzj+agMJoZR7vf7peXu9mXl61+cCrKEv6
F/T2sOH0yd8yY0ZK/RGN9QXtn0ukgzf2fH8FtKwhQkR2GNEWB0KykpIqJ46VfQOE3g6FZD1Jk23V
Ui/WFlN63azWDNo0hp+kjBMOVNdnpdU0znSLDBo1OAZDsWf4xqVDRW3bashH5Z7Hvk5H4pZxMRre
3cKmhCDrRm3fP/KYtBTpVNT4dECkqNOPU5YF30Fd4hf+5Wu/gphXaRG+fwlEnrRjz2Oa5ZgjcAg8
xsd9SGyAKFfI/1SjtkycicjTD2taoC6P6WQYOfaOUwlkp7Y98AFgsS1Yi4Ldgi79jbu5qG3KYFkX
GiBCKikxKTiNmeVCy04M7roS8QHdczFjRxcYo12tAbbcdiQjkOrg0XKeCXbWTef6xk4Lmego4ufg
shibdDb4FyzHYnMgBahiiOkq9XHTpAc3Ktc767EWNaXjAe0Kl9sP8jGvSwUNmFmtqjxjPmdaykau
mv5y49gzgM2e90MIeyDl3biyIvvvhCTstm6Wo76PUitStkIFwhTbd7vgD2E9oMkTtEuGPk6z9qJj
cdUWfIkZ36yuSwF305f3lOB0hv8zzGZzKyTrUs3yeoDw8hcO1cIgIDv0OU6wJ3vNHVQeCGSecq84
5mbFtIIgct0HKVqWNqnmglhBnSED55McmZtb5RgsAFmbHr0o/HilY9zGPM3p6fzjN4L0Ajc+b5M2
zcU81VNg6N/sxAG5MJbfUorlZGszD2Xmj69bHfhzVJK3TF+gxa6CMMplTeLUN3XFjDWQlD74NYKr
mkt4tRFwLPzGxnVZ7pNyYnCsLS36vwZELHAJNXnjgDiWFGRwZbkWBRDa3eVqBkb4Q2K4wtGgFJ58
yisC8Laa1sOTFHd9MimNpr+rJKxHXWO15pcYoyGSQt2Ein2T2NjANF6A38htzDpf+vMjEPX9dzRB
NayartkAFB0zokfWEDX/VZ/8rP92106FPcTPmbQnbv+WFtseKnpnsm+3QO3/piqC7YkujrUl+lBF
mUfW9XroGWZSLYdMKhiWsbpR3QdN/OTYhRsVES5vFkKOQxFUpVaus0sOhihKl1zMhw9T9ecwq/e3
NpsowsZU2SgiZvjz1RA6StV+hg475WdMf0aODhJpUME5byymUSntNzekH95AmwOW1UUzC2Hgtf3o
BuwiAIT8TtlWTZXEwSC1xAw2HEaWR7rIxF1lejw1jYvMNgzDccPe/yJodoo9jM2MmLDqRkmMrofA
LbzETNUqdMV3MtR3DqV2umDtO2zGlEUlHz1yDS8+wN4VOH5GSmNyI+M9IsRD7p0lIWXpvYyQcIej
K8i6F0vl8OQrxRV1z2g6ljES0BdkUHXQVqV92aLvdq2iplD6MK9Bc7fGhWEcSjEvBMoBh/QUkdxB
AxTDke6nIwcrnwXzlMODsmwHIN2TM9gHoWJ9s3iqG46KhK7c3EzkGOyY4ivdFPnWExaMXK4nzFuX
IwCSSY/nwykIQUjuGlUcC6+rkD6OWY/qiEU65DyISuqZKkzYwmx0TcsOMAULPviFrjwN2dAylANi
T4+x2OQV61Dz2Th/VqMqdRCDPV8F2N/DvmmVui/j7l32YEUA+I9RBBQA9dUwuOE8Tolaq2jsxU97
u/e/RUQEllbeIVgKsEg9aAYpUwcjrGz60H1ApqE8kPM0FJfccpqwSEGisFAvRdkbsouiSBiMa6xh
tyXIckFMppUkybmvmKnTCLxAE89rnxrM/xfwMQyo7BB2h2j87sBIUTvf1hmb14PXNTeI2zKUmo/v
vTun4VjiiUEqtGHvalMHr3RL7rcTq0GyYJOM4KNXVIyxHbo7VtMhRIJ4ESipP5HKZitOa9npLPPu
LL20bfXRqI4J/cEzPMGRxSif/j8hHikHaNgvaQAtaWEMUkXBiW0xfHkowL57yzefAMYUU7eIhiYK
pMKcxXLF5Yjh4vbK2Nhtx8zTGyFEQ+NgiHWLSMkAB2uIotTLpJ1CYX0/QHXa1hDn/s0IEMhnWZq1
nbN0QTsnh7lstS464opsiwYP/ZhmbjrQvqAHOkr62UmNzLNKc/T2aQ0OJWyIZTBzwEULvG6wYVWE
IkPpdx0Ub/gUAvNKDy2pYOmTSLppNYwTsB3fvOr5hNV19zG85INYHGflALrZqvhc3OTHBU27+xE7
xkFLqa1qpTyDG4Cp4zk6dIcFJL2PBYObPOW8bdKPTnObrrqW4yUje0gJiNrBF6iMSFQHDkRitVmx
dvT7vXz2BkrYChDN5aR9XFDyg4kKT4zkR7CGggDgOmviEgHqGQ5BXiq5F0q3ulVdZ5r2ua7YaXbc
lxPdQpi3z/13SM+Vo95Stztt10MkwPDyZ2I7z39MHf4uh3ZIUXjcsAhWEvrPrNAxwNRAlm4Oyoqe
XqPcbOiSf+PXq7AHV5Ua64TVjoPBg6i91kfOjCJg9rii7IsgzYnI5I255ifb9f01AVksGORXJLjG
QVPTlH9HnuCqaedseF5ukGzdzwmNZmy0ttN6O758xZT7Bgsrfbu2/2/po8wsAd/D+RAcrAriDbC1
1vx86U4d9fI2yXA5GqU/C5aGzU5G2q8mkUsvtS797hYm7ljuXCTM5TocEdOFThva9Q+vh4S1QYAq
tJFyCtbLwMD7jEC9yyLKa/m4yjYzUKMxJOWYums4Suyxu93r0KJt8h6nIN1WmS0MeySP6xcNm74y
shfDj6uOKzFVZYwKu8z2dBNFWBoP6FzLPimu6NdBpDHKY4hpAjkXIM+9H4LRFErhfpEGFTlr6HOd
vJ3jJoHfwozhAFttpaNvNE5+MgHdAFRnlVhHqyr7Je7lglFFk5M7ldL69i18V10Z7eq5omlepqTv
YL4Ll2SVFkLjKFm9T9TWJmEaeWxD96kThkPjLkvh4cgiZywS/hF9cgR6fVuhZZcSvVnPGSFS/IIt
VXW2xEwtv15A5ryyXCrTDsSwQX7oc1wP36iMck7rDUea+kC7KrLrH9FuTm5Dc6cq9tdYvICR/ieg
o7sTWOUjXE2KlMxinYlbMGjR1Iq0JMN1T7wr+uMysNSq4PV9e69bFhg7ALJovPNv8+b07ka8ec/+
ssTPMYqR0GVbw8uRa46/G3bZIhZmiTvtpQfcoA/bUA78l0oElQfX8M5aiFN2RtOFC61YUrsjRoAX
f437CqTabpLY4tBzvJenc/K/NcNBKNMOUYmCxEvoqnJwC2n6qJBXC998D7wRue094APNn4UXolia
tAxTDuE1UBW1/WoGckSVHeLP6PBm0TV+ev4LO97xVMLgMW8f3q7iXMA1aHDwuRHf9cSRT9GSwi7o
7Qr93rwQLH4QRngFhkonHRansdsiocOFYQMf7AaKpSt8vUvA35Y1CcHyuSxCMps/a/qS+0lo/KSL
LL4nVFmExBjeq3JvOuZjjRR5mWDoHy3/mvJekU889fWH6lRNjnEUXw2blquu0E7KdQmWvrkSo7ku
iN2Xz6h5t4uQfMEYBBe10ss+VOP4OgDqpUHt0lSA0G9Ss5XMq0cxq/GvJpqoJ4twguuCWqtQQzqT
vCID2nAQCWs2wE0wjrMIVBCDbn1DkpqVRdGLnjMg2gEiBJgBrNku0kUmRlxo1yA5h1t0KxdIm4Bs
Jmid0mJqpdnT2d3iUNFcCAvzPWZrq5siT86swbKMP30xwkgD9Ibb62TcoSHdZ6rLfx03D/HgoogS
rOjks8QXf7D3jmHNSxCeivMhsYuSE+pwkg1D0YafrGCJTpMlKoHxiMrxyTW2Y1GLflphxYcvT9bW
G/Gvlfq2pPsYefKmfR3FpRCYHTMZLXWKJp1pw6wIfbiNCyrZDW3tKTDZrtL3PuS7akl3Ei77QHNq
8dEgSgc+a0aaAVkhNHTnLqKuv42E3rlAiUB72HaDcCbHXTIzVFXb2l6i2QhRkLkcuiWzOrf+Bipo
UpR9bxeZCQcy3PiWxGJBaHrHUIaw94HIimjHnkmo6JCMk8tjA0hsmPJ4jGsXq5pVK1llLTW1DtCa
dAUF/e33JbQyUxhbUtwaZwat8gTPMQnZYqRAknz1TW+6A4McBqT9yNVFeWEBMR/TjOs+1aFYZt8w
jRgGgZkNZjLByKkxe7jDeSQ0TonJONeYrPpk6a1iIFs3DzBCjKHzmiOn0jI+0RHUIC/oeKswuQv8
fo3yKlko7vD7Gz/c9tXKe8Sv4YiZGRz/lFIrrIBcVpOQHFmp4h7tic/LPRjgoyVKIvv6tfsLXzhu
0sd7fxCP4C5ka5xRp3SPoAk0kba/4raBgrAPtlQKE3IqJJYZbysYwNNvS3IbdWQVGCq9dixwmqcF
DhkSNFg0gGnnP5kjsMK0lGzWEL1IiNkvspeT/i5hbbs/VmFIuH4B41kAZkSSA2Ckh+oHVtuZSsdc
ICBLfDY0YVSf+uB7xsF1s89CG+5n1lv0nTW5P5bP8eGPJiRyI8Fae1m5dM/zffCJGmMJZ5qWpQhj
D5os5dT3yJN6M2KKX6UlZA+4goyEbJWvsvOO6lWO80FNKhWsz4mritoU1ar+5KF5cKghg74dnVOE
omO5B/JrJpGOJ6L7+K3ShXfdwRKkrETFcEMUmGDzZPbZmBjH4UOc0fOeMR6yx2g8gDVI+58jS2PI
BUwjdvy1/WXsp52lNDVzPembwGUYTgnpDofz3cPz7WFlcRcZj2BilCkKIdWpE5eXnZ9hVarBxKIo
lC0zl4W4sCTrmTRQQf6jKbDG135EMpp5XuuJsGyrRu4JHrRg2SNDA1ZhcJTuYlUPAr8+7I4n3D8y
xgH0z0ygF6P951cmqZsMzxZfKT2eDUuHkuYeHrfWe+e5n6Bq3TE6A2MnIggUkPhU9a8nwZiBEKtI
j7tEGzD0YxZ8CFOWLoMLr5kLX4AYqcUfeIEjuB9HRjyxhU+ApBZkP2hYaQeqqkaaWP72qTafhT80
61jzTSR7nlmARn6xz1ICTiKqCA0U2amELj695u/ZDu+V9PnhXKRd/4i9dTEp9XxCAY+6Lajd9A6T
9KIP+DGqzF9EyTxrdmJ3VXLSWaZ1tMPZBCQ9Sb0MSfdpstsNmWESrkNstDXQeBmrHE7QuogSjRNx
nX6d4mW+6qS3I+aGZzFY+9wYaxe+WTAJL2ec7oPZ7ka4Pgd7GnR77IZJ0n645YDvEASMGuWKM5dV
ml+7NFiF57wppghZsMJJZFZmIZg9DMpbJfNNp02Zui0Os2du7cx0ts/WWi4OH+Zef2P0qTuD9/qD
QBGDkY4pmF5Cm5iAkaw37OCFTtBIGoRTgYAsU2JBrx8w7UVaQhIYbt1W6lgr2o752yH2UmhS0yOA
JorsQgvIr6RsNnFNbORpYstbhHSKi6pCswJejzKGSO7P24iLyV+GegTq76M6RN3XDWxCljwb/2Ag
KQScDUjblhX6ssOvdSe9MsLsIiL0p2YCv8n0EPc9mAVzs7r2bryZK6GlnYLy+kO8T1aWMaAW7Qx0
p/VNJSfqB0XyfJuyC93fQ0d/nXQEdFMkIhEA4t9SGkAJxnOU06kODwkAdJVb24Vi+I3qDFEKaRLh
n7mfFh71gw7aZ93V6Jr+TSqxN3zswc3Dp4+KqEojQ5fYBrbVOTvHZ/+KehaLsrqBAofjKuwitf9h
G/7/OFZjZmhQu09lrKN/jMy+gmxX+C/ZFBu8e8tYrnnhjJ7Uvjpc+af/9UDE0nflk4WGw6uoUf8p
4E1FHep+C0t+2ziRYA5rJIa6Xb0NhdSLAgEo5R1OwaTFSjpVvl297ebqi8RwXnyuCtknQNEG1Mlj
TkUeGC2fP+RMxP1NbqzpGK5cvcX0v6K+GQyj9fzazbQGXv59jR6rUI+IVWS7TzR3g0aq405vzMSM
g1i1eanB3daX93/+wQRPscRy53c0xG1OkizFU7ODHvK0+4ow9KPnbKdwe+oyQkGDJ4XWKIrKYDjv
PAJND5LzeN6+ukXOziaTa5KaKv+mN1K+odMYalx89Qk7S/i0FV75a+X0AZS3pxw08Zo4ULKtUD8m
/cmF9cFHOZ/2e3nXwExDeuyv74R5LKarXyzTzShzVqIKUhZHfSOupu87+sOkuqXRixbpoTjF16yM
+UtuQ+QUBSdUFK7+Qmyrn3NOOydPRzaEodmG4EISM+yUfz8TM9bhp38B9b9R4k7v1/yYDct+lQNU
3PdEYwPGYHjRUcSRatNyIPz03LS+PjWrr9IU6TzqCUr/yStmDAOgBcHLiADNSLpzwkmwkwTTa8of
Jbth7LOD7MTshLl5bTt5No+bZcnW4Fgwub6kurLVWDjSaBXwsRNdVA1n40OqZoqsl0j2yX10hr5f
pT/lPrlyQI1IU/t8SEQshK4lDwgFGSmSAxu1FlVcCA4c18kP3eR2vXKJE+5k+EMq4P85guMEJidk
jOJpPtvcCl9H53QRiV8l8Fn+i8/Zhg/34l1CTF3W+7QM66qG9Gb1/ZzPxcSiI2QbdHd+iCYXR1u9
vdfd+ylct8gwFE8GW1fQ5/vsh7HGuJDoIqF019bA4ojGylpnko6G5LKdofsEyG96cHv20Rjwg3Av
bj3CPoX7afBfClN4q+NkYz9wVIsT5hj4RwWv4QwpE6tyxgXq1CZ7ycBMzVWiC7dSlMEUSTOV9oSU
AH97ShfM+KQufphkau/51Fnk+P8NDLMG9AXRvApoBPeQxkYq6VqnUOWTxAVtxNWYX2FdH+mvWczC
ZpmO4bPAEQBfhsbAkkwAJf5pR0Ej9TkyvCdAsh9Z6pxwPGsPuC7MdE2iHzjvzsjq80GLR6VBhdIi
lzjgtP2tAr+oOqKRmTcYFaYd+FIhut7NQk3eql4dX2Z3dlqrBTLV6sdlJaodddMPrm494dxXyOP4
dPsZ2qxgxiX+bPUzfp+NgVjY/NEZogIvEjgWBYLMRNQfhAaN7ZYL50VwAWwunatpTd0uOwOhasKM
acuc8PcHnqOG26Gma4jZAwxDR3RMYoGIbBE4/lM9zPaRWzxMtUdkkO8uqc7ntim6ktA2NA1SH49D
HGUE8xvTuNYKM5EUS9MudYOKWZld/UZBiXrxGS/IOuIY/qVLOIYTtTJ2agMz8KetmpjWKoh0MSjN
REdw6wJTCm17asu1i9FeS4auv4ST+2WbjZOXRuci2J8OFEH0i59V+M5AvGISAYMj59nReEBWF96v
DLEc9h5uDak2Mbe4l4wjpOOZ6AUGE/P+I5bS5I/U2670R8fW+ZUILGAoOdu2Q6LZoEsCx3sVKWfC
S1wMadgDxAkakO6bDSCK0tqSIHf35QwDQOFA2iSvjQdPNJwsJH95PpQyNw6M6gd9RM/DwLOz9cEt
Xsocn0GSvMawTCZrubTJE4ByvWChDHD4S1WBY+vzL6YGt6wc+B/J81BK5TOtPpLn0H1qvKU5C76I
9e6xX4s81tpWKDNPAzk2LLN8y3xlJ6FyZSJuufRAy7LWqAULURbhR8riaoLwRpwkH+d/q8YvnmJN
WE60xIVO/zkdoN5kOt3VonWDVdS+TCeNwOZf26h49969a6smD3FVtck/5NIsfrTouRDYbfEYDZt4
iagRhKcQr1tCLGAbipJ8e+jEvsVYWdqr8KRQ5wru6FkAN67NsKYOQCkJZWVOBOURy2DjFODpIuwT
QNe9sFRIhDM++acdfGlKiGvGNUP1B5vwSOAXl1wpP843h0DUEQJGo7zl3Kqhzf9w0eNGZclgOt5R
HUve5YMiZIn02xhL+duMMfwo19HVOdUEuRBbASMvJiBTT+Y0bl7fLb1W7cKu6546/v6WK2P4V9id
Rk9F9YBfyfhDxyR94cRz0Zx35GIME7O6bMosd+Ba5kF2jCqXF1jDCpaIMyjUCpsREN00p5jEU/3P
YGP2jM0raBiGFVkAK/8UJ751cRrGbtfVdzArek0QOWfelqwa/bxWazUTZxVKadXv0GEU8IjiRvEn
AITwNFqzVWtM6NDZ6dymksO9WYhkhITGoGTTTFhj/MI9xhRQvt45tcuGb/ETLKqNgKzfzmCMoBru
aJnrWIMzwZeIz84/DCIKQ43a7bthsie5spi1P87SBG5iLMd/wbU6vn4ba8/TjNigVPL/hcxCoX4o
34nUzUM+HOk7WhewBNXaYyIbOn7XNpASjhCkqL1EH5mZSasAAHF6mUqHsQrAtmORuUtrDEgxMeA9
5tTDUfeZkIgd37JCpWt8hkPZPJPqXd7t+7mXGzOEEkuVfoyCwvo4Ze0aOyzYz7XG5RnVUZSQjJPi
sMptYMFIb746LXeTIEoWR4ZxS68lt8T5E2Q9O6YSSxxHdvPVCOoyXjYwDHsOXPHtSSS6ZW3pyZNw
XrabY7YLPRKMusDWUmrAS0O3QmX539srsVNo3WcGKK59m17sUIf6ghEi6IDBEjhGiY4rPBDBqTei
SYOyHNGYY8fbVkcmkabLzXSEUTEmTnED9u7cg1LnRwLBvMCalPwWj3gTLyjk2SUMKaTPv0p0gBFR
+aLweJCU9XbJdiJ2ckFiMIqGaOJvZ2o7WazCvLuv/e00+olDWYGwas1Dxy1KLC98T7Y+Wn6zl4Uj
KnttuHo01ad2KhIGvhahIYUKA0FwKL3KwoZ4SaoDAupeNO2CUtEDTVWfRGkJ8RGtMkFbE4BzlvTP
2oTR3ZwFinZFvekV2qBjvXJr+4OW07Wsz6lp9tUi76GoWJVCOLBifTiYY97sIqH+PmYdRcSFvovI
5K5caq91JSF0oxTS9FJJlpleAvq366s1XWymGb6UfmQ+1f/rM5q7RZ2m6V6aqcsku1XfQj60e6vQ
NO/fGDNnGjKGtG7OyxP/xq9IJXIchjSt8QXK0Hcl+wB3rBfL22ZVSIg1St3QUgG1+heAiPxrLeQv
XYFKUs1PfbaMk27Zyt4IC8Yj880/b+snoz7nnKOLl4N88M+RMSknu5dj53c9zI56qI7Ody/e4FfP
nVamCxZPU9888g/uMQb8IArhxo1TGRhORq0OuBhoicJe7VJmulC0xcFXg4KF1sQp8Ru0gXlhSeRS
Nszo97X/6leWr4HmLijbO4+q1Rm0wPEDC6UZPOjUNirSSdZKxpOQLU9+dO0jw6wpqQeXKO/QQKOT
BM3ATWysC7V6yayGvkiGHX4TPPw2mxnsm4gdviATbwa5fLdcXV1gmHWpeQcyydw1E6i1Vbbx1yGZ
OpfPfVhdClm0Fm4vmeKImRkM2GFkBS+SdQzpiZv+LJ3laOFjGhXs10kfIUwCzdD5NOAB6QpFYatn
JaNf4mmZmnaKsRw+rCxfyCxqq2xKC6o3pliJwhdp9RuHWeRY/sb/m+gY8FIbgTTSuwPv0919+oJJ
gtaq5+fjPaO7QW15iLoZpqco5CMNgWduMUGEn392S5QvNwjBbI0JhGp+REjQFUkOQIvBZJ2dcux/
bmOc5KIw7L+p4+wfos2y6L15yu+ox5ERwlB/RihHHKOmPTMGRCBNYweB4DF2T2b+YgydVkWqsNdK
DKD8LqqD754123zeIDPBWazikTo2CKuyp6SQFJHzgkrXFOz2whUFrtfvx+l9K4xuqNSSP+TjSqXO
O8BwQEtvqgp/nEsMLtLrUzNnynkR7RT6F2NE48I6WoysLXzdGWTSrJ3k6T8kRE5Nx0IDoYGjzQG+
db2AhYazzZjYAPln9xYOmlWfboyrdMJQw/17TmDF0Z0CGo/SLQJJNJ/l4epCRGQ3nzQ/aubqiYQ9
B3hGDPlZDQKp55UALwhFS/7VPkc8i4U6RmrlByO4Kna4HFTTzI5Zea0WxbuIhCLaqi+hff6Vc2mt
I1rq7L+p37NdpCNEpF/wz5R19YsSl148mI4lRTPqko69rIeIr6pVKRMOPHgaKl/D7zQToMQQHfuK
OtF8s5tLIQyZyNdKL/9gFfdEKGmAo6LyaPfACV6jUJBy99TCQRFH9SyhX3f4kP5awkN/kHvldYbX
UfAWiAm9i7wvcWj+Spa2Ihkb7efUl5kSPaZaZK55NUp752bYRnefNnAvQBPtdg7fWYrf8lXvbdc1
5dx9JcgNtHSC+YmfcMNyMa4bJz+Tw9QhSfapmOT0V6aC+zDjFcSN58DfPLSiXfBTDYNbt3fM54G3
Tk9LXvKzxu996dQ8/isd1Bj0EN+BYkmPGxQyLB+R/rnPEjo9fk9z4a6yEHHHiFw9dlF5BsiDXORw
+XnDlRq5ZLSm8LZr/8+gYqsfPJSm4HUka3CHT2schE0xJFko+JoUHpAfZUpDhDrTqfkqswH9TaV4
O0oyXROYHNKlDWZZ/2aHHsLQprnHIR0CUoI+wkhrzBOner75xNTBkLXKlmxEZoqCA7/YJOCF7qhG
kst1C5DgLtOyEjg4y49MxEQl4ZT69ZzTH9pGTDcY7XLn44hhYirJC3BZJJvLkECjHn8yvHeg67Y+
4oyo1PmMwTrkbvtOeYNZSD8O+w6SaGAqT39aOXdWUJH/Fvfcf7WrxlJdzCvg3KBJvRCk6kg29XP7
nogV4OZXAgMrtIS6ohp2aszbLpDzkbXtRL+oBTr4GjP/w6AB+yjNCMvZnkn/a+v0RznQZA35fo1v
AErgyrzoNML9EDiBL0+zALfrXT5iE3mkAC3gtTy/9xVYTjs8+yKd6KuKFZh6SM7RhJli1+kuHzFm
DOJQe8bbb/hv0v8ArvjImh8sgAYWOhFguWAVr/6Y2Aahre1UKfWMl6FCiZyyOh2Kib/J9JyfEG/K
pn+MHu4rrEZ8Hoy+NWCmYx07CvHQQUtj7EsNkguP1lhIUpUsSk8AscVvaH/sCS9ecoOSUgiMiaoL
KNKARu4fmgu2XnkRt8u0oQxFtbqK3Y9O2FizLXoABLVGdVQMION1x36yBLLO8uGVgPPb40OOtD5W
KLN8i1ikZgBtId6BwXJcjnsX8n09W24Q1vH8CXGCsV5EvadIrNemK1f+HnLlPFV9Tyb3Hwem8YJI
anvU5Ki4GelO0mWnEKkb6Z41O/2YLF0cOt2+sD7LXLWk76L3N4nfSxkKZHfPjXmj3CCOr+aGrEs+
kumAtpTJ3cTbyCjkrz/Y9+ipm4F8wJhEeOGYGhkEB6kc3hc3Ww7Fh8/gTtO5Yi8ynmEJqVD9srvw
Xo2hxrrO7NNngj2+96HPFIxcG4md7Ie7hK2szQ0R2l3tLmWXpyFXqITn1oKAjz8qY4Pqp7hMrvTC
SshgdqsNURvOUBprkw8kviwx5J6xSg6NmxmViDVIGYYV7wVvFM7M4E0dGsjRfFHYhcJIfNsWKo2Z
ijqUgUNnzzmXCEdUqMzFpaBiU9MTlboxyFbV48IvKw1IfBWfmqYmT7iR5c0rDpa7nYLrhRvRYSBW
w+a+ReeFOMbYRy8ozykzWCHkHKfd/engNK/85HYTha4aS5DzkQCl6WcQWhXL3SIKRQUhCY0Mhne2
fokJrlPvrf2qQnBdmOr/PF+UFkc5UsEqPtLbRJGzIIQGetLWKcjLJbBnk7RTGqcuB17pElx7b99Q
ZWNHV3i4Cyzg7LQIGQoOJgDCOQbxyrF5AfD8EE4O0UT3/z1mGMd5LmbfrhB3NT5V7zSwGgFyoiUr
FePa+WTKJnnuSvvaOcf2GQGAf+ZiabBCbF3j3UR8Xj4wpvv6j5aDSUbJBgOmDPNdcv0s7EMU3X7+
URpcM8je16f/VezDLpo4aKqR8dKSfAZ7tukst6QuG582YkCx3J8ejmK1iAB/VcIPW6kFU1Ppa95b
IYPOUsz2h3/xAm8td5zMp+EGZBETJO2Hsy332iDyUHqUa7bYC6A6Cb87pKESPC9GnZbHunNCkv1X
Z4ZZ2Vn/1KkwP9/HwGZVfAv9vCFT6ewTYKr4bu3UgiMLNHynd0YlrN9STEuM/YqCFk+gCPMebu1M
PQJ60vItt7Xf3w153A7IghThefPsdzcOj/W42HD8KRIl5lMpgIl/4T8xk4imb8bFbUBEtOKc2Rhh
L1jhXq9B6c3NGX46FOoCb9zh5wm4sFTS7rkob39VLW24Rmxg8vbQVnpsvhkqnNY+yZX0wl98Gh5i
OwenrCOiytWSPKG01wjmhSXKwgEc/iecKy4utpVlhsfhYSnoB8dXNT+Pwi6y7SoiByfZAB1xg9jO
YPkaWpoyuRBYJzbW9lxn/7TSYh+gYc/eFJnrwoOAhzhrUHElQlJOYf0WislMcPtAAC/k2l0NW79o
IxoypN1KB0Bb0BsadbBTWF/0Hm2eNOXBFvY7nN323ryiOysU9b8ikneg9JY24QsiN+Dsl7YxtXy5
7nbLfTBjmZyy2C5kfW043lcoQgJLg911QtZMm4jnG9CFT9WvsnU4H382t0fCGHTGJYATqoiJksFA
IfQjSuYM297Y3VoGqu+qgGdFpwIcOGjf4ASljQlVax9PrUdM+r5vnL4z2UtK7zRDq9phhuccm/Yu
+r8rU5OrJaw8+HKbe3eM5eD+xSHmizDOyRSHVM02LOzk1Xp+t+bM9em817n1H981kOu9eJ0nHcOp
gOe9Cw3kpxosTKVjRJky4tNKaNOwzmekh6JhJA4Lh1dSQwGbASyP1dpcItU8hNaU/EJcedSiMg7K
MA9ca+UeOc2LBrHEfyGAmMdycZI+gw9VkqEvXldTzDxzoTkWhhSpA3g8K3YKemkURLg11Rsrcb12
L8ve6fq6nwUO3kahI846fMx9cA2M/V/1Aeo67deIQumLHfuD6LhhRSD22W3vbmbhyj2bYnvf5SIf
OT1M80IHmZ/k4k5BszBivyZ2gMZjbPZ5b0WbpJZ5TvofTpbzCDC6lsM9OFLFg5JZsXV7DkGMBssl
Z5hOXaiZdApDhK58lOaMF8Yl4tuzOXubksLzLwI0fZYw4jEBHLIVEJDqZ66ZojpMybhRBkExQL8u
q0cTWQP1ozdU8uLtsFJuwrflKZBJnS2GKh7Z7R4XmgaREYTx5diAQoI+XcypzX/aXBjsWcQyjPcB
GbxZ76N0TUYulSwPGy9g/Ry+nbw3wuyWO6byzkquhWqxqDABBQKkiDR0JuTO1Vqv8apeC9VK48Dw
I5HtU1+kcpajqu70dodLVNlHIIQgBJzQngGFU+zKes5pfjdxFe31mxMxewSsqY0Edv4Gf7ITjRfb
stHWFbgQcknowtD7CLRbmwx3nIKSuBQAFC90wcfuoW4KClQ7KRQvQzuChcqo86kdOrzkzvVSAt7g
sPXCCeV1AKlK2BJOqGCGRIYcwdK5eLXJi2eUh2wOdzlyVY+eLfNQdqFds/qi1oXvybBgR7HqBx9R
reZBPwK21b0vjgNmi6YjDoilvq96Rbu4HS9zz+B/D71zgir1qMeLnm43gHaAkMxk68X8/MpPcFID
iH1Mw7JhpkwGzi6OE1h2DV5ZSAVlYIA2s9RyLUBWL877K0J8bAhWNFa41Qe8gNPBXDq9JeqqGGB8
IG+UZtN5q4RDCe4T7wQJsYfiECB275x88eH47CD4j4lUtzyRq2nabySrDyzfgcV94jvQVBq8HDK0
xv3AVrIA2KRRGul6NE756s2JiiKFuQ2WLGxw/mOu1Nr6LdpiI+AZT19yXLw0ZK/qLhUdenwatERm
nsy7W9frJSUme6Y3RkFeLkWqa0PGRqOOyA28M6w4IVAYsNN3chncQSNMPx27GFdNSMHhCwrdJMb1
YZxo+PgxiGOwyXVb9D9NTU+6Nmm/WbPxs68eW4m1D/epZ4/nCgc2eCYJcOYsXtCS7I8s73pCGmmC
ECdZ3cK+DUwgsOHdfMMgIqAQD4snvRxNpS7flohJbuPde5Ap0UjPu+nE920w2u8fWHSD9Fa7o6c8
XVdjIYn9d5V8oxRRlI7kJ6FJ8MS9gzoqFYhw0Z8071OhQPXXa1LSx4SHQoAnq038YFcwKwndVFMl
KObCPa5moy1vcj0cH6+OKfTeAWjdyOv8ab+KXgaAoA6St0Ty8GJAObhaiPiCzIIL8cjKJGZ/xfbB
As71wHBNWbUUuXPTcvQdd7dps3CUw0Q2JyMq2kHxTJFKxlXZNZ/P0tI/VnRk+PjYigzjgbYUsACB
fkLlczEdwPsVUGjeZrYtIVw8LfgIm2bzsrV3e3RRbNNhaWWKs/75T7+L+Zt8Kwgp0dhz4AvNnKiN
7zcK4Sw3Olonbp73FhXYmRTnxmHVzMrVLBTFF2z0uJKDgUuyyk8Pb55OuxhkmMa5WO2V5kKKQ2F9
2bXW8XBvwDPxADmARNXVSOhMIV6kJJjy1Ovt0eOivCSL31jRcjwkgN8XgTjA+ik/ZWG8lCBPsh8p
V6AAIpaUTUZRflpXXeYaPogomraEmdktB4BkEeoi5nGq0hiYTbMoJuYHTMrjCh56L7fifAgJbeQL
3gcenH8UG2az9BC9p+wJ4HrMUe3RwZCfhdgHgpOA90eoeBXDT4nnIUFQeyw3KmLXHUs+6vFG8AK0
NSrBElWs6kNObUEjHJo0Ona/fudbqV0Zanv48h0Ul6QYsWbQ1wT9UpeaEojDCu9INseaVIR4gfQy
4gah4E8B9oXF+w0xZSM8/eo1LWcjl48dYETbuIsWVFHFVyXZAeZBhOFLAagw4oxgGWN/VDZIvjST
g7IvcTYh/rW1d8MLMMVVKrdSL3qqYfZMeBo89ieaBg4bR3PK1nRJsHSdXwdYt6sOpgMKhDngxlbg
ogwttcAxMOoGkt7oJkkVTj1I9YBo/kL9McY8mR/wAfbdwvd8r8XE1Nb9BQczm241eB8zoDfbKo96
j0Qacot7vGSKSY999x/ODFxLtc4ggb1F5am/3fyxQ3ibCrRk+xFBm7OtHXRrvpIOW91c7ZmCfFQm
ZLaYh29gzODaH8kvH3iucIF7jT2GM2baVhJjEHfufNyqRBOPFKyZHCWnWPu3ZTPZONQOZG7gdm92
DKoi/FF/XkIq+BTe+ox+gWpv+U1upjaWpXIc2bjLySiUhP2D+yLt9zQ1ooPNI3TGRx0aLXRdVbKD
Zv20QXR4KexGo9V7zP+MHx+0n+M12yF8YaxBSbGua1KgB1sHRuDY1hJjiH7CrWEOurYCK2NNmgVJ
YWNo0xivdWQ2hRqaUFcsqvu/EWbp5znKj7gxUaP7u+xy4Sfm4DuV+7q5U7BRdku3R+s1BU21cczS
ruuZUbqVvQP+/kFQ55PafxGMxR1g2eSN+jouBzuCU+vhsc/VPLptCjIk2XkpLuExWqRvpjm5LKam
VNV+JusmOcI7PETA0hsq7qo+tq3pJuV+v8k7AJ0DsAgVVdMW15HEs4LTvMbaujTXzR+OTbECkxWP
pDbNheIaBnBfmSCxy+TxUWNNCxh+2BbiGnhjXsP5UKGi+0mFXOc5iTvIwNIszIcez5j+DreTB6Nx
2MmVE5Uwn5QGQrwOvxKQ5TbrZvbXr5li5NPM8EaZOR6++6U7OyEfhvZf40P2UVC5caslHf4GrGgp
n0CZtaAXBmozfwDHZFNpzcQHTmflEtR+wcreMSJO/rZDHzreHZdX/+sfpUgCq+ZDvEks1Bo7GmK9
ZKK2wSPOLsMn2Tz95hvXO5Ar6cMU3EaY4CqE2oiBD9SqdPexkX9JKPyJPRgYn+KzVnqZyWFphZWQ
OP4roNMHuvp+ldJBrhb+mLcaUisPBJkN0+J6/tOVtR5oJBdPa7IvJFyN3Xh7qb3OcLLJv96y24Z0
/lICHoqAT0mHO5mp4V54FjUkds8yMrlqlFHXNYB02cB+ueeipSkXv0A4zyEcgSPqP5NP1Patv1N3
3xvqUFj0VdPm2lrrBIkg6VZeQoUxUkI0nGVDJNeCmoh6zKj+NwNr2AsuIvg27UT1Vo41vrpi1vaC
mDOcTKYbH1MoH+QTZMuE856Zz1TNFiROkAdNuSdPY5k9RehhXy5Pc66veCBCoYAicbdb7NxyLB0v
4rXDlRnd8uru5mp9mJWoWlSb1NkQuh+JVjobIw3nSf4rIVg0pQswhsjYBrBVXRR+bdEk5I12Jcu/
RjVPPjkGjWiyX6ZzwhWuSThSGtvE1KXsP9NXu6wOou81mssQ64QuE/gqqochQTPZvBmYF7rfifga
GAdpb2j9rYj54u8bOEPeeZIWLx8Sk00jtjaZBFFpNXWf+8dhhmnInQjExEMObjWUpVyxylwscFGa
CT0iyUtbDj2nflFbd6PW2uDIK/OdkM+rPeqqCE+0XyobXxmU7HxETvgBkQE9cnxNuwehAupINr2r
O2scVbLc8lOg14VvtWIAiNC86DAxX82icwq6b3dMVy2xoRI/f6Qo8iBae0oXtoUCrSaxJFuQn7wA
Ss8JSqxvjQ8ERLztNynd5qew6CcoW18vb6XU6D6Gy2hhmPkfNkP15jnyM1wLBKSvx84bXifPLpFA
QNWH/xewWoBWLB+0w6Q9PDY3T42WeZpy5NpZJSipLcUbbvaac4TJSCfJIAbWep0BEkYCaZw7TzkT
p3XGpye9cqE1V3PplQckGiOijT9pUwtIjnDd4EnBV74FJ/RNgNjQQZzSFe7yVXwGm8ngqLFSmxrb
8xiEPXqaPvWfhXnBnF5TRF7eYRosbeAjhZ250z2m9Nfu97XgVW4qg7Uuqxo8ngqlVNb2GZAHWnDo
toDK5uNGEDC64DsgPjDW5/D9H1Mewc+7Pc1HG7FKPg3BA5iJ0af55jexjf3sNPVAdQmEcgfsDdZ0
gUGuHDKbr1+jn6jaC8OJ6QJcUPHxBdCy2pLvoW+sWnI+jxQOqkchCobZrA9IYzMHkjN6ELHd1RE7
nIX0edE+hbvgZ/l/gmKtqJ9szDQVPHuBkwV0nyk8Vzhq1lH8mzrZBr1NW6ULJdKe58tVLHvKQ2vz
wOLb2Mgh3Z47T4CPT+R4XF1vtuy0jFBlUWoEorYsDkHGs8yV2KJPhaaIjzwVQcpn9c4mQN0/5fg3
328rYGcvvsFwLzbetr+v51NnFbjAyhovf9XM6pbFkkfudINI45lhajtTNiJm1imrte/TfYsGKluL
au3QF0wmOCa1JKTAA4csXw57V/by0JEKrbqWQzITGJeKk861NJoQdpV1NcO8+mto32n9vc/a3STJ
EdYXLsh4Dkd4VuEulSng9mbWpY1XSkgl1UeE/9yYEqS9or8y3gFthMwmn1HL63FjfT6jJn5GaMhv
FmtEOQHrR0lRgkI5v07Kr6FCIVvJSFus2mHHWb8uqAtDzEz2BR2970b1C64kGIUTL7RknHZ2+a41
jPgxDupBBuHvpxf72kKDA8zKTRe/Np/juwTjDghlf3TjBz6TkZpqGQDtWLv2rhpmeI8h96CwBklq
iAyON7VmmGPLbOFBCuyQl5XzbT7nuk0WqYdfe7wj2CvASD8AKdLFiIJ0zr9/6TzNwDXgrLiykRch
NB82HAMoNq1Ryqu/UGy9h98XiWHu+XmgRbnbW5UNBP5tnnopCn/nXXSZEOFm+fgnn8AbZieiJyDJ
6ihky2A1xDGyeDyd/sTRL69Ut9NQYUUXn7YEa9cMpkYStCu8jAf/18yXGvgW4rRrMA3wcKo+DcFX
0YR/+ZtTygxPCr6kwuIg64Efgdy3zmV0JBSmPymJAHDTOibgetlpJVqR8hxvgGlDOQA4BRq9sjxy
jTeJZ3e/mK00GUuNY3ZhOqvYaMU+kWZL+OmcBt/zPcXeXMRlUypcuz1li7aqrjGsmmIwqsxN3pFh
b1qEgx0McWXMH/3YgWLYmPDPuXk1yvmtbUKo/FEAxogUK0NUlUPs5L2XYXOBq54afTjjS50EzYXn
PigtgkswryFQILgVOMRbTE8rjeeJGOZTJU5y3r5zBVpYPQ67Pb74G+C8p0Smg27IcAqdAknHLSqw
T525OFRSLmhnTbBsTReGdrN5aVehacEg+IOEGe2+W0637MP61hqEeEl4QqwbgBAO0xOBVBO0o6xY
EOU//44w4lp3shS8s70KY5B4zXPQIjt3UwRi9ji7e2+32w0eKkJ/mNWlrNqLcpu5s2BoR3VeIFx3
sVBLtCWpsdSJ/e4UbrZ1/Zb9wrdRQjwI7XImcv9jyCsmqEFYQuq2mC6p0DOH4ksu+WIlZ49uwHT0
a8wvjH+vNXJGcmnJcH2bKI7rLmdVaLiEMNBtDMQwmtHfNJxioSO5E+EVyzyvHoDTiWvjsc37bi2l
KgmXKXK+GFdF9026U7KdQIAV6f2A41enXTD1JfGSadGDaofKoTS2F2NZziXT1aH9qOrwwd6V0PJk
GPINQkzdgMYpu6Us4UEM9lfkLQHGnGMUFyHHSJqCXXgD+4YE3Ab15FOcehR4UH0mQ5KAqjbIwo9O
U1inNxGCFFgZRRVhsiQYnCGYwR+AeU0AB9E4XJzRe06/aMFkdALPx8x5kzvIutwFbvA8zZDPdLPB
d2U6mv9C+mc1jRcfq2cvtBHpwrNj2fvaspstYU2yNIs835SSFPlc+SQlH5tYlf6eoyH66xvGGfjC
l0eoRAPNsxLiVsk9O8WtX9C1lvZIaov0f50hASkf9V1BuZWxJpL5JlEBvRfrKF8pvNLA5gf2XRw+
HP9KoESqJgXEdBpgX5ew8fDD/NMYAZNmyqqfDc2s6+geIPJxms1fmWgLWRGRK+GyHus6Vr81Cpq3
74ZpLcB8jT8Mf4KH8x2gUQOJdbW0+sDcjC9SEOK4jji7gFGUJWOugmGbg0BX7q6RlrkxEVi3Mp/V
UNAv6YItAhWwjXTIEV2T6gQf4hntTq+3oQOwiwbQtQcQqicinDvnWjkFxwSYfENw9IHgSeSqn9gB
Kx6wQBTh5rf7Mx4u3lSAU0vsUo8ZgC+aquOZuwQTtL0S9gEeDLlSzF1IchZ7hhFFFl+jNVEM4Qoi
WyZWgLn6HSKYvV99q4w2TVAgP6HKTeSDtscvTNscCcagE69t19Nhah2Y2r9tftwsdrtpqOmB8tMP
ksYHEGrumdGGyRZCMczebrniFbKWmqLrt/CNPNClIZFgqtRkW+EfZ3xYcY4Y3kx82CuDM4tzEZRx
QIAoOf7onOsTMHuXr4UBmO13fkNIrTmnPBu3FG927grT0euG/XqPlKOThylsTAfZhgE0EH4Lrlhe
74KFUkJYviaumCNyS59kf+f9cZyTOk9DevNQhREDQb7Rkvb6tiG+ca3tKUtqW3IYsIba2bY6nt80
Nfu2P2sGyhIT6db0BevQe65r2wGPAkCbejtSzXKUWX1uNv1foKE8U65AMd7QQcEVZiDP0Ky7rWyM
ca243tDRVW0AcIosHK8rvBNOfmXlPxQgGQjCyRbg1ISFdV/NeEqlvSzsLxyuUC184S1sf/pUxbFb
4ONfgINSiWBM5HxDSK9wyQ6pg4Ad6GjpAgJfnIJnySIydibIcOG+5XBFLy1iBtoogweH/05/Qq2d
1pt8p4BIoMtzYXFIu5qqA850qHZ4tvVXX2OiJWrxVKhF7LiIXFQIOcw99jJuqf9YKSdjyZx6qY0E
dcw8+QaH2488+hwxx6r1FnfSS5Q/8myr0BWNaJhIgsTrEppJSt/FlYP5Dr+654Fz0tItqI2u2me9
t+R3yDzG6vlWgrCYBktmn7y4AcLW3Jkmmu1JdZqCT2n3H327Q7f9q49J94uInXbvysZyorv+L70B
pn5zvuNFwwwsyPHJwXZimiJxU9VodZipJfspaXjJQpKjMb1lB2ruAW5jcEWG8OAmdprBlo4AHEaM
MvONTb/Gi5gfM+Mm2E7/kzMY2JlwYROkquyUvfUbQfmApVnqeDn3Q7MjYtawzFbBVaTPlVTclQt3
D2908QA6lkU15JUWhUsm+raia3ahZa9XbWrRsQGbl9ha7oH/ismZL9jBRV8+0KJPkcr9No2J/bOf
uj08Nqu16zbotLlr42tOg1P5akUGgidXDETh0qXtNbQTBGXNd/L2uU6HsIA3Tj56p6+FjhCNrdYT
iBf/Fv7mM8gn+mmRHHdfEEQYbsvlYyztumJ2SO+0HN+SQFxgPvqVwCF0pvWLZrdbTN6AXsM2yCXI
qPRdizNu0CB0/Wcme8DnyJ6w2SToGxdsMQCP1FAw5qEVb1NigWjnO0noKB8KF9dFIEGNd6I67eQh
SZNExembDPKFKSRD/Ys/r38kQQdLeyiZOXQfMqcAro+HUmlJUh6U9uJJb7Qvq2/lQrKaSk1loPNw
7zh93X3a77hyVcKPAh+TErwNuovyMJqFqMVmN9Yf4mfD+Hdnki9C1yAY05Q7ZooNQaaF50nBUwOD
g3fc8FDboQ2tgUIxuxecYgo5D+y21lSwHB6N+GLqrwSl5cy9mzq6n7KYx6xqz41EyAuxvUQpA2Kb
pJEJFDR3wMYluHF6bRlcJyNUQhizM6pcdamxRHQaJchva1/ajF7wnWnyQMrYGZWM1s+Jy/5zlSoA
3b5lOJaV0ASGEyNoQ614hdCIYZW6qzFWhCH/3lLHLkPL0UCtW1+zGZChPT/N/F60e8lJWWq14RoQ
0sv4C0ypjYvpAzkkYvbPfqWpPj6nev4RuDD4Zlxy2emZJzS9EDyw32Xu+wxXtqGLbtJnrhhv6ykP
uBUcY+P95n44p0sw6neJa1a16Gveq6buJsGpssdLV7MuHQvy8h9w5HO+tjy8yn9hrguPdSBd3SuI
MI28U5A3Z1MC+xSBp6nC1H3pV8XHmDxiSrZRaFGrwmz/ELCD5vMYXU/rFaQ9wre4d2JBSJXEdP4m
Nsn1b27Ntnhcp5b11A7OTpRFG3zEKJbZhmKzTOPpXURXB1/SkwmFyQAaZJhYSw9ATAIS0nq5lHQ0
PIhcxIL8WOzgVArfR80ErF3exqMYnxktTl/tDUlC12Xs8SBLmxWjTDLiadmMIneeFcr87ppM+jGv
kbLyPjRO41byY7q4oNsT9isV+hGNZxp9hpNMJeah1FxOVkw9Kbc465kzLQuPBUZgZzWyCf3ln3nC
h9L6i/vU/e3uLWdaKHaiLztdo4+qNYqREFG6x3NdBGrL7QpnjGA6OA3pNCHbKDLDlK/NEKeRN80l
TXP+ippVsIT+VhO9Jv7c9NKEcd3hjN4U3pQWQQveMMIm00PESUH5zNfdYjNgG9zbAnKV/qJDab1x
WPFOCQgwncxXjZEQCbZ81CVcaw1juvciAfD7X4bc+cwiEfv85H1x+dWDLnaG4/p8ZUA00z2PN8NF
F/7hltSmP+/9nhoiS11QVIg2LLA0DDi95LaLHTQgikVFCwtjBnlIhXeDYk8J1QF1yBNfYljy4rFY
600PxaGnImUToR/2PlakkAClI8zJ3GCrvHHtTn4j56rV9YT4flOeJyctWE+OHMlpa2Aw5VOPBD7A
G6FfKpPUp9U5gjla3APrOCNKyC5I2NBvSk8pK1McZa4mvrFAcW6sFJjZi7lIJagzNDhqpPW0BGQI
QALyv8a8T7CVDVvYrUXrZI3W98oAyQ8+qHSPNS97kzVlwP4A2vbXkXLYNxlKdegH5iCtqrXtbzPo
Yjnio1Mw4YJgsljEOEmcQqNYM1mACUf7VG+LNIsRaQuhD599rXF9rOgF8lNas+lXAwovU4gILVRl
oqcE5B3i+qr0Dmi1WP6qRA9hkkPTlsv4O2bXOMaF+PHHVRwOdKUN1m6wMdU1zXUJfigZE1dy2A+4
ZERk9U+ZSt+tVZt6u+ovSUuDh9CAJT9tNC5v9DuIuemoHQ9JT0gBvMrjQ8LhVtspF4uzTdlO4KT7
AsN97QTxIBaqdRBZK1wsmBT2BC3ywq16N+ssUSp2RPRiZzuOVJVPpql+90B4EFYsAQMrremVqRnY
4bu21oHLZHxeVpUfB2F/wZGtU5lY8w1VuNE6lstFshfA61pgF5ucWP6Q9ZewNF5XW0CHyoVWvb/2
oZxDKA4HVkgHKIImXtbwoMW+KR4Y8ay8kfZM5hMSiQh9CUmMzJ2BmUnToSa6MyOyTjyJ6uigWUXL
NZEKO+LoSDjAE0AwvU7VMaVhe5xaqUA66DOAGLRbaZxjcmLqnVFpyiV84E2gnFLq2gmex86mPcVp
bgIcM4z/57r93ht2Pd/hAKWz8hyNcw5YH9PYC5j3G6XOcPB54qP/M4SA+8dGaLqHF2GxRUUsJ2eS
NC0dt+ST/nc7GbtOdyMbyK5cKwREM+tXBD1VYEfVGD0FL6iCE5fuD0OfWeHdKukEbSnfwlaSTGXy
pJY/Lw8GIrUT0OIG2n5B9D0snrZlZKVU5Zmm9+P0XFHRVKMA5/E5AqkY2yxwDibcumbNAJa4svX2
++UbctGH3HoTljuP2ou/WINywKqAeAXy9bjrbvenYB+rU4P1N3JGozjHbru2CoTp6wzj2QjVGs2F
H8H3+iBQ6nkIoVVErkVz+xWvzlU7Jz51j3agah3j0Ykx4fHHfTbThEYVm+C46JpBAqldv4i/E4qa
fnqtFVeWLNrlGbtsJ6R7F+nIPVMkQoR1apZ2873WGy/wcQMijQKRNhqcdFsUBnZm5zhhq99fEvro
s5X1jpAYbcaM1TgDzCXbOTJbRjDAQDZGKNf68j5FZN/+RhXbcjy3Ze04iFUEJku/oYy+vrFOiuRC
RtAUxxsv6vOkowXfVF4+TJNwwUoc6owzHqRMZlPBCXL9aRCIRqUY2HUT8Cf+8/2Xy2znChrs0vvF
tV7HNTyoALj/zr+ikkh9WrHZilWpUdLgB624MNt+I7Eva3I9QINiyRsKnG+T5cMHj2nQnaAiiql2
QonL8J4+EJ2ghtbrUhHEXemcBaMvfDB9JOXjPjwKxz1L0Bz/8mje5pA41zE0Ry7pTFqn8ApuZJSu
pZzD3DCgzvvMIMAOnl6oqeGMBjAHyZDf/NmrpeT/4bjl1Lk1sdkFGyLOi1HQw4UbjqLAZG7mK5Eq
TeuS7r4vnxAomRPmt4B1PnamWgNjQiWhoQeDn9Oy0PDkW+pkCL7ILo0l/DQYha+CTamuTjXZ0EsP
+i98ibOz8d1Kv0oa8Sig+dVGJU5bzJWq/2yCS4gSrqS5obdE5apWp0iItXoMp406gd7xupdBAyDh
UQdc4v1F9OluxiJ/oUbfUc+dat/CxpkAprL7rdYpfLGGQNQLfinUfBoTYzvSd9fnPK9vIn0XEQz6
NqYwgUaMjvC9S3q2ozFaL3bFOFaqBFqkeLqztu/hGvQhYk+4cNWfO8yXZoNHXCjrnOVmSa0l5LLa
cU84PssbyElLei7+J6d9tdOaKggoGjw0o+iGV2tiK18bstqr9z72Elfv3vzJU/pedAeo79QYmc8L
6zajsfFjWoAMfbfa0UK8aAGaYFQGEaXy2p3U3NTnlWqXEMmFpjSz5s1WoouIeOuDhhJ3FDk8/m3E
8J4sZce8mOmG2xBnjx3hz/NODlwxLF3jPQPldIO6dmHfarTXw20S5Pa83+Q0p+cK249ksFm3LBE1
dVPwdVygyVBCVAPpQXVRAY7vc3tLnh7okhICz64iuzx3h4aH4tuCjmxCXNt7P5afvQryTVXEFvUn
gpxlkbR+YuPxJzQlQUgUIpGTpQR8kbAEg3dBabpq/Q2B+sTvuzistVBwt+TV4K+cOSTDobsFxzbG
o0bcGjnsnXrNmBiDSO3gYef9SpRCoxCiwCHiXx7BZEiTDrqqH7InZXPfAg9nquCs6uSwYDAhbEC9
J0DNBiqo0JcBSpFGJqdxL0E8OO1iE4InPmWPe7X07h2EAoV0q4DixO5560/1Rujvd0S4wQAK1Ju1
1rThlA0qyhULFDfVaCFXsnpM8VjDmUTYb12RI8oob9qEY1GoT7h2o9mnMB3KMrJHvCAux8A9yfnm
3CL8bjvJXLdKHXMejCCpdxB+5Gwfs3nZ0Z3xNu43SuJKv35rvlLW6aSGhnpf8H72CCpVIkmzKvJj
z99QERqzYxU5E1PhdhWP+Io2IwzIJ9//gVF7f+YEuaJ1MZ6enOuETRlw6M1V5N5pIfwiaWCCqvsL
9NQyxlvnmyhjrcq+GAOBL+hWnxZ/Zq4LBkFctje85OkMtnhpcjr+DwVsy2s/o65RlBN6QzL1iGsm
a2WbZPTylbgWWk6VQ4LxhLhepQ6qjFaxPV+on77NYDPVltZKdHLTXOI7saDG3DYi+DMeEp8hP6If
+Y/XNPE6g2s4vJs1Hq4PiwVt+Uoi/637TavVbvZ6zKZDJdF1kBnYY/pXkAzY4ukON1UbTeKCcxQo
O/wGzQGim385aASEhWNIUdwHlkwbtwCYvB88gdV4G83eWGPh09NMevDRNCorPUDhIbshzfD4mcxu
4m0ysTvy3skZ682FBmpxtXZRoXxjR7cnZK2hO3nuTPaW6g05Q9VvoiUkhAjI3VfYvf34dqHM4LUb
Yda+Vhe2l5LSNm23sVNrYt0g+lKOMP5HFkdWf5gf/lIXu9ykW8takDTYfQbA6mucREOQwcPZmw+b
19SOscrDw65nSVCv1Hv4pK2jjE3mudTcW8W8Y2dJF/x4rLi2G+pEkdeaeMtP60p7lDfmQT4jHRCr
zBupHW0SwFcTdrrvqa7hJeufTzUNxz5d+DeMKlvh1a6ePajEcWNOuwZkSsYSUCwaLeCzDZkbKR6A
DAE6ywpyqju/pi5AUAc8Dsp3/cmLqePwGG2yuwQjHDRHr/GJ74FlQfH0N5Q3bg8AMJWF+297JNKv
CUej/BhtWwRu2sWL1UGN/3+fD5bhr9fY8uk6zrSDVOMAITYqNSb2FWzVwbD7LIFhn2mende9oSC/
bzyuYchzfDyuz2D8sz5JLCVchFk86pv1HUSUDIlZoaqcKtLY8nHa6JhLWKV4/6nE8AOfLvYyiOSC
9aNdQLgGx6BarVimhs2JdQydZmUoF7GYbZxgbekwLJ1BMtcQgJV5cM7pqr5mdMCDFW5LO0Gk2HeD
2ko3AjW04AZWC/ONG3x0+0wMzo/KInJ5X/0rASFrlIzQdY1MXbn3TgafR4GRDlFo4/JYaKrOIeRC
k43vab30F3Px58OJSszCCrR4BK57yf6YRyCNLtC2UdwXPGN12TlXCFgn/5XRle1jTcvfiYi0/DyJ
ALhKM9PScHYL5eRfe0akYZfsMlGHR1aOt0BETPTmsE+Dqepy1GbIjwNSf95sUFhcTZPK2Jt0JGqR
ZV324E/LHYWFOf31TjTUi/jw4P5LRKoYVSQ05mPaU2aFgLxlqGSOpEot82Dh6PFLRQwNhVNtolmK
9C839pD/4KohnQ9CetisILsY4OaE5/KdAEaYJr6O03woV/TGY9isbI5bmjyoZ0rXGWyG1UxXDF/p
qqF05pLFTRzGrefo7nnXHT8Rfyf5heArL/+x6gtitPlZcuqj2iQSoda/3tChII/X0ZlrqhkkF/oj
kWvm40kfosDiOPY6X0LzLr3bN+AIpuH5clIMXibTXIv+vVSLyAYZUrb4XK0sDz4BSgeCMRvzecnh
CuX0yrMxU8MnMvkcP9gfOrpLVkSby7BrF4u4+WIyVWc9PbwfN+ByVI7e9bn1RgxWqOR6ifR1VRRO
EfbNSsHgCQ6+Iiqj5JUJ0di1V8KbwDhyncZ2WhckQkXpVuxBukA+IucAE6Tm4OQmjFr/bGe3owIc
FiNK9n0A0QjJ+kP0j+2x62A3l6903gPY39I8cbUTOhDTYiJcc9MW7DykL5xBKYsNd8uNWb1rPY9X
fIkPZ7R/zHb8NloXtOL5iNIkFGxGFi2ONIh0OzHrdU9r//hRbba6ljN5oR2G3kJIAlDT9r5z3ult
y5P8kfqZP9JJoWkZzOQHNHKzwxea4NztHL/wlGK/Lk6gxy1Ogqkgp71bq1SCAzO3fBgwzM+gWtZW
UVVXrz3Wg9yIJM/S7OwxMxPOBaFYDVgcpobgsAArpHLEyeFpyaJk4qhztlhFD6Bn02piYIC+sG3t
tpaRznyepNnbJ0wlBDf76K9VYWmVqNYMKyfOCX0eTGeaRZLYLeeMVCPR4BRSuK33OaHBXEpk2Ugk
yQaIwi3jiGWj1/vqWUWPk7cNNtfBpIqci3IjYjTphoOgaWSFTrHiIG8c+xEXcq0Ja1wBmhK5IcVJ
DwQtOF2sYFYyOIgABxK0a+wH12MC4J/SMSn//X7tTmMhbkf4YpgpSBpYz5Y1PLUfNIDcerzkM5w7
22yvtxv3GMnn9JaH80Ea4k7OOS8zRNUb0PgKnTi7q//5ozEVy9TC4T2cXD3IjzUS44IziFruV+jC
SuPtTUIsK9B27fk4Cy+V0NIlcBN6exOwR2ETAIjCJDpa8oxAbTshMjNs+EmUYQLXUNb7KIwwAAYP
LZ6YU62MMAna6yvscvR+Y4/KzsA2/84OMaDZuUcZx3sdoLk1emtEAYz4Un57wEhOkC+W73OnFk+g
Bgz7jcDsP8YLm+9LVZAnmUJ6YUX+HSQ7BfJSxrtRjT1KDC36gJk7wYidYKRIbZP1IXWa+wGtx72D
EpgHgeyj4jYpKtmTYUyt6tYLBL7JaVhLNSt8MYzN80/wI0NotrclWUDORUW6g+ebczbpH0qdu8su
fuqCje6+Pjad2vrs/9U5gqxXKkA+uPWZX7VeXyJqCT8FXZwTEA0bxlg2U5C8abFrj2hvVoVs6BFu
2a/8vZjjWLwosze8f9vTr7/onFGYguIxql8FEBGKAiDjn/CCKUte40WASZq62NthEsp64ev5Eg99
QNnCdQ4a7Hp1iLCY4T0K1EIDCujzAGv/XQLtvfS/Eg4h1hpkYZyMiXnt/yC71D10isov6bezC/dF
UljHiHfTpfSaZdcu0BJj1WB3gW5A9a0vu8yAWw4QYsIo///Z3T+LWeT9OvfLVUPEhQFYi3HN5OK8
NCENDozVDbV43p7oiwOWVPFPN7Veg19B6yk6+hZA3a/CZUyMa2/ghvzcWLjp+QJrI4Ts7JIJScmB
su0H1mo8A1gC0NqgEclAGNjmi212lwcocO/pkjy+7kfxE1zQrY/rEQiK/8ynZN+58UdMLnwFS8Fc
2ufVV02pg3TlVjWQRQ07d+NyA3fTKWoD6x9RAsyOlyUEqXRSNcyAdg5rvTZqMkKMBPKn1N8JX+9N
T59XD7cmfVMhjrOZKMLu9tnM+cMpzIJtsR26hSxfbZ+ZqcjtX/z/FQ94Fo0Ywz3CB1e0+ieq6xcf
g2tXf+ojAUdRifHFpEI7Xoq0xqbkDYxkq/Hl5BM9F+acy7eoySK2jObvC+8GYdHbQIxthKilLcGX
jFsqXxcFWiruzmCyVCtc3lH/7/VdyrYBLsYDTyIABAu3M4IjrLeaC25lL++Vzgp7YSy1esVEHYfN
ZqS9ga2s9TMa8EYPmNGcgh6/TPpHIzparnolUrhv4PEURkEjvA+GFyvpz/hRiBolY8HcJn+vSXBY
eEvvfM3MvsMqo+QICA+rrueHtHvw+l3InAajEMITgiM1/cuyGxv4F2Z3qWMNgck7ZVAj+yU3Ah+A
4xWLG1lGC7TMfRn/XRZ3uuXOknXkyS3h4OwvVWbs4I3Us/U9rq8JC/DmoAr97u68m/kMzWwzyKCb
DKPUyAPdRjy3wTXf95A+YX4FWvDUQxQ4RV7g82NELDvo5VqpkOkKkBZxj15/CrdjpMUI4jMjz1bZ
132dGl3iq4p4hr5t69Pvf52916m/8ai7L5eAZic2plhO66JMiAM1ZCavKz8qn65z+986UlYcUnx9
cGpCFjdeemVromGLsra2FTl0QUBLuMxnxZfv5qLPe3NeGHb9a3jGuAflyAHkIX09NiQkATW3nlEQ
jo2RefKHEmCtOiy5Ao3b/izIs+1f8+WTbzAtfv5b2mgnh6gj7/k16D+Q1HBUus90xem3sVnf/IJV
GhKTueFU3M82vKhW6UN0jw8gXE9bgQMjeh74Bkkrsb1+qmthNrbgxZ6A0R1/euCHnHQIy9Uo6UmY
EMmnkNcSUMxdiC697GtZWUganEXVKy4hX3TDQJQwCfrEBzq9UEvS4bgLD5gcvmboEDlJvrAbm8Gr
YrPmfBFB5NNpfZeKoXiZbVlsIKpMJlx/YBu6YDZVLVeQJFsKR+gxsPTm0tFRNyUaEJ/1YZKU6F7X
qfgd4SEPTb9FYKyFqjtAT5ZV4ltwCsokZxyPULbc6o+mta4kS7VfA12lpu8L2YWaocT0xf29DjIy
4qZMVS3q7yJvDaWNTcTuYRgqeKp+j659eTj8q6/yueWgIywU1QJnUWVRzqTb3K52gSuPf4hhPROJ
NNKFQYUd1lTuA6NX+GAGK2oamVBz0h4IDbtITwR756wElI3mHzwkG7BQljICG+6mAzibUrfc4Le+
hRivgZ7i6oVIs27lzHcA90MOOquPSDWEvEbbr+/W0nCvDIUmrCE0KYdueB5sfWuqkVzqaTIDIwFI
9DV5N8B3pe5+1BdXlBse5N71QkfbzJFYUZSpMrwj3kSh5z4uSYTkAjNgzxKaKgiZm9ARvbKQTHxF
RpvaJgM4FWRdJW1lRfHWp7vOiihp5Ozg7ASCOfvTgQx4VWpoa+RteBlcRGzw3EiIVih03tuni4Um
B26x27Kbv9lNaKfRxVb9opok3E2qvTIiUeaBBWZedp9DeuNqZzoIBScIhRdqFeWz8k6X2AaQXaXG
Prrxv1wF1qaU9JMA9/B/e9Fr8FlXlw3wU3MBe+eG+4TWYEg/HyxW18+LZR5jFOse9NpSoL9TLq9w
GWjuh5hOq8xfIYnCz0EEd902zDmXGkf2PvhtMJpghzOy7AGTwUbvq+FDGglY3VYLwlzwOrNiXdp5
qAIdWjXy7yL+UFlzRLUsULS+yRkeRrAjsmA+WhpCsl7KW2kKzolrrFZbAV4gnP8s6gIFtXk7zzH0
358G+BPzYYWyf1NSHGcQ3pCR50qCMGvVh1l6M2oTgmPSIiur8H7kSGLY3bIefhHis6QH773N6czL
k/PwgplHjJhW81OxiOGBbOTmoXRWEQcmJn7mFZjMmrMLsKG3iZe29/0VLeue3Sw/rdyyKLozYLuh
LznuVInhOyDe9NQlZxDetB/iu5BvDunFPXHABTdWNSeVJy3u1tf0yKQZtwW2X/IYbvSFFJybWjnU
7Ck9pQrmUKfPqXE+WrdBG+YgLlitMW8mr4mIVDLvUiQwbqUvaFn/wlYZJ1yIDC28nlLoaQWDonfp
H3uj1dKh7nZjJ0d+ZkW1jKlFCRh8JLl3EAvH9MzTRHewPuBvDRCpPFqhaJZFQgKLUrDArLdugJzc
C6WzvJnvKn8yIkmcB9TENzBQjBGAOMyjfQeqDCrPC/1dxWYpoBITfF+yW71hQmxs2X0i7xgrU9n4
+bHX21mCd8wYcg2ZpOHYQtw8LblthyJhBX0qmbO063TJFSzmAbn8WqRR0kI2Olr8iGjdMJRnBvWh
yXuq2DTjH2PHiCrFTUvoCOMYq0fG3BMFfk9P4lkfeBPq/wuaoin5N272b10zlsk4IkCXoR6DWkUj
v2coqHxWCoizSaJsd7DSCnM2EjWdtvXmbBfE6xi0xJT3bW4JzD+ZEJzrgjWuoAwkJqqkj5LUI2iR
T8UJ5ucn4JvbcJexFNO+GJ8g+fE6Zft/Tv4cV/LqWx14+x6V/u26GQ0z070+3sjscKBjvfL2AR+T
bbh6X5YV6rYov/Gl7jX6WF+uo0QArIkZJcJqglhym02i+Yr9sa1SCPu21A7HDmT/lLR4p10G+66Q
B07c5TJKsjUhKqe0XypF03HTafDttxrhlec3I0tcswGvFdpUEtf3Qh4yQdlRv6Lvwz6fY1MOpOWn
bftq9GP5/FB0hBFTMJ8RE9BwBR3ma6Nd3+WneAD+fw30F74vo2fCzXP+6o2ZqvLewdogKQ0fgXqt
4TJtrx4EKzy6rCYtZTF1eSrlHMptrF+d2p5qOjwsoYWapgLjs7Zo04k9maPCyszIdxiVTUj6XdTc
xYAfOHFmAXaB3HbG89iqJGF3gDfPY2BB+HaBuWVuc6Oosf7+QVBYpCW4Xyqdm1wBoure/JyEDSsb
C42HdfZYjtSNrF/U4SSlz5u8NgevCEACglPvts5kTdZOg3nPgnd7rV3tW3sAa3nfn8jA00ZmC8ol
uJAWcXHseyUQOtIM8wvEWWNCB6+FiXoaL8QhjkOWwQ6NX6mU7eFCDktoj36AH4jptY7oz01A4WrY
Qg3ccEKEwfAT3WctzZxlGRXMISqYzfp5DkyBvTW3Mla5jaIQD8zBqu3eg665glxp87BAE0rzn4nw
fardyK5sPfNtHU4uCmV12H54B78m5S7/J/TThx+oBWfRWyL/BlPKMnrblhc8orOCBMpdnO1HUdG0
PdDqyt3I252G+mFNX6OPL6bYoZ0aTNyNysh1z7K2eEiRnqpjb+H7jughadh0cs4R/R3cAiJlBNe+
JDSXGCT2vQsTkm5QVkTWcLLACEWl7u8OVlMXcpKtNksVyx//4BpZu3uYt7sm6K76SZLsWl89+B3g
y7Z2ZxefVycShf6M+gPxlZC4Fihq80fq2gLRqY+pshRf3xTt+2ykiQ7fxawSqpUcBg+bxnzjGDXx
SeGRCclajROj5IN1iB6KVrcSA0MbCUHvDc3i59zteefHzyzEIoc+OYtjL1j0jpq17+jNXjxzSB3B
a4Z77Q7KL9PX+9dvbft6c2xWv31HQAzGNmZ9sarlZwnqpxECleW/CwP9gV6jl1eiG4hp9XNdhwwg
ZbM9lSQ6QN9JezAUgMUwsRL1+3PTvNR4YnJUjWuZZJqtILvhU24/tOXvLg2r4G1gH2P5HDKbdbDT
LTM4eJFNcC2eEP0e2Tkg4C9nXCXegpUC3NSaSWVlzJtuM19EApLeVJs+CD8/UWcKXP3g72lVE9a4
Bnpy8ArypfRqPc3iiVUmzofwbzqOM54gBzWeJdj7ttJXvBUtL1YB1MAop3hqjZczY+QU/c+ZUP1I
WHC6DLencC61TruCcHK8ceklHdfptVv2jPthGNYoXM+cUkZOO9PkFAEnuOCwQiYj6bCuQUQdD4PN
DkEU5CHhKkGpiYnZzMAnKIIMmjImMJeIB8T3gOzxNtNgDkCExVMXF4Ss2XSCBPuT7prxaEdfK8NN
cak8QE2V22JcwXLouxvyhc3mMM2e7fz/TBzJo/jw4QjndUJFBzg2yLJXySxLpI9hy+AlLKwRi/PM
A8eDLF5XbZHPVLPtkCMr0XHSaFuwy/Z9rIzY4sM/WmfQuH4q5Lnhjwzx8usPXSd+jfe6TIkm8QWN
AlsyooY4yiTbOpG4JT2yod9sfOPIF1mVDrW4SEsA/ydY7YScpaxdb1LFmRmHlR9up9QchqqGvZho
XLE7GYhj/+mME8+XPoqB4Ch77oxA7CNskdEr93OynrYmRB/DQiUfjSLiOC1AQAqfwlCtzx6ShRe2
XLKXxDNvee2RC1G4P6uCEsDW2JQoFw2Y27nm88YsuxNlYCQfpAolX/QDVmzNnXxufHdmAYTKCJKe
o5QpAbhVTc3B3XSvKdQgttOGcL5us65QNFZl0PTu0Bnv0Mog/8tzX6I86axY496tTAstkz/iVSHW
i/mfZpoGVJC9oPC21bxkan5HnE8pXCLqSG0pXXAqJn2Rv0MXMhWknv67i52+1+cAmumPkWCP6Wn2
tn5cUIg3F+UP5OJZSjOZz+JSUKjkWBa0JYd0/qHGm+R3DaYfHbsfEWP7fybZFAV59AnyWIA/Xm3g
bTzMyu3m93QoJRpof2u7TnzjQKuj7KmEinbvYFH3XqG1Zq+6HXodEdTm7OhwbHSCa2Aj4Wer59lZ
GwTQPemFcFCoJksDUZ4sbUIseAZitkRVvEOB+3DfKKTgD4hnEf+s9nQkQHq/6Xznz4UpvEDJJ5Al
7ynljS/9ZnVPmv5eSGzPAPuewBEfXF9myBzQ7bu/IBr/kkvZ+bnLiwDvV3bu+1p2ELnOfG2MfJ3f
9zXZyPC73oq0gSecqLYwtpixTLfYpdsxYXds93NEcisfBMGiciJnk0EEy3CF/KZXSDaW/Nj3x8sM
HpK7uD34zkMnNXE9LKQDDBPj6ue9ee7Dv4gKHYi76AWFKBuqEG0Up53KB0nB5/vHOyKa9L1UrkS9
JL9DcQOigpMNoVb+R9qktjfwSsyCFNqys5Amp0X+ploYNIyEBOrPS7+z+QujJYtmANUL9hMvcCfm
hV1KciugUK2uTJAJ365WxFbBFiVpVkZIEqR6vptSkGHkyDHL6cQXtLgWxAkTAP+Flv/SfvA2HJ0g
pNQgFR03uYy/dnyGPg99qBbriYfftAKW0dOepixLIZ2rPZBesvsLfUditI6/Usxr9UD2Gofv0TAk
x/9QgTGm5gMT+vT8aPfCbSbKcs3Z0sxZPxHanM1Pi9ixyh0sU2+0zREoIt2DeuKpCohIqPo9W4ef
egWb/Xvjw0ds+mZ+4DfbbUDK3NZOLain7MWm2C8Ix6ai7bPALDvlsyrO1QqLCmOmTnIifzyQYUp0
o3if6gpM1RIqoTNvW93N6sXzsjbXgbi5XAZ9FiWtYxozvoWP9cE0Lneg69d/CB/eg32IyIOnt0Tc
enATEG+DOevesd2zwfrpvW3iXF8piNWEiklTdJgd/1TBc0+Ku6V21dY5Z2Zki6MZhm2ef0zAo8d0
cD6Ja2l1k0X+FWL/bbvXPYSluP8vhAkcBVvQ+yH3YNnmlcHHlc4GWhCXs62DBRJXFwf1PowM/c3e
QtOwY/e9Yb62E7abNbwpgD58lZmFWajbEKRxYkZ+Htyrmx/+kVwNwq0EQxZjre68qynLPNh13mSl
lvP7fVjypxWhadhX+O0zKvFjJjGSMIdGmQeCU/H3r11x0zD1tdI9c5N8ZmANSgPy3whWkcVyZBe0
ORRvLiM/4tt4CCCtyhNt1wbWt3RVcQGUx5nC7s+93lorgEWBkb3UF52EvY6aYivQv+3mjRcwjLKr
hb+k3/pSQ+fJ01XwTHkFk64XQ8KoJSfKUslb9Sz/5KCRTu3ycoVfwvR/2CFXLDqK6gpT1TQy4ta4
DQ3PchJ+e89Dybmp5uiPNMlqi5jM033sch5fVXtVntcdW85Skbs0Xdz370gicvW1+HQwwFUs0aDW
sx1J4o7FTllp6itOnLOr7MI3bTMIyZKp1u3yklt5xXqaeUxgJHzUr2YPBz7tJmc0TWClhQmcICUu
W/JLA8G+btflirgK8dxpq/P2Km+2cKUJw1YltqDhItMQhoikZ2VJB0cizuluEi6Jh/rEhb/i3vX1
b4yXq6amwZbEjouyjK4NLZbTnT5ZTJ5NkUVXjHp9Tfn0ovGQdQ4vvcWekU5Gx/ncgNo8AOl7bJMi
PPjKYWrp0nl25467IGLIPilBVcLxxcxvTa7Ea4Id/uhJSrnnz8CvSXIe24OA+MSw0mEauAcx0rDc
IkgYSyw2rE7M8tVyCUOyqnFrOrLYhmS5h2p+i6cBUSm7Mn0XHkaKytvCHLAEuFLPB2FFNh38frjy
0pfuNwQFNF2WfY2PbCCSeypF9b4IdjSE3Vydadctc7Ve7UNIg9eOu0jPX5UL+3X/iK6PEIWENAcm
8+p63txd/E86a9kg/Brb4/+f0PWKWv7CNJuV4DxDw1QYEtU//lF8N+ToLQcKuv2AARpUkvwsxzbh
ujvMJ7Qmwf/lZt81Uz689mf/6LzKKYr9uauNosSFJjvwBVhSeXTg9+/lSrpQB6dt56fdc+RT5ifU
Kx5JO34OUmNhCfJHMekR9BuTFex9Rn2OSLUOJvT6UbLvpmyegX1rC+D+Qmmh+U7+JvXWqdl56iyP
G32YaqTDrB0c5DJZWJfPg/ATfmFxmzwQpYOpju/uSw8NtqPEmQFeZMl3YqRYW4ThkM3/gudH+JG6
7aGPtvMSSXVCfITWGK/BXhY3NH9lMCvhXPnv3dMXP5/lgsa1hkpJ9UjfrGDqg39Z6ZuEFilgt9Ab
5BHmXN8wessT9WdQ2t6bRsrtj35vyQwSO42w2NHEvHuNOJgZE99wXIc3Sd5R7iJIeNQ2RPcuT7QJ
HUwY1bC+p+ubdDkhV2+DVtHFwtv3444PCBHHi97n7LFCg/wX6nr1k/GYbKFiprMgyXFsQkbO95Gx
97jZ1qx5Y3wr7kiRKiCPGiTrz7WuyC5Mq+yJzDc7ntBhA3KfagsXoiOmmNjSbdLlUVUwAI5zv+rZ
TL2DbL2R6e9KGeVNzlIwovVLcM8C5aDCad/DXTJeGOiQtq6w+orqBkEQGeXgza7TEMUVhmRA0aLd
Cd3gIRRQLAkjDmBaI6b7AIfPYXI4i2ETXPTWdd1IrUQ2cNXwV7hueZIBQ4xLced42fx43HOGTbk0
knF8IHIs5tccWUoUl/QW/OhpIGCIA9ATtAQ8i8cDIE58G1P4JycYnW2Vm3zbF9lB4iKDyWT70Id6
Wl543lifuVjV2DCVs2hgI6fbmieC6i2qlZjIF3HzDaGo/Q6ns4hpiI5YK2/cCX8y/owIqIj3J4yk
aWeA2daGt8ZwrqwakBwxhRGHdXdF9+dQAY1UsYs9mT69+6oMHG46sR+2x4Q3GuFJNgoVvpvYP5Sv
rA4WprVubYsI+wnZBV9bwosXNn/0ePRXXTkx1fljulFR5PFLkePsFVB1eQ/bidrrQDjLbkz8bWLE
TmVlpdm1gCdS+DjKMp/2rOQEWhyFlr1gKplAPqgR3y9bkOLXUfGX0M8WSXWuQN7x1oglFftFI1zS
fQQ92Wq3RIc5Vkhwvsjgnojlwr7k9gHYpRyiNcZTkgpVDE7JSTRAqbUbkhF6nuTmDIsef2hQhTZ+
ZIP1G3DfYRHFOGkQ8+b2pxos+aOZ2HVJt1XFQ3LT+bwhrekSPO5PHtxHBYY8O3znlwyhsn3AxWSL
ZCZ0CxPUhojX6P24lEsQuHD4MhkpWY+dC+rQciBhFCXkjchbz5WrTRT5H7t7Y82XPIsALN8MWlSM
CffeA2QQdOl0knU4es0iPRPXAXz0Up9LzTalY4MfPS2OoEs3W6Iefn0wDppodrWXVbnXakix4KM/
YSbEqo1TWo2NZQm1GuFK49ZUVe4fekrHLXUdiZYapPLsZmdCMSjXhmsMxMG9l6uohii7a2J6rcWN
0u+oGOiE6WTasfbtjtzsbO0rGif+n+9qJ4lzfuzDMVaOGhIXrnU99Y4OKENmCqifY+lgjn6VtD3y
4NhdAV8JEWoIgnavkl7lEAYEPfwU1DT55Q5+LGr3MBJXIwM/vIXGrdfpdSxAckxSMYTDK8x4GIvo
IAE+L8FysEx2OhAHxuHfKkLJC/bKQy7YEpFwHcTNLxGxu6xPfFCo1HxkVm6gFFYEwDk4b66qGr3g
l2ZN60IGT3TrGPg7e7Q6VqT66aRp9tNWFpjx4A6F1LtSF0WHjfEehaP30g6ZRlq/T5u2w0t/S3E4
uE1wGeZFG7glYXRSJtqzdGahgvwivdzXVXScDZuAX/reKfoyrAlRrfpUWAKbz+Hs7wFLAR0Eo8kA
2Ra9WDHMqrhO2lQib6c9d2GOvVauYSF3U4dBF78ldr6wcMwkhu7In8oqKFpFnMgNSnTCJ5a0wuuj
do4LbtKkI8iFj7iVo35zyRBZigNLrT0HondEGUp7JkyByrlg5PS1pCPj3cOqUAXC+I69DP/52ter
Ng18TJVTPUjJBHj9mT+98u6MBMTDiAaq9p8SySS4cxItDaobG8CGvHFJO6YbPvoC8izcT+FQOSuZ
UjVB/qwdOeNnS9Mhd4NiWadAVK6in3/ZlI9jHjpb0IPpTOO/Xkg2qQgK2Y8PJORZ9DJ0yQJmThiv
j+V1h0tHrns/ruryyWGY16jVnLSX9kAGfROqjeVX98lGKCz1q+Jg6QQ5FIPd8ObN8dak46XkTnxj
OYuR0d+i1xTHS8Akc7zji1qv/UMKh0AtoqurFqWSWZQBvVA962hHRstAa00JtT8Pb2nRkk22qRAG
iEgP2qOpXtg1XoKW9Kt9HRfN18enF6SI1TaMHOyW+507QieNrNo+lJmn+ZmGknL1B7WiCi0ocuej
m55fCXPN9bgsNYFzBqRbch/m93bBCSGVZxNKZ9BBAre/dfTKpTmbvMLzsJG864rukxUW4naPr48W
r2XdEf4vLrfenWTuipqi6HEhXzZCoHLDtEREp30YsJI4yhC0oiMThcKWR28ZnsfCFiIQC4bVj9Kf
34bsPOVInth8Pv0cWCN4ofwOOxCDLYPW+0LgIPx6RrJV4hItAWNxvw+LmlcjMKTArCEx1L7T1o/6
CuNiHHkeJ94nP8ol8dFvtgEKnD7jFCaQAzonP/SNa+RkQinISMr0iPTTQMe+I15s9KEcKSRb6p0w
O3hOFI56Ji+01dVFKABThyM0OHZZuL/mstfrXX/g6it80lJdlZevefkuN9i0lYCiT0KqUS0+BaqK
+5LUCaA7ciOOy3vCIIAc5n0g7qv4LkZDp97uTFrUnSf7hMkHNwd6ouVSGM5OzYtfsFah99ccYAO3
9Rzc9Z7mZ+7mjG2mZh6EJ4FQdY7i8LGDHLh4ks4VsZ7ybl/un6mzWelu94BlqaZrvvg03GkD7axT
ZwyC62zH7iQUG8lc21yqc6Gaq9wISWvuzSXWiwJJcyfau67+kKdfXT+iMSADZobgldQibvNhLOyR
sO03AekVjV/S+p8aLdgr487sgE6LlmMt2hacbWcMcy1wZ6nYEAx0+9Vjj/QFrZ5bSZfCSXcCC/35
3DkpGGEHFdwGBwm/0NxQnuZRMSU7SETYgSCWLGUbm+i+u26gCoIkwDavTlyD3ii4axypPst1QNoU
hjhuwfvEWKTU9WdsC1Qa9KZzwucChynutLnIE5HhL9SO/Lx1Wu4X58ZNOBqPPlo+APh2vTbXL+tV
IQW2woceIzrlG+5klMWZXyXITDinY5MYVYoCfgJxY85PbXrSo9mCLV5kdOvYcusiF/aHZIp5DPwC
/9wtsExZUhYGW5Xv7c1UohSQn2CVc+64nvKX+5RG8M5Fsr+D6dn6LagQPkU9nXpTEI4TUc2eVLgA
0jmyVrmgjqHIMEWHMpvv1rDZtKyTgbva/6Lu4D9XfKGhI59KEuVOjgpzIg5lIahbNEu/74kfb8FF
wOUDIQzeZ736KAAiX/rf4JkJJS77ySIUpp74Oc1oakS1mNfhjA==
`protect end_protected
