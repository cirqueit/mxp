`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25696)
`protect data_block
NLrGrNJwqR5HfD9a6MY6ymwuE9vpCdQ3ZHSm0JANIWU/b415KOTE8ICWCGY8ReQ6RcmVG5gWlz7e
hbRFwXdo6j29szpyl/xB3zcgCNJ6gKCkmD1K15b7s5i0uI6jqrWrful3ZtzqkKJxUg8DlTgu3jy4
wEbsdudh16jrJ3OGrb0YQCh1DZVAf7n9V7Lg0hzKu87tgIT0Z7pWLi9knQ13FioB6oTRyXcf6sSL
IZJHkzBtCp3MbnKwBNST53i8G7L2xXHDnCiXU5vRlUc3egH/COIxbZ+oRnA1wHsYWD7/iOH1zeA8
x8oKBVEctSYvpe2e88W9I2Ax02GdtNoweNXiLG0HG83mt1NqQSP1mUc7fNCCFQXg+8YeP9z3UVHH
iAOIQApdxmTPKf5v+Tgb8alkR2xNLDKH9Df/4MiaeoCJMh54HD0SKae0g3ilWpv1T6YTrIbzwYZg
u0X4tVqTqEy4o9R21LwufABmPudkWvoIrIxemo5Ri8UJceMQlOT7napJf05TEusVpWrWOJZeaOPD
FQd5s3EIeEY5dzpqoxlSZszyWgbTRj/CEMI46Y3KOAwpG49A9hmvjhcjdZks6zPUda/aEarqP9xR
+d3M5xxyvByZ8yUjuDtsR7PyAe7Htes83Ij/blAb9RRVG/icSw71Q1cTwk2Xm+9NrT1Tt/+hUwMM
njTWrBuYLrC51VDnReSdnCgow0TqWFXJ2HInoFlNrZy04b9uHwpoSHo0yKj5KDSXK/vrmqxx0ZfK
66xFvG2wDS0PRrO9AdK9XIEIDJWAGV2PEkQdsvo9aAvLUAFPTtzGm1JbRiujrBho+M+nTZvKjgwL
5Zt2E5n7/h+vlE9YTtykou1GS8VRoeOc9Y79H8zxxqdq62YreV8ASucGcmuPxkPASwFQ5nz+/Imu
vIBvVGBWdhyp+5R1LssxschUm7NpHQEGs6bvq29EGV0X9nY17DM49owTD8ghoXTv1TbaMse5uHyM
XIWw0CrGv/4SksdOgvmM5F0mvdjlE4a2zNtwymcqPSd16wnsuL3rABBGT7wPisJiSlNI5kps0sAv
GU74Yh49AWn4yC/BGOh7lXHFe6KbB6xKYzh2+tUy1OmSnuc9mAICKhT5bEFmUJZsTwVFXiuHpGa5
a7bGRYduiIn/TgAzdpEUYN5JQZYhj+tKrsrat4ndZfX2C6yDMnVhT6smPcriAQbU2eL8Kq0EUu2g
J+Hsitm8I1oQTZ5oBxvndxgY7CybFPr88a4XOsNmcX5EE3C386//nPjoO4bJt34WysBaD73tFM6V
8tRwacvT9VqflHfaZbqHBKQRQ3VGz0vTKIItIHCRk1G8wb+TDNhiTyjxgSIiswBes7g+Uho3u/CA
XZ9SN44C7QhkRDxWAxWrZiEK/Y5Wj9M+o8Lz9C7d8W7hZzWdBQs5HeqEmDnIbRWwMYocGFlHoncv
WniA44lYL1dCabbcD8C7OsyAMIgvz+3yrUgvJ2FDxk2rzZ5YjrDps1hWhMBGX2O4S0K6XUqPR6Qg
hnZrKWS3xCL+GgDpu0GG7tc1pwsoFe7HHXZJ/xeuhQNMvgEhkXVeWZ8ZbcXEplUgDWJ+pS2w/Riz
3Xlv13TwTl5OdczhKG9xhV66ZW4bsLVMntnVzN4HZjWP7TbnH+O7GnflL7PmOiZB3emkkph55dKY
/3ttHWWoDHbSl0ijKOOjS1kxalWn5plvtAtFA/sahCIh17HUr8QG1/LC8IycHJ37QRx2YxwITtaE
tBsM67wwKGf1zldRGX1Rb8KNj/Uv/tYzTOcLA2pWXRRa7uViLoWgXy6pwMehG+r4+lKcj473P5Q3
IFZHV+WVxaoYGLxRhs3Swrsmo4DQFjqd5KR7nAtMz4WaHhIFXPkAVZB82Ahmr30gjj5VhvYlK2LV
oDui6XD3iBEe3NZfRJ0M36XKn5KnCZ51aDif0NnQ34quak/6Vb02Zh2gom9ahh4FqUP3bFRCKyHb
j7PkPB/NhSYb7IwGs1d7bgWqcwXaUL25kKtE621CymjYwVnbncFiYuMWgL1uP/ExbKmWxFfA1qhs
fsRC4B4vTSi2ivwXmL5QqBY1R/WMNA5fz4NGp9cR2BqUnJc+9rKJs3yXnlBPLIkTc0ZoBQVX/sXd
s5c6lCaYAWNloihFtZxdhlSzN0ZovKrja0egtXobdxhBHcGHj+yh/Mqz+R5dt8iJYCUJ7uc/HN85
CrvQZd/a4G5+SL+rEGtBLJlZzHtzC+w4x2nGa+GCDPTOnQIjuTJeOEpU5FTmgzcungPrzHZ4pqXo
jH6qcBFQDPD/ADw1vwBZGP2o4stHgSNTJLbeMICR3PBMmauKu3xbyzljl3NMSgBJOPlG7SJ23Oyx
qIIfthOXdwNwueImOqSEuBr9/XeyquNBeDfGE1Vo0Jvign09Eaka0Se1R0dIj+a9lDdvGHgR/gOm
R1Eup34qZqIGgjfA+AsE6mGEyr3a3h8O2IbfPyCyVj0atALr7fhBU8YCNEa4WsZmhxiUlNk6bRa9
o0dCiuFF/ikYRxd0YDj0ckOazx3LTNYR4BTRHVP/0d9WQxzd3DqCaYYei4XexybN9Lc7Mpu8dhuc
rYXKTnfllZY00VKbgiY/TmtHgCZ3d+MxPIZFVP2xl7wgIoYkEF2dET2j7ywhzS1imnqCPwSMac5I
7n92PVtk9C8emMJiPoYFsvA4gdmfIptDPGCCK7LwZjL2OAMc4ezYlvVwDrOLR7mzR1n6LX1TYt1n
Stvm7N2/vFhy2zj2EqK1UPjXicTH0bcTY1f5WcfAKi5BA/+5O3GMAAbM81UOkczLg8VA3hc0MIm6
q7jbrN0sUuRhSVAnai8xXSVUrcwV6+qbvaj9qpJ/IdSRbWok2l0J63nPc013Wj4lnrvXoNdnHjEB
Gjd2r8pWEtuel6Mff2d92bRr+HsjU6S5gY+tKSk+eCyiGzCCwPhUkx3uuiT8luIesqxJ4g8y6pYY
z4szU6YoXTgwKLp9lNzdvxAPvEq/ogXhi/16XmpaqBBlKOGseSHS8ozrN6q1lPKry3zEAF0pNvM5
nQj6RIR/P2N0GskeoeRqhwDOtyvTr5gdeezagzNxjpHM1BSliE0ASeOa5sp6DaTTwBZVPImmXADZ
hd+b0RJxFLH0jfjNvxC4SZZ7QTq2ytO7oTRVsxNDCzCM5gjyZXHoHG/dRYNia15fReY9xgQnb7qo
a7tE1elfuZOPB9rL6ZaIfouf3ZR/1Ea1Qp5OUwTeLb10BCcHU3iE+4/OCgr6jNtdwzWShFxdehTa
BrAdikZNuwL5qgR+0SZsGOWBp9TYE+1PN6uZuo60wXSE8rYkqQoIa0w3RGKQUro+nEIUiK1pxtVV
miQ+aZ8oMydRyaauZHey+5mFMuEJwKx+Qp6n3IK/T47/l5Xqy/QyPP71hyUTS9Ia7v4SgwajFTPq
x5wR0WLwCbUzb6NPxdho6Pwpg1xfZtOE3hSWsQmgJNTEDB08NmfDm0nYIGGQBfNWoccIF9CBMrPb
mwODn9HZCtNxGcxFI9DfQx+dVFmS7MBBOPspz6hV/hlV755bepgeSRHRxWf3eIm3FPxOjEQuhhTh
wbkuBIsa5faYBW5u/n8pCfuFB8TpbcBeaIsb7PEtF3uqLeyqP+AhJRxL6fLbMqnjSOglpeHcwEOU
a8srRDNQUB+VWdf0TRGrlFmjARGKyKJhWBLYI7HGT3zXs+uN4StRyQoX/783KjTne4tW9Dxb7lhF
2XkrfuMNYZWUGSTgk7RiYxNe5um6WfsxXNuyah7IRrPT+ZqIIts+xgmJrh4o7BhWE9GVGedxbEbu
auAczkID0dcSckT6QMKzVf8jnFfWQC1pDjNqfDmb/r4Jfn8iIQGEk4A9MJbaQvWwQiSo4qsWM4n+
V34uRbSkYVNhAdynT3hIx973XgoHJPsV8Okvz83J0u2nwleQ974mjUFnQEVosHzRhpNfP/m6aj9P
oHvsXh/XgqQ/8Ytp8K2NTQbo1tzQ1PMclLx55oETX/8FskNtvDjSt61JWhjDukMZoI6RqTudu2Ho
gLrA5+jSEC4u4bFRNX5ncDslY+A9Hx5/FSSxpnt+oN5w86/SYLzHwk1FMXC0630NXiKWWig2BZAF
cc3plgSUWwVpKeHL8bC1VphdDOO/2z9XPPmUGYljgqhhbiXxR6eK6lO90EM4Qo5KwOYUNmJwQOHT
u75uulF41fcePimYRsziw09+t7D7hs6FfeV/j7RCObes4hsVDii+xeDC2NQ+sAvmrY9jS+xYRprw
8XwH+Jf2m1ao7TTxVTEoAztQj36NW0bXd/es4JLxC7BURHl/tIG5U5n0NJFHe0csN9UfNCMGs6EM
OYn/5fwTXd7WdFnqczgtlJ/vcnAb7+RoNoGEOP1azu3iQ5glUKQKmO7xYxIWHiL4ahSvE98TzHcp
3NXUyByHjSlxRpWHTs4kPnTJOWDgze7H6P5Id5WLJZUF16sOOTfh9vl8Fo10iHFk9L6HhGATf8RQ
AJKD9WkswHnKRXM6zLyP5iVwgqCeYXMphXaxTl2b0byEh62nA0sThhQhIkudiZHRZ0LXYZfrERLt
mhTB9Qxu/s99hS5Lu7w9sUx/KZPOBMvlzxNbhFNcTWIPf3OrzXo6q0aoVWnw2ve4qDM+QHKDIa4O
V4mNckuuCackL8au+z+cvXBEgmXOuMbM6v94I7r9x7kEJ1BG8XXkftSLdbsquE14fV+oejNdeDLi
JRRydr0JcJICDD/oJKM5UyfygalzuMR5M+8pYn6YeCt9fmPYHcB9ZO+vbaR1CIWFdzTqpAYkN0EZ
JVNfG8buyQ+++iGT9+l/Cou0f0hUuqWEh/g7j1+dR3dPgvXWEx2RTG4sPbulikqfv1IcYCqXzL33
zBKRYnrGGMcBWLjk0odqhF44CEpEVG7SY8V5yBkcLyyQ75mkm4shnhXRh3MODf8rSs5oe5lnXT0z
l9A2RO7g/rbL/gyxeltZIBs6GVOPeBpNDZjBBD75Ge0Rdl7wot2Op1SXXAKkGGW/oKZqfGED4ol+
8dp1Jv9H8LCWPkAEkVyu7HPECcZbjK33jtt05PRVjYuCWeGibUnl/8xdCzDKGn3NsjJd1VLzdokC
P8/qyiZApO4mKzia8QWSH4ssJQ7eZGKiTYLhjBT/PgyZqn5DOjMdETqXgXfbVh4OOrk8KDaZw4zs
wG2YUu0iliqoGXhyCk2qT8xHGyBgoNDajFMRvasFZmtizvX/jsniQ5RoU2DD/9u/z1Q+a31ZKUtZ
SHfnJ5VeoONwDJjJXizu8nARAFE/weENWTpLv8Yo3xBB8r+nRnq972V35E1NtRQ9liVCYEC/gcwN
Frv2zhJef/eDhi3fguRNw0dptimGoutKCRc7UZNaGqLSjQ3yoZcDJKnWV8JXFxPyNMhxf0NNAh2T
dPnh/Q9R2wZ9ee87Rwz99yxYABwre5E/3nmvncpDnNk5BUlcw8rQgIUDTQQDuZq4BuKkaONOY/uv
XHqilMkwAb5I/a0JHoDYtXrFsIFNa5hNfb3CXx6QM++a5uWZARlvDD5qAf5et5zus/BfFVdhp0mN
WglqKHdzOBqurilq+qMIf1HSQ4E2ClLkbOIFQy9KD+60Paq23Oo36A4U7B0jBRghalfF0b5ne226
yYBwm2KVeXZfcGC0d6/9GKGS/lHVTYvn9HWC1cNRnKDVNU8YJ+2mgVvbFvaEklX0cTJ0DCk/nWY5
3LNAHbSxuDwfcmUArvAYinCr/TF912U1oarrb48QttJIt8hE25RB9BH/i4JaArXFZMHqmQemeIyt
PKGV5NPOmxVFZH7A0LBFS//vb8sMB8sY1BnG2xdrB0TEatpq1p1nIfN6ueR+gW197f4Fz2hdCKxf
NnXhbvlh+ywWrl55WAqaL1wWgeo+7KhHp7t0QFaMaGc5UOhJUV96La/kymCvG9wLxpJUz+nA+pZZ
bYc2yGxs/Ng+eoG4YjokWiW+H7W7g2j7+aJnYH6VEP9BcA/mKSR2rBWixBkPBCnCK7XUNM2W+G85
sFdmjcxWvDtkMkd0iyVqoXnkhCRYWllTILkv4MTXAimyM5CtAPzrFbu72juC0vTZmu1OZfGZ5uMO
brFmeJIQfbytpZZ6FJJbK9ShfQ+9ho2CPpVVbrhmunbWsCvZGUqAJ6TmiQukCH1rjLnO9MJ7OZ+5
FagOiM/fe9TU/5oqQ7lx40pdFmZNpeUyy9AzSzVHFWIEFc9Ju2f4QG3xjrwfyykWOnkRfFKRM7Wk
UPYRvl7BHQugd+9L36HTUJIHjFVr8u/cS+/w7mqlj/fMkWpGGmmfG/RXs3jBxNro+396i+07lJjJ
VQXytLMXtkfXZKlaU9OOS1O+Gjy/K5ZfW3uTZOT9JOWDxIHjjv5wD7JYTb1aULoM5+bYgqlTFIbE
ENo/vnRoJ0g6hlpNkUBQpR3SYvga4h8dT88epYpU3kTaHIEufNzZrs94b+kAAga6iFkuQxbtxA9T
oTFD/2HoNxSy1fbP3LUjGlZi1r+q3Z7pp3JjH4odkSeaJg452Xf9YhDRwCde8/ORlSRDJtR5C7mU
MkZjWj0nk6NjBa4RHcZLvnstC+5EVhaUZmPTq1goUlQAy/ehXrlfWjvO62Yp6ODgGLPv/AJ/fxaO
UTALrmTlDDwrJ9bBayAlqWZU+nvT2X5d3q0kebQ3MYhApGTKyVCkuwzpM5BMVOp4z8DITdSL3rpJ
K5/MJSjNAWRG/MVqt2DVxNhx8Y/L0tFQSH/az8Y9t6FbOwISuHAJFujNZOUAP/44SrKlvjc8VNf7
NbGTubNkj6hP6Vo4rFX7+CZ4aMYIZ9klWDzEt60grPI4KUDznIjzuPtCLgqI6Hb0mxBHH5hiU1R3
gCLwoWyktlGLqBjr2yKtPw9QW6Si5hiOVOFZTB39eCWCJ3FQ1Xcw5l4sDxar3nAmwSzvTL1TSOBY
iU01/5sn0EKraZhWKxXygVzS7DRXpzRb0j5KNSOKIkoi5/7BXmYhlp2rhBuZ6re3LrMS89dy+bqO
69bOOrxTqImlbnzyHLUSAvNxs2Z6rgOvvtGgWbwWsD+/ttg703G+Qw1MiZy7pWOFT/Fc7HysX4Kl
Z9Lyd440cUZhYyzIvUH7PrSwl372/3xkEoFzTSr3131QjMRK+1ObKWpd6WywDPLdrA2TTjLLtyMP
bOarL8cB+ekh25IZnkAhSEWn/m8mV4cb9VOimvz/s34ffyh2hS97imLf4SGQFIOQCfxdgssDli0F
Uk9QjuqLW0JP010q1TsPDzUFliK5yCSTiMlZ9HpEwYkGgniqgp7LyzfyxfXcl7FDLWGuVxChwech
e92fyhbKNg0O6E27hMlC4Tbt6WDOagxAPoZH4Q63x8R6tCIWs/Qj4vbWTPHS4WCeEMZtdKFd9z5v
B6Rwo06Dx3CYhlt3v3u15k5ogNnnouwa6FhC/HGVQVY2EbwVTkCku2Ld1TOvnihVI4Lw1+pYY3zF
eiyl/q5mCtEe4Gk1nZZFsk4tmVVBqc/fdo8mucFzuDAROWbeq4pHLKfgDPZJ8iZcI1QcWkXIEIZU
lppv8yDF8Jrs1Mjkp76USQzTP8fiyX0+32Mlpw4lUAvPYYBCjVXMU4NP4BvdV3x0FRmE1n6Jx9wx
yIw5r2H1k7kbec/9F6FRp5oSAX3EEIouMk0ZK764QFFFemI7df2aEDl0ZmDyzXZfqnkHprKiBnVc
OPlT8eAHT3PYObPgnw1fmZmidmBs5kDzvPHfCjoTkpVkAhHviCiETH7IYRF2VEBmz8j1Rv0Fw1/Q
UzKGDXqiGYUz1WSJ92OGKX4o3usSEgiKS0d/4WB02wi739PCBobw47C1whBzoWRMlj5SVqP+NdMw
JvkbJ0r323C3Ysmt3kfsHs7yJp535zmnh0JrkCq6g0RHQk7TlaroSZL7PHgkvS0kT14Qfs7JQhGf
jaKbOOht1Xklea+oir9QnM7tvIX6mqIFYP7mSyfC+8gpZEfM5u3muOVkMZZR8x3T5Qd6sBb1Wuas
5L52E4PADJyYA6l1FFsmV/k7icVclOcww++gq8PGbq5d/KIsl5NrpZgch1ULUxdD8vRTYZyr+JWa
BhmmH35I+qmmiNYkh+o83iNn7H5E/myWZIR1zyrTLUQQyhiMw0Jp6yuGvWNcCRtzUMtBtFqkciMb
GTeiFmev3Itebt0vyjhmB1wDo8HG3y50yivP6XYiUCc6GtxPuQop3YFLKmB4rSxLro8cYiaDrHy3
DyxTSVssoy42xeNtURSFKUN6Y2RLllsgqTEKbptNtWSOM4tduEMccsams7pjTVb2EekPtcQOX5mA
i0WYQbDfm66nlznwJr6FolUzNBNwRiQcR9h72COhb5oK+nO9TV04vAsepqhJTitJVd2wlBptmsDt
ou5LN7tJDrK+JpT9bo08ozC4XnBA5/wAjFSpKLMcsr2y+OQllyGnqM0h/iQuoa8Fo7q81a8BwP1v
i245wauzo9KICf7Wx0Gf+njmN+B1aolL654M27iFoofECGKuGwle8mqsinYkpBNBxnLQ+rMK6Q7K
NbjQDSounvB8e9d6TutKSOWEEKcP7o/yacbbkVXekYIjolT1Z/WSz5RvOwowSGt0lBjX3flO8vtd
3tYy6Iip5vn2Z98RzEJDmhz7e8zPfv3TzSS/UjJHxEOZPsx7VKj22OuDfLfgXBmc27Rso7oGIl5K
LOzfnHX3kEwhedNMBWNuK/4hTavRWDpJxN2v0ID+4sqng1Q16nxtFtueOpbFMeukqsGxJ6yXayAx
4L6Mdw+Sjs9712BnIWnO68gwaMIbAbIaiYOOa7VK/971qx9Kee7YyQFREkiSsfbfB3ZKlgj8ZMr2
CITE9ZS+RcHlRbld1i4S5PwS4DBCzkGh/wYbJeYYKq9rm3Xt5bLQa3WHtb0WQPGGjvVsbUNybW6n
eZMqrTnQYrkNQnGGZPw4tHfu7Ytsk6GefKWQKdH9SgC5qjSdQ0mS5Ozq6HUZLiWZeoOkaXE0exDL
jMCkGg6TjjRsh93Y20NuifmwqcDDHAWrCMooz5KrQEobgajOcOjq92Te83zya9hAyVEfBcZ6/oBm
lKDPGhLg+9SHS42BHYJY2LUGwifUvwrQAFvRmySTe4LzrcgLz2wHAWloaAaCD9OoVZEbhOa1/XWc
U3IIGTeVU8YabI0pbVZsHeesvaAMPON35nepke1Mh50h27UFQ5/vpg65kqAKXLEecwiH7lxQ8rtB
bE7HINh1pUjNMHYgLSKapqMFn+Tu9GT/FebHvh1DfDchREVwkWYd+b8ZFopEC0MosvUCQXbU16Wr
bUx3aR4XUGhutNbkeNqH6WeIlNx4MXJVZpCMsk1DCkoGd7pWUWbL2kDB/VwxUybJn6fYo98vktye
U5ygLfdTS21I1ruwIUwwXnDyilW03s7LbF5M1Yi6wlVGqdi+lN816S2gphU7y8fWZ4aBIOQoPf/A
p8UWzo2yphq6DUs7I2SDS6zvVaES6yK0bWuOzJ5/7aggZF7P6s5whl8GuA4qbtlCiKh5tgBZgf8F
FuAqvOvnted8nL0pIjGuQT0vAF+p3dpZaiMGbkV6Z/nnKnD4gfTCvI4+K+6Qs8Fn+bM1OXAmPUnw
UcwMtdnIitqGuqe1XOm7IGYDy4zCaYLKuspMoTEMFTIju/PhBf8pUoi92Hh/u7D16Petv72QQWqE
/CUQ/K23kobT7h2An+iWLdeEA1evf9GlRWRa3+2fGaqtskAWS5EEDcOKIck7dnKsR9VYaesMXOjy
BBJH8PvOvs9MmPOZTDxefjxBBNB6z2HTfoGT+GIKs2tSo4neBytghOZsT++bl+z6/yuhz4Dfybde
S0imzwedCf/BzBX0gPAaG0+J8CDCmqyUjWtvOmo1lAJfWfidYPDMHWHgvdZvFoUR//1h6bvdVIPj
TRyBo1bZWSbhjpkaERuX43PfTySWL3P6P9kcH9AJiyymnHjFMojjqQqg2YjKMsN76HKpPktGiAVT
jny80mGS3JiviebwO2cHTuovP4ZnKiLbQh+uI/Ejh5+0DNW2afRkD2LNFcnpXlX1LI7o8MXhttE1
xegVD4OGgyynVQOax5NyvY8l812Gd8nW7baJGyRrEeEcQemy4eHzkt2r39azABDTfNFi7V3g8L1x
ZqNGPpWQ/hU7QC8cyV9TiFU1KIl++9+40M3DtqL5ka0+1KPoNmJ/an4+unNqgupE4wif46uxSIlK
At7X64Cs8yc2xI7yCj/ojYf9JwkuqIZcLG9Rzo0M8vedl5I/CHnmomDrTLKL+XF5T6jc2g0aLn8j
KuqzqbZP38r5TPW9nAoFyzwksquRiJY+zgG/CZwVoywhYZQN8HCoUNyNmzVHHrvWl7AlITRgsB24
jsdd/Pw0CKpqywWXg8v7a5+pVSWaQ5m6fDmpwFSTCVbq2nJoGGDVs+PpyT4wIe6K5qWymajbnaBn
qFnx4hEhyN+9Q4wYSqhHz71/WAzqK+zJnU92EOci1S+cJVNOC0prv0zlnpaXzsdcFqnWU2QiWE7I
zbFWHvQnWCzdU/HoqnOtRsVGVK3W9v+itMvNWfPQV2Y2ScRDkmnqGDwvlF1Wq4ukppnh7s/UCWgu
c0JWQeTncjdgdLwz1V1DDuL19VDxrM4OdCjwFCeLnj+xF0tpTBzNnzT9yPnLVzkXHhpfLurEhX8O
QcFhoqqM1LYcOwDwIdZpC6/DY1u/aARbKVuHNrfda0bEZYG/3I3RDjzM2FEcvw/of8C9p44VD9HH
a4b0jXNiatDXor3KqNipErYPtbGimI6Dp86ZccwVyB7hrirqm0R5PxWNO/EOpQUop4xmQRl+3U4H
CLv7PbPKfuI7oYG2px8OzS3A0ltqNXPXFxzct8QQEhadjygXltFzsrQfEDx1obBCweq0G/57YzHm
zMwWWI0UnWG6ADnk05f+0t3kLY2BdJK3nEvR0OBhWlYqWQz7bSK5hBdlNBbemoev6ohPQLtAp2Xb
7tebUSx1H9KWQOQ/8tpfCMEfAi8dl5rw2YV+9aCQqkioEW6aezf8nGbvo1rikpUHGUE1noKtTQD1
B4y+vt2tQ/gfDFVPElSVe22fn/FBY5o6p2uXXlV6SCz4YHZvE0JiUSQFhtPuQMQpFIQ3aJnkSH6w
ad6QNWopD/cFfvHoN8v2nWZXaM3sFk+n5NZaFaFw8gs+7tmYS1XpnJaNdZR4YW/T93JEJ5uEXLI6
R3HupmoP8vFHdOG1RHuG3/IiBu1c6fCTiMAfuQA+X4Ype9IYeCgof8aA+tl6Q9Scpj22sskzD1qB
C0M2Z0nLmw1hFzuPX+7HCJYmDj/L32zIZdDHcwY+2yrYCYvAUZIqcMmmPeZJtHWrZ1m5uaD9IQSK
+JF2fLv7DZ1TnGRKSI36Ga5BYFwLdGM/+Cj3s4QkpCZv/enr1oE5H6q5ykumVtElYtoft4Af+uRV
hiFarc5u1ls6GsqmoPLpoX6rahlproISUKzwPSKg2m8iT8DwJZxhxwGW8jv+Z0AiCFqMdPWvt6Z0
h7xJDfoQyMC5AHZnkk5ySUPX5br1wSBcQFpdDqrcuDZHg6thKVKKISzy1fvj8pfqmsWsNICCZgLa
l0KWSkzZHnHmAKzZ9jLyUEKHRhB6++W8ZMWZX+07OtVM/3y7VI9b7zxU9H3/RI8GKpZdnmJ6pmCf
NRrT6nRUBZ6bamsVm9OLPi4ITu/xu6vXzRLWZcvXDaDhtt0bp7Z9nZ1IVyl/k66rkSSG2SujfE1A
rOQGOVGKDXdml/tmOK5uHqQyibkDoxh32ubt91p/H3XbRPoom9tL9BwNtGtF5UDc2YVHclC8W+C9
1Q/joDgmATC6GxJW7ise0fEBG46Ynu1+k59rxNDAQT7NFQEQVPt+SiBD1HFE7m5gOZGYe2OYDV73
BDxOkl2vq/kH/kQEp32eCdSqQJNxCBfUbzXR/J2gxLmfi3FdIcAAUwng+9qcQAyRGMEIuFzk5t7/
/3zdXXfd7QCTpargFMVEYfisvAMdw/M1fESVXgDRpa2DA8UD+f1kP3HwYpMIXKfx2tdcJUPKxims
HwyA2HlToMpnkzOnzovk2VQVVtiXgt2gdYGnp0SYYRCNClZp5SUcMCzm7WVLVVn3EKqGGa6ZHv5j
vAvvls7FSTc63LEjtIYYBQllb23H8xDD2o1KRZCEkiFOSLRIgKFWuy3qUVStIx7lRHbz5MCsxuB+
KIoAVj5v01VYoMI+RP0fQhBhp/PFeTinJNkoWlDOoLdl8tZ00iX7ATWdOmEqgCFgjjuBy6zdlUTP
DUyaBQrxZFUZvLvFwSt2tco5Aaur22D04rkZ4YWrUnFShq9+ICYyXrdZEa9azCNJEjQHDyDypDCI
WfH3LkBQ6J3H4cN03reXa6AlLbppiGf0iFDMDbvTB3TzyODyrv5o4ueEjAJS2OZFPtFbKyYq1XMZ
M15PqB5Tb3ZPwB32AFi++fLl2CubuIEUSTbVepKWfNO3TAenp/1/yV8AyoQ2hdezoqf1TzlT68rh
Pd9QiBZQm6DRjRd6im9TMOis+LwxBIt6Upf6EieywyAp/DTpGZW48gcANrHIGLsHG+xmrkDwVUX5
aVFc86hs3XCqEAe5nJ6owt69MCUOEO46q5VsN2bLGKhYr0v55yF3caf0Uy9NIMwh8b6gzfaln6Yh
2rEus8od/ROQuBakD8+vjktmQ5iH/d2ef+bRI7PyiNDweHX/AKshka9uSV6MlWMoAZrUTJxAB7tN
bnM8dFSllkdfj/MD5whGDzZK4H/rjALZmLIyWWQBgBPYvJIhcoKf55+4SFF7B6Rs0b0WNR5Kn9Y5
3uhIMlBDr9vWraWwQgWoseix/vRnM1Yjb0daipaFqPAAosqXNdWYeOaQqepNU0E2T/20h/tCg/1g
wv3GoV0siczcQ/lbjNiIS4LZLxlhWjAjbRkewliIOYUmLdn5NlP0LvxHpWa3rgRzPvJ3ByISh5AX
+DPRCizamAVwrxO1TABCmnRZv1LVaOCCRzAG963uJGIyWopR6gy2mTW8W1vf4vfPi2ntnr95cvlk
D4LpnbbKiOhXZbfwTKdcuv+x7C6+C0qa+cwdqwYvfM04ze3BUSaxqRJkXFUIr+6Gu8WU5hkOprJ1
l8I6q0KVAH9bb06QRKYZMnQM9ym/Dsw+wsf77lSXPrWRz2SKU12fXCtTHO+aci9sRSEcNumXmsAZ
vKlQMIw0/HLmQ6L3JuP5aqOWWZv6ipYi5gly2JLRyTf2u6kJRdz5F/y217krUKqn3kFlUnQOe0tK
RUovi7S7hgGxtpjUPWBYybnxYv0uW07ahQDq4hqiD5JNzLlSvHIbot0r+RmP3ZTFYqjmewdi936l
48dGbeEoIZZmkJYLRYZJN98C9t5f4OZk9juHrN2zs58oVzsnTWn/eXEHTn1+MbqVuFzxeaWoQ2X+
JydZJDpBvuFF47UYfTuxPp3Q9rNnMKiEXAnDZyYK0cYfC7KhL4175QFB6YYgEdQ2Ek4ag/D4pH0l
eNbtE4wYUCFiL4Xz+KfxAVwuoZyuzU0dn/lp7oN+1a2yQERYVOo/o9iTL2OwdXyRhVRGQVFrhJ0q
FvoswsTE+M7E3QClYXQM6P1XvBw1nFhmkmn2lRmMM842AJrUG66QZjCqRUHr2eejp1onsKBo86k1
OynVffZDhUq/JQxf85aZ6BlMrnObgnkaEL+GjsLS2RoICGRdA8/9O3t1o9assZEY8gJSNWN9PIsl
vGIQDU+PLerFrGCljFKRkzkgIhnlx2UHdg/FakZnyS0kxUGhoScaSeSoMAu56V7HgC5/Vx7JIZo8
7ZUT7eDXIt9Ba+Ga1OeVC/xkU9mBzPOr4+XwE62RvI2IRs6dFft1dpfb4+acZWTFnP2im1VP1wNr
C8bdLiSrPmRBbaevR0QRnAHCWUKXLdwYxS7R2cshKc2VXXQhanOdi43jJgLBJzgokzIPPZ2P+tr9
tSseq+396Sxte4vJ2HhMcWd20XuA7tEUCvmzDeykDK8xOSU7inTO4IqSmZd3+Pd6G0AnBcqHCJXA
qDCf723JkaHMK2zxYd1MZttB/bhUfDrTgbHtIdpCIKj4vUeUfzreSs09L3OcHgJ44m2BrZxdPFwd
u1bUxSNcUCd0+EbVc7ogpgtWMJAv+XU+MmATNQcuGBrXiqkGkpbfx4kVSBDwOpSa1dyZ0c5jirNk
bsJP4Ow0WcyrQzIvj4tuLJ266bV1GxDUkbMtlpPOZDwImg0PUXpyRgeM3IAv/1sjMG+9WJT0j507
rRo38CkFhaCxZZkcgZcALWv/oCHMj0oEfVttL4FSQnVbaCjciB0p9AuU0rOhoJseM4PhaU0dov9B
KaEM18jkhLY/HRYbeUi4ydgrKj6YoXcW8mOBGXSF3m+XGnHxV4tsA6uv3WamolyNc0yYmxqnEwqS
sEjKiFSwBau/w6UeX5kW8Mv0tVmhHPOA2ZIvW/NF0HqFx1pJZDSzb9ftW28y/VYMm2ZJAINy6auv
PrNzEtDdwKlVIixtHQ42gQ+aee4KdgOc43G4153uWCpDazamPE9j2gYH2fcUxJpX+200iUZBuD1r
a5qKKFowEoF1rv5NUBDfF6dVrWhbPTWHt12yDDZuuoSW8EEvnhlH9jphQA7tCQv3oHWF6mAe+JGF
ZRVIzM6SdaUA8uG5IaCGeX/EkwYByfloeK8wALlOwcO/YSUQccutMHOFEdmjsp+q7rDdGzQMZcCy
oScUvEok7D4EjMNC5KS1TxZMVh6aJKPPQbkL7THZlUB7jKAxGQio0NeOSPjHiFoSJt2M9AaC3KUQ
251e0RMjAk5204F35dkRB9B/oKE8DGxNjHoHXJrU8FeL20yGlSgVsJlWLxgRrSVHJhfWgnePYwMW
LhR6ePH9TU3DbJlAU2kHRnz1MPPLE0HmEKx+N6ws0Ba+31KIV+ok2jh2Ss/LuuROnEqMDQ8F7x7e
Xk6zZ9/AQAn6Z98e5eZiSuMf/qOQt9UOUYg/GRCfVqQFNpg2r3Efx2NrgMoRWH+iFeYCUut+p8cx
gs8kiziA/wQZwRvZsyCeOrrUOjUYJLEx/CTTnWwZ/HTVm8OK4neoFQRSX0uXKwgeSDG1FNYtMx0k
+UfHSHN9IntTbJZukvYNL07UCMjEB0XKBerhQyr/c11TtrmWggjPj3vyXyDrJh+GMkU0uUeTMhT1
Q9r2qzJsy093oKkLhOn4BoK/O7ITRrFM+gfDQ1A3PZW/Z/0ZGjMj6KrGQ0crrUvtrx0lNUIe+HGB
3pUiYCiz/ETcKGtVvtFrW8ZVFM0J05WKhvQmOTb/FtNB8Rihht7kY/rU31ZI7GRsWQyFrRkegQsg
Hr8lPyzNdh5NaFlTb65FbTZ0JWHLUCWwvltAA8LObSRq5KOC+g91AyJ0rSExit9MYjMHGe55L9B+
DrKPOhB2z2OAWOrdgjF/UAHipcGSGttFcyHlEqYNjrJuPbFbCnE5iuhbpiHyp7TVFOQq6KCArm1e
xCPdRw1+hgqLMGOEBv/baoNp93cIOXgFRjOh6AvQO3GLLMB6Cnqz/a2Eztby9a3sZD/TWlTaUDnI
Lyvmfm9fmvxDR/Ckb10v/tje50dXdIgTtZT9fx241BlFsTIoijvjU89JnsnQxTmCqGw4IO5ktGoM
yLEDiPwnd0IG2jCSrzqu793H68lFu4mOO+C81n4NZ4Fxm83fB1kQxLBklHB8QHdPqsx3hT8AugFl
lZLCbL/S1pJX4fDEoHKRn52FSnWt6xOGT0aMAnsjjl0GQNsbV/qkLKrCnorhNRQAMNOiCtHQQvwB
Gpc0HUoL5b0UWaMYd17XK+FvrF+0B4qBFvSHKkAlLOmFlSDh9qRBir3TGNvZU9ADXHfztqe5jGV2
NlCZsUhQbUrsnjXSM5jSnHoAKZ+ZSgDUYDTM1cwtfxfTdg0/ZiI15fDkPkAMwPHLu4jUrCAHafZV
c8zc3w6XnmK66m1symm7IaK0mg4swHu6jTehHqpZuEu0rGsaZiJpdvYghyyJTLvVG0DY2JnvDRzq
0hrHw92jUjC753uVkEEnzdNP7IyaKul/tMx0FORFRhRMVvUtfhkvVJ1VxQa3ILJa8w7X/t7QX21Y
o2/HvvJgywqA7lt6Vq+KM2e3AvcBsMpDd7kt2b9gB8CwfNIXmBI9H3EWQukFUt7v3E80VTUb1WVw
RRY/gdjhx2eoCWNd89imE7LzSP9/Gkoek9peAN1IAJwNS89ofoXl8Gn8jiX5n85cMbMvFK3SOmap
t3xoNfMQoBNd9F3LABDpWA23Clf/xxqmFJJcGSCtSF9I7mpc9GoTU11CE0UyZhJGvZ9AYdzT8Dum
yl5vxhv1xr50aecrjFD+Eqztl+egfXNZ4Hg3neonpgM2TWgdqQL+c47zuu57QZUyfTiccWmnN478
LzGeLK+AJ63xmJ0AFJHgTNo/kSMBijapxtJF/MwI0ZbMwcG58/ohaGRjjUEIiYiWF0dppHevqt95
i/ifXYSbQPE5zCkxPVUazM4yck+gxsDONzCcPTElB0zJXbOQ1js24uDHy8AItRdMXE038f5AuGNV
iqVBwdNW5g3b3EK3r8Ov3rlOKkftxP1ZWgZFZIfzAja0TopahB8FfzU5OY1jYfibI63hL3/bclF1
77SuouC0xXMsnzFgKLFOEqqeYk5/iY4AkK6mK+ChapOjaWPYj22OPIpKJmvQ2TwKlLEgKgPakqoD
92HyCL/6C9NiA5ErGIHgk9Bf2ultcjYy1pGAltXiiqPSEpTkePD6vsHVT92Pe17Z1G8pEzcUoumH
NHzXiS/NRhOJNYEfMbmqfQZ7gxrfCBKv886vkm646tinSreZ5IS6++vgAVBBI+UfRzNrYUo3zKdj
rbkFQx9Hjzl2R+41lW8oP7h99J/Pc/tO1yeAm4Px+Py9jcp7cL5IMP1oCra8I0osXny1rG+LOGqz
46IXpwwv4WKhrLQdO9uLVHo8j2iGjXpearyEUxllu2wSqMzUPKPowicA5jlm5QdP6pa9ymg+GYJP
IWhZF7FnLhsux7FF7YRc6C2fgZiKmdZehJDTcusEXvlKGkcomWCWopjyc0Q29+gsscnmyFfnFM1h
rOjhBJl+aHQjXpJEJBzS3SS2n+cg/QjsCIBeBYVfR6ICeWJGtn+D5i1SiicVH/KD3fMR/koU9P8T
cXR15NrO14VEo98IsT7BqSs+M5E1l1zJ7rsm3KOie6Wiwh5b31LEfYvdt3ZIAssgPBj9UW5A2Oyp
ITnTpsRNKXykorUAPWVapNpjsWu26B9BDAOBIoIa0Z+oBIU7lub157VL/BQjuWmJkgoT86YHv0nJ
C2rpg+3RG8py8Ri4xY9Cj4gSdmOaW6QBaRX7MA+FRyRP0bz5Hf2lDLAdTK7gC94MwLAK4EXJpReG
HZnmRZLbIIDvJNg6AYNQn/w0vBl4Pix+YQGRD+SwvvAvHltv9y46nfwkzCJTF8a5VdQU2+myQr/w
an/8L/APtLYifd3HoRpwy8EoQg0yHvDrBvttIxQ41WEdoMm5f4eFp7MbpKgUfLkwnVaHvZfBgjeM
P/xaWT20eZw7Urq5b/Yeu2qkX7eAvx+MFli86WhlQ8pxvOKKXDNCdQPzaLs907wxvjQXCqwMjhwh
vmBCI1C0vUbqZZmN4ZpNsHqE6MY6g7uc3zQb+azYWhCfvuzndnhHqx8LD2NVjaBLvWypxl/8PWyR
HSj1sZ1RDDDdJBoYDSHnaKp77fbF28iO6KRR2Sk0E3pKqr80xYwnURMY+KKAT2FvuFX2c4zoC3+l
Sbr0bFen8eSI1HBLE5pu8nJ4I+hR0Z/fzrJOUVCRwCIa6NaddHnR2KJ2Zf6F7LfNfZ0FEcg+1DX4
laBI5vhz0JclQxYqHMODVXIu3f+VlKI6aS8HuaAtgyT3TO1PrJg5u2JYpCRxYxiTEXY7riHLCtF2
f/9fQF8Lb/A0tg7fv3kyTJA7Cm+Wzu+L7qZqhAXGTVbZQdhIWfhNP57z130nYS6AWVI8ayQW5f1Q
VFWmIAmol4iWhtQEjlzQPX+v+Cal/CdJr2NNfh+yLGZCxmFZb/aeHJjI9g5igcbOc0BFMEgmB1Up
JjAz3A38VyskaVga+NOzs6NTZRPvIQEdwdYT3n+rq7qCRwrO/hqkzitGaCJQ+ebXlDQQq16Vut9p
44D4m+/kZnTt4lEgaQTLAgbi2gmaPF2NScl7MY5B1SlUx3lNmE4/FFb1ppRp8DBLr7a1UwIbhDfQ
ncCkKuw+UwBRA24Ew9POTp4E65tn2znrYO+J4Bz7zbsWI8ou84CjZ4k+cE7/PtYbVOMVxgl4wp8n
XvphRczC6ia/dArAcqxJrAJmb6And/+merV6q59uIghL74QrtcOGz1pSdKnNZgTwNgxG80env1X6
Kc2oaS9AgbIY0tBql4cMNz7k4Sw6K+W9qVJ6vwoLim9eIPOVhYGdW7h4f21BogxcJmAIF/gDk6dj
cAgM4N+LwilY5J1tHFFAlm986PZMqoceJ97tLuabV8wZTV0qkQ7oDb3S0GdDie3YXBe8+LAmHNMx
46z7eJ5FSbwP+yp3bX3Hb9jg0wk6jdI4lHnuvGTxJZgCV1nnfP2b1f5qKnYr7qnj30wExHkDJSop
uWsmDso6ab3IuqJl8wW1D5AUzo8oYYjKJ2aSQy3096D+n1QNWyFXcNsOmQGjePgXEUzZlqK8Z10k
oddwtGcBbyyLbrXaylYbtPqGwyV+lESbjrX/DxVv/fMUkugXfrJpuisnv0tLkxrroEltU7sOrXIX
KjdEOeu1ZwgsCqp2EnekyN6FCT8ISPuK0YeAZLuz0AqTXmWD9Y3Y2BW0zMG2Tt+40ezwYPYHo4o6
aTiJAjcOmnnRctP7W1fafY1vx212XrRZgeuFPoxTqL2x+SpoJJJivIVZypS1Z7KcCj5lAJVOZPYB
SejDsZhTe1g8oYOEtCBtZFHqlYEWIumAC0Q3IeYGnMMm5LbhtefKCqq+ARmXQZ9j039pd4goue89
RhAXahzATM8vuoIlI8JOZ3EOC4DU0b+/j1Yh3Dy3JHoNvrJmYPv2HBEASeaLlAVhkBMRbxgpa3Qo
SSfpzeTtMsIWSPhMw+2kAK9zsah2x085g9AOVsoT1rIYaX2tCRcNOQAcOag0xV7aD/ESh9oEcvRQ
3hXoh8QghGwXtkScDyik66sB4X5qY9VrjqPwoX81uNwUzmq0pvDtppexQBDL7PNbPyMvtoFJMqlu
/fIYFddJSJUKOSw0WRIl8Rg3NSswlohQIYPreeYvsSR4gpjPhVJRqxpyriLcthaEA0woqdb9cMX9
kqPWSP6NGFYCcrdCD2ygNYh2c4K9uO0EYR6T9mCDNmHxVbgCOM3J4tFsf4mrQ+mqX3WOuDhY6Xkq
OaPZ2dUF1JhQd6gIfz7JG8yPRfPanQI2qBnWl5UPn8TJZfG/94uZZc1vjcYSJIuOgCN+MRsFb+ZA
epMK2iaJxrSWNvKHPwipcfCwLLSwxNKdL1oHvAd6gsEBkw1jWYUw+cNLkjmkaJoTcg74JwCMTqT9
s3z67TSkgYWam2M/PCehS5Wb47tvLZuhn3nD1XRSU7W3QbUqkViLsvjml44u/GKi7qPSzqnm+mNQ
W25nG7Xnr1cOJZ4apIZnbKWDh0hrrTiH7iZ3LnVfgMQjiYPlkJ/8eDktDitoNTFgjbriPCi8jVC5
8lm/hHVKDubXgeExoH15PWJnVhnIFDHUzwcakmbh69a7taBMAkz+8MpzT5zLeqNZf5+ECWp5/0e0
WzA/74bY/52vqKnvK4EwCQOxxlm6ISdXAsErHyywsXcU0pSNPw43a8a7iLvGWEldqJwVww5nP2ae
HW5McWiBTM0n5+YFnbYraV39I/YiE0HR3XpmsIUJm8nS0qLF9HM8dUNlH11PQcXuck75Tv1psoaq
hm15m24mH0TYX+b48ImJmw/1Le99BnZBeOS9TU1oiKjM2QHb/uzIxHvHUTUj1MuZHmks8iIety5o
V+8OL+tsqpnNzrhUTX0KoB7MnRRBH6A2/yQSIyXlzpxb5yfoUdBJl5W2xuDIQ7erbOsG0+NNu1j0
WesWk9CmHkcD25uuCq9YvP8tdf+rkLerN2I7WNajI5stUBDLRsA1Urm8QcpT/z09Pue+YjHbbfd+
Ztlb7eQzNfp+llVEL21rOwHdYc/AcKxjdnFnKU9q95eeZa2Dr5oArd7j6/QKP6h/npo76AQKe4sE
Y/6LhNtwMhL+qvj8zDkS7BLP4TVkLUP7vE9rHYboiurlKyCA+mukyU1S6pzgUPHRXxvo3+jHjM5R
Kop3WGEpUVVel5DOCSlKjZYbcZTN4K4rY64VKrLIlLwe1n5ATJOfXSLfcOl2hQYxAPO1GfulqG2y
hFJ4p9YsAL+AssOAMUx1bLzbTA3H1qK/K6xJcxLqDBhcHemJ4ZGLOUdsSaup9JZnl/HrfATNQb7j
KH0bSBzDHPyx1HDCvAQVnMH/FIddphEsAC5ozDoSV7qBPsD4UM/4zvK+mVqSkr4L290pPCLrwxH0
bI2nNwmVRQhUoZccWkwrVR79DjWw3oICWmVN0baKXd7zi7U22Nn3GusRVPBTBsoq2mJ3MQgqpaZN
b8Ukz/eZQUfn+fqcUG3Hi27Bc67nibizS5Jo1allFHwwQSMtxEbp/kEIZbF7JLW4Vd6cN99IhDM/
O1qqFi4rC+zutvxy0WXxKimjbiENSQzvmE4YsDwII94PGYDNw8867F/Tb3rjHl3DbRh1pohcfBd/
6pfHLTl6t63meAvFd5MvBpdWg8L7L2Wz5u7D+fs4quLHtHB818dd8/0W/YmiFr7/ZoPLvlTR/oED
n4OmN90DrBDkw/FQ22IOuAdgG5zcZUplumsWzZsDcSI6k4ONpLO4C5pP8ub4t+nEtbvMRAp2EL/g
vRtAhl86JGtLvuMs7jL1D3kwy6ECn4U63yI5tEq45xZD+8nJUfyhPiTorufd6Nd6enw2SxetDbqG
RcaMCFegSFn89/bUfH5MCULNVeOEtS/xQuBzmN/+Gt7z8fXG0Cb9M8XfIWdDDYj0qNFBJGMQ5AWP
jyzQnEjoNm99wrREaJc76vuHsTuMxGi7JmlFFQuj7tKijCXMUpz4z8nEGaDsI4F/b0A+9aEKcQjC
4UNfjavBqghVC25EbsvYvf4Laac8jUv11t24uqYO9SVi65xEzV29nxqq5ZAu4MbregyFwF/vEZNg
l7nJ9NySXiaHKEhcpB+WgrtDw/gbfCOaurKLkg/fPMiWXBBFOESpxWRumGQ7HpFjtu0CJdZaemFo
/T50xd8zTq1nPnnZBFjMxtzXp/1ntnE64fm11mB8Og4ndgKxYHUbrMW832YI0R+WajV1984QgYwn
xhqR7WeYFylKg9Rw2NEi0IVnZ9RhzrhP1GbLPNwJgFanypX0phEbkQQ8fPON2DyogPI6geWQtLQ5
dZf2SwhJg0CaCvS682kMKErJ3ZTmZRlRJlYYqE9YzjujDtb9suDWUkaYJcY7oLzF48+8R4NQrHYt
Spo4W4bBxbkALkcZHfmtqR9mGNhdC2CR7beneOfUKxLi+oB0bbZvx7Cwhphn6b36eZNu6eBNDCg8
gGM98MyvwhhUwlWcnt5v9wbC/Yyd9WUs9K8q3GpOOEtBF8yjWMWvMYjQeeglpImmeV/Nt3d/SOgB
dp8wtat/YSrtmOgX2TUy5/uDy+am40GsPbocjKNFFPj3hi70dUYyjj6xVb/wGVi+ujKxl2NVPHmH
LWNI1dzCeIWmQG4ejPOVk2fQuX3qC96BULHelMKtTBn48+RHRErv+4ISSYDL8Sg+ztBIoscE8qFi
tPffVpaJ1GwTbvDtV69rtv10tPFupvyJEdQL0QgghU/PagrPmGG6fOCIfL+jOD3w/AKXWCw+OP+D
7k7FDcH7xho5TvQDngo0cH8EamyBjPxPCJTP2q2JIluNEnlYqqV809Pa1L0uOo5T0cvtJIVqBHvU
cD4gmcMyKA96T9qk3N4ikAf5d8LAinHDl25FrmcPH56SSkoOlr8swKl5jmfo6y9KsgECqfnSJyGS
lCmM1bl36yjG5McRt7gdxd6R00zLhzGvg68idWo8pE5EXLrM+hZdLXLar8WiKOR3sqW5j7zBkDn7
aNlRkO1QLcitbyrXt9EP9AxisixWilrf4E95n2i8cCq9yIOts38TI0MmbRO9tz7UDdqCVquco3kr
wHqDYBA0GaP9G/IEyR7zI2miqqrCkGbi30NyDGYvUg/tD/XsxHftgXs+z1hqaFgrS91OnMgBm1Lr
XIFxTgpMI7Y+I3BTxHui3FwFKKftqEv2RCLHPlRgdvbi0RU21ExQFO02l39L/+d6/JwXK9JrWxZ/
fu0XzD9lw4FuEqErbcqFK7YrEkKIt+vcseQ77gAxkp09diLiQs6GHWVOQVfjBORm2S6XEfKi5oTb
7VhgnOHR3PMHO8AozquK0ed/SnFAk0e6MURgIITA3Cs94WkcBxPZNOxbDV9vDNqbOeSD46k7x7OL
Mp+4YLPQCVE3ADsk+hXXru9/TEWjfVB2Ty2ncqryo5m7PzpJUZqa2cPXQ1vaXlDhRqanxvn+fgby
wUB/n7R32ZCoHBdyKAcEG2Xyy3hGy7Yc0Ntb2GZAS8Xh7wKg8kf4KBr4mCzhgMbJmO6axQr8MCno
ILUjZaJ5PqhP/779hBbMjnCEQJmsCE2fEIKtKWI7Mb52bpdiTMLdl+gx9QsrLW50p70hfJ9/ceVD
O4dQYq6vZHWluEbEhrXSY+c4yp78JAAM+D0yzII/kqUf8HKBSoFo2hIccQJXPE/7JMqrfkxGYLM9
R3sRn123TmQTnMLu4HXWBmdbQnWwostkCafowgnuUuR1whJstSnhVdEbGWovS0ClLWaOpfM5ENdL
dgsfk65GGRnNsNxvG+SUZqw+SWJ9D0NeeEQECGRvL/D4Lnq9GlR3mhYt4KixyXWDB3IKfdCqlQ1F
qtkmLfi+/s/ob/UAG0Z4vYVe/elAp/bM3fT/2kbkV5pk1yBAJkdJT2DfC2dFT50lfHX4JXURg6mF
N8Yhy6hxw8WiSoPgWmLpwfSxgm/R2J4svr0eW3x6OZeL3WxRSQQ0gEBz+7ULZz1X68UeGqF/2xQh
QyTm3LB4ArvWI/LUVlg8nvlXXQaU7hd7ijXxEQK9jLWkJh4cBehndAqnt/nuycSmtIu44qczz2I6
Ladk6EeI1kmfGCTLEs9VYBvNzy37KptLRAXhdKQY7aQmIyY9vDBIxI9H3ZENHbjON1kGdexopQ1d
hnc2DXLwr+rt6fM5JAC0hknvID9K8cj+n96KvrF4+JnEKN8FGfjykiOgclpy+IPJbuEb4y/+b3OC
aj/GMFh52krkZcXd8jgrFlt+WE6Pht1c7Tzci5owdsazKUJ3jIsdn8xQp4xihrqI58G/24/PVsur
z43s0v1/35OqZBknareEGirflm4uweu/ZfPuLOOxw9zyByPqdL4eByeHTCzc2yb/xpzxtLuY1ND+
wQ1soQhHvNmSSVu4CI9X0FqRo4mprxLWZWBf8hkA0OMrttX5ZmEQu364aEKurKURp7UvSwZC9WcE
fB1qMOteHcI3CravGkxrpBKNKMNfPKdmaa+o3cdf83ylyo2lfiAdCfZlkVG2DivWLGtRGNY+xOnh
y5bjrgVNV7RL0vhKnpvAQG3D6en6s1WHn/njJkZEGFFCmAlhqbC0ll0NjPq7pX3mT0l52LIHqg27
bQQJoyT5pbmTe93UeKxcs64Rg2DPkW2AWVgHyTr6Wg48TJ5bGV33YmUmPtEaGW3fRyMgav33Oc3T
S+h196pohzr0HKSRCRI1+Gw1hxCXzh3KwzDhQzPZLL9QcQCuWCzbPzSloBTa2BvUq2lr0cWnll3v
Dzt1y/gXq+bKyKzsUkkrGuXZtN4j9h2P7vz6WLkbX3S6Qj2qGOO8g5+bbGVIkPQ0hxg5/cyYXZv7
g5e3WYh9r64EPih4TYGhnEmDPUlBQr05ZTpXM0CqtqO23EuokU8xFqoZOkSW1EraV5L13sL2Vkgy
gqn6E/d2Fgr2h81TXZ0lDTG3ImPLozTJa9L0Gw7XUut+RThSBoAyOyRxCuuHGbcEMsCQiYWkiLdQ
TxCMukK0cXLuDgMiTMGYGsGGiEC42H6ReqDo7Qjl8b69oAyTXLzR07MphE9xl+ZJSAInPvfudEJj
0DdG2s5nFTQw0Rapr/p1w0+op+hqNgOp8nVQcgrpnEfJziz3bW9IoTewqypAcKhjU6I0sXgIKVh+
Hnlpo7d9cmyDg9vetYgvFxAZISX2hNjwfipzsGF2eJcIkwA8kojAzAF3ZueWRus1dER5c+2fUgFD
hsf16d93sfDerGzwG1O9VXpEo1jQZ4mOZjoxI95pYn4NB5OI/lcm7yYLvzHkSuYy602jXNHZtwJN
tHTYI6UxfxIB2rNFa2sF+8P9Pv9jv9I3hRBE/CJfuTZERF8/YhY0rBgSf1bB4QepwNtbRIUyHP+K
GIZm0xEXFUlkcxrqWSBnONQ8MA7qlG/RHmYCd2ZkyqOKOt+oyC3Pc6C9tgtVB0ojN2aajfL0gis+
2GwbuWV29t5Y3ePmAWmrvtn1GGbWMoUcTjzk2+nf0nT5t7jsnloKe5wmCS2CaFbToHRKjcSjtSvy
zKIg9cSTtfoYJddDYWGzBtRpwhIC9b+/o+GaJffzAiL+luoy4bhB77Yf2umR3Pn2zbJgCu0kce6n
MTbnmM5RQKeWqDR3neCPtbBtePne3VKXG8ZM5zF7szr+0N9Rs7o7OmfvhE1tPiiEsFhnU0BefMOU
30XJAv3O1zJ0rBf/RQAzoOJhQ3f094xszVCB8ySTUbbAnni7/iLf4ofndFOjUyvB/C51RbRCQ22c
H2RrKaDcHPoTBVn8FX/pFj/hgkD8nvG/aS0r3Fh+XYJh3di+5vpiYzOp3xbn5M+uVsneDzs5Pg7G
ry4MG7apT9J2UjtyfKsTdHoAE0SDPZuhwYW2Oy01rnuvp9Mm9CQ1O6lztRMizQ0pFXFhL6PqT/jj
g7NirXiqvy35Gyo88lq6Yix+fgc6vGXhgHBchxPTV0RpJpw/i7h77BCX2IuaANkkMGwuwKqb+6uy
spH9RpvWIE8Cw2bra4w1kuQY5lEFY9CRBOUlTxvuUZ2XUouHk/NX3WLRX1LAR3cd2yLrW97kNRpJ
zoVrdj6rlYUVAJSreF5tkKLlR0uVUgUsYc0P4Tyq/zmPiWFnyw6OwKLKHprZ+lJGya3tSVl3wlbL
+DXXf/v2jC7O4rga1o4SY1+7q1BOru9DFgZGX4C+Lu+skLtB3fl66F93DwaOHxlF40VChTqv/xJ5
iLzklasi9F4JS38JFBrIOqks2JhUHaaHTI2BhmSTbt9J+TUvkEKi2C5o4ebOJUbIKljS39lf7NqY
hNTRs5C3H0kcxmbO5mK4wB7zAeV/oLLnGwgg7DW5O/TpKZpyZASo0S+0UD8MEJCwJwEVKuSZqnAt
cvZDdwaGU66FghrS8I3GExCSsvXckTHCnfzONXHCEDa1Pb164R08XWlvOZ+VwgCMqJB1O4LK9LMy
ZcvieXAbGQu/l+uyvzx2A0j1CGLcOzdt4IKOUqf3O/p/ujmzNYcfdS+d6oDRDEvjGO9Jxz5UB1Mv
nD4cBxFfvjYKzOhxReKwToU4LWLBl2oqgxx9Eb8QWt7KdDLa1G3bHpveivoUKtUF5KKzUhM4cbm9
xAy8UjsB+0StPfkKEJY8yLLMR8ByurpLpL4mmg10fDViYyVC2hGKk7JdwyZKG1r9uFs808NPxd6x
BGKZp9lBBlBd3tDOPe8JLJHOCc+pRjw6vr9OOQKQyrfZuB8Gvxc+U1onx/hiPxtDF38+M9YqSXF+
qi7DbxXL78pgS2fOGd8bkYwufRSYwFjDkjTSckzkScrVzS7v/b7ztcIUQVHGi5CcBAksgU/17hgR
CdQTFsMg8Ajwc/SKGDnPO/KcxUK2/1k3oGhPzN/6uIy2bauaJDn6Eg65YmQW+r5LA1zIwndRnISh
Im3EMY08dhQTX9PgTO9JLPTzKXhJ5ANwypUTdbRkfmRK+1mMPA4AqLK4iPcQr0LYxJizUh0SsPtX
zpdIe2x5HsZDIaaXXCCY5IRXmes9jLZgAtlAQKoB+2TsW1+tPUzEd3mxBmXWcLFY8UDG4p+O+IpO
4Gz0ECDylAJfsc5WMwKXmScy8pYn3iso6kcUXpO8ABiomIMNT0c3xFQDTvSBdGGLnvPVQ2va8zVP
sGgiVsa1vbaOhtstw4OPDtSleS29ztCOU9DDCvGCBw1H4XHjmFyjnwRc6dTQNJxYVqhB2y5h50pR
fWdC6PPw7b373m0Thw0ms7SaQXuK/VECqzsvKxn4jc2ACUmdGm07Fjx3YfVHXR4r8E/ZCJeTU0T1
c7x+Kmb3pCcRwVjZn7oF0/jWYzoDxbdwwZug+vrpJjnhuYB/4LQYl/YaSoxRYHm1Dnk78ipNdKgU
FaTmCjVN1tT0/lXfah3kscVl2yTY2ug6BPUhK/BiNdmDzeRs+v1syyCrlFoy4ZMXXmTydyrhTAID
+pvFq+toYTFMh3rV5bfboBruiKTEo6JyhHEus6FoflT7RfAm9BxapN84RQfOU+PXZ+dr/jvBQ/1T
iAOSzFozDgSCcGjlPM/UXP3nIriUyLCZNF2wG5tWd08lfXm1XOY3+IT1NGlYKHVYKakiqZ55mo7z
Lmqmo16EC8yxPzIspjtNx43vxqru5xjY1/53leQhahUIUucklD4GLH+xmiPs/TP05RZCl3kEEb5m
lK30evvPyj9Bm3D+EuGWFwkJuj4mHWQQfsuf2/znuhSPFFmhp08rYLyl/XwHFzMpAwtTnbJRQjO9
IBPynUBTpYsy9ODOkshLP8SiFOUgPbfpIw9cQEJV/mBejIURZs+4g57b6z8QoFoa95OjYmGlBWEj
wvmOBb49GpATVu7P6dOARQLqeFHZAZ9NPurwgd+g8D06CacdAKbqhuHMP0QyD8Sty+22CD9saTIG
y2C4JOobCKZytQUzhCjNifmJfsTyAbMkIjDXGYxUX2IqjIKusHyN6eUXZZk3WUOv5+9pDfFTYv8Z
cVgDh3ar35uDbeMm3fbMnUNVmHlUEgokFsILtLW1V0HBO+IAB+v/X9NRrV5p5pVs+qJIz3HnXJiC
3DrVQGMZUOnSW69EC7XPRL6tYdS3vYSSMDgBKvATKaWlk9fFTdH3BeaSjaIHRt71wSSZvn0uN45l
vzEKbxhoP2uqEIZIuR9YPamveUYUA/zC2kljLWnEDUuloZgOxxP8KQdCKytcsNYwsWMfuUVedH0N
8nqSAchwx6bsoTEC/JLa2fHPhsgG1DUbuGkvYGVEpmm3v5ICF9XTB5CGJVKBFHnTcyz0vWy+yyTN
uw/+mYOrem5qqg6awBiXubatHR7PuBoYHIY4kwAjR+xETtUgqlWhPJqDskLzR0DvedRwehUuHUEC
b2YA26i4IgQiO3yErw81IgjkZb7YrId/AZBl32nNfo9h4FZqsh8nSS7d+iI2BHjTdfVqS8d2gjdF
0Yv+Tb6DI76kKcIUjLGSWWHkPV6D2xTEzwLmIcZz/wxxkK7ApGrzFP5cux2Q/Ii5ywZtTNLfi4Ll
Hw2j34jfpfeKlaNeExWWA8/lo/nttAL7Bb00jpTVhrsG9Rom3bMKeJxV2H9BQ+0DBeQ1Lm0SARoE
6WERenL1QigernNVMt4Ba49WW6T07T88biD13IHcU4tJYR8blCmrXxgCKwqjLRQwv7WrHm7ZEv5D
6csYTUx77Bfl1gZcwV6iKESKC5TKKlerDKKCg1SxkRAnMFaV8OSztF3e61iLTk3nNWCpU7GIm/QP
0jKjgoce8hYUvCqLjrkTrD3c7Mwp1pwyrEO2CifoXbV2qvUJ40Wxvf45kCNnOyfwcDJl3TBDf88p
sHCqs/xv55AJuEvIpK4+FF1IWxfxI+4PA9I86z/+0C0xpcEqQhrZ7F36WwSymMdGx0nv9DRh/HlJ
a/uc5yWAkWEdSBqFbYwFG+vNXCXbO+c8TpTcqN9nalQ5OPHkDyCRiugyvbF0iXwe1qIPdXTM5SY7
ugy0XtmD7G1EaXAElIDGwY8a4LFrML73KnVFK+zxxrrQ0FDazK3TXVKaz5yrYOKQmtl7EN5PmG8a
+q0aqNcrg7KaJtVVIPDS9zZrt96e1YX1HB2gF9kEq/Aa83o5ROFx06KfUV0x5BF0ocXfnxk696ox
1bF8PxJEsHfEBaJN9yRlQIdlDSm/DHKOOy4JfA0fI0W6Yzpi3IJmQ54niZSR7aP7kRZK8QCpbEyX
T29i5yER3TnvR4V9tbToKR2yI9UubMs1Js3guUx+bbW9FJNOWR40uAt/krF3S/el6xyyrJA1hXgM
YUCFb+En2tv3P9+4jSq7P4AqQ3LAuXpfoXgkOTwgSDaeGXVDUYd+47QamYXaKMX7Sb9oUEL3vbp4
bRRUSYJXvi/uOrMKfedQCoeNKFq0kUqtbaIwe/yoA+lNkkGR70pdKNn/aduScbJwZXEBM6CbNnHO
4f1zAL+DGvJIPLKg6eD0OP9M8XNpgBFKDPbVg7wTZIiwkOXAwv4ErhxaNs6SjxAGAyDouay44Qfk
2q0rj2VxSUQkDj/90AVJtzVMujA7phjmIWl4ARisW1zdXuhT7Q6pF/9yQhY6yH/QTCyH/P+ln3iI
R20GsbN3CbGj78nWm5SMg9ACsw3XmhSY+Lqp6X4mkZhchme2xjC3d14ljzjimbJDmKTouL1sIyvz
qPGv/HjV9SjVYS2WJzZFU9eIVYhPGj0gj19fREjKULQRgS6tIB9YALZ3POtjpOaKXFtr2HDilNr+
CQ2zUrawFI5yJcg/aAkw/9JrIEXQ6YCmUbL/pqEIr4ZnkVc6roctgcHjsiGcETyvimyE+Jd5dO+P
95WQGZhfIayILCVSd++uexbOiCdQa6wUvMVbmtDjMrOsxK2ldNUyPAPrV0gROoomyMismtA35UVs
Wio93SeH9cuSWtw14DRpw7QQ/DyvakLATWeZi0M4bcjHfPRrr4WhurgNeal9k644N92VoPWXVyf1
2jEeh2zNB2sTvdeeVIWLiG9tXgLyJXAIFslwsUmeJd/5n7ywXGbSAZ/5KI50UOgDsERSl/JVrzli
mD0E9xnyntv0ftIpC1AAkZf11WD8Mijkx8elpxeW6NfZgfWEzWdEnB6vBwR+t0r739mbQsyiD/pa
HkNhAsqi9ect6ObhaE55E+0vr2K/gkCkV8srYC/ZOskw05vYcOGo5oBvPxrLTKTan8TDFsInTFOb
9DdJYG00B+gva4DzGJgYf7/SGqSkj6hPZLxa9g13/3BfaM41m4uvh52+ErLeBifJ7GLy0JuOa8d7
b6gN/gkNtBVpnPWL7SuuSqm0S6t6VPIJG/2V3//kcpQuPvVmHuhjgcB/PZeMXBUuKKltHnntlQvt
PluX/VKCXU+mdev8Zcu5xisRLbqeIC5ulGlyoxLAP7BSIuCSV7RxatyzucEjDHHi+WhC2Kt1OLQR
MKACpCo7lfnce5T4h/rXxhLzuR/6msdJgX2NqDTJmEkyTk2WUSjWVQY5UPcQlXGISDLKbrI0bhk9
DgIjQH8OJT6CFZyEt+0tNuRiPMEFe5MUVpZbnzPEBbn3cQNTnIWLa524pBjGMbus2grN2hYn/XZV
Sn9ZJ3mprGPwjTRKQvYwl5rMZZXihGBw8QVh740yV4XtSLSoNWQ+OBIQUnbxpjcDJTfPY0pn/b+t
GxKMuiCREC7oeDq0sjK+EukqnS1IrsxT34Rc1uosKhciFq5+qB3LEWz85y4avQUI0yjsJ48ibAnb
pUCD//pPNbEF6F4r7MNqHp1Ue7rIKtIu1N6gj2E9eLL1FxQRTkQji5tg5iFTRUTuJcnyoTDoZPMP
92DxYmdG1l54d9HKg3maS0vbunrA7wAZ26lm8TAaSNf//688FNUbvuSUxeKH5xq66GgmW04226vp
vHQG2ntE0sO+VeBgq343Ps5m/3waqk0kULlT52dmG/7RnRfC5/4TCXIdnQubxIKUztYww3g4LkyM
SI7BILnGF3fEwRBWDXAIHPFr3pifGqkGEdN4/caIRlP8gOtzT6uv3m2t5wJ6I1d5q9QroSmLLT1P
qrm72N6XK8F+DFOYeSsLO392v71AVoJEe/kFMQTLUk+PMSkGbGrVCkHXzBra1P5d7HhhLMdKNrrm
ZKuU//G8Aet1a6ifo+o4rFI1Y4hYvdq80FIDZvHg2aqqpn+wNpUhETquN5kQR8CSf9aTEC81rYHH
SMW8ye7Fuo1W/3PP1vvgt7L0/jdXufoibEyHbXAfkxM7va6rJoI9vn2sEwnNtYGxJFj7+Mg0pF9W
2vf5uhBizbGWxgJ+Wnqv3VldENdwRTnraJiMrHbNPx4ZishkDXaL0pBDEBIYM83KnXaJZPJcDZy5
LO9qXm/1WFxE2/sDjsoDYEkkOdhthixppakVDG/fiZL4ZGaHnzxyKEz4BQKfM/RQrO8aNy/RLZVa
MQ/+uIaKraHy8JsMBEG6rvqyUIooZJosBllK6Hh/gjJGkIUf8Sxtv+GQCQ5iYFG3SMME+6Eg0X9T
0Wz76nuLTOl/1x05BU3PujkXFGeU0uhlumELZXo5jWW0w7nKmKJA9WxgTKsC5e1OJOIe92jMevol
/ZLQZvbyXQXtlnngbpVHvQmZ9a4X5w1KsPAnJ4961y/WNKFYOXVGUljJtCtKFzW2L14smmEUvXE4
aOvcbCMV8DfAR97DvY6bDBgS+y06cTGqJTHaytSD1Xb7XxDWYLzYyJxc2R/T9mzy279CHeq6fm4x
qoc7/DBeBV262o61uFsthnbyoSKxN2SNd4xeL8WbDFO/BrdP5kdSEu3HIEeFBqT7u8OHmJbfZtFW
3oOEgH2CI5SKepYDB2QI+57UErgDFBzZ7Ti3zZXUASvuO4tOWrlJgthHDa0JcF+N+UFCT67hKFuS
9esuzCyA3Ah39Z2ZGXbstgugM5XyZpUwb0AHjejUN35/5ZJ/s5upWyygUI0MNJ/sP6qF9qP3vtBu
l2ss24ZOBmAh2/IoQeOQBSNEpq8trcDQAoVu0nEzNpdyZvhP07vlfB2O2fcEpPA27mRinuYmb0f+
Ll7FI2oEwR8CAgbZRiJnDqs//AhhmQkV1vPhDGE9e2He9L0w3o/sJTOmIwZlwBHpN/WXNxTyi/C4
piUgBZL1b9cpOUZD0MoN2CDfIHAztfeFFUgVzi3G6SqAVPitBfFttWu/Mg5tl0/HqFDMdEprDZtm
MUCkjF+cOzBUG5nrWQo09VQL3oyNWn/cQ/ma9u331gfgoBG2elX+cEhlBBWKyH/sF/hgZGGHq8i+
XAZmiam+CGe3N7KXZNVWIfZRg+0Fu3YqAWPzQ26MkEo/dAfj14C9EfnyWyUexeUC4+7PQBL7q2UY
UNbfbJwtgPgWNHeZugNB3EDiKIFIRPdzjOyxT1DBPoh5KXPilPzSeVj73QP6FYlTb/+Pr0QmF39u
nlSuwZlwP0hOoH2lYLImM/VCthnazsmRhPybIRE+e4GT3XwWHJ2T/q7d8tbJqGVuDH3cmCEJAA0+
8/YWIKjUwMBZa/DXpu5iAepKqzKX8j9CsYSeZbcU3nW2qgy6g/vjs7qaXG7WSvLZO54OXpVtOZKA
R5OSTVxeG9UgTyB/TYo2uPkgzJxAqK2lQ6J7VWQa1kpJ1NIFWYDLHjilRVsBWLO27+a6R8etdrRZ
HawFgzToKUNA8oqpNjbQrcw0cXkYckVkcDrAaFencQ9hCBbwHceEbYrl6TJBecMfpoQHSeH2bm4f
GMQmeHEjBSnKkdwsk83RQN5sxAxfdQmCGrdshq3q0W8Abx8BO1eNyYFFtKBGfBxwT30nOO227Nyp
ZIC4a6YSG+/HjkqRh6DeCEM0E5J77hAO7QvPfzvBo9UNL237+tQHvhLffnZ0M8DTeoufJO8jzgdv
lGqtCXSbuczHVdqndgJIBWPppWcQUiV12UkajIRb3NaQJMYIPmDcTwqUwGofHj1m9Aw3SXUwNXZD
f2+357CPdD+MnHRf7M8rCOi3EZW99mhY+SVEsgLodiZfICb5v7RYUkCymYBy+JLtrTbMyvaGCEuS
aMXAKtiVcTYPaB4RBNxssChxi9fZA4770E01u76WL2OUEk1jhJVaj04k/ITLNmkQhopW7TPuBDYm
WnPSsopI9C3FnZrgSDCUn4hZOwlIU+xYximmGXXSuxEcs6wdMWClyN6pUXdUte22rqF2oqAODZdH
6Wg0G2ATYshRtcnv4WUclNXchC7ZKuzBBQ9Y5wfqAuVvvLFql5KPU2j/DOZLIl/tytqyFt5PrGqv
K0eNcp6RyRt9raisXbv1iJJrxhpTDCsKoYmw6jGc4cxpNQXvKsZemwYeUqoPjogGp1L8zrR/a8ur
qdxzJ1PvK1ojoA7LPsxz3rULZxmffbsDSEN48O+DtJu2N9YnfDR67G6M8gVxjQapp9KQVQhf+cP0
Ixrp33FOD/lSOKhx57Ser4iouQQ26kw0PnM9xEPi6QfqQh+5ko7fTLum4zFX8XSj6eJHs3jBC094
ryXCV40UTLbTD+C3QdB4rUFki7KvaupiCgB5oT3ukAHxHMLddrP2sA1fkgeZEN04TogpIVlmTDu1
LmllHjukgOwj2m+JOLMmDgzOKegewCsliAOzkYEM0y932lQO7+w+TEouTltkQdsY1qtxdYwpm7hk
a9NxZL6Lu4TMftV7ueia1VbFoKu80zK2F0frv4I7wDFTjLinRof0u5+OKIFeh2DdUZqm3XCHMVc2
28/LqQoqZYQsqQP80PZwi2zrPhys2YIdu2OE12pTXcX+S3zvrkokDWungCiq008b/RCQG+hvG8S/
cB+nd6SELrdwMgUcM2Zfq9fb3rPjKqZmgLdy8O1QSBngVsnn48Gc73rNsCFDVOdoRnKJhr8ea+bK
P2J1oMvR0p5ZGeKJk3Vg0wUJGcr17ZcopnTUCQmUGi4kc4HSTeuy3hgjCvpGylCBmKsTcXeLqBxp
qZTupIh7dL3KgcztlMQLkfCJQv9J/TD9rdVOmUipwYXNztjm1d4D7krhBR70IQEs3cN7sIgE8iMe
rLGrNKmrEDF+1jYyYkSlwpCPjkVzmwkaZYZc9akD7ddepGMlPX9wK906w7LOlgMj1NoLSHsWhvxj
GQX0KwLJ+Yig1YWMuwjLCbrYXV7DTy/7XaNSN6WJZsGz+YVVco+1mncd58FEqfIGTJC+8BZ+H4B3
RNO9UHt6Lwfindw/VXYCnZxZzczCRGNl215hngb6AonYzcga+QY+F7KUw2RCZPS9l0nKrhBLMG2a
1RIz1zAaoBOweV6kqFSAez2iNX7zuBKA75szN0XWXjrV181efnSrl61QhXnIGnPJHhangX6RI/8z
dMdxp6ngqn19QS/p/95t+4utj0QTNEstenWFZJyY99RvBo+gV63iyYo7jtMwTx18lS1NMwd5RMCj
D6irR3dk01b8etA1YmMLgbzGzARqQtyJbpl7SSDx68Ug01d2ksJ9Z1SYh36+vVrfU59RZ1YT7pXz
1exmPvMA2zM6RlEOQEaK1yZfzPfMt8wbg1bWVDQQf5VqDKxIvGTkYpXHMAodYXNI7yx893wJF7ag
oABfhuCYhPPPEqj0vpkj7d5ssA6XQFt/pdJRUpGH4sAxVhMow1Pnrx0uNQBazg+zPgKCr4QFgcRx
z7DXiO3QbR4E3wp191Jy3FovNBGFT62EQMZX1oegn8mb4S4WNVCjsYPP1ZZstaZahANjc0HsMGWP
//NhhOgntrFwRxkSuhzbVAxqZBnhYgbbfJH91xFP+2pqqi40NmR+tDTWeQSSbD8o6SB8duA3Amqo
sGpuRyOj13iVA0WstqD6TjBpWIS7xi3OVCw/J7gaXZHXcuMoEBwJHb9mN2hs/7SvoaQ77gWZEH/O
0vh6Lobgd03Kuk49f8WL/asE4AN1v8mUMP6libmCRPz+4guAMA+LXkFiiz5j6tZe1RXn/Fqut4c5
1CtLWVJPkFDYOjIdkamsbwv0RWz6cA6UdxzxkIK0OVS1rMraN2Ogv3DkDWsT9D1KMJX4odyyEMSd
Eq1zCaShO78nBhItaY5ePWmNQOj4kvYDXXqBtWtj7B3pgNJXe2fvxTrQZGKlQXmmyezfa3xZMqDU
ZZJaOR4NRUbNGVBEM1JGqEcze1tErtiCkEyIHEsw0HetmGWApSTKspw5dDxV93vDmTdggE/L6eUz
x3LptX8QnjlxtUMDRK4FrFBXGTIGMznHXLUI+8ZIQhI/izgVZwXq966nR6gACsj+tj4KGkRWZeR2
mj7ISJMQYt/N4SPgEsSXo5g1wduH1wyVx6gz+RucjhVHqDvpmYC3vRXPzjZrUA==
`protect end_protected
