XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��rBڨ��mӆJ��M�[�a8����y����B�iI�8{�Q����?E��I�pҡG&E�a�1ñ�D&,�` R��Tl��V��4|�����vN��UЧ�t���w���3	 ��@K�K	����8��ci,:��@ ޿qp����f�SD����2�r�~X�����\��7�Q��^ Uˡ��1�Yjqtv�:�$vngo`�?��aۍY��w�=vǇ!Q1O�t�ơ)�T�p2O���L���B��ݞ��� �U�.�Qk�J?���$3��ܹ�������8A"���p�G��mN�+U�96[K��N�����ȟ(��'�G�T׵ϖA���.�Ϡ�A��
�S!��M��i�ƴ���xD�s剸ĆB3�������:�Ί1�^zUH�+&c�[�"]US�]�����n��dm���#�Q�&�`ߪ�3D��h�L�Ğ(��/ZK:i�bHy���[���Ӹ�^�P���Oc�Y�����nr��lܣ�QK��W���� �VV�X-�M�0-Z݄�h��l
܄����h��ݹ�­4�E\�ײ�%�h�]�
�d��.G篩^.d�寋	��$����@���.��n0�]�c���<����e(%]J&��o:�g�+rK�t�?W�*�֒��}.��D��ƳD�D�0��-w3�+A���0(��։���<͒]���3�WHU<���X�\-�{����zNqa4h�Nu&haz6����
@��,"6��I�XlxVHYEB     400     1a0|���ec�Fz�l�5{�g��N��-w�w,�&�r���Ҕ��^x]��/+5�@6�ηxcb�����nϼ�OPƳ ���H�5ӔR7*���+���������.�@(��m�}���_�	��TS��������=�Dm��1)<�ܦΆ����@��X��Wo;�@�L.�M�᥎&|�;�v�n�v��HA��*��(�Vٽ6R���np)�ZrV��e��U�����v;���U�$p�v0%I��{d愿����E,������]���uȿ�S�X|l3�Ҳg��ݤ1��V��'����4f
�a��{[�	ۘ�������jk؄y�IE�a�(�Բwy�_R7��g��Џ�֎J�<s����@��`*X��[��~u2�7ԥ��
�XlxVHYEB     400     1b0�j`�D���4R��r�-?���7�����q���V:s�
�B4�$$��J|�z�����d��N����f��=gj������^;)U��mK�������w� !��)�D��A똊�N�"`��U����9�>�צL���w,�G.\^|y7�]�Z�ŀ�S���V�;�5��
�Ʃ����N��o�B���+��]F��5z�j?��(Uf���/	q!�qLk�mˤ�P����yl?K>*�ͼ�6Мz�pҎ �g��b?!��J�U�6��%�M��^��)rr�/"Ȃ�����n/��n�(�#)u`��ȧ�Z��ZK�-��p%m�1���XW��9�	*B+w\�/��,Kv�	��׵q��GFJ��,V>?�B�wY$!�ޓ��(+�χ���%�
�+��x`��XlxVHYEB     3f5     130���\�5��FU<� z|	V'<L.$�������E;ڪL�����7�Q�����Qu�7�Y���{�Rx��M&%�.�����J�?^������"J��`c5��n����b ����^�������J��M�o�B�Ab�ZE����lqG�b׊�����s��I^��䮯yq��~~AVT�/z�Dq���/hDۃC�*�q����\�@c5[�	��5�-�~�X��"X(�@8���l���O�F*I_�~� sQ��׸��	��Fy�D/�!|�m&��4��ݍ�ߝ�F