`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45824)
`protect data_block
SUaP+dc1a46qZpxp//utQkiXV/tP1yBKQprYhR8I9oN9knczO+EuB4xA8zElruh9fthXWsMqUiKX
iT5WUbARS+CKShB2aSVQW4R432RQ9VCm5+NWBFp3LpIZWo+pGwPmqGj6a7re15OkNVf0OBe9N/nA
WsJKxR8CAhhkUWHwWrlQpMfwh0G6Vt7zDMMJp4f5sMJCX+r42NF+hPCVi7p1bptCJCPslhUzk+N1
XhNYugnrKY9kBe2xaz/e1dH9tWYR3U05oFPcOt47joNyQIGulBo25epM9JTXCdp+UTv3yVp5n6vU
cGL0CxqXCVaLHXfz55SIKxlaXjZJpQyychzdw0x5Co3kOAPh4hruUPx6MXmm58Q4Ow+7EH5+1IxO
LrXA3PLD6FCCu342r5SW3YarE7tdBJUaN6/T1UquV8siXnVg4ZJkKBHdnYj+xM9C6CKaB1Md91YC
WRrVVvUlnAmvS/EdXz2CFN0AyPQ2sOMvayBxv7aGQoycrIrJYqDfo/lzguF2WGjAaM8GWljsWTqm
F+tTjXypqPG4UsYWiBTBl9vKH2vJkx4AAZ0cBvXfRCANTaV+vl6V8wZpzf3Vfquc5tGAHxyx0+4f
aFHpT6eDdIMFdXJpjSVyOR3nCN2XwsMhN90/3Z1zQcyxLRE+Cu3S3z1bwJJmp0nb7Z/g7VarY22G
vi2gw5UISgvdMA3NSBpQYLVWcm7+eYWDvDkXOiqD2RVKM5+8YjoiQ/jxeMLgH3MEgOfppgDu5VqT
yuiGuUYDIYvV6VReE7gE3umFcqwVafTJubklgGjr7Alhm0Y+9nAoTyP69JWz3mdGJEIarPK+yZf9
r+ongQHzsy0bjc5u7AeFtZMNtQWiVv9yeH/im9ohe9PlZKvV72tWTvmF9UcBQZ693qiRGI+h8n0/
hxdr2KBvVjj8P96hNCWBQVCq9pJyRVHjvQvhino4No0kCdmwY+khglw6w6GyZKyUhTyUxu12pmGR
nPG+H3FtJi2ilhkWRQjbPvf4+0FFBetO3I0nTCKGBX3sGGHcMMTqICm8DDpzzw3nTx90xdR3engT
0nYVt63taFIzcPRawk4nZaalqd/UOZr4IrCNHYj4c4e6lzLEcYLsnL/EQpMH6CY36JxV2CDIkrP5
cKWEysQM7bK+x6sTr0eANFHR7GUblqlXvMUS8O3nBSDSiQLPMgAjKc5jBtclxXa/vY+IVTVcfjxz
zW6qwjuM+bAzTEISL5cweV5n4f5GBP3GxeH3yjgRKJxUvvUvS+WsE6gpXcZoc9SLs/2JdBiFWxGI
E194A+yZYPLNKQo1LZMJl2nmf+FJDKCJxGGzWeKwVuqSLu3Ns6LH/V4BMma7qmu1lRyweVEVEruo
nnQhMnv0PZ9Qnl6evLOyEY3u70W3CR7Z/wwtJ0z6I8/X7tBMeS36L1LGWjH4o+7emYggLanv39l/
SDTXkwcyPg9jyjZacXfC5FIgIUY00B5LVJIcZ3u6xtwGQ1Mq9NqcJQDfIEFkPN8cHOoNtLhYxuQa
tuYMA22ZqUOhFvLfnnAaqI+Qmho+4dDCTbrsOct4suH1sAcDYcvGjoEugPCQkSrAS59A4G4NLB0u
rVFKlRFoA65mQMZtpSSt5Fi9AFTrdGKAcmxSq+wv0RLKfr7mC22Vpk+uC2j8zzeP9YCtSV55loLp
jqbbAcZSgvSdyok0330Jcug+FfhxdGlEjfTgHryY90GNYwp2XQogppael9c67fQ/6wmlk4zCXaxI
sSz5cOwmRw0pd+wOlLYc/G1ItCwtOk6pL6STKvcF1mm3mmUHMB9GfvZGVN2A29I2ckP25P4OhAV5
ACK85mpwOdLgCJJ4lsuCZeRSTxCqTZQ+xHkI8GvFVzkpxUE7+eka2W+3yDHO6u/NMyxU/zO3B2lg
XUkr5uFqkRGmSRLrtGKocxdlnxZz5z1KCOoO2PDHW1Fu0jiL4/J8VA289MrrRy0dV/gNE1998Gbx
AK4Hntw3kbsZP0abEExzGj4hL8OqIiWDmMB8Q/5wzvcqpFVWs9Hj5heUx4fHZGNMd9tphUB0A4RA
smXKj1ZbOgzAa9k3klLq/k38KYLiPyiSU1vKVYJQ7qC4gnZC81pPWQwDXDii55pZ+us9y4ULXROC
LbXVBUmACEkjYfISr07KB+AfuewHEtIdjDaNuJTXTXe7Ekku7z6cE5dkiRhIcgWaG5eBDZeStaJ0
hvo1IeegBiA4Wrlfzoi/zWMD5aui+TBo+yHjVUgoWknDYzMxy15QL5tqakgU8ie10kVlQUgtDdNE
osmoQR8CgEqbko8ezUQ1q1mgmx//Aom8pf7/1Dixs5tIj1AxkCz6hpi/MZNver0NDqdHrxQSyyUa
juWSyWr2lqX2KMb8t2F9XLbMG85PjIUbTuIkXLyl1RFw8odgqvGKU7sy5EsEXSIaHjYF35cJzfIW
5TZktOc98n3IkV6emFLJTtPunlbscnDhFdt40YBDyWRv9I3c3OfaTbWr0aniptCouWUHsTZmBlFZ
xYAud0DN+Yq/9KqYQNbL2PX7BepWWCWpol57ylHaOJpxLLLvHcDzXedIiEJxNF8CfX7OoK3SajR0
5LASV81mWN091uYpiptzH+VP2XQxmGznfNOsawoivrGHIxvQ35NTySyWVT0d5f3P0kaOMzW73r+8
vUExEedKk9O6uGhDNOndYZT5D+EFOelGequ3wk1dhUeHFtV4BL1s095nNiLie2diatxOEu5tGEg5
Kg9jgsMqfho4ejYYVaBhD5iB/hutvTxsAzRaSvDdRQOOw9RTY+lCBh6Ls/o+FrPxqYIrZZsMYR0b
vzrtdswTI+6/utP/pjZUF3itsi0HmI8MUF8yTzmUUWnWr2XmkSlIaTubp0Zlkb3F9MvdxONvQIYA
l/IUPmsuj7o86gnMErSNtS1li7NPg9TTp4KqemupC27EoTwXV+P5NeiboIZimyBh/h6u6LFC3Odt
5Mlq2zU8Zf7EgXFPp7EOJOqRNn765vuyDMM6ttSvXqpXspKm6MeizonJiYvULLuFS7RmgMPFRPaS
CEtDsxVINCpXrOkjy2pLEvOsdnh8KvqC2mT9GX4q0AolTV+clESaOBg9Ci9K75yiO0z9Ze5s3Ag0
Riqp4oQImW/H/IhRinciidGfOFKDqd8gRUXPxNlZtbc5V+K7lEeI2XCG6lgDPSChXAmVuAVPQLqm
zCrdsqE9rkZvwGnxvUf9y68M3hjhOIvO3GSN1Z31hv1f88GwPKaqr0tgzvw97D8lhsT3vxi5+B7U
+hh2YWNZa9jvBR23AY4Y/qh154Yg5xykl9NexfPKzACXqDLU+ZTgrwES2KO891eOxvQJHMEwTmJM
XE4qRjW4ZWMiccalBF37UkDA02xLHzwc2E5vTZ6BRv+B644MluTuE/HCEV0wm+DZOxrGX+QQrdy2
1bYPTWX0bnQgQ+l/HzluyZLQbKBFLh7w2uoEMwbpnBmaBgB/VtFrgim3mC3V3HmzbPAZRBlOc1VV
nVKJqEZr6MK9iLT/F7wlYcPrFToozYSTEuKGci4dvr3cH5gFrVvueT4bcuXqcXWUIhrYpKGkISNH
7LSDHJOE/IyyBgAJvb/EzsFvBO5BzhhmPXhxDUBnF04sgLZhj9gQIMigaoPi02+Vmpl7DaXlYh2f
3erQIJolaZFevvzNeRc4qYfBrHAjiH76N1hE7xQiTJxAtkQjAjJzn0iQoOc3zsBoe0canPTnu+v3
Xm5qKZspjMFy/2MMB/z9a+EzzUwW+eQfG2adYpJ+/GEL2kjg2P3+ICmC8PRKDJFiCoSByPpMUj/b
H3sJBQseTVaK6pKMIYFlnH9yjXxKhVLSlYIrceW5qY/sddXdYRRrgbmr6opagylDus3Wsi+jCdu9
G24lLr+vRDj1Vf14IyDp1j0ajDqCvygUXbxxSjA9+XwpnY5sSCa096grdoulZKAB86mPxlPEMnSm
Lu6K8ON31FtqMnwlBRJp0xUgJWJdV4fFmNa6ig4OwNrEun9g/qid199354yios/IfT5eEnnTQMjH
pZcnkdcSJe0wTCiY2VEQ7pQKUyCqYWxBu2mCL20dhHniuWdMV9UKCZlQMrynruwHTPu12d6Z3kcE
uG5BWlfhoq/76nSDNY60JYy/UAD3DrZwUfSsoRCDLUSGSJuBjaruCPf+cW0e5a59ipTo7nHbqbE+
lW2OKVSFGzBnb+2t+GIzr+qLsXAaKriRCPWMwLarLs+Uz3STrwnRlKvWxOTp341yjMpkK+/ofheK
5EWN5Nm5aaGRZMweP6dBDC/RRGDVg8Z1eafpO/QHET62rBn5AFnE2g/WCixtH0S9KzqlgICbDq7z
i1cgpAAybPAjjNYvImo/E20rilyfMpHj67tvm2Vh/4CQ01jq2q7taM42t2bw6SePYz6AJmZ2w4wB
a+nxCH9x+pKlYa2MlTDQDGWtVxv2wiE3lkb9uS1A6ff9keoeOPsQ2Uanj1TpkUAx//lp9ECxq2L7
7EBJYmhfT1ZP5Gbdkt9/nc2r5EsENScHh1UN8R2la08UwSZHKFIzgoa++iv8xkCeWKv8G/6QK4e8
mgRtVzTOrKhjUQgbaJQzKZwJfMpP1QqSh2mqnTF34IY3k28+FQv+7vus0wD8h7XC2+9PtqBzWgs1
TqrD576195ekz+gHGK4W7RKEayKolGGt+yk9ToAg1J0f6/5piVKEAd3VEPisnGDms7AmBFHewsxb
Mfh563jK/CoBAA5n1anE4fO/fd1nXOmJ/eAmQUKJRr5P5iBS8agKJGXymkX7QyKtSHDITmGL4Bo3
zlhRgQ+QNRTHGD3vej2hog5XZlxWRhX0VklKV+A2Ry/O+GPfA6lMFdhBAdtQNSCFbH+2kiCUFuFT
D+j0kgfyyt84MruwQk6+D9EmedQRwhMb/Lg+zAkGvaMmuHD2MABRzNFO7O4mdUpegkVYl8Eq+Vtr
x5Hjx4fFD57OSloTJ9sx/PMm+JCPt9p3Mh214vHA4v/1v+YmYqzpGGwUFl+JQUzIgKdAQCBNB0Wm
AqilDIVWTbYQPKd15/j5ifV4qG3K73Q+ElynU8WA5JHBtodNFQTXow/OX9prnEOnfqqyubZeS/Gf
rZqeH8XknflU8sIGgm5P2UnLK2d40ew6ynUy7BMy9ykN5Sw4bCGcZJvBLk+zHaGjfoQEHZ9NwH/b
tZmCFCD1rZnwOeofqAO3664dIRO98W5RAM921FqaYq+xeTgupvHDfqtsWYccZ0VHLcS1bJMQrrHv
mScNuqeyg77wCgldHOqq6fdITyQgeTt0Tqf7qJFgG43Kp6WDh2JE1sa5WdMpKXsvtutRoH1c6zzd
RICTgsfaQy5sgP4DAN5+9KAFYTTCXzKCofgZCi7CvtwQphPbXg3UK1xu4wSDGaNADV+IodI1p/v3
pA5XhLwzYKPOQTzj3MOzfrAVzQ2VKs2Na8B7Pjytqa6Dtvk+3W6nkmFK04mYfHcnTIl8QJfO4VsZ
EEPTTTas2fUws9yHIfHHLSM5XI+PV9S8NpEUioIOdcNzQb6s494pE05+6iALrWLEUT//pRpAWF29
0tLKfbzDlBEfBW6CvbA33Q32at/s4weeakvXOsytdRnITIgWTfQAZkaNF1nCe1jSVeAVE1cBFBLR
cQ47G9pOsqOTiiRTO5NN0ZhUCeRwlNcyQqL/fsiCrLatXH3Kjw2ODhBZcJ3zqfwEQzgr2HDwQmAP
Lcjn+L/TXodnNrF5UsSL4mlqUBPdd6bjaCwhvIc8AKYiN6TS9chPh9jy+iRM/+MkRd2va50vY4S7
iEX7v2ZpClkhsdSlq8MltF2yJqGwz9XMUGVfHwXRZLqQ7PBtbwwuhMGOyqA2Qti7D2uopWLznqpS
j+XNvddDxwrRFsitqUlbHGrUYvExr+Ilivd1xMFalGc51VO0q8HKwe2g7VgYPsgVN9jflxHpLPds
zjhlrCAnAQOjFjAyxpuniMRJDJdlpoxfaqbqWu1yWEXVVXpibqLSVGJiIMm8vEF/ABE5HwEjNtSs
9DWrgampQqJt7S624FI85X50XhKeylqgK3+2zkFexPubWyImhJLG/hmLtpAsNqmqjbnMto7c4+Fn
fJr6ZBREODzq8lX+VQRi3Oxnl8/I2iF8/6liTGdi2F9CJ/8qtisupQN1s7ePDaXrxN5EQ87SmGd9
iAV1N3qnoOmr/yANdZSc9y/iTpuXRDg7LC9un5yA48DwgJZT/NbRbyRfXaAr2Og2wKtV7IC7eXHD
pNOTVjQtmFWjMIOcti62gEQNuCadTwDV66ykZ/aSvto/CpoqlATDH3FI3m98qsak5edQmj1buBif
snv8HLa0A3lWikYRKn161vfAfiHJBfLpAAyxJGwn/FAlUSWZGBIlEcmj2uNR7Rapoclqn5RC9B8x
yVCeLRIGSnSXEmliMhGwTV6L4bOYqDWU9P0Tqo9SWWQ6FhP82B+a1+iyzmnAIhl/cD73FJhl5vlu
cO2TqYXRwFGLCrwlaLWerPmmK5jJKXkbYE5Zov31TUVgHcGlXwngigukNUhtm3mpCJttR9WS8apj
1LJvaFf4pT/OUPD8OE319gphJFkzgMVVvTa4iNntU5KNTz2561v+d2nwDa9DzEp7ym404HFPJdIP
N+lYkWYqWWgvYsAdaUt0tmeZzIsefVLE6Hl8ePe1f9jKJmv8ZFrweZuDnvgBrcBLA6ePuLIBz2XP
9XVpPTZAOn83BgFAuycFKuN+zDTOQcmTf5nyy6y+2h2A66XDTejX/M7Y3dovEz+KpR71ge9n0Vem
2ogPFDuvdUNs6fYARTlSNevn4FAYB5dJLbJIQPInUvYN3TWVPODegpZl3Aftn/5+FJyAWg1oqu0b
QZHWw0fEg4+RM7hKaDQgsiXdNfhkdh4DOoa7svxiEy+7ZuQbd+BeZhUuDoagHKUJMV1fKb8KPFc5
TpDXFzVlM/3lmMSJIRPMPefM273gt32u4tHGNzroEY7aE9SQktx7IKNnR0WTbpSuYFGQb/DCW711
/g9ZxdmfR3p1gmA5h9HZpO4X60uu0POplRn5U8j5lBVgJPClebUpaBMU3o7bv+dbyyRlCQJCQj6T
8iH4cWk441LdtucKPnum3qLrZx1F0KR+3MQzuIGH/t51KKN+PcW+nd/WZEvwwqtqj9+0ZdQ8x2xY
l3YnBdmaY3joRj60tnpRMEub3Y6OQuRDniK0SfGdVrbkrGvyJgOQKh7Sz+1Vzw83b81zZ9JC8okp
aaGYyZEqD/IlbJ5Qg9Y9JLvrQA3sM46c0DA2ab4apdLwg4CB+C+bWg+NB5rn5L0EdqIXJ8E7AQSE
FZEwFoGxdWaD3V6HRw8y6CRw1TdTMPvWBay6CQfmAlwp/VLdXhz5bxLPd+I0wbz5fM1ffEfJT1wI
Fg3qPjlG8fn+rL0uUHMOqEHgCGi7g6o+9o9LKUh+xmxYL3KqZuv/15O2H9Hn1eNvhNPH8U9U2QB2
uG+WKCXxJxVSDGNa6MdwCUSffUK9A8Ls6YtZ+SBlI3b0pJRBmnoTqNgLn8IOl/SNRKSWPK9LPXFh
SY0ILr4TFebNTSmj74fmdtre+ig24UT5AGZBzAk0qyx0aPzzG35/4xx16Lc22whZL4kkbt/YNW2K
aCASJUj2LnduxB0JaKETRiLWjLuY7ast5Qj8EQyy4OvOgUWz+zmUCQRfzZkEoOj5DO/6gIN6jVq2
ZH7EEdSmyt35VVLHZSOR9oZjltnVwmEutIUbal6KfMKZSc4VEFSPoW+ujABC9ov7zqKH7A+C/XlK
8M+/lpZX3WErvuj7/3ZLw1ms/UX1dDgILl3gQGNOh6Ib8POCpk8CatyxxnKKvgfADldp+V371x1Q
Q9MsFrPl4gVqMcNnzA1ifnCh6GHfFJ2EXmpawjFRHaIAYjaFqDlIfkvcGV8z1/3l2WL5QwKmjtaS
xgoRTZ2SE/ZvvejZupioXYpBERi8NsnszmGX44mHJpHLBoLmFVY1bcPAg3LDV1XSkex0aj7CDelv
rdrv6Uh3TGwiBTyUNBtgOBIwa1pLYu0In0yhuYKoEduSwQlNWCx9V96QJpTmSAzJ6zbmq3U5lxTm
bWtZCxd+H2wpFJg4a7vlgb3rnrOwtPQZe8ONHjwPvK3BVSVK/zMFt76pLl3YU/KSRoOSDdbpxutQ
fu82ah278kSC9fNeeMjOqFjDy2t4kHqZTlgxTbi8h4aRKLyt30Rc3iZzP3r3edp+qVw9V1GJL+mF
SsUl8Vf7aN5psv5Gy5BjCHa3BddS6YhdDNCtX6yqAhbVk2r4mb9LVfjrrRvBa7rE5eKWsIzS6zcY
cxI404Oxbov98m612buH6kgrQSkNKsmEJDb/TaJaR6seHArQc+lE16H1vW2WHEacS+YLx99NbTij
0cQ94grA4Vqq78gZo2PSHYuqsEKDSgZLTlxWav/3BW9o6sogwmaF9ImtQSLaXE2EJnUgR8VFcs9R
T6SmhcsxHOeqBzi+woheCmcoNCB4ofUpghxt4hpusrkMI7GwzIfMFZfmEY8qXBATQxM7EJ+b7p2v
JERR3P95vaffNydAxZyXydmz846oAoimuDYVRVMWcHZN5rBly5YQSugM/zvq0t7cQMoP2gCXwiVG
VSHucDcn0faOfyzM5gYZuRNfmOQrgrLEq+D5LdAfQJRLB4n4XA7bmYKIYiv/EUJ/vhIvL/oZ8uuJ
DvIgp6sLQSmiJPFA8C+JE4COw4ZbvboSJP+qOhbU0KKwWbYzLdnJgY34JkOZjA70sNPaAeE0C/cF
zD6KIBIiGbEvJCYS/w9ofiW83snhm+ekvoahEuNaDlDzDbIiQTG9wosIx2IHgnR5T8WPpTFWlNNg
j4bm1muYrOWuN1mHN/SUMS6MJ/AI5xsPqi5jtCiCfJ14DhY+93zwyegSsdBqY32cxBzMtYW7ghcN
jHgcLzLTyzoV6OLLPi7cAmEwnAl3JteH7frUMw+NcDfqYKgAl1aG2KRJffK2XfH2CdJonMNE3IRL
9Iyst+gfQVaeM6ETdIVqkQsvTXWjEqi9jhtC8QL6ruWU0Kp2AqVUJIJoZI8cRd3nF/oInV/Mk066
W/0RmWl+WIYDvKVMIcvoNfsAWVuW9uWC/Ny+AT7z5XV9CCyJkmoiVna91itQYRoyNm6Y3MYZ05Th
0UHR3LiFca8RTObrOb554/2RdzW6mxH/OBk37EaJuTi7WtSpH8a1+KZ62CNEUGl+M7LVGu4sWAHF
tjUtqRhMnLbJtYnahl7sulkdA19MGNCtqCaBxZhHstMVBoRATUE0HBOypCS2Tkxxubi0K2uYjxto
G4LdLuIfRYz54vI5poTwUT4n9HGoRAMkrK0vUW6pRQHzTetYwH/Wvxt0ottKncISxeeIxQ4BiCa7
4+DjBX/9IazuTRZZ+rY/SJKiajyO8aKow8i22KKq6M7td6aIFL+9CY3ryCC6WnpQDqYtQr/2/LDZ
t1EOZh+otKs8MNKnl38eLmW9AdTy++SRmDkvAoPEOLnTBKYyPF49NduMHPySXodI85/DGmo6vOXd
U99KCPOZy1NMTlW3aDQH57DtVwaylpj8GZfqIK+d0ybDJEpycdbjS+CmyAA7rgiEjMR0svG695vZ
wdJa7NX0mZ4gYZbyYlUEnlySYCGb2omt1UHHx1GJCvdVcQTP4rjfaIrQLE8G5rhpaeflIC5PZOMe
ehjN+JQyhjj+asd5RiiAxeO4gr/yxBwJzL7fEoa3zB7Szk0rmP/Gr2Cz1SVcNP32eReUjB9WMoe2
NLfg6itPWltV7X0EU716JVsXoe6SPZ32urAC/lFh/RSRZpHMUp2hllljapPxI7ca1bh1CmtNVOHT
lmm0bgYTukHuE4mOpEOXqYwHRr8l4OpmphJgEF1WgJ0W76vXbojHWYfBRc6qdTLg8G2OCH6dIiYA
i1kEs+m2gta/bLqeI2f+bxxZtKHFFc23zixwrRgU+s9WY0+qqjeV3KYY1h873aY7mxuWytOaZ71M
AXYxXyA0Ap6EOMw/qV35LnryouJbP9IDwFiYHtmFZhd75Q+lh8+4Cjb1a4fQkIpAUJgEpMGaL/66
w8KtCKjm7WurgvMQunqNTha1FvMh3ESpR98L7ZhoUV9RmlFn/u+tgEadsA+H6uLbQzKBKaex7EjC
9Cs/oAS77dLPBp3o8eWWz+Jn4LruUtXJM8MqEKDdGN25UBNI+Xjz3hSGhS8Mndg9Kj980oGHfHKw
/LFt/B7ivvrPfLwhZM3EFRV/UEHYCx0b1dWm+bqQ/fw4WGaMqgSAUjIyLqGPABVyZKPBDx0pXJa3
aLvscRednw6zd0wNV5ijn62kshQknc8YsC39T2BcgHOhf00HduP0jg06Ey2lc2H2C5HYgL+kzoxk
T4qsQWQUiP/UOBAHfqmxMebDEuYR9taNZiHXxc2+hD6XIMAdw/jKgPjZaFXB5DrrDFu9afS5STwK
VdLGRVz/YQiSMKsheJM4uipFf1pw9FNu6IC8gvXPTzfzF1pCfJVhJveuglg26yP0HwV/bPLMALn9
Yb9/bfzdHmD/wRPF5SO+n8/NVpiiwATTzUKEnhIJlcDX1fUl7cl3RYNkOibfGCUfbiRLPzPjd7Lq
dpjTNT3X4AhSqdjDfe+9y5UKSDU2yI0FLzIThOp7gbuMF1cFwLYXqLOZcY8cpyLZ8HakIKhbOSf7
vmGpOkFe1ZWe6vBjnfyt5S/bwU+5QelnVmfCi8jrPqgxgF6NjnU5wsvgza5g/aTgd6sL8VsLV1kH
gaDFJu82uMF+jXgjXsLgGXJsGfhZjOcIBUcQrrbs9S/3BaEh2YUrZTVgKnaVTyeT8VJcXojdE2Qb
sUs5+ghaZ+qndOksaQKpuKtcywRCg+mZas7CiOzUBQuhvc/eLVq352tCJBOsW5zR+kLtZ+sPCFDt
Y9CepCG5kOjytXngrGtyfb04W1lKVb25GghRzbuxBK9ekQLao9SXiXBo0XLAZu1jSZJSSdr+Wqie
Iv+LxeGlSoxN3grLj2btnv8K0WGyi7eh+pJyy+DMAKe6visNdu80aoa4pAkEHeNZm3pThpVOJbnD
QnwJiC66wfFQA5NuPnFJ/6A5keC/SSuAV0JNfA2UyDBLMatdt2kWHP2uaIlIj84A5GQVpFkVIjHI
LwSBk+lzceFb8xdrvkLmPXWn73lRLJSXaW211fqdpWDrz9+Nu1+txhyXK9Ux+fpM9Vy5+Ol+CWEm
VzhXJGhEFt0BPqCz+xkH7vxvq81Ws7LxwrrbjCAmKNHBHI543meuoqJuwptNHk4ZiCwiFW3GUiAh
zKq2lPl/LlkrHlJEKZs+cvEVPc3SpxBEbGDftZASvDbwVTPTjR+jV9xYWzNXPuUoBaIqKNXjOG6o
ir73gHiZluyPsBzeyea85rWtW3BOs6huQWbmwXx04F4bynQzCMfIArwJcfeMBspMLkkEbCqbluxT
nzYKFawatl/xGUXakepeQcvMPGdHMqefFAkRZsbUzOQIE4NnLbsNhOnf2z4dXTCLB2L1dT2UaqnW
FdPuvDVFrhv1U2AB3+FxC/Kw5FKV21G9h5M2JAp41ouRGH5SsU44zVXo+l8WaywJ+DuVEx6DqBSj
T2/cWGx338jnlKhHJT3QgKP3hBRFWnsv7amTTQU9bl6jfPsxWGCOrxLgMf5j0MlTG1q5PaPdBDiP
trkoSnt3hKxUWN22iRMd/5h97sxTQ3bAkIj/IkRPQ2vqFDX5jVfANBsrhmpHZmtHnGILUrXGbq1I
ukYWlQDr08s/SdEwjewzhC9GBJmn+lohFbhUroopH0uzrQbAVIBTKvz9sb9f9tZSUAEJ2BiyZixh
Ex2hmjg9XmkmCmdrg2eEu2dvedpfjvSzcGz5lPfWocRR5mDvuG0RN6sjCOoPLYhH9THClFZ31jnC
9zyJ++w1nh6FzAYCSkaB27Ib7JfY+Fk/JzRDUk7HRKbNIL+rRgt0+FAOnrdDsiAKBPHpW2jc1LC5
qHOkZmglYl80uXoxQRaj59yMZVgaSoWuxwyZtLMUK2qPjMJ3YcOwXen/QkPcS8TY5YE/ObmZWoC0
x1fAMmgA0mbbzGz7FdrmpJ6l3lht8IrisOThEyP+P/H5GlE5F9Q82y1MQ1AFSwD8wsBYbtMP+abC
gD5ZLNIOEsfrhXNX20dV3sxwns7LcHb2BsosI7NzIZjTT0IzX9yl2It8RsGJCByzvk/GJ8ec0hxL
cxYLbIIBUdwWuREV5ehSsISO6uw0IcV4YQ4BbR4ZbhLyelcmfMWJcU01Aje/iAS/oybkCSWZEcSa
Khfq5YKRzd9FVzd9rVi9JYnH2MObcwwdsNoiX+11Vxdv7nN1UGwOLHSTDioU3s6tfYxYe+VlwTrE
cTmoYgghNUeGEXWiwO2oKtivQlbXiXFzY1/NyzH/9EaaaELhJXrk9fy3w4DIDnxtNkoicUIyR81O
rJRfOxkUD88V43Q4hYPd2YUEgNWkMcD4v/0dJw+g+d4B+bMPGk0DdU53SnSoiSu0vfOL52giyCI2
nLYXFZ8/jVf5tXeecVg2JuWOlXzWeox12bTU9ctV02zv2F1EJu2QPKozmBdSYkIwNqqa7HufYdx0
YIn0Tijzmk51xjc6fSwQrk0ODDNA8z/jURU56wtSAukzqErxCk2B+3llKFC4p8uAg122ZTaG+7T6
T6aOI/kY55Ua9yihG9Vncfjt7VIdjeyOVFlK9kUDu3/6kuWhCxPVxRRXh3UqLCJiqHYhIcexdFHc
YwKeXnywpuQ0/9omySC/Ww60gZyY5eufbUndC6jltwiOtLHsSCGulTRP+PsIXmR52EQAxlL0oh5L
6bDNNbSF4LoK83iBoLzKUZD2/3W0vNCpmTAe7AbLNvZujVU5EL0DYnCHSikUWPKIN+C5A70Ktwfh
K0bPU3u0kLRisZISp/I7jyxn9d1+3sEh9ppjUtAzPRjTzq1npXZaE8TRz8r9aRTu2l15OPmmHaqB
eU+k1gByMqzlE+7UhkqNIPK4ko+jUQkyoTlFzFz6d6XwS0Se0RvGxHsFTOj9jYSWVPXEjMHdH2QT
7eEq3zWwBSoEp0yA2b22+CY5Z3AOUMsj1lJB7PyfL9AvYqHW9U07tAJEXYq+w0h6OvZpvMWi36kt
3UhZR5OTlhpda9BlycFHRtFb673tjecbJaOYpDSiGq1BOaXp6AV8w2QhxwM1GltlAK1wg6NK/qWK
kWBhlQd/4YYjxVIClGsVEHIEC9UA+ufYRkd1Xx8WYvGk1RfyYCdkJ/mGKccw37UHNzYQV6PN7NEx
QiFfSArZua4l87ARWA51xKMBsxOdW1gxvS/+tR7XmRlYQUDuK1Sbj8sLGjUjbkdTEchDoYBx6VMF
zCu31Qyx+gVw0bR7gQ+zW6I0xO6xsXPCop/lFrtAFp7RSZUA3pdafDzMUsnjAQeMoTYeAWCnX1M7
+jA8lTSFE4Mxxu2Gm0Ltcn2krpe0AvjLWjVbGMPLT09adodlOOHzGl4jLamjx0SIcLki8lFowoP8
MY+qiDj20vno8h2rU+/qgtX7PwzW3mwUlgBaMPsuv0aocfMvknXmTvBG/UZgEGdUXV0TkH7BWzu0
S2hulFL4ttzR/qPS58Ku4TCn9r1r+1XA9Rn77Ym+fCO6sRsNW71TY2HWWoeZLBr9BiQei1s+ks/6
nFFZi/cerKBwQaLCMKUjLNS/2R6LdMv6HMOSP68+B5ZZSPy8CIRmRji6Ce58mwrMqvGL8LCJIOBT
YIEABU3Hga3r/pJ3RpkIHORshfTY9oB/V/3LWeB+IxUUpWNd+YOKlPHP433NsMVqRcJY1OB8ghaU
tcsSp7wLX+VwpnG1GUKfrzjpN4lAqGulxJe0mqc9GMDpXpbFC7V6Lj+HzVlwEAGCESJ5KhdVcKIr
OewaE6kJXcGr0tfpd0Ln4zUm511T7Gus/6TIct5bVYlxJdmMVffG7Yn5WjwFLUac9YQcTJB9+dSW
nN6AhWm1VTFqywGhxpr88OpW18OsYwCvwMLdxXYEU7NZSJGP30FbcrFa9oGe4UKzxAwJqnkXY7LE
GAgWH4Mv3Gq9nEbyxCeH8e5t+kMgSzf1YCu9bX96/ln5gzyUTf07V+LMSFVauSz7bqQsuTVbzGYw
IQ7C/9PmzI3ELebt72Y+uEWeEHTUPS0xeS+r+pMg9gDPAdxG8AP8IYrwyKOLXoXADR6XrORytU06
BOiiIndhl/gmBDavKOGPJpr/XjIpqPhhjUbwDZ2CEIpYbOFdOHGqbszFfn58I+X0WXnW/Uiw9CP+
8UihNrd2ot8ScOM1mJID8gYJCdHJSN82YplAA2BKoo3cELIu9z8BpxJcj9OnUQfGKUEm20wYZ8hu
ICbhCvFMSeWnMJs6CdjYw5vxFBlXBPwQfIcZyEBYqPmE57VFEiiVCbH/V0DQki7LhFruQj7dNksf
5plyj22pJM6Emzr+cTZQAd+KJBB6peW14v6X1lt/Yl/MmWRSdl8FNPB2x+G/z2rgIgQ/uPp0NhW+
R6yllFyQCRFsFCdz6u6iyUPrypV+cb/eBrapF1TpR9jdUiDYEBwjTbRkFFBDlaMgyq5HYeWuGhl7
joWzKJj/GeVo/i00H/puw+G8DR/XWE+ZOXG9Ad4TF85XwjTpXRwv0mCp3vF5MVMZfLFcoVhqxTu+
WN1soaKjhulM0nxkJEkj5Gs/09lRmpa2vuUPQ7UHtcwuflnvqJ7fkLLU2IubR2hgKGACYy9W/ZqY
tNq+q108+yTPBEADzSOLUzHvLKtDLtLlLBGB5jO9vg3lNCSwlHWibFgtj4velluId00ynPIljoAs
xftjuz89oLXp3HyzT4cHhpUqo/W+CfkTqN1ZMxK6Ao/cXrQjKpDTd8gfbf2sDY7GEuryclivmM0b
1qM9dXGGCH56CxtmRyJvDKzrjmoHXZJUkQ734/WKcqUFuSY3uqGntWuZD2+pO/Wy3SMuUwgcHl7U
XLqow/pg7x3TaJ5DP9t5qUklLHmevpw4swL+8znwcwlDN++a06t+t/hKVFv62aGAKfeZqtK4Gtpr
bmDXnmG5ykLmW6LJI2QwTbkz6ObCgMxLSOgW/Q+L/87OL/uV0UTcd911tD6/t/KKok6pffxB1/pj
z3FXAr9Za2jCJYaW+fUmk/WITRo5kp94a2fe+sSVX1j8RA8wAl/qUaP16+Mrvh0iWA/BAnVopGAl
CBJsdUohWacD2q4gVwi5t/9my+Xgu7aEZdPDC0A8gS0+Ee8koDNCXv3SnpwLQrXg9itxFcOdJPhr
9ez4+DDJjt/PQTaeujxj9g8BBRpaRslI2ZH/p4daH1sW6NyLn1Mx/3E+dmhkhva/OBWPW277cPEG
KTLlLq5w0Zz0kcvSILZHSVdhZXaHWVob22X2HmIz9fbGTcy363HLn8E5OtxlPQHyrRbOm2Subx8d
MZgYNpJmEJ2l3XXQD9ziySMEiAQBnM7XkupjbjL4v1/8pbpbisw1VxIGkJ3LoDooZcm8bLKYCKJ6
iVv64/8WlPfeQcUEYdryK57VWMbCJi8CwXD7y15gyUMZEhvIQkcpOZej5NQVhMlJmUZGMQFtrhN2
5VQcNyXvFgTux0vWPkIq8xiIhskXnbKcMN3S1K6CBH4opFDYFjsGmUWNIcNJR0yUs+Cl8Z/RFkMi
ZCS7ZDEBuK9FZy1Ee4nJvaEjzueQHdhtS0HwmZARsWbDP7OMkwmhKzxrpfd6R5F4vsiIyadsHsXC
8Sz30KJObBDOgN3bfYqngYmehx90fw17A+oYhwupn0f1mgGkalZY6VqYGflG+hhizAFevvZs+WtY
5IpjhESYLgg6AhS+jBjRUXloSamOYcrV1wZUAs05jDVLnV9Vf3FfZtND9MUSUWKB4Uq8yh/jne4l
WT3q6ksRik3b5cLK0k6igGksWr/kpExz5QoTjhGmGHu/zdeqCY70cNggSW9hOgoGs6qiKI08uwBo
IvGapFikhensk34hDIlsn+BEOvPR6j2uzJ3yBxgKCHjvyA8v89g5JjurKp66ulFHjTDCf7osTtQw
KyfTrIuhaRggVIxdjSJkAke1jCU9UsQBkaJfvUcLJqFsl4ObSNbLtSadNe9EVH4paLZzBcKIJHhz
LBYuhMiZIh5UZmo/ah4Dfd14yj54ydoU9jwuB4oMe26oUmr3AFaiAElMmCSQwU0vXdlh17qTr/dx
LsuSTK8OG+eqLI6OjQzG/G8Frgg3clCpQja00Qpb/Q2k3a61CHlQKDowXFmDm0/NjklNoVhguzIG
P+As5TrcgsHxr6sUuJCp9ZAiI5gP+wvNlNcGMd3VqDoTt1X4oq/8CO645Kvf9mwTNeThW5O49mjl
8VpRk6cPQMvBlfhyMd5B+eRj8KkrxPfytVcsN7/P6dbD5XpCE3/RP7Y/GAMV4sP3YR4nYiJoX+8y
sqYWsC9kUFoIg0X/NdnPYA/R7CxMxy8pCHOVqFzNl5Ve7lXJmXcAcLSHsmPtbNipC26/oJxt+x0K
DpeHsYZoFefuBxdUEp7gDh/RusflcDBLM/WT0vfo764DgSmEeCwNuPv5nkYOVp4SYPm4RlubDaxv
jZEIrzhLqN6jo8rgL8i2jBul51jaaJ9Pxrunf+QlTpu0GJV81QO9Mq3nit0zp10uV0ujn+VKEzeb
WGavzoeMvBo+LyuF37E+Gq3/6WjhwkPUGSRjApnJCgvczVHS8Id/KJ4PZhLK6tAuh9BWBQ4hC0NG
LUOVD4g/rJ0NHnQkdHPGTU5pj/HbA8EGy7grfuLUL/+bF1Q+S7tEVVrecGK0oCQTpvAj3TfMqUWF
qJSZVZWIJRr+ymLYQae9CykeeLw4+sXfyU8BjC66AmN45DqCwpbBmCR6sGH4Gs7GOsce0QTTTzQu
l99G1zau3yP06GaA2xXSY5ePG6qup+bmdTURprl7W174wr3z3kQdhI3t8ovY7KUqXZNjrtWNzMpX
67EhZKX63NopXUQyfTkQj3WIpLHYOcc1d9U1ws3IwVECSXmHU5pyEvtOY8RmrUMNds2me6RcRDRh
adJ6TmBtHfLAEorzKUjjhyNySoRIBfckXL7qBYD/9ghTVRwzi1S39u6h4uge1czepgqhngdUo6HO
4o5UR7IP7rIpJdUuH9uQWLlmblmCQRHhy8u1BEOG/Gaeyk4plAfEBohfveNY511gqBf2rD8ul+9i
ofKHrJMOBcHojJ0cmxazWL3UuO0Cy+KU+AMBeDOnzZ2i9AmPvGHj8nGKZXItueHS8qPnSLCfl9kd
XWLQXZOJC6udi7x7hKefAU/HUBPNgNMXlcuO/7PMhkJ7n4hq1KZqQGi14fJwpJVmyRqdxC48ZbHi
P2KYxSwpSkSnkCk4KpXXdfrqEbAZucjTF9pcAANkWgGXTuhMczoJaGEjB9gtFxbHlKOJnjyUXqzp
8nmLGkK2Fpqo9m5SIhQsfkWAIrQKIq9jtdmlW7rJ1lFiFJPFvu4hzyzx4FpQeKMNDBLlGJoSqWtc
QWmhSmn/byMg5uNejlbIy+F6jsT16Q/xubdoK2VuIY50bxM2CQ7ThGKtho/iYtPXU1Oz7VRvTx/0
SKnorVS6w1EmeJIbxtnVb0ib/k7k3RgbYOVmMQCd0eUUArpYNunOBr3mo0qbp0k0zM29pWtVCjqB
/sLWd3AyU0qARQrNE27HgRReUojwmqJb5nJPhMVR5Ffi+L+vljumSEjv4HKtj+E2IoI9SQPlxIa2
x2rdj/A2XkKtJ9d8RPRZxoO1Feyjr3RX3rpCVB2bnYzZFD7GeQ8239OwDiv0x7g4t7YUHW31F/IA
wkRny8g18Oc5OZGJaZfliFq88exWIZV9xeruFDp/97biYJPkhvSjKiXhdhs+4wTINwAT22zoveFY
86qO+HqOha5GdUI42SNaRWTEy59b6SHcCpr4Nhk2Sdc8N2FPFMjLMnwBB0h5CtUc+Bh/QRv+rl3p
T0zr14n/Fup94t+qgkTNAhhYX4OVkMU6IPcrIgC2ZjEIjtc89BZ4Mav52VTW6y6mYv77Y3K/tlNk
NEv7KRMZ6LCbrSWPcXxwdzLftMidvP8svc/RFrPhKzbmBE1oaMnpeB0Pm0hjDQGIb5X+ZcchZMNV
RglHAyQnjx1KiVshMhXRsqYkbEgH0bwIxur+bsQ5pPIu5LyzktTMFRnX+utb2klKazYMQEVEWG3B
tdWmTAtRsRmLMWXYRsnDNhmqVTSol8WxmZTs8UVirX5soJCf8jqzooJ/NmZ4W9EEcNCi5X4VDFr6
yEs4bmWgqqMvFNjCr3aGYjaRtxFUEk/Xbv90s6D1FI5ol2NQY1YYeTwUbLK3XuLhSWgDUHCLub7Y
czuNKKVUGoMBouSdBVnqNbKUoh1FCZu4U6iJQwF8rDPpNrzH/D0EHE7zIyrlK4tiaE48HWkE+H6S
dXMOjoXqSkQhol4IYaGzGK8nf0IfZpPLZ/LZGO5pdn8OnQUd/4OCoSyJV8FLqRIFmxhC1RBGrHqe
QKTDaVaalFEFo+f48JXjBR5TYKHMtGjVovcBU29Znqkb9R5MLLc5gkI/jxdVWmFJXFim23cUli9d
ZKA1MUdNMToNQ3er930j9HGsAW6RIYjshltYpSUaXzG9EpDANbHe0s71gGt8dx3J7KApmLmM0pY9
PKWIvCmIlDQy0tXq3BVlV1v/eBtY8YhIw6/3Ya/nKbfEgY8h+erFyUpP2WJPdt6NAR3vgoso9DBj
6sXu3DIYTUwr9ibadA+cHGI+8QFlX7H2RxOVqotzfW5z67DOHYg7m6iOLw21RnrcTBgARNed1tlA
dZfiAUDWQkN2O5/GRR485v8Tj1ZiNWMk+mLucl5oXswlm7rLe82eDEBopNaGYWlPvK7e5Jn3feep
IiYDHct53ywXQCerbvcXQl2ajTpQf+vVt7eGYSUnvRJmPS+yjSdTDLgYuXGYCRV8C1nZNIztq2XV
nD785P8CLe7Lvb1tGmRKXghNR/KhFCP1WA1J3tDU2hJ6+SJV5hkuBO7DAxE1LP58lOvBWU1w+Bhe
t8RoZInLlTyyVTdsBt46RYhJHrg+HMtwGFSJlhiaMTr9qKMccIFQjwMWITfqGYUITlEmezkYLUjd
4KVlfvkpJLZOpML9sgXz1AGNMa+WzWTX5y2xKEUNMgqzojBjrAinYgby27schvukOZ3ryiPt7tHZ
Lxy+qTyJfXny9bHFuBB+UYs4f5YBuqb9l4frpeYZ+q6q+fGAfDPCOXlMaitw53fJc+9Ai/fBxWKu
m95tYQTO6IjnnVg0l5Ht6+Py3LaKPKX0ceDvO0IUsUhzhni2dg5lajAUlwocMohInrosSQDk9QEk
6bsWgW+n5BY1qAuWEy7Qa+RBA70kQq10a4ITkuQ13DI6h6/YS3RJNEH0uZg/wBFlOMcEdz+QuuYk
OHCb0WqHamRpEazXlpZS/pDIKXOuMZu2KcPap2r9UEi0Yl+9uTdkeHRV9JpdIn8FqU7GUk8ph7QF
BJIqyTqVC1bzOnj9kstdcww1KYye7Ox53kNo3neKUZBSuqTLzFjLRZQIIgMzvWJS3ILwROCc4ITf
Vaa2XKIQrDfJ9fO6J7Yz84In8U3Z32AgEu7pJNhUoqetNtlj/oKEHjqFgC0lEyOZLF3SoB4WiOEa
IbjekeIpbvsXVsmV0E3mU4TvheDdB/tE+Q4Um1heCODLnoGr515TwPRBGBeRdiwjJe/DU+0PDt7G
Owls2LjAlmyvvDuBnlKn31VimATskLMYn6tKpB53GNTY6+Mnkx+qiIDE5A0BOLf47rCqpDL5vSHA
d3xvvGnW3Kedbb2QE9336v637Mdylx+sFLqCzMBQ4Dnpj6r5b91APaEyHGb62StKbCK/1RkN7mBM
XtmOcdWpC6h7CiqLxlAmQPDQgHsz6RdFx065thJodXPvGkwkAK2/Mv8uapQbv/dpqxMUqaw+snct
UFSGyhWDvEL8X1J08mnFg1LEkrdgZleZfZQ7Wb+kfJA62uFMd5QV+CCUhOaXtIvhpI+ZXzWz4wz9
nLjyEPCcjUbXwYr6nkEqh1osm2UBMluF44rexT3zTA5gUbTDPwrNeTK9r+DS3DDdtz6kzhnUaPCq
rFTcrHH1jhJ/qeK6sUbOhm1lJKB0G1qEfCCgUQdiR0TaVuTAS9zVvQG+Dcatg24dqthb2SorlmmI
VXPwK88tahfFPiBIkJakV4owV3bO3cJ85DyTsobaNyDqWFrjmUC15EJN1dUNWR67eXzzXY2O2hYy
obzIuG0d9bCMxW1CbtzeS2spXkiGA3HGgX8SYGq/NwOvk/1gtLqExsa17kptcm3YhqVtAyJok9dB
T+NAcrT78Kb4orhP2IaO69ugmRuyGF65CQGTcYEhU3JZGW91Zz8l0M+yyiWBPJpHHN2Ux9/fw1MY
CDRiDHYSB44HkQjlQIf0EfMza/lxFUSefn0RNXUSFod9+I5CS9ONDb322HDCcA/wCKG3H4uCIhDu
eG3SGRtnLNmkgOEU0USclNW0dg6wDaXS+zuX6Djv7gpthKiYEQwIzTfjfoG5wHwpsFrdzXqT1lgC
QFRR5PG5UY0xxgZEAlIzQ0hMRpIuJeKpHGnSZnUn/MG5Z/NYCYf/rT3o+4sMFkQAyFFtUp1cWk4P
LQu3Yt56iK7dFfiPOawOtyX9H+K+emO7UAYMEhr0s+I3M2Z5D2//KdMKUkHuydAGeL2SJTclvry+
e89lu1ZkpS2fqsE0MLcmMhw038b9OpXy4bk+7X55jBdSHETJAyXr6jij2ZPo1qFcVFs3YlbbvQtz
kQgU6oWTR/KIZvgdHCXE1ef4qxpTImUv2sQInElxl+PnBteYprGYBcMe7vxZJybSobq61g6ZmC+6
wFBaCWyzUmZoB7XqCjloqfnQ8fnzIGthkitvruEEqvwekF/ri6/bLkVVUNxVWXfp7Sat1Yradsyq
RNtgraor9n8Q6IaMlpnyaeNZSrlUZEATP/wzvuS3psLRdAiPDS0Uu4NIhJCqts40Ntp3XVW4zzoD
QTQW0y5Ib8gM/cDnRAOdf6BE2xoOfRrKqJCRCQLeFRqoCK/OOlPLs5u2ToUE/sfrmCjlRNR0Abk5
NBFuseoTDBsDfr00cAsop4Ml4gOK2S9NAyJk1Y25PlD4rTyoWqBCyzpVVRwpRj30fFA0Biojph99
M05Wb80kizgTNKME3Y5vEPlYQuvA+FEYQdUaXZ7nExu4rIEHxrGaX5w2ODB2PCWjJk7OT7ZX/KWg
geca6YhMdOAQx6F6X092PCrTiFLJFiKv+FhRJgYKZRIx68Wz4skBWqNzXaWMbKSNjq9Q0hL1CgLz
0FiEn2eqUv0+eNbhNGow/yP7iQnlZvAR/jIw51O/bvGQkslNeCnafpDUxXDOclT48ODowzeLKM7H
wwPrTC7nRZl5nWFAzH+IeMNsiHuDZ2+WtYbPrGDbKwiOugykCE2/UXpCbIqmhBNM+Sd8ZmJ8o2VL
25rmlHv6DMF0OIIRAMXvCLSXGd3qDGqLAA5zr5vagPMsKq8Z48P1f9SDDRHE1MzLImfANztqkwrj
6eAZNsk5Z/4oYUH5rCZsBLOodPNQnlz0Mxkrdv2TO6WpgjRulMwh/q//lNB371d3Xf6X6ReqtxdH
8cm5yQ54NWqMHXbN7kcFqoWLX9Zce7ewmeFLVGzilg9NlekC6pQthvP73q1KjbFEKuMgEw1vQEDd
4yTD26LtHEdqupNZdEVuTSLWD3pfszLsmrnCZxrqAtibYDHvnWa+uFaXvA4UjeywKeO9oQ809lCB
Cw5uwTWU5CqFSgKUo4Vl3hjFPfq3ISw3EL0VqEZvdzEa1ThxKKTATtLGvdg5fnAf3vWWqdpu03ru
QR3CJnNKRgGBBW8g+uaq6sHsoc12j/Jaor/hzfrw/8Pb8TsNyul3uQ/B7CqvleZTs4ziCyMQk0XO
Yi5xkRMYnJ/nHyZqfwM1mQZHYnxlaCHOR4rkwpykGktznkluNInYQEMqciE1rBKyBIImbMXa+Clp
L/Pporxi0l16GNpYlrXP1YFMeetD88g3i+/A5MXDeBViJ+Uts8W7q3v7CvcdbAWDYhCj5u2mL5YW
ihaIGmg/0ctdUD3Eh8a/OZB9Gqt/7uHiEnj5JWFovc12Glnqzu8MUeYV3pD9ZWQcRGc9B71M47jK
jlHd9rDjQkKWMH6Eg3tozNTz1LB2WiDAHLwpvQb6KlW2cQv3bvCIsYyYb4crAcGnpfiixA3vIUlI
JhADq5ZuzCL+p2eY6qFeoRlFTOUgmnQXzb42wxs2VXjH/xJINKKj/Cqe85DqC1CE39mwclktqu1f
TjUm3aGqfENGn37PR0NVzaaW5z35ehEVj8q9FdMOPLRyuOk52Ktb7AExFIHpR4AHPEBCTrlJAIuU
L11mhonOXlRdaQQBX6u7EohDmzh7scgyyc6HFPUg2qIR/afOhk3bTEa0aF3hmMu059Y3d7G40Npp
LB+TbGPuFVFCbRt70XlHM5kU0ILhBktwEgXWbRPsctT+jWWUISvuBdhSdlPZjSh9u7UnbtiBvKOg
6e1M6/wBYLwaIMoeJeTr5UqgX9mR4tu5UEwtJFJNfI2RftfQBC/Df0CIeskxBAkqMWxV4kU0tVka
8Wgp3ytwYmHuVyj6iykYvs/x0I9yGrTJlg8/X+5j6FRvk7D8Z3U85Vmla1XNchukHrwAiEe6mpDe
SoKRVnbUiJLpxOSkmRiBFXGF4mYcUlksKL1mACyseiEj3D9yaxhfEKQZjU9OVEJoQnQOK7Y3UP6y
1noqdPZcvsBkSBCMmFDxNDl1eenw+5szE3SnUqgtm3AfgVGpfVQsE4DQDqcnOW83WRtxsCSL6rCY
X6D9dxQElxm1Jgsof77tn9G9Wtcyfjp7D1AvjlUgavIHYB7BplyKkso0Zij35kuQ5Tg1tJmkvNJV
XMp/AAzoClDSJ76P/Tri+WQwHof/m78k1t4B3xZ1nx0MBaS8rSdZbRwuVbW/jx5zpWm06x7HIBoJ
aNKb8qKqQvAtS8ekgP16xyS66T8Cf6p3pbw9HtfQkUIm3rmKo3EZSSSwOQUel5aJLLmXV4UuIUXl
tP6wKoCqIWV3RHf3rR56twAlguKTL5obssfiwYewcVVC7gdcpFBS3PQ1C693lAqtX5+H/la5JIzN
kcwweLAe7AEU0U7gnGmHdZSjm2z05kAJqhSPJ2Ll8BPgLkieF8gHRBnmpdTKwgugXvBKlBneUvYZ
qyll9+GyAe9YYM34F/a1rOLskbA2K49rTWnA4t1XAzJ9im9WWx6NgY/anbXgIUeWvWzddJmKauBC
zS9KphisPn8OfivMrVQbOA6UhFZVKYWyVKO3k3i/gG9mchHdSS4BGEqIh7ShceDtWLDMU8bHW2to
Le5lC8v+nF+EqF6zSsIpn2pjzgXJmVwyUzueSOfe3if0jf/6Fqm0TK67o1ZrUnH1kFJWY2sEzUhB
GAFrW7T+i9A0tnMFxUKE9vCCVO7Iq/2IYS4iZNonN9YWYHVzLWEQQa1zJGi5LFZSIHPrUFFuyYB8
v6C53JB8FqX8Fm4WBh+kL2k8csMNObcos8HjvuKsuCHVNOK957nDpSIqTtqUcpVaFd1FyoEHx5f2
AnLB0tjjopR64mETg/ayQmyXHFstXtWKxNJ8hVNRGWwoSnJcs+Rm+ogKnigdqAoDkNjWio0FYhim
+JIKGSnho5isvEBFFUGmYvhCoB7Z9lLnXn6zTbaxUJQMYmAk4Ez3INA/0HnvFnqSEtht66JvJfRX
Lhp+Gve2+sFU/YB/zFwa+ZIVQgrvBCGiXUKIGpOJNVNnEJk/qPQqsJVFnRTX6OXx3glo95ppG8YS
KkBU8EO3kVtA7lJ31zsgXI2DFINBAakpflYtqYptkrn0cwxTEFwppO2OyV8phY6BaCHBl+kLkXFq
Tv05YTayKx0ASlR25IMFiH+v5e3ezAE3iTVZyD9vZJIVSBfM5TTFo0LtWY1t/mhg+oVOmFpOgFc1
GjsDeCqn3lFv2kzLka+07Z/Q8pDsoYD9beiONJApKJ9Ko6ElaFdAm0EnwtVsfpTe/xgbgYeqo3O5
2tX3OJZLBbuv+fbdwtxi0Vfv+Pb4ZEUfsPhfZan+F0+DA0dZ9GA+1E6yQfxCITb+OU1MlIHVpDqd
86Bq9fO+vE6mrZLQxlLaeTKrA/EWXgtGCL16uhQ3z8BhvVfFQM45KG3K5xVXz4DQLm2oAFCXj5MP
eLfFWveiwBdazNZJZZah6dSRneAqGuhgeLZG60I/NV5juOW/swKb9+s03PtRs2hLUeTbYpkQ6kyo
NJc9G4GxUUzWC2oqhJBRBEuETUogQPIaYaWLgX1jFA+mCKVdxjKG2RZi4QmU93K15ADoeKo7qNKT
RP6OegjzRQ0YbA3Jp8mrj3jBhI5ChTH0Um4gGbTeNBPBMtsF8a7s20p8ipOsL2NN62zVAaOCY2vc
rNwL7EGWQM18oSdBYDhxG6d813/9IA7Od3yd2tr4o9TsZ5OFfcfi7gn+qqMas6nea19lLXyzMHiv
w/2/Ig5uW1Vy3TuPe5AtC3CNQeoFJA+EKHZ5LvzMLbBC4k741Z/+CtFTSHh0g8og7A1sLhRED5Li
TWanecC8Xw2sej1Y4AsFO/5p7qmKSC2k145avUtRshY8HkbXm7UUjPcXT1HQ9yJnK1jWF+wjeQOK
u1geX23Xt1M/DL7y5Sq9rIFSfhHqFIIaNC5wBmIRkGubDcNZS8xlacEn/HMRR2VobCyvM8YVpcsq
jXWATlcA+XDvDE1AFgS/cKGMPt6gPjLfp0a1xOgagei1wSegbbk5I6MD0HNV8MUOTA8MRp4kY5j9
D23jSK84QB0ywGH8zdpaKICP796QzvQ+PgT4DpiTc3jSZPFRI3E6Mfck10z7ZXV4XaKA5tK87XzF
s1SIEo7WOQmVl3LpNkXxMRTSvYP6h3mGy/lfVK0JOQdJJx30dtb6fWHPsNQQxQnS/L7EFpI2E9FT
qdrlBRSBp0FhwoHVpPb4YEElAa+UNRS5bAmm3ihK6Tx7RjZN7yYrThSP1OEKMmY03TF/rfFEr6mC
ZoD+wOMAvMPo3RJPvhFAPwaWDdrFExfXifjSZ4Vppu16kvTk2eYDijHYw4D/cq7h4tDu5HvLnpx4
GhQ33Mc41ZQdvMRgI4UGBVH2I1w0boqUGjLDUp8huBeXhxOMTgUUqjukHo1rXrLMrbYEUlCV1tJL
RGGfb9mbMpF5b0aI1CwDE+haDDPrYUiqDs/8Ev05/z6uin1ebGmf21LNZNXkjO1fuHWEqDyVlJw/
YcDSgvPtrkzDnE1Dse76RBs7sdvE+qcAYvQvkZtCtreRzN+tqX5z4h+2inprhNq/BmQiAgWtKZRo
U7cwodIewq07fYMTM+oXr9z8r3RYIiEa6kxv5mnIFhRJ5jjDzJxJgDiWyE0BmS+YvQXYiWI9+seK
mVd2UpwEB9/PCbt9dF26p+42KPG7wdrViWC/panUZBZnlqyR4Z6vW8iOGg9QL0ZeaVWhDArOzEsI
A/oFT8TJ+fhFVjpEvHwrl1HcaswRsiI7+2RBKOAGcCdnrkUaoRYxu+aQwR54+7qDof9NOzqiGbrf
jZF1P8IHNAhcv4dRtYK9U/oEXVHBXwL3E83Dkiq8syySeFUANiHJV3iPEKaYgJZq432twjZaxet0
KZwKZscM91/VXreYC3ObPrqN4l20C3rlKIasIq2FO/bWgx7vknMyczxkqYgz4GiXGm3EJGx9FrVB
b84+IyTn2SMGd4yc2PJgPaigRV192XzoPbPNs+UzXKQD4zwCWmt/5GjnD2IO7S2HccHQ1UV/3H6V
kgh7wPenLQMoWPeZQODeTvfxni7WT961TMU/JUMolxO4pADKX7tLLX8FON4bceOs+o4E/3a63qsa
jK3Qc9ugaIeqFmCVm/I1FlwqAuJ4AIvWI6ZDJ7Gp6AhrgNHm3OkfTrkc23X68xJ4aM6qmZ0Bva9O
OP3/CddFqBB4oEnOHBax09crpm/On8/TB7WGus+4SWB2j34nb57H4IlW87AOf8COqHc9uJWYb2BF
S++UpzZzTucm+PsyL8/KQt1z8rIEo2BKgSrg9+GBEFz+rEnFQr1otDFNAnofZGZQ1wvvQmUrxU/9
u5yEtg3d/bwYpZTAZoH2nh11eX8K9cBOlt7kUOjTgXKNGZas1stVUdaNTKbvp8kyhXc0CHoo+AKy
xgoLCl6YvffHgRaZfhPg+ezZnFbfzAUCXcYsvynOjJvv+hrM6kxmEa04cTdPZdA67WXuiL7RAxtZ
9f/TpbRfgHatnnjJeMFjTim8u6f3JYwSbERSg242SccQqbHDQ6gyBej7HkYPnY5YodCuFY4OnDFj
VPpWlxB5OeOVugeTudJSEJhnXQ6o3DRG/KXJui9vJAt4s73gPw7muiaGywTIFwkEthYn4WExCi+m
QtNfhvZHzfsKCuPi72XnQg4XCGKrgWve03udk+I6Yl9Tp4NKuvsYcVfEZPwH0+0rmrN8Qcz6ekc5
q0FdqaM0iT6PicrZiy1j1kvrRT8n/LNnn9sp6s0a8W8CUjTxQ/0v0MGXSIdv8XjMD5N2WGi9m+Zt
/0IZLoL71HWGzY630V89LpcYOsJK+iDwpl9B308HUC3gLDOTfJa6VfAryhsuQ4shVzXKqaMfCwC1
uQqwH6VJEKEdk/umnH9PNGK0fuSFqLbmYjRHONqMjIGgJ3qViWMy5fing0eZVxcIGJ1iRoRjuHYU
o75HtNTP49JcbbYbtSAmmvnHvsscM0AUZk+XAuV6s+XVgW3mMU9wppdXg6K3aL0Z829XLtFzS62N
Ki9zVQV6NdmC+1lTVPmqlbJ/5ICKK5b4AR10CKOiq8GmBp1zCqc/OxXdUtgLG5W3YESDPirtygaG
lOrSdyhVwPj+4IJUj8irGPbJsAvq9Dpmk8JvTw1o7BHQJMrYkQ5WD8z8yB7qeI+cXICiRUs8vZsk
/rDalLfHqHRK01Fe4hQV+z4pIMqEyXo8NCMY7t89uGp2cTnjjik8xKA8gKVJH3Wt58hIIdxqf1ve
Kd/vyRQVGv+hvk9peFxUvM0vgWIXyjzHYBg/0xpr0OLqwvILCG851u53TVeXEI7d0W2Dw50fovZb
b7On2Xi37OGTuTbHGFxVb3RnV2gXuGqW1GxIDgjvjU7qmc3dnfXmAFQpuLpYQRkwM+CoAKq/SAXi
zRwIXCWD8Y32k2iXbZIZXKsFldAb5ApJPomuhDFK4OnIEjghrKNctqkWC8Z0o1yXZblVK0SkkvJg
Vru0orHxOPCMiA8uXuDprr5sRk3Snx434Fgm3mrZmtcbPqqha2EMvsRg35i5zALaIA1oMzsWay6X
CyJqDLnQqbD7xHhEfM2fTh8IhG/i5dZ8VZr7J+hqkMkPxK5KHUybXuA2u+zbUaPno1nUACcN2L2+
J3T/4Zm653BR8NVLuREgHD3eB+vk2vBf4eXpZfcispG/mUWHHkbp1pOmJPUxzxv/jNV2jJqaAKYT
C/EHNvXBSmOvjqpf036AOvBBhng/w34TTHA+YreqFmDOnq7pOnXqkAby4bEQyU+GUoyTKdBUe6+R
RIdoDDqtryivV1IFy+/OQldb0psJOhnMmZWQ/7VBzBlLg1jXD6FIbjGwMHRHBfGjkDBmRaS+oFt5
p/IcPBIpMqe1OT5THIugZGafuD5U2/CqtpT+B3gQaoH/VbItkWh/UdrSPgIuhEl87ucpq3lTp0XW
5JH5jcbRlVQCuaPvWU3EFpZApEk9nHK6aawKQEGTvrvJqawgdWdpdf+gnWXHGlE5HH93yD8GZPK/
rw1La39p1Dya8dl9O/NH/EWCxRFZNBGZTqU0FZdjJWfjrghh/iG4v5fipvl8M/hTW2iOsoHBcdVz
Y4VfxxcdnMg66MOgEEQarOyLfoz8OO+Z4KC9fAFC0wSQmcCFWP3XX3MvAyeDTv64MHbBSfP/GUpV
xOOnxjL6v/2yrBgQc6ydehZ7gFXSZhcHtSCuSviy9vNG08irsgQy24G9U8wRy4pmPRk4+4SwmKqa
Dm9FujOGqSGNnhJfFm0PIkmu5WZ4BVDTOW9T3eIz+QPvWPn1d8xNw0CO2KgY1mlhnVrLCx2zjItf
t+4g0+T3PbWZduv09YsKj/B0HjSuAitR29D5G6LTCK74p56VecxEdGckf4Brod8y5ADcUvQC/21B
EhuxYFVNLAOSxuZTtDIi8921q35y9b7eEfRHTxkVW7XazoUty5KK4/VxD/Ww6dh3maoCfJs5fj3r
vuxCuDjZvYG0Nk9hAQPewR5YOJ7VEh10ZnWpTSonzfo/Bnp6hxak/uXPNfrIqvVDNwwXjOVqb2Mr
+IE1FBKJuNqrdTYTL6jkh3iHpZtrvbR67pFjXqei6HUnMS92YtYjnYjxq+7AEdNTy1LA1arw9QGZ
QvL6tcA8RBqDobBUpcfX3NczOL9320SqvPveMrgVuZyX0on04ASyv02H7rBVa+eNjD/RpPOQtnvQ
0YUgRclFkvb2rK83NsJ2XoP5xKmyN5n0wLZx60ajq+MbzfNNeL7p5EV3GgGl15/xWOcBzz3nfWGK
JX3bjGJxJoJhmFi/qIgBnEPT/U/lRo1UIh1Nh+BSmK8bde3WLqhTjQxSlFFeodB88q+Iqh/5ygsX
eb+Dwl1vvzYs97br3UpgkC6edk9c1dGJZ5ktpjoyQmZhT+9JQyPH3HxVgbVXnsYpbaCK0jJrCP/Y
3Lhf1mrDuadWXhTzZlPVO5sqNImbGAL4n32Ka2qe924h+XwA3Ptdi+2gaQbQPpCZi5eEzI1h496/
2vAnQi55PS4RTEqSEcoQf5RtkW1XuvevXz3F11GlkBtdVCy1fhI8obmgrQ1OIJ8SPwRQGsOc4B+r
VcbY6ptBAEDzdUNaDZZkCW1G2Y1zwhuM49A7axaY1IRwZh0qSovO0M44yE449vKJyC4C9/ec/Ct1
2lF+YqiFWXLQdXtL9RpLqBE6bK1FlJo9y1FNw0JKG6RwkMNjfUjLzCu4n1+whc6swJYCDK4GaJsV
W6CciPsdMxpKZbmW+3KslGOfBlZgNU1XVS9CYoy4OgtdZeGilBudFk41p5nP5SzEABgNGIoUojpo
WN/DZzP+hBTM3I9QB9uYhcZuNUOtuZ3PziN125k1BiR6xRPvZ7HJW6V1nIQwxepBq1A0GGB9JSoI
uuO+n+/LQ2RLEbN3Sq4mk9hK6tMcdBye+gYUYrv7L35fY/Vkkyt06FPmRboIqLhTUtPgpfVwA1Pw
K+yA/CRElxo5WJBBtvUygihyiC5MuVLWi5nLhIDHNk/5M0Bcvu41ICigWIXU9fg5+/cGLHIp6WSO
Zd9Y/i05d5gqYwY1wIGr6K6j50/p/t1yIcmUlhYLwWzmAziz4Rn4oK4wuXygCJ1z1qpfiaQG8Auc
lfW9wCp65YnRSlxNsssQToVhHZNRmVG1aWcJimQre0KbIg1cRuJ3r3AakTyfRGWaHu+0xGAMEnQZ
DpBLQbBxBnEz/CORHVjDe91O5nSqwdLS+q1nzCt48pWJSxcSmZxHndLGYM+LOLNTUlBkcZP3UIaa
7gb78H438LiPpN53DwJWLxklTNuwdQedvVBV+Kz93ewQh1UyIsuQmnzwyVNVeWNmS0AV717V/Z9x
nOMVuIvbLIH02t2PVnFdJybcuJF8Anyh7ij6uDCZflCp7/1FYBtxzP1UIy+OYuK9R6jFJHZBnI3g
Ue9T7XMxh3NIvL66uCGR2V/CqtcgHGKBIX1QgYHXTIgfmNDrv6Vifie2Io3W4hS55CTv/iFlOIQf
yrrdp+Eq+SV0yTdHetGtF0zzYCsWPZRHlm5EbAyLJnTKzXaK8o1uD3QWypS3GF9g6JaRDojqWchP
uSzUxFZcHtFDQ7yTavlthLOO5/Ppj/JdkZJ7XVSyaDewMCKS6U4PVDRfvIRy0kFUoda31wSiyD0q
E1G1X9pdh5MEIsdaNQemSWUKcxwDdwky+SkGqGO66cjzridWKRptYVRev2hEk63pD2k4rgUccHBk
0C0XbhpQct1Ydpsby+Dn23oj9E/unC76PD+9lO9BygXSMCEzTsKLmrJL3Wcd4wpUHBGjlrQGwrKo
uYmhP6uQS6Gq+QQl2Ac0xrhQrwVOsZV/WTJbwCqTr8J2XMIJJGWmUAnjT3LVbfH4aiMMwDN1b8kK
L8M3m51ZK1zn2kZKGoKvHQT03Lu2m/3/HAuuIMuoBgpiZkQFeJAVs+xNf1SY14NKf3n/dpFBcIUq
RRMi+tZpg9d1G6iy2/9Fb9Ykk+Vgw6BP/TUFeDloNMMv8fC5t7QPkXEU6C33pWe1D6zeUiBrdJ8K
6H4Ij3ykquRZ79FDafNqQVMSUBrrcWoTvuwd9gVlxVZz2mUOyY3skS3sBBxqQmIjGRaQU6jxRqlN
V7MO47o9PX3a1jgoEKbwEgXYkET+MlQFsFyJUAuB9AX1Cq7wjc+2S3UGg3bRM41DqdrOlUM+nzhB
gLtljx4gXaDxunue2NMMLz/yqsU5DqcV7FxDg2/YWckYAOkV07nU5BOZBLyXTuCw3aDpjanRyta7
w1l+H2pHcXVorHGu+5xwI/Vx8iHxf2uAyWiCemUi+Ayf31kousprLNJDQNaXx//gM/MTBCz0dLp4
aFzWrrkCxJT1ZeObCru8u9JF9/VzQZs26AdqZBWSM4tvTtHDEP6XU06cQHjyi/wOb4OP3jwQxuOh
148uMW+VmErwN8KyzZKQ/lUONoJMw4r67LTu5fMsvbfZVDJ3o93J1RAqW61OXHuZOrMmBIXWLunf
XHQT0zmDeufKSs+p2MgTTfOc/qICEFsS2o+df4iLwWnyobuX4jQfFLuJlAWUSCTg+cu535DAm7q7
4CgCzk/xwZX5ihL0vFk1zqIHgA2eR6DbDrkiPKg2S1fIYR4z3OFeppKBJJ7T6Xcm32MROuVUcFzn
y9QOACV09gILDrIcEK+UmlD5FKYjiQ2D2lXikluNrlzTp9KEKiSaGn7AxlmPD1mskYM6wuVSgS5l
h6MFiLPIx8kEcOiq+0YrIjlEgEufRSP/wPvAf0OdsBlSEvhwijVOizp0YzM5xjrAsE+gBz7HEvZu
TYRbmj4R8ijwPuQhS5+JiAaKYHOPWUqkANk7eiTqARNrwyrIAjYRC5O6KmNBCSbl0Iu0P63XwJUb
Lu0d/RACLRopRFWXoGYrAEu/pNuEWYTxeRIa6Nb0Hl3798yo2knYZF4w3nRt/C5Ekk9cciX+TdZK
E0Hf4D0Z90Oqa8EZxRv9wKaBrhudYQKeJdropejUbH8X4fNTF1er5eQNOWwNh5znbJmJ/03Bwocp
oamGG//Rukbyma3KdHLry89CK7/NOJFciwBj5oCxQHDVc+7NjwqBgJdKkAIKYIe5nK7g/9TA/cs8
b7ua42X/1K72KrGXRPWYPYN1dtiX3Su/KjRNJXedYY/FyGK74zueP/kOnY8Jyv/4D4U6+UtMUdX4
iGnacVgh6ewnDFRmpbW9WORHJCYZZ+8/WZDR12y9eSmb2q5hJilf8A+RZ/CBX+tq1vzySNxw9JYf
iNSt3cgTiaZgtwidzcdxNsenkWeSTnko317+alI8lIuz/FgkE7tN9vaUkhzHsxsl75pSuIy/vKFs
ueiIfkeT7gnKlc0tYAdU0JqE+kI+E7Bm0rGxkJKbhCz5jkBopTLOIYHGpHxWMbGQBj6Ky4eNZdpN
8+8f6m5BrT8zj38EIFr26Wx+4vKty3s2Y2sc0v7VwWM5C3U1E0bqIUuAU3JO74guOyLgCnsXSzOz
0syi4D1p+MSJzXcyPO9Kvx0kp5Au9IwqLHpB/zKSWvY08Ad+N2a8IupaLg4l18I5dKlk4k0AuSU8
XiSlHdhN0xR2+6akWr21DyGlBJL3U/0ZcCJpLv7/1ghslBowEKzfMZFrrYmv4huWb0SornrsFzz2
OO7E4DVzCBK6/2IzcvJRzcwBYlJrsVm4bb7G8TzNttD8ZXXm89VI+Mo970KxUB9df9F8DPg5cVBd
SjEs6vxKJuP3MmkcFxmG6EV1WTYZ53AB1phrqbw0ZqVKKh4GmOvulo9QVUVSF3Ns+pSjMFLKKiog
Iw9Zs+8JwZeicnJrZ9y+aXqK5CYzCvy3DubPY429faSVecRhXeeGA5st7Sq5cO3gpAOEzv1jNXnW
O+0EOsxzzJZEIPkRihWt3VpAns9vW6UELXvAx/DXouFz+qZchu6n4sUrAzMXGtOv3hhZ0TQzegI3
ttAk1kWqYFJSo8RjnvKez++8yJJFrkc4iqkRUqdYSRnlqyr0e1tMQ3sXhnzUhOSqMc//DCQCvKBt
uU3MasnNi8BvmRHlQ+eTWM/tnGVGerNpDlbaUJ84vj7C00yzNAMch1DJJSzusWRgr0jkp36QLkzx
ELZL0kbtZTVpvBkeFIhDPc5iiLhpSyAd9zb+lRPHnY1fD1392MZhggj4ePdUgHP1mDYtO7fi2k2T
H+UKRuo5HWBWy466C5vVc7Z31U9sbUEDYnpxIpIZh1M69BSsku6mIRzRPh6QmKl1hDcdcMqv04Gn
L4agvqkv/eXkN0rh0TtTl7yx9SOQF/Lxmgc80gIxstScoFcUdWG6ETTviGPB2wAqXtOzL/7pcZRV
qFBijlDV2e/tv4Y7yx7WJJSHBlOn6iubHDo57yzVaHyZ9RsmgY+4b1UwJ/7hPHfhmgsXH6sSP9uF
7UHI2DIp2LDfbzYzuvAC/fcXo25g4KqWJ7sqh2bNzjM0yBtDsBPymsJI58T2PoUqC3fT1pEqWRFr
si0cK9DQHONR4IzcR/ODO6iXRLI8H5M4aZqlaI1//ItgrutJk5eb/K4X088MU7zCPI8F7o8FkzyR
Fje9SDuERZbM16/FcuMMGi1F/vdt5L4NtADvQCvK9GvEMxqbyCuuqRPg/FrDCJxOhNKSpPdLmrvj
oTuM+9GxYCAfHKUY/fehq5/sGs4TCoJk2NuGHeBoCuZnL5dS8eazrTidlTSZZygQxFr6xWEw2Qg9
c8gFs7/ihcnEm9jWAWdKa4Xs6k9rm5k/w1kjx4LgCrCVgBCQSH2S+EIXrAFPJ95KAoj9BxCMZ+Ob
DqKnTMsF3qrCd0+cUv5A8UyF+hqQDxxvYmxM7niwqecdYOy3XHDG0gBzd0WFSKKg1XeWtjTbTnSB
1rzdFjjyJtPUd0V2kUaSxvEnNLberMAY8FclMGPHHPaIn0GDY6+j8ret/nack9uedrsM4bbDPTBc
BiCQm09TJYURZqw1KygSiPQ/oIJi6nAMdURghbrI6FCtx4FU/ajwQk4VKk7VtMMPTE14XTCS2qhf
8pIgptE5vikqzblbfNT56eis0aRRqZ9S5Si+RbtTsUg4tm10vBChacm5hoUjij4SLvi2mbhRPI16
UcopArsRtSK9dhGpzlrVWlMkFdUc9GiZdklfw10Ug5EghEWw7tsKFWML0Fn6eAbFeWH9Ivkk4HID
WxClCnuelXdI6QWiV+dhl1WTm9LCpaq5J8zh9vZ3aPjDJ1bHqH3QbRgC3eWyJDBX/jkHtrtB6AkB
cRzX/ctcfeWOoKEZw4AW1azc7MBvlowzu8PWiekP3/q8CVPK+orvQRVV8Tuwzbv+QM8a2q6Xb9K7
qqbAL6BV6SLQZax02ULaDwvd3HITjIvptJSBrSatYYGS1OeExaEydZ/ahrAakxsik8CEjYCZvmyO
q5Z5GB/0BBUOTUb6pR0FC1KmKZH2mv5tMJtkfJfvFqf0AoRbAPcnLC6JEfnmqctrj3oPK/+zffcT
Z6f41R49slfz0Eguc3a6DO84hLssLx+koKd02z0/mAhRP5anpUAuFZTI0MhFlb2QsgpoHdOVENOo
bHNzxXFdK+mwAKUk3f57h/zSDJvuyrvYwsLDRdpUMYJj2gT6mP5catikfycpVjgH8jKf1bCzoGTv
qMiujypj9ci3/XoBKJd8iCM46q3I1J1CShg30okhPQ8lI0SJS6yTg2Sp/rlD9YfSDP81S0kxjTqr
C0ekUbMbWjeiB08sfTi2Cx1kRMRDoP9ooAZoLs1ZIBe/s5sHG/xsXxxHMyH7KME00gSx+TCjgJrh
5QT+nQT+cJIdkf84etmbrOy4fIJsKAq4K7P3T8wmZkP7L5Pdhxs/RwzxP7gsOZeCw60ShFy6oUvs
zXWRfLA8jznVCbtGEtQj+f4Yaae6rcZrHLJPd6FVWdpxDS3ymBWExU02C99Q8DCU6ZDWGrc7SVki
vMq9rDTrm6RwSwG7SbPa+oeG/Idr6PIwjlCDKowYArA94PKb4kmvl8fygKFHBEBQFIV4oG9BD1sJ
ztU0E3FCBJl/KPnVujBvbz60S8GVD1N8Ib4K8vCivkFYhqx3jDYJb+UwK1vpinfG8UCfQnG72XXc
y96eJcp9LYjwOf5JcqdGuK/jvvt6dWUuW3WT35a0e/NS4BOXa0btQF+ys08FlTcqcZ7djJwEBUs5
Ul4OpLfONkjIIZBLaQZzjuLgPrVPsfaHQLVSoLyXbPI8pdZAGJatHlqak09UmjzFTKTPIqSS+FQR
zGo9Dtn1rVoMyKPWHfoegwiUhcfa+1DLxAHHCcmRsYJoFK2aN3n8yaiiDbF0IS+ZeyfwtAd1cfn6
+xiEKd4xiRti0bnlP8OR5VnKltUCWRxQBWcz3EDnvyVhAgbdRw/hasmUqiX/d9NjqALzeD1dvDZZ
JKOTv/MmCxPnX6v5bA6e1sOGNucbTs9yTcnnWcUm8xWIWpVYkpPkci4dgMjYoP45IBumc35XsnaC
TzjfXEDagjrdpmxP4on5iEOzrU9r+Sk/htJ7NuorAePN+gp279Ry5q00m522d1dIHuvp4xX+VbO/
W9hq9Ij+1bIcfvh6xO9s0lJO3af35riCQKEuka0qAYxLLQjDh/+QN8dXjMypdCfEKCWl8zjpQ54t
hTzIv4X5S7YEWKWV8shfa0zLLFl0FBUCIB3bdcbcbC648dg2cmj0RdE178fsqiSblXKcNEX2sq4i
Tzot7eRIX0Sc6Hk5kVj0U7ggQ6k50vhY2KTGV838P9ePkVGGZ0ckctqgrp1tvkIvb6EIFVHXzMc2
81a8nJwycG7KZcUuF4VwCaQKqqlLu9uRcc4kG0KSEoN2Gg1OEhmrTXshROxqe33ezi3NtIrhGESZ
AyAorNcbgvnq3s3Saf/r8mINvvus8cPY4ET28Ju3iXLn1MOHSmI1/9JseccX8y2C4JkHcZrKA/br
IXDipUsqWmtWbBBcikRPd3ohjt7HLO86Dio5hUe5lvWZCVxw0hHk2dm+44b7EBwIw4aexsqlBndj
ATkvd5/lEz4w24VXzEMuwFUafwQDFGWoMIlI6HgSrKdbIwBYjOlxRf4d+B7z4JKgDL/pIF8wTpOB
jF3xjn8rx/ENVheQ097/N0FRG/dSJZefuPqLyeSDq6MV/ZqdM15eeQvBiQgvevJ7G0PGeqaHT6ms
fua0mn58Wjc3oFRaNfGfcdPKq2EyhENNE/ONedMp4UkcZwlEEJN5Pm8hVsA17tzCE3XfIMRitS8P
gr2YR/fNt4+k+DDge3Rt6I3+l55hUakN3wM9y4tKp62uWScT/XmgrtU/+/b33vpglioH9uZUGy/S
fykCiFMC7ioaK5jhHYVJB2RnCqNDJG/GlXMJTdC4nMx7XWX3Fz8+wCExlNnHRY9xUzOh5USRU8AY
z9xSTy7zj7SJXm23eVNCP7fWvDPEvJyIYZx/5/ChZRHNIMsEf5uzgtiVDWN12F95Y778ngichudp
IMRQywwZsaK3xWtn/T9r+bdajIypR3Pkj6DFWGZCqGNzdpXa6wIMVEUeH43d8CxOQFay9HcWzR5S
vbcWZh4F33MdOT59JQ+Jpl/Aus8Vo3eqIoEjhGlrwu8qOHiFyLS/i2HEI39jbE0sG3KUAg8B3nCy
lRpWG7cqrCzjBDLXVeOMxaAEBXktCW2zQuw5WZoDZD1Qr8uXORpyMA6Q6DSRn9LIFvJwpuRahFJh
pBy3l3gV4PR8fHOT+piSvHsRmBgldDnw30UkRjypOGxLb2UTBqD1FkxccMvfzZaUdJtqO77aWosH
cviBN+5XPdzo8ZCX8O7QDRLH8l3jFOCd8hBTGI4LQlrNNrE+tD2EmKNv5MsnfdW+x1kbx21CFLA8
3UMD7TLQbovw1gNGclsaJ25w5ovzyDWBSKj7Y5izjLaJvT1jBgjE3Qral0qOKAtVfxTAvNNrgG6p
luZUzqrB7PufyF60lvGBvdWJEYypxNrHdAbMRRs9Y3R1di3+8IFqqr8Q7eL9HERhETnEvmY/14+o
ssLRTwFrpAwuG0DTVBI/3N+IsqABVzeuQfi2pDW3RhLDBJgvMGxE5oFaLfBJx+2C/z5Tqj3CdFA6
zxgOYkyVAP68uz8w652M7YtUemVpuLYlalC9QZQQs9yQdniUZnM2haPSPIdpq9zMat7J0Z6UkQN+
dqYnVej66ekgclcDTbGmM1OVZ4GdpOHPo/0OY79ySVo3R1h0rTpxkqcRzClpoKDa4V5FV13vTf80
j6b0M161KjCCZsmUqid9J6F0AOv/HxpcTlZcSXY+6hQYwRSictVZUcBxjboa+MbPaABDbXaRPwkv
jd4Lhv5d7+oGkHrOYxK7ULNTCVPebAbyZErbMFY9xsJAVNtcrbTW4mPit9jgmdBTAxqMWR40BazU
Yq7/LNu65I/lwxqyYuU72dxf6LJiJdhPYcGylTtHPT9j8rKkWY282TV63MA6Uckr/x+cFfMQHJ96
bjgvyKOw0Jdp1Iv0HqL1w9Zds2NdZ5GZ2MA44wffNJS0qv024mN6J4BHM2qY2DCOGg2EhHh0XeyU
lJe2lbS3WtIXGhJvEatU79UiRINM+nKKLRGtFNFWSpoWDIJllNP2JiyC4TzfN6dCgn36RrhC0sCA
oPAvEOLXXDqodh25euiKZkczu8yX9LWglcR+Tj0bSz/K+vbrqibJ1V7hzd9VSAYib8lfSsjubkgH
+XCiXvE1NlDsKPZiJr/8z3h068zD2AlAt9Fsta5XVwnFwDcBxqr6t3bffg2Iq5/ZFRYBh88ypPWz
L4KNMoSUkhXOZo70W7Q8W9xenuchswAvWPcwY9BsNzLBDMXgKtcZN+2MuuxA/jXvOGwI2E2X/pyQ
FLvQT9aPIoC2yqHaP/oFFowU0PGTKRmjmh7RXFl9IRqQgrrGhX7Ifglc5zECk+iJ7KlTk8y8c1np
g1RJ/sBe+bNAiCeSRWJPBt3Lho2VwPnuvi/LHjTuk4JKDeEheJ+S1rl2SebKQtmhYUO8sozf4SrZ
pxfvKRnm50hbVxTQYtygaNQoWDt9sq4IZK8rNHys3/oH7gfquBYex+mQOzRX8mYEzf+f8Jri2A1h
NS02NleRvUtL/CLRxsyZ2Vp5XP+dOdhbMCVkAzZSoeiFbhGZssI1Tpjt2jrfSIQnlN3sLUIH+O2e
Uqu1LaXuzYcmYWpR7kcXOpkyFDDRSRebsXowTQ7Ysw6uZziEMxznaA9a3N/k06JN1Kc4ojQSvF9R
tu1fG/TgNJ5US+MTDPpe7t3/ez2MyO9FMyV5csmneXeJ07PYI32TKwAUq4f3VG/e+TdzkDrvFX8W
QMtUWN4ge89EtFMUNgP9LmuDRcfnYNVjjv4qnQVuC0c13K7XcXmqxfAugf1FTiDmUHIRxSZurDsY
y3jFWHERXiyMJSgD6EGx1oAE3dIhGjPN7LNkRyjQCVGd9zKse3xJwWGtAmyldPmEDg5txrhSMODv
83Nm81NO54JHX/ipsAbKObxKcVE6GnkySqRJSX7ET6Dt3yRNoEmBLa9PYqpPs7XOfgxmiUHyzj37
DbcufGKYnG92FD3UQ9bjleGm48DNP84m/r3s0WSicUN1+zAr+R+mhLJXMdRtRmwGWOkWSeSqM58O
CNssM2CGsg9e/Kux8EzuLYK5f+U8ViRH4eaeg2NRM0R3HYFmbVSHik2ARZiZP44Dejgo/0s8FJid
3icW+Sb1sAk13RVMZO+kivOFQruL9mW+ZTW3CYVyPCALRjU1CnChjlRxCui5UsNPKUQ7WM2XNzbE
FJJSCI/TNRfxHYY2Vm9w9dGEaMyIdPOVoSa4I7fgnixJe+Q+5YOQqnw3V1BFVZdQUyq9amz5I1oz
mSOANuTPKhmQIXRtEknpp9mZIY9dC3KZ4dQfJTkc58TepEsc5kczJehkTnJgGyQ/tHXUl/z/X+gr
paJ8KkZIZWtTDnqX9O9QdqWHvuloD5OU8yK3HZm2sib4lGcN/riCGkfRHrow6Q99hlISWoYh10Dc
VMhQ96y4RnIyg+P3MpXo2x/HZxfc4aEh6XBQ2Iijn8St6FNYsrHRTcnMdqOR9ZoIVhF2FMdC8TNk
bXiRyFOPeU0E22o4d6fP/CN/qbsuwPMNtY/oY4F90OiPtcD8z+CcuGpIWrjz/sMGtc3AR1qZnznq
eoJ6vznARWtc1vhisTxg74ePRf8osQ8iZcsTYPlzRS1z1Cz2jVNOgcIQ/Rx2DKzFV9k0p3c1pjAl
O/ciqUx8u9FDD1G3jGOv4APaZ2aVvG3Wo0XRonLCmwEKjvn5h3S7sc8ciwTE7LZ2/Ag4WPM86hvp
UvpM0F5S5vtN+iUTExy8VTktmWka/0TOHdTXDmzV2cwJ5vH22sWL9joS/RpR6piBdWg53FONijZp
fqBM34u9iWMdIQux+Tys4iVPq3mp6ACSngIsxGlGg81HRRqh3TCa7YxHt5db+IzrN8oSKx377qKe
2Y6L9HwUjT79yMtouHa13UyKispc3eOg37PFkLEQ8L8xenHm9Vr8yI4LV3R79/MT13kuwvnWKRYC
VkmWY94l0wBKJmyKQJoE5/YYyLCmwLn37eWIBQTIjXHyz6TUrw8e5i3HYNBrjhr87s8wmbCjvMZs
hYs52f/24uMFA5VQSDL8kwkNBy138Lp2JEef/tEN9h2uYtJUqvfOZvN5ZCmQtvDixz+xFLu28PUN
rW/2NLUaRC6vFrvAXfoUclNtMrDRqwESR0Xc49LbAUmbrvLp8VjeqofOaLm1b42TcqwdW0sOm45+
sUSaDy+cfJpmTPPXfqAVFcIvt3BeYt6JFGRD+DH2H9WyYU1UocXwquHWGVveBVpMgzx3HcvS1+i3
BNtjzj+ym0e2Bj0imtII11em1mplVpxqDx4SIdBCpUsV/tGcqyj46LFoLYWL4QogyB7cyYkjoojK
ezTr2Sju+wzGc7kQqyTLmZgfMYZxyBsky3dRslIV4mz9HwUqvx1TV2gfHN5WkljGvB+2AuV4pT6p
G0E4UVZJBOAk1K1KnvkwqHNw2ICGeXrmKo+m8/UQyt2rTtxH4w+qbym1ghkclaa60GoOyQjtwkRY
Dffhcsnhv9bWu2B9p5jL2pUK7I/gkqensWWMDIndZtR835rbUA3iBsggu4pi3ZLCJy5P8fs6vaxo
kVePQox+q3KAS2HQEZnoUIMXYco3iu4Sw+MU15DRCAk6/8SYMtJ8yspIdD604dvosWHPIcTtWt7T
rniv3QHP751ofXgs55EMy0D0tYJYkOMNcvYh5gUlijpp5GZBUGUef6znr1O5jgHNUUW5WPdMfo4p
30Y54F2f/IjWbuCrSkwbAGFlX71Aui53K+Jein9o3GoRMpZ50UZ1vyx2+OJqB0IDsXkv4bX1tSXX
Tj+4duoURyNB/OQ8MP9hCacZ1no97OHTL0wRMuE63Bxf/9CEZA42phEUEA6+F/smgtyzDADoJCPf
oFPakWjgfXZ+8MshVCIAUnP183hP6/Lnk939YuBh2jWPcG5RGAaAyYKY76mn7rMZWoO3/z/rjbaB
ZentDOOdzm9ptHtn+xuziSYhxoRfB/mV44iwCxdOZunT3IWQyfKy0iWze7FbWTn9THSgvFqXC5qw
qvgbkJlOEFuWgnhkd325b3ESRHtyeRlTpn5yQS5goQz8F+EA8bbqJ+m0r1AlpEeqTagnk84gMqFo
3XZG5iJKbBLBleUd8m+40H3a3t25IdzmLZpd6WR1NQ1NuMPJJTbMn0gEw+lEAB7HzZ3WGJqHPf64
aaC2Y3dcMuMhFYFRCxSbOrBxkyrxh3OjkhEAEeAvUsxtE4uJd9E8R4UhHVgS+5tnmZbvz9+YZXFa
Ii0tEbxh9TDe5ErOiIYVBWg9ovutJCcA1hzdN7tkRY0JzT9uRX+GhJConRN2O7xn+uOJP70h05hA
o/VgAbyjKWmTc9dFXkt+Zaudf0dmDSTqadjqOOKzNLtXG8/Oa+tmg/1IRlJ131HuEB3SBu4ffhYM
xJlvZx5J8ZKP8IQU55k0m8iIUOyjtNiZNKKCTNhA2P2F/YTVzcLyvyWKkn6ykSKJ9w6EWniJtgkf
GpTFC6bbUggxT+IXe55Biq1ik9mrurS/in48BpjhCIaPehXlifwcGlhn7SsVIj6QLSb9Jom3u6FL
LPu28oDYXcY+Ln5lCprPe16X5V9XnH+5w59uZA33JaVF8gm7xlmRLYokxOxIQyWpHt0Td77ag7q6
eSdricnvanm94hPG4mNgEppmwYz4cvToWzmsR9IPqqj+p+DEc8AcVxkCnx0mNLh7ziEAqfI201Hp
k+qRgdcXdDhC11DAWpZXQSdno+w0Sg86XpvQDHv3wRb6FKLU/0TZcBErdFgUlrgsMv5UaszcCK9i
sZZqP0/c4Nr3+yoGlvZxaxNmaEMidJYJXB2Qi8OYqtbiMRE1CTN7Kt2wqituAZzaEEtRIKUhFsvd
hbaK9WeDAFoGjQuwASjO/OmFHwHCmIbli3eqIdPi9MWoAqBp8XJF6k3vjU76Wf0i5DU3zxizoHXK
xOqCdUjrbjzWH9rmspvSPGzmpeegtl5g1eMcQ5TOXjMmeC7ZksSPFYyq6CaPFYYRZsd0Eot64rG/
z7a9PfPvoNcuLnjYDb2H2yXpLgzPiKiJYocr0R+kC2Lx8sBxXTobiM+qU8bqmI/aAX28Up2Yg99d
vSKug1zDw5RSwGfMAiMiF/HmF0A3h8ildY9kvhhd6Fikq0MhcqTHp7I5187P6dAJngD4IdyKk4tp
laBts7ba+BythTMkLaf2GUjgQG6vcD5vp7K3nnu27GW83fgBtbxtBv9/lkaRU+1KNdDt2JOUrAjE
ezbvfEQWGCPujP74pqrpDLlGcKhAYoy1s5USfSCPpUAOL8wyL7LLwlmKLAxqVl3qZaBVpYWs3sU5
Ldvd1vXRkZvIHc479MG18Vtej6NKGVMlabaGuSXHIGpGOgX4MJ1fOnRWFY5uNkHKA8FnLiqWGyaE
ezsA+R0UY8GXt5c0WmBAgVkMPqlevvMgTqV8mKR+gxoN41qvMsJguG2ar/h04LeQpHlUwr01nV7W
yI22dht43i3x2DuGFZlm5ykJSSHUL/Cr9SAVoadUGcCHb/7FIkf1E+6wFJcajSAM8lyfc01ZZpSu
walIYlBpuT/wCIJ3JCMqLMUBv4rAsBXyCbRU8HAINtA+EFQq3hl426PdSczaNgSYHGZA063y6HDs
aaT4QZs9L1pdXKGf3ayL0jaOxF95tHTt9dr+Nj/xy2Xam0k2UqirY/LB05Rp5v7A5VdU5ZwoB36s
/klcihMSu1wPrAVE/jAqFM/02tYVwojdrhXT1J/GXNXUyjCmxYlwAuTDmlsNNxOI7e/z0Qirp3on
8YXPcC9IpuszeYvFaKrEtivT/GRVM6aQBzh/N8ZRDjD6b2/vethLwZnjx3wKUyzlZPH/+Wt6YIKO
3viF7JPMEUjbV3q+drrhjuB7rFtKQqno21EOk6wTOca6VmxA+HOD3EDmjWRVwYs+/97wdXbt5JfR
awJrxAKF20jcKZu6/HC8zLzOATuU48fGRjL85j4fjqtQEECi52XFpPM0641wfX4fZJcCd+hb2p3k
+JQNAtGH6czEwxoCaZqTL4h2BjccdoJ/9mKy39EJQ9rZHgeMjqWodgbZSuhtj3bdDXo8VWqUlm4t
3qfPJ4LYkCIiz1icDiuGX8n5zTtXH/P7yS/miA5qHyJnz6ucocCcuYQrbPZP+fMaNDYcHAjFSgCs
ggk7+0SuH68cwDKeC1azdmNscrg1MP5DXIGZ0BjyLBIk5d3QnSG4z7k0NIc3WUQhHCym8MjnbdDC
RhagvBgJJbKKeBwCCZoapfUEDkgVm+Sv3+Q94U0iTerJ7zwpdIC8cmQMjSHZrebhrDRGcV+xYuXD
a9wfu2cjaXw//0+Tbyo7TIMVOuI08BR69f44T1WaZo/zV8mdtjW1nGASxPVEYMOh6YTcLNM93DgC
82VS4DQXERx8iqEB8Z5sZxIlN/2Xg/hFn4j8ge9IHcfyAs6a0BlIIVqqqWjand5ja5AUa7TeLrng
0KG3zOGxWB2Me8uPxIkSuOY0fWy8zFSmGnaBdKvIEczVJ7o8xPFG3eltOaTboNDGLq6aCAa1IUeo
19m7OX0qNtj+/8j/AxaJ7Uww8PziNCLlSSyZB+Rw5cJ5FF3+t/lBwdf4jNyZvOKB5hd9HX9CwRIo
FN6z3ImroqeDXw6p4vb6L2/8hD6YCanIrxcsfCUp/dry2WI9iYwX+pCdh/AVagot2GUtk/fVZK/H
+koizUx1XgMD2epL5jJjYA7jbjqxx30xyGJYFtJNK7ddFFRpMrbCcKRsebrhqVfyNwksputvAoB+
Hz1gBSp/j7HuwxJ+Bz+idTrmhQNXuFx5s9lyrC8OGwVo8Ce8Hz7Q/7JXZ1kxD+mJoKUlQuGBBMV8
yq+cT1/4woiYwcqwanEvs9NNm/bASiV7QaJu5pSzH4LUcogGjykZSmqcpjkGR2t+q6spgkJitXZo
z+WgewpRFv1CndX84UKq8DTFyvsV/4LtaiR4NRoT39gPKZO1lwRt7lJIaxKEEscdF4yrA93zFUbd
TMw8Xa2B3B/DlPkUXoJ9YEAKl9rOmNRdOegNXHTWSah/AwoFY7FGROBDxPITBeiXCcr0AIWNrGDE
b2t8QvTS2C45LdHoq9MZJp03WoKjCNYZmdN1UDaxr67LenU4PlmAnY+mLioJEJ/lcHas47t+BaK2
YZNO+o7h+y/uNfQu75H78P26tWS/MilGy6dxT9hZUUXZ/Rf/JAWEnhb3Jr3GMazNPnPPUP9w8u83
GXXH/PZ9790mZ3shdImfRAZQE1OV9DRN9/qj5afh2oy5Fw0XG8ZaGC5vPMqB+a6c8DIt3a7YG1Xs
+NB4iV98z5+o8ZGVYmfjGn66L/jqU6pb4VcKqqhNsD8pJJGkDpqsgmbKLiI3PskcwCuLA3Ts0yuy
SufACYQoSaagKxMc8RFPfVg9pJL2ic6zZLct8B3p2ZpzzVI/Xo+LfKqk5nMQ9gvYxtb3x4mQdvB4
pzHf/8Q4dqMb2KOGspXLBPK336d6m1fQwcqcmz+efw4nNtopcKnXAUTb4FoKg1grqr1O8SdEL4FG
0l3+8I9q4ENl7GjJ9qZ2EcIBCzQcwU2IYxQL0RE9CWlRTK671LUSpnp9v8u2JSijmBeuJ085vRT1
4VqzI2UU8x+ofAdFQmzkwS1DCJ9YdPVYZwU52+elZBNTdHcc5oNunzC0ubm0jTGheHtDt8ire3QH
nrKRd4RrbLMF763xheG/M8F/UDRKGT6fYDMFr7Uwa9E/4KcmTH8AL2HwcZnt0/HBxhGr3kxCbLz/
Fgy9kCqVqEPVWpzR/2kjfvwl2D9v0+kpSrRPqpFa+CtqTiirrTqFnDVHxKEEu7ezCJZGTcly3pcE
zKm0uQckjQPjj7K/i+nWI1DGgPvL00b5mIv8TJEkR7HCgCtmk0ay0/tsJg9zfuXW3quP5zaOubJ6
81fsChrSh4Wgwg+HFaEeYIxHUKEDBFU9tDlYAn5thYAuuVk/3q5CnIGhHR59owgk1RWAJ4yzhrum
25xrfKcCUwPAdrF0scEA0ZUPuUOKIoTBW3eBGLyeFbHSHDpZZuLrtUsSKZn2RYRw2oTFeXjzHsOz
nN3PvoRMI+QLepD/fl/id8AZVOGZQ+wxSSF/XczogysGrTwfEp5LNFcuskFhJ5xMhcAejuqUBdC8
vwj0lcGe/xI4OYflp2SKDEq8AFvZ7il5xHqe6W5B1B3X/LHKyHCQRlv8rqwfzWJW/JE/J5vgFIub
wh9ohGnE+DZL5hsbqoph3aqo0FHZNffeVvtxeNS/bYeRgih6tjcWkd8EqQSJSkvT1oWugb/2wKEA
cs0W8ZobrgFGC5M17LTC8/LWP2S8SgMNatzk3WGU7R7sUNprJTcLHdEFH4vQv3kC8d5nZJGbnZG8
axPD2DTMip7y22V05wN1uZQrFXCBPqAtZTopeTGUUu/PmxLk1JfICa/JLO1lzk0CGIZl3BWapiKr
weU18qBiWEiaCWD8YA5HP8wbnIO2na7bHvEY0uNaRbfgE4s1pjFiK6GB0QBwyJb9ck9nIhSOI5pB
rEuuaY/5dbzY4ELepeBvgx937DlK9qmRJZqlq8C4IFc7n4C43onL2/nbtkW1IWXdV3bM298jm+0s
XzSfyw3zo4ZD+e16mP+5y2ekIX9lFbzsqE8nUXjf9Iy183fXOqLBVr2Ej+HwTS4e1Uk6syOloQQr
swpZvp5p9eRFxdIpBVgecOmQ3o8/PW1OD107KN0SYIif65CGKx3MOVBTCLmwqYLs2ShYj9v55k8U
p/sEYCTWnoH0WBKlZI9ngHZhg88RC3BrHukYp9QSVfJZDJ7bI8HzCE0YCpyWXbYcjd5XEAkF5ffe
O8o4cs1s2TfJxpwFyiZgZRiW/wLCZHITRmzEE8+A8BCzUcnohPZt7AQvsu4CuVKY7CpfogBs93M4
FZ2L7rQxYdClMDBYzvIN8u0Qs8VG/J6wdkPhHDmQENUb0rwS6mw+IoNZ1bJLHoIU5sUp0jIDzho1
s0P6fTgYFIAktWi+x2VBazmhBPCieFl5DUqkl0IpOfTtcKIybwmID+NrXmOwcqdyCjox1zzfE9RH
qUfHcJ/ILE9ol/nTDOa8oe/aEJO/jE/kXUMlWlRi+Bq5BvwJHyX+KHrWt/vEa6juJmPZm2aY9VjY
6JoysJ+B6f4SMiXszUejveIef0yKGqprB4oWxB1w+8IXl+w4BnekLQ+CQ3PqYeQyep8kXAGohOJj
XiJBOq1HLfnKsEI61G+rjYmEKmZX3Ld+/w6q0T0KPXnct79t3J/M4knNLtMQ/XO0ROCIGzPoHkSk
XtF5X7k8KQ6lc28CWBVXXB0ZqIspibUJ0WDhPKAhTZ3tmkiTNNpMmJ1nPNcBSLlJCSmvXbXWeiZf
22u++3l1nQTGa8iernwtd8pIxnDn439IUEMpQnDG4qObn3cPAJwGgY2UjYkHItwFr4zGEQSKHdSG
CGReh0OHdul6FeCQifxne+WU0mbJLfo/2bKxHzvJce7lKmZXqTMfQhO9JPoCKyDzf75rQ9QP/1rX
0x6iMXna0uvXukzrAmkCGsu48yUPN1gUg19w623WRRnwGSka9lRoYTJAYn9Sfg5VANh7rE+OBGmf
+ASmRa2PDx7o05ZEzwUYzRGjMG1vKcWbTKP2J9rAvcDR3ThbmBwjemPqj3Ni1zR2mbKODuQdRr3G
ICLEj0JwoRluP9LA9dHXdKyIYfyqXzye687aamyDTAWD9xT6Cv9nwTX5CgWUKa+o0c9ppn331Onx
wuVlveY/547FZcnJlsNMyofMbwQR8jc8BPmqr8YKRS5jDuEY+zIWwEiIXWYQpQAyJ8GWdLO3IKle
QDHgKj70aaaXxtt0JlKOxDeEE84HhO4GylW6BVVTuoxNXQj5co9YKYyuWb3Jk8jAhC6YMOWWCpvx
CxM8c9vQebH6g4H/vWPBCNgQfSRErKafO+FGyJ55LdokZobT5ZRkacgI8CgrqCDRIxm+0glx0dMs
H325XWuVZP1ZZj+3p5Q3WvULWUGJ9unCjLA24ZV9fcl161KAKcGB682YxPXmVxGEU32xzLht3q0D
HsAb2Dm/YuONcymVsZ5lO52JvacwonAQ3tjQJgSLfdlLMhDK49hcjPiOywjl6oPW0O9EXtDrEbaS
2tx/HrcbE3tgVLIQkibp4tUFMCV5/uUlYWxEVCNZDxZfBrBXTgQ+DQ9iIb/GJdQkBAEhX914F2M0
mAv4KOyXvu5MJ7v8dcxyQ84mIfZYZewsxx9OSf6jSRgqNAvKu61/wPmYW0RtVSNyBSkHMtWcM+Fh
Yy8cYGOFBh2QE5kNPWU6Kgo+1GWwMCtVVpuddfbE6l0tOFHHiPkfRas0rpnqmVUGjfdv0w4tRkUU
3x0RvhKDn0XyyY6br63LB2bK0Hp+adSsV+KmEKaxyh/I/uNOocavfz7e0U6lzKpm+T23EwTveDnM
pT0r3vWIQIB7Nrq1d94NfUVt0boImdQqigOlKJBAChUn8R/CEOn2+IJmhUR4GncIMRVJrOQQaO0p
eqMM+2pFGwDO9BkJRZWCk5wSP9V/UCWttsNVMn72tnYZcAFKWPuL7sjNS2VYgiiHkNUBHZHtuRuA
XfS+nKFwmDsRh2CIfgXiV+MnLLdvwfcBa89aRzKTczUShDL9tt4vkon9S8yzwLIoELciPcr9DeY2
xfDwSRZjhuu3iVJCnNofx5Rr6t31Issss1ii+tzMWLp5ZdrS1urEripq0UgKm78wve9tY8KMWdNx
QBWBve+DF6oDGAkjNy3wuH+KKrlTIojgEyobeLRpQfmtoaHEKs1/OkA8ohRijJtKag6UeLcPwDqU
yvQDegd3VsiZmTexHVZkWFy89YEqWyqFvEaBnjhGLnAlRsFOk2TLEPAWJ0BoeBBaQI2KWgZkEuTC
4Uh9T9azlVjg0gW/JPGq8Qf/AhZWDe47wGQxbmh6dsLFxuuLhmTUoRumIgGqjzqgIUdF08+Lvql7
WatilSAMMzc5INqeIPcSoMBYgIx2Bm8fbBm6Ny9gseESE5Rwb35bjL7CtaFBKYSxBpGkvKNbOzMq
z0kEqqUApWf9AjGW9jTdlClvpU1SU2r8OSNPKBOg7o3CNWJvpJ1uvnZU2wi5+2pCTf9emTmeoWEC
1F0n+NEfjzVYrGzlnxCwh2DqNGVvPudDz9lqm+FJX2tGKnrGMB8xUELXBeDDhydUdHvQBek0OBb/
hPRVHCw1Zh6wTv4NRneZncxO5AxpQHaw97VAZHk9U7CVPqMst8S/YEBGb3pbQU1kygM27JVo8KYo
VE7DEPvrsKksk52jW1FHsHqPEVvevnaU1qYHggrehT0AtMNhAee45nnwnEu/Mfj+XjiEPsAXcH69
sN4bq76353v/EtXjnEttztLoOLOC2lh9MEMGzKznq+i8JjVIWAw8QXLS5dtJiLhCRMfbtqz2XigE
/HYa732dWxGsvVvmBmN7zQOs00Rviy3xU0kmwiE/4X2SbZF59Mfwh0gCa2eMuM8ClO9TSJlacSZI
UVUv8bN6KXsOGoL9Tr94CEW46PIA3i9dp1+IwP7XqYDkm7Tm183U0zAVOXWpbtq3ucS42r0AD8Pk
aerlWV30idRDfz9yD1DCyql3pSRwPzyeZ4pp/1LHPn6lsvl5Lf1+gXVBMwI0psLwe6A+9dS/rvMB
/D3CWdXQQXQuk7UuPdOiL6scOsJpM0UmzDiEElUWE/Yv9Hf17MDgNp4ccRUB8pb6zbi3cGgaLvT9
ySbSRKlLK6Gkmb1xRWUI4svF2VBHwnIUvQ4qxOgiiVgLBqG0ikPP08KPsY6Iu6Bk6VMRdSTpRBT7
KNTDvWe/EINeG9HSLaBWF5Z6vCHFPjG5EAvbjxbFjY3nRPMe/XQ/i095FdrW9VxnZ6bp67LN/G0k
a0Xi9tynR7wJpFjUeFp5+MskFoNirg9WObJf3kEukMHI05rQkcSi2VsRzUutMvD4Ic10sCvPrPo/
SWYVNQi/pi65m18dZjVJnnHFP7oWJ7G5z0CPTP+/1SlwGZx0jAbSrT8m9baQ5kT0MrskZRBa/rLl
gAYU3iOUEPIOEW4UHZ3L+98YNml+OITfAm5qkqVkNZuR5Yzcm00J9bbc+baKvhWzTfnNB9zKEB3e
4lBU4+z6sNPbYWdhj0P+qRvLrqMT4W1t7P/tIq+W91mfUSHGiO5SCvWpiebPr2u9wsepJmPf4K+n
CsfF4K8rY+9DDImhOjs8BPRj5CQkQgfbSGLAyjRO3u1H4TaGqjFftzkX9rBtuk0+kbwAM1X1WVnQ
rXk78E8ddHOl9Uimw/b0EhW6M9UUf/GPM7eGCH7I38IQkXnRB/0gUcVdmV7NYkDuqvdguQYN9C3o
1cwfTpQN22VTFKCLsdFbEdWwWXvfUUjxHjME/cC/yA+IuWRMxx7MmHN93g4AnC96jpct08uiLMQY
3psXmXemnoHpx5Ris+6QqyKaTxZmmnF19YycGN1x7OFtzL5rvZj8tjgbiN4VqJRNB+XJkL9JzGTB
KtV0eUniq/kw2iUItMruYcXLsV7sJXof9Lv/XoaklIKWD/vIceEpiRYWfFE4MRQD4tITkxzvcOoi
XmKLzSb3pKV5IY7EHzrFsybYsRB4+CDBvgg22mf2YanbfOKN8l+zn2JzV+mI1kJfevmhuuygBXFO
Pr93//YokQK4rj2C67d1pQyh3oK+eSUFYGZZAU+kuX6LlbIXxMkR3XLdKWSPhsVgBfeJAPRhWh3V
K+Cng/P0qqB/DDQjDJ2AegFDhqpzXIDfj+SYYZo3/CJT9GuQYCakOoatw+QbMPVz1k0nt4BeZVCf
24qqAugVg+AAIOHodlBw/yTlIxH4OeixkOiX/RnH8cV/eLIDfvLJSZwA9GvNUW8JMWh0sF+tdgxv
IRS+T4CgFUhSmfZroDLvK+M5f7DpR4Rlf/YeqJqDzCZF2Q7G4ztVLxPii0ZM5KkW2U5Z955z0k1r
D/l9PQFxN5F24kx/YHhBaL2qFiGm2u5t2LNBaKyyOQS/7MnYQ7Y6MvtfYoRuwhBS07MulSakCloE
59n/1Opopsa9UHkS2ndfvlX8qSkXQxonncm34FiSu6s/nvoUvJB1EUC4nnZo5fTj215sCt3eJFRB
gsvBFENTh90stVxQvOubnTM/rF56A9heQJMSgS6Yef8ra9bmcVm6W08XuG9PkBLXSnLwC7xjBwHD
ICpERzueEnTVeoGkXraz1PE/mMNyYnWNOUs5w9t9YmOLPaNruu7yMrqoa8YYivthrqyNyYFSKovD
giecRmOzVeEPJYwDX0/ob2PShKpyMyS7v2UB/a/o/h4n9woVsb4jE5DHozO7zKYQjsg6OB77rfO5
VfOGXAaIwOe/digKI9KYmPld7SIZS79dMcl/BtF8rzm/spnRs+Uc4jG+xDnL42bNQ9tl3zOvsrP6
5AbnMCadLlRFS1h5QTb+W8HQy+CZaSLf5uETOHfwQE3CzO8Hp68Fk9D1PfW0mJ9g7440NmIOGc9l
cXWGV1H01FwyOdEAiZFIOpT/5K10q/7LW6wlrNgP5fMKXdy09If8XR0PRoUsYzB8hTSZYekJYda2
sUVUp9Yvp5npnUWh1FiV4cPDNAamkY+o9u1ueQVCpWgvHHdK09ZoH3r607rxn+ebSOy5mcLyyH8C
rUukhdJRzNP0QvymsAQbMqhsVBrJZKNtvCmEKG+xA0W2/gjoiZE+m3VY4VTENtvX3NASWZ4N2HVU
1T4GC2IS/pV5hVkMffanT3CN/ZwXjDSkfm5GGQ/lGuGUKVkMT2bzzTOMH5hykv8ETmibVtxtu4kv
MK6N3tfGdQWZSsjIflyyP5MRijgrW/ZPmICYmIQAvtMal49YA38wn147cz4q0LrHi9HdCUMuF9Sm
GDAZ1Afm0QwJ+DtbusmNSmOFbGaOUNt724saV6KCLUER2zIOH/GxAc1/a0gAMXkDXXndxlUz79St
zKoYokuS6btvwp7CTtfGZBbC9qjVP1b6+fIqJHgpYd8bkpx8x0VuXKDS6zxY8DP5IbqlWBSNgam0
V/OAH5aY9qrO/xDosoBLACTorhohI2Am4PQN6ju/I9IBneM7nGfFUGrWi5c6Hh66r0PC5H6OkBpW
b/TMLvY7qnC8ZPYjMLp58pqLMRSGXAojFM843NVq7Gbu7w6eAJNC5FMbTfJ1M5uPr/30Px34N/41
EJjw6yyOYLC9p3WiLNSp0XXq4Ou+LTfUNhp04MbDYd0/6pX0KFxhxdM3ELBVWvOtiJ/i+4+/cEUw
WT4A8JEofBkBf03XHPw7yrhRdzab7EBJ3sbEnKE7Bw16q2DOMv8H2Ugfl1X1Qqn6Zs54eD0U3BC0
zhZfwrE1SU3q47BJFN5PQg5LIsQjqcLk7l8xqBXtru31ZJJjGQFAqEGB9CUPXfd0jH7YE9Q/N1C5
HmpEn2WiamInIJ78ej5KACsXigBXazhXzQmk9JbHzr1k29F/UuAibf+nhNEuE97L22lzDX5GZkHF
+emDzzk95tyRUSG91VtuwQ8wfAGg/BU5w7TK2Ti6Kay1X4Jy1ZwQNDxzN2Zu5zkE1nhQFLTQ0p8A
kvTg9Til+q1TX0KvrksaEuRVR8Cvm1ibAX/EpjqdAeMOeeT56CcgnrqtCjvlk2WOUW51+ZgM1ceM
FVoRe3KqGH2wIVnvDMH7bAOaYoj1EzqO4f0rBoMoi0II52+dfyZWnhi9qeFojl4SmuyGzu2AV4A+
byNPakgQLGIJ8FTg4jcTLfEtzFeu72myf0NJ7vd5ZBcB6u/qaD4oMwrlXnkXeTOcgm3zHN1bRB+v
07ngL/HApxhQerU8oGaDXIafqn1taBP6jkLgTCXRi4JtCP1xpfJfCDj+ZNaq2pKg7JUroeKzokjG
3ZnR6QZxQXHYKbJtymdDxcvraFsDCiUGRjQYWGj3uhwyI7Xcs1VPZHjrisTUrEGZYllO3LyKFJ3k
hGIa/jjcNPPSMwjTgqUM4QaJ/MVj5RivJdLF1jWOcfPDfffLUmar7OSyOnclbu4CwMsuDPBpV3EW
AbyeQAO0tmd8ONo22k9YjRqTshmQ6MGFoCBLChOubUcwMD7JyGMhft1Ve6/H2TSpAp29ISatLH+Z
NhST9liIWPoUDNn6unzoKS2ec/UbUvtPcpiIePvy3P5a3NhuBByxX7vKYkR/kRgqizuA6tMddr5h
m7MOmbkDlbGSEWyS/jgl6kI6vbt0bo3OQ2473eGk22Xoftb6CsVRs7behdt6bOHbaxwsee1a9NkP
KCs2g7flTgkorV+QEh6Jil5zwL7G6LU9tdkxvlKZMt7LHLVvTko/tKDQPBG56xEAGPAmBRo3ofoV
YVeK7ODW5IOELQI0X1gERFyBYUd7/3rM0RS1WVSF8dOjhnSo/MUFg9k9YQkhVXdvJ4gZnrW+ob48
4Uwy8fnVjaEuKeNUYJCczcBJldmn80LLHGfUAvtdEcU90mNmAjd+p7cAn6u/EM1nCYHBAwMI22jM
e/xOuDufUt0uPJN/+nh2KazyBlrFm0Qu/4Rcde56WFv6VbjomR0mC+oH67H4d0H6ZRBqAL7yKfDp
IA7F+CZ/fJ7YadTDop48x1QLrrPCkHdquBQeNCuG63CHcxGVBRJ8cd36s2O6+E608x+4fzC6M9aD
w/Wmyf81vd/1L27KrOCLM9OsQFAbvmdUmlWeTPMq8KoKc59DUOa7O+o0pEp9EZuDiJsbeuoldpIN
RBtD/yU1gagek0oTn3+L2OqSlZjH946q6NtYrOHUs18wrZQw4J6ZCocAH9b4cbxBVkKVbFkviH8F
9TMce+QIklYSwYfKMz3eItLByJPyBYTnitxz5rw10IaIAPZXUsMhyuk/NK8kEuxWTy/7TI12M0gQ
x14YNNcnDTnXGMb99OeeN4AEGNWax52QsQ0TAHSDFHe7RtzA0bIMgNMTrY7XmqklBCin5edYOVS0
KepT9vJWq23WNxc99I5lEvLLHtHq8i8/9OriAlxHBX24Rr9ObwNOJvR426GkGSmjUxNML5B/YWc4
zfzCdN+lwCkzQi2686UuQtLXM9Fmg0Tfctv9fk/WvgQO7zxOdMP0tcMcgBg+dBxQTcY6qigKFvJ+
p4mzV4qPn2n0PHB6fQI+ree3TeBE1yklM+MjyeVWU5/SRiaaqNnvpudbAfbwgQMqiuOftwS0kfP7
xpiZrMXwE/3y5cDfItI/IsDTIXixA2IukZmj1ax2886OdG2i4frY34wrM55/NLq2D9gxcTjHVLOr
oM9U3Vqb0Fa1iyaxPksGNn6Onst2rSudW82GYdHlZd3Ex0fq3FTLEZHx7sxeGbFTiuvodrtPxDr4
gmBtKQO5CsC3aFx/jf7bMZJ7PdwCUgmvPU3NOvKrVBH1DW5f2g7JI13ZY0LSamItXixK9bBfwER2
xwhI1Z7gPDZPtcw8bU+5PUaeTOn/S6BYvci/9aPQh0ZsqMwWB6hqRag8t9WBzSx7EPRu8vQDMRlH
nHeQwnzmdADpYYLYiJHX+X69zHic7vrt/bSvN2OrpELds3RENjSfjiwD4WczDGUv4IipLZ8dTrCq
GEMlb4n2yeDd/2vxpbE5U/PCixuBXDJrCs81MoICGHMaz9NQtiRPpZln1FY9+r+mDgQTvsvyDQIg
dL7sdObSCb6i3MXFCBiR8CccYjx3LgnPBlZhzdGIqLeXsyJ8DNwBajww6hyuBF/gAorTEujpnhR3
C71D9A4pCcwiLKC9LgAeY9izxv/pEvqcw78QlKvUKWY7Xw7SCWSWTL6ZwBYbYqjqkLgfI3mjhuMG
QeGhtSBd8EPY6r80qVThl56qFu27+Gcr6fNHlIMVhuezRvAaaigj9qdpFZ5ho3ssUcGMM5Aofa1C
JZNoCx5YM7NFcmN8OZPCKkafR7MXr42OFhP/S2zbFYG6fiU23j/HKrS9pwY5P4/1dxIWG/Xc3E6t
qbPSmgl7DKs4XeX9OIfHToNxowZkXqkZNZtFCy4Zi2cv8P+zpbvv6m/jGbD+VLhp37PWwscdbXpW
mupboUeMgOQ99/wFEpnVwUX4VZ5Pjm7mxunJbogngcyAf+HbIPZ7O+fVFIgZJXjVmst5zxMaM7ow
hrnlgI9W48pMi68aQwjz5uObKM8jsMZkb2VVyT7hXXg6lIKH+uVjkb3tjSQ1KvCx+A5u4kgltLcT
ZFsEQHFKiwWDVZQtM6TkrtZA8cKcQ6TUntb7n9xHaK0AJpAs24K14d938ePEVrZiXo7GERhegpsG
ZYADelCh+6HMdRyDE9GaaefE6d5u8GLE2gcQV+b5ytlr7EACAz7oDTLi7YAfLF1WWnHHDimUgCWW
iZh+EfwgjGg89HGOEzFa7Pjrd7rk1hohX3WFcuhJ3TOJnbcLl0LxjLt9wK3gz95W/gaVLhWmkdfT
uWyK968Z45LgSYm1fVAaXtUyvmK4j+O/989zppaJYvSN8UlVmmQyqJNdu9is2/5cuMWpOYo63ag9
LMmd4bLrm/bog7gngTULJ9Ppdd6adVnGU4bEW44iGxdtumBCv/ahekrADbMng58b/EwDeG6fQXtG
tgAG6x9khykPIGoRXTEQ7uyHKoURgDeZAsYDQvge5yaHU8/1aemSQsHzyUCVlIQTb0B5POeizjKg
FmKlJM3KrIPM4mO2hcv1wBU5QgncAZze594D43tLl0t03RgETD59yZ00zzf3FfUDl5fw48EZJmQu
1GbJJzljHLKG6F64RNm5NHIwCRD06UJ/qIT0dFpBNPgagm8tYSQjLSoxEjihbDFz9lHYLTFswW9/
0fzprM+l5SPv85g6NKuOSj6dlySQd0MaFLW9LdQt8KzUwRFCq5/2OChFf2xTpyfbihmv5sXsNkKP
5JVC+0BTnxGjoD/ckAjou2rBUx2EHQWaLGImzSfYTwa+hcPdGKXQU0v9RYcsHHj2CYMs+CbxS4pA
mveUxQlwZcbvmPf63c0SsuSWbG8gpHx0AqSVx8GjUs7BwjgV1GDoLuJ29jCTcLjyCUY30gHKNRd7
5iX8w+eEEWCMuZsl7BRc+r0SXKSLzh7eUxVtnJCpZr0+IHB+EwotttLqfVLj/izo/E2COyLTfOfs
mkJEvdgDSLRbWkDAuthu4SOsU6H8VjZg6NeLO+EMiOT0KvuTphHsxM0k4Lmd5sBRN84Q180T/f2A
wG2SODe/Z6TEv2eQyYmllxe/iHQrpDw7NR3xWVnklo8L8uB+BuIBAM4eJFAiaQLC3BW72WP2nP0/
SXNZLwnkrx8/Jgb5faE4h8e2IIsxu1bdmuXvzI6Cn0wmp97ZFwBCujc0IcHuJst3hrwr91X1zZEH
TC9Dkeh7rpRpsPNNvKqcwQ8BoF3bdOUSMLQqao8c3F7cnFAxp9+hJqi/LDMwqJdNiS3RFR5elEVh
qEfDwADQp61ZJ5xhVtN/ssO+nTILkr7ZTzG5T3bIKkJJMoYOn7IGi5wSvAWHpHOC36fgeLXe2y2S
/Tc3h+co/GpA/Sx7cf++zfq7DWsOsKDsQ8xGw4DNUHV+4vreGT6WZ7dEH7vMXFHjmMnJcbp31TX+
E3d+tSsjJaycd3sI8reY/5NZ/uxEn87ZnV0Q4xwH7ujbIVyR+vjiDjquiR0eBKDqzVqNtHWYT/CM
2nuSRjFooAuhdZhKUM6c/CLQoia8gwhkmXomVrNyDtV/V4amizUKL90ARS5TfrD5uNhZuWmZWi0+
Hq+siJctEdbuF/gSXDQzQRBCIbATfpDZ9JtnuQBhG++y9eE5iJAcEZmywLexWPfLGpqb21QoIucI
NxhJ8gcoJ0i9p1CPinTUGce8hgAx6n9Jc5cwyWxUo/X4sSpvqwDN4hEpbcqn74hTJqA4lfMy2cjk
MpfhiLOAeDnUPjTpUOcSDDkCQ//Fz1k3TUuetrM4mHSELZHmMk1qvokz2cw8qr4Z8/lAghvf3OtX
PTl+st58UjP4NVsEVav4VOeooIX+2X3g/1YtaKPSy4RBTyKrnVCZIeLjqnQnOp5pXX4t6YXrUqPt
hDwb/IUzNcBM0Ag/kpboQDAE7PqWdSPt3EcSbtq8CKKBgKn5NQwJ1Zwqd9h6DiYjg/jRGg/wt6Qy
P6WFVf8CAsx06baR5HeO6EXkYGh6hXkAgKvAoJ24lQ97MzQLpWRehAmI6/JPQZXxTRUu4nI9Eyi6
Idf1PKJTv7geICR+vyjmjLYV7Vx/ab67nQGPDpDRx54qxQFvRtJaX4sAzCIhVmT8eDF/BXM6WmSo
zCYmDkCwtkhL60xiNwa/bTuvaroiDr13FsA8W6PTeTdCTrQxLCF9N7VauhjzxBnuo8JZGXAPOXES
lXuNXuJSxrL0oM/H3jr82Ymd72GH5nkL6sRttQQbrV/WddPrq6Y4sz6Pw4HWPUOHzVQG3pnoN7b7
O7cCk6YIm7zEVk2X+5hbkQvWZw1zICX2a9AuHlnxGiqkrSBZikgocr0Vz1WX4B1kzhbrb1HLebpN
VeP1Du3mQ0VAPqotAgtVfolEcdcigYSa7vckCKcQzcWq/hpNvgyAtZtru7jHEzK1ngxTG5zqtcyD
hOSBrgsbAHHTzz3zmrNkYCifJYuu6tfb/WpMxPQdZ+VVOtrRTr0hhauyme20jz8NKNSiQLDD0pou
Bmpz8Er8TxMxP5JrkGdwe/BKXJcqsrlN900Bf3QFS5u8hzgPoK1Wf5Zs6RlKkMAqwbeRQ8oQGr7g
CfugkYhJpIjL4qZf17WZDtfdcFzWpnRH0bkZl5sxz9a/gz0LN7FlFYCi7ZCDnwA9yw/dKLVn3QYH
aIhSEEGZsAuxWKDluUSUZoEqHTVvAW0ahUe1ZnkvY6Y2nHisnd0pKf/XbbI96XJcC9sEoaklXwiI
himjTOc/F4SrkXnJVR+Q1Pu1YdvgkG1/Y4CAbW0tBf7kILIsZnrV0L491F0sOLD7Ng57XkkJ0ZxG
8HS4zvFzsO/ubAng10/eJkzj4pf/LovECA9wezP0UJCSUlR16dgZmwLIDUmttQCFJu68S+GHv4LJ
wDG1dyFjNb73AdM3ze5M57ZuFKTI1NZh+kWlkykEtDGMq6Le27rxe6POePhd1P44MVcyoEtrvhl1
cOgXZNU+leiIEJ1Mzpq6cytUe0XjOtAB9HDhSRXCZd2MFNUqlcwhem8MMZnWelmO8AAmPnbIEDq7
w3dY4p7A9uWNZ80bz3HhjFzU7pUTKGq0xJHKkX2AWp5UarLLsS80aZkZSMjBjrb4CzuAXmSA3Ldx
8WQqf3OD+tKkwiS/dv4yazwcCgyx0/vtJ14x89jba5jFDW2MYIob14G1op8qlprlWWwj3lRkKP48
Z35ujr5+CBlCWu/268L1hrJhITKDiut9MBcME69AnPmkXjxvUtNdNLuD5oXGU0kcrEiAJvTIoO6G
3LRUxLhokCJ0ltNMZ9q3N+mGHgs9xh0PxJRwzA5Xuxgrg/8wTVs61/YYudXpmBvulFffHJUkLZ7V
tz85zYyExQiZwOGI/+OUX11rOcFfKnjrzDdWK6BgbjraxH0QQQ1uFywa+23xfAZID+VsYfHqggPV
loOHEaaHplWoEOSLZF5zaSkJiwoA7i5hM/mXBBcTwIwIZXWV2h8tCpEYABjEeKwfWlmEHTs/9FTb
Z+S74v/aRhsGa8eKkraVfSQgHcGkZdn56Cc4KFSfbT7fzuIex+RHpEFsf6f2ejOv9n3Sr2Hy1jiz
+7fbPBaYiQ00vsubu245XFuYnG8YE/f+zTZMCDmELzVAboLW6WTLJprj3igpaBguvKi3BwaeOEQd
JSRwl8R1tTkuXQbs40L+HwgtCQRVI3cwqvknngO4gVmsFGHD55MtwY1j3VqZ4mL4XuT0+3PibWoO
Ww+jpjW74jMsB9iNNc4jG95UsUbNUqtAAOK/pkQBFNPjTAk/g+jmtclk4EBXq5Wp/9chvr4BP8/k
RqtkM2yYOIgkyTQMH9BUwm+ZGe93CSr7gjMvR6cqp+pyY69qziT818J+/jphVj4+psXkSn/xJgsy
pV6l72GJV+SEwQ/i84kAeCAsn520d+x7uB48uzlMY9cQgskp8xZ3FitDzOCLVFgQoFJJzMom51zN
cLL6F1YKL8x1NViuUgW0+u4vLrFWc4SsCB0lpYWLJNELTCZOuddCRYJVGpTadYl5PlG4nxcLCrfr
2sRj35WNaVypTGewUGRqDf2DZ6xhFeTC2PbNZ2f+CDcWURLnpSPDWsqtD8g2ftIfCli3Lm21Fl+6
4BgB7SaRdn9iKb5g4zFiwsRNzpajpDjHOiuGYM5V1QWccCcDxWRxq9mhn75YwgAINuzT0QkFTSDj
/aMuEQESgHk3yFJ7fvodg7WYe6r3BwBE7zWx5D92/m4wOMWdvsVvB2TdCg6QdGl6cJrviRQfBqJ2
0OSvyaMifGpTVHzY+OOUqG4nGHKaIyNXoyFRww1XX65CRAo6YRWXPqmrU1GSbq9ACsgMvbLJ9XIh
8Gp7Jv5wmg1xtGpHz1GglFR739tGntamaxLxgCp4WhPcZOxWnHvhhKgPHlaO56rfI0nUvNcJ1CNu
0gBzMuZ/jj4B+ozxWR8E8dilKKklHQF23OBwuQTN1hQjvN4F0vjvVmz/AEp7Nyvyqtye/DT0v64C
YxYaZ1VpzdWzV2CvyYLr5/RdNzMID7gi3le4u6OCZh9QfQ1gLv5KdptuGjYzagsWQeR2iZCL0xJ4
E/aZI8ZQrWvIRv1HtSxkMGD8xwTdAtmLN1LPLJ6WJ9LbIhnXSzPqeVwmvLNJwtU9Wp39Yzt1+/LL
FXUmZNN/dDA3eL9EYF/b9p+FXEkV8t2/QKfNhKsj5/PHNaVxe7BZXRgrfvutUXxH7p/U0+Ib3zgm
ewOZuXC0zx8zy3e1gwxikWKRg+nsLJleSC8/s9thlimUcGG6LMGShMWpVzw7d4Jpo3Atf0LPBwYx
fh3BRW1VZT1MG9BqIFy3N/lZAG1CSbxG7wAvXq6EGc5PY/eenwlREIBXD/aNYkxZrdDSFT+wBlKg
dS60f2jnc4bIp8KdhBB13Mrd8iZlmIUH7LMrE9OyXki8Dt/xlqGaXcQyNu42ghNv2/kKujwNJRA5
1Jl+3J45O7fsxoe3Vo+DmqTzcAWhYRcdTKpIDnE+jWYaKlRgvT2ikoQzZxjVF4kqXZWCSbO6DvXo
r5lwWinhEuRd4U9jvrG/aCSYqU/pTIZREGT9mUfu+FJ7mbv8E1dx5jRrZ+Pnx6JmBpKbSH2roasE
rVxUHTb/wPaBnsxXeQYDgUbPpYtKXL+OLgKFEQeHDqU8k1NVbBHMd2CWuwkL+SHufNlgv1yx/Ix3
wFzwJ2zE4pN3xpMHU7RQ736HHybczgCEypTXlgof5f6l1yqQBvUegYgVdlO6smJsAAZZlNsBno9u
51UMbB68DqEwgeD8w42SMTGyTNbSvpFpbgRMbg1fpyQWdVhr0Apa4JLMJQ+5TI4XVzFhNtGxuLl+
8r6uK8zCFzevgmnL9CNbGTn6MhJfyKexk1FAB6XNtKLQw4+be8g0RfX5iEM1pUEfr86XGUfVjrBT
ag9lYILCtmNtKgur5aAenYFx03WtqNOGuIrSRNfBb+9NCOY6j198MJ0joo3b6GSlShWAzPdamHSO
k+0Vg2yFwxygM/hXgAf7fzO+9JtYindNki73YWEQL9lya+L5NR2Dbqn+5rWgf3wXjDbjEf3Sgnqi
Yg3P9f0Swh2sTWc0Xrgb/G5vLgpzDMCj2veuuhqJdZ9AxcX5ISYETD/YtsJe++U8v7F3V8X5NwAg
g+W2V6Q/wSaIk2xj6EtQbp3TjyBsF7EtX5obm0myVBj5WBKG+ljdTlXXzUJIGXqz7To0p8yWxzVX
49HLjzBeVVR8nM/emLJw11w3slL2qYnyGQFIVtzU1ACZtr9Zsst35ki5OZZi0PmZ5NSRVQP4pLy4
qB81hp40Aqwu54AuI7sQBKmW1z3sjrr8jB7wz4GsQxnKnexQkQOcmLHQhPs+bGBaMGCeCZBxNFme
+W7Og/UobXrz6GFs15rzGW8TQUpMD0VePH3FWV8v5uGH+kwd2GSzkpZKLhjVfS/wE8WLvY3cs+YD
Vl7PcovTymv6N83Ujv2bHmHCxpsiUUGCYFsMZUCuzRekXSMFzhlUwMX2BQyTeGzSPgn/tXJdGAbr
19JUFa9Uxi/ExFRgXTErqqJQaIbTGC09Shau6BwuIlhJOxV6pnT2zDY9bPdcdUqYs4afKkXgxxR0
JL1vMIg0wgVMMtNLwfjKE/CsH+53laxqEOZqQXl6O52Saa1rEJMUAPhvMW3yTo7Mr26pEufsUG2d
dsc/8qwB+MpOND0KzAT5r2V2XVJd4O/xrJVfXRP0XBUhIpj8ClWjnB44pC9WgbERhazDfCr/bhhn
o6O4ng4uPwI9cOhB/TtfgufyDAd5kECIXwKISbuQeUmBGCmg8IWTuJXrXgeFgMO/vew9UAqrIpRj
3W1DfB5Qu0k+rZ+quWM12GI1BH5H8XUrfsovLNUpyXS5DbY2LZyAeSNbT/K4g2bEwEh3uoL9hVJR
/otC0R0NbAiURz6YEl+TJxXV2l8IG1416HnqbsrLyeJ9/zhgq98Cu/oH/V/Wtv62VccX0BEs170K
VvUUAReoi2YG8OmIv92q/I/CJ4dooX8QEGrtDo0scWCX+gWKdZdnDBdLZ9kXDPpGd4o1dbLdgq1r
fKMlIgVf7fL1LyShpOb7X/t/pwVrn/yWHALcps0w9wIEY+01kvW8qzRgEIgCJXT52brXNdBmcfKr
pH3qoT11En1j1MzeWOpAMKWErTpRC+OWMfsKMXfmyyZhJq/43Kmua+39AkK3/IxtzArS1b3qfl6A
/a6F665iaGUiDgy72hX4pSW4SG0aM7Gwk3xo9O1r6S8RXv8yjMmidBp7OemtttsJcaPQeyIrONhR
5+XHFeRCAqZyNdppLHkeGW3v4xvsegVR7XZjIHPi2WSJJQQkP89JDOhh5UpZMZQk9YGeQEMYf1vP
y3l/b6d7u0jWtf5IR8l6IW3HgfATV4ywcJGfyIIJSS+z1yQjupdbymorq71mvqUbRnGKUq5sMnDC
8yalkS8CUXwiarRx4c60VWzgeLUKhm0Xa+FhCOWpkiR8kwv5/PZS9jT43wuUIDoMFaSs/KNRyhc+
hSbqqoJsyj0PxcxiIFwOObasNx/ZKdF/+/ZjXb8FsEvG7ZCFqguMRx1Osc0CXhyRLIpdSkx2m3IX
gAz/B5Jq22NT7O5Ojqh24PXcPzlSN7HufZL12OORYJyrpP2wSCGNGVZiv1Uy3tyb+D2J1/zJviRb
tOYDTzzL4R+a5U38t9we8wmzRoVyQZGzlRyV1ZcK0Zu6krzoXN5f6tMEv7Uc5630Ec3bxwFIigV5
lbPhg5Mb5mpiF+LA8rAgpkLJ+SVAyVSq5g2yDOaKHkgBSAup8mIjCRRb3fGdNhVQv8FKRXRSNNPA
ajPHAbL9hmg9AP4T7lWhzuJfsaz7vcOPyDwD6b6FwS6fc/35Pb+wuK+jznPOlY63vZctA6PUbMGs
B7W6d1gT2TyDanPQKa8hJrrNN2UGuUhYSlIC5J6GYcpTFq0Nkx5gYJ6skJ712lplpx/VKiVFPXaQ
yL+2m9eQT0a6ULNaL0Y2VIbEvyIh2O16sIp61n54hSIa7/CuXwUaF91GTPkYPljvhH7PFrGxqLXv
9EGF/xbI86ay7jnDKkWrI/dTQ3KtfHQbaRNgIR6fNHTawIbJUr0ylBgg99JbfMp6xhhWtauyo/oU
KVXRSIOsbZlFdRPjC7u/c6MV0XFBbp/JbpZfTw1NGUrpS2PGa4E7kG6rIs/mm9Iu/0jG+J7zuPLS
IAb/5Jj+JCJoYyoMpvhMOKNGU3Bd46EDaDGmSvxuTCokgrIcXDKyiHSuWxAhXMACqJjb98XS8U3N
piTmVJoQrU0qoSqyduh0Klppefc/DZyON9b8tqXdyttmnG8YeCsjSWyYyXXrR4BjgnKbyQiDWwgi
JU6oZMKzlxUq4PipF6q7qiii4nTeasl/AyLiO4eL8Krk5IL06ZCJqnq5v3X7emXEdkWLDyXGd9tG
r8VQ5myT9XHUCvdiKB+x8BpQWmpDai1GJhDUSX+wwO0ysEgIFRFcV58tVJ/NTNO2p51D4qXvM6iJ
y3lwqHph8NIDUbC9P14MHPZsbS6KxdCSHyVCg/9Lv5nBiJTfZvZb7bT4F+ufahFkOdMo9DOSujIO
M2Nthm4WDTvhgaBHSlHLsmd1t6PbGiD3RTpvOKICIt4zZhSCnQYSWuTWY7XbKFavzJkfIaKfUDOn
Hmus61wW0tw0oeNRKYHpvnymAA3EW/HE7zz3BWUdpwueUL6Kb6PEQUGzH8e0hWuYZdS8hdhqaZg+
13W0QsFXba76RU0Vt7vB8j5MZR0G6yQMPodjP0UKV/gcRCuYpQ7I/nQx1tM4jOztz22LB37/jx42
T66S8jmjbLRC/sSdkfy+u62pTr26jzbhJm9qtArs0YY61ACQHL9UjSsE2B3oqNi6Yebi1UEkP/pE
nzfKlLwqQYwj8eRmHPerO+Gufiv+o90bfXl2PsnBWq9PezllZ53P99XQzfBtPDo+wl+VAh0=
`protect end_protected
