`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12176)
`protect data_block
LqyF4N/Hte4EBiG1kZRqN/Jj/f2vsSDkWu7sk6tq2+N8LVcUr0VOmlHMSTuhxeBm+fK1KM7REfIz
KlkNXX4aZcqPl9DOvGgsIvy7XmDavRqXxKdNyJgHHTSqRmpn5M5/bDOhB5yjN8dnMA+86yD/VloA
FOxCk3CjI3WPLwV9qJFdg0YkH4SOkCIuoNGy0iA80D/ONdJtYoeJnNhBsLBvDx3fgI0Qh2jLVPVR
DDbE6WGLcUufjV46ZAXb18y4hUNKvAvU4DNjIQQK1tP+lvfjbJnEkJlQCoBsWm6FbBZLrCHtBo1l
wuZ+UIbm4JAwI0JQ/70s/kSLFT7MiKOGLIIGr3ootEBIntgUT2ie2qogSaLLdmMV3nv7AntHBCN7
hj/gl2JKIWlVzpRJkV4XMU/y9J5WWy5pVgLsd/XWRllXBpiiBwGFZ3nVcRl1gY43fU76WCpaKBpu
B/HW2ASDRnzDwI/t75DVzYqLpQ/xJrYSBj1RoS6t0cg9KTXOhNsm6RqaOddDRselTITqcxZWnDqo
INnjB1nyPk9xnm7uKcmaPDJv6STeIM9rkK16XEcBto2TfDNKhmRdept7Gam4JOhbhTYdto4VLadC
M8FC9VKlWtNILFpVjoMjCaXqCD7cTlNBD7I9cyGwWQVHBj2gtbW6QLihYc5BfonDecmj/Ge6CGVS
TKiH2BrTa1sTi/3yqshes+o+Ycc4FC7jN+vGhPChXG6QOJ6PUbjgQX937siQEgspRdicx/bCpBRD
bbEu5lRS7WOAQyuOE+3TtzpDfteXJjWH51/52dk+tImr9cFAy3PEWPfhMKeKBTH3PbbpyJl/7CIs
1F8uAfL+36NddtVMqMEkRCg4yjACPt72w/t1z8vGtR9F6Ws31/AowuBdUzTAWaam++yCkKNrZ6Hy
lyo9FrXbqH9fmkq1i0GaRFaRUX8FRFFspaAEvMzx3iQ1Glq65bXNdpMl/9oNIPe6mYuWWA4ETg59
RrOv2hath57z2EoRUMG1zKeBqmQikRS9zGKGFFcmrbEmfuJb15pHEJrP+R1RsP9uhmrJGRgSD7VA
SIXYIFpp1uVlk3hXLouvPXv4pKsd2rOdQJ2aIq0mYq98KhnF2q3yyNQCbY+1BkIs8JfqgQeaUgIy
M/rHka1rg/tjiw9Lq2rGvQCCzUNrxt2OwJtlj4NiN3cvSf6995FNx8LsO7ruo5GLolWi3G7Q2EA2
Cn5Lra0ZhMUyFNJjV+l3FkBoKkYERuTqs8JMQb9BT1LROO4bhPT6jNcxKtq2C5rz4TId8dA8YXLr
Jlich7uVRlHVQXv8VogF/vTTSb09hjI63X2xWdzas3h09t1bPY9V1taJlsJP2HS57QzhVKpzWpOF
F66AdnnrTxcKrgObnc+EUupQd5O6v1g3/vJBxjmTRc5mFPdxuTTXUESBgqe30jdGkUiXczkpVsyG
34gcRVScnNRf7OUKJ/ksTu+kk9GdZzYbimcs2hq/k4orre5OX8v8Bv8kHU0KcFm6a6za+oA6cCyG
xhD7mQDnEGbWapZR5dKZaNOTUQfr9ClH0EhxghwKokj197CSWzt1UCXFBbsTootk5XZzO/378DPL
VhmL/NYn2T5Wx6uCEJOvlCpXGoFBCVKk4Sr37+rsEJM0fdN7YPkcztqzn2UgWVACjfxBh9sj0WuY
n3ZqH71PcRu8FSOOF3Bopzg7RIacNOvmRkgVxm3IAfT9QRxIAe9ZlfzV6pERqg3lVHEtbW9vCDjD
9eGSjNKHEFdO8Su3rQmPKVG5cJke8a5d6hd7RBMZKJAa5xjNTHTODlYX0+1E+bd+2AgRaVfYnWZ6
HucniGSjCkLE2/dCC6z4ULXo+tCW/Oa3wJL23VPPNMNFi7IMby11jnW8/EuFd8JSdULfCHlpJO1c
WA9ZDa+dljF5P8aNwghJgfawt9zVNcSzMbjxTMrnZgyl5PsMX9mH8cHqBFi0R0D0cvLUlvY2stKk
0CgjXuSukrKpleQFx7rkH/mYgcIRRU1XUCvYj8m0NrXukyOvtCOojtP6G4dUb1K42ZZDDbEfcrDu
BNZhsTFSigCG93BbNtHLxarLo6vjwEpZNZJbO9ZJbkjEVrbveNWh3MOoqmeAnGd807qFivYKdpYz
K0S7LFRWAcIixWF9OM+F61Jl3di1DZ6lUJ1Ajl6RbzRjOfpndaihUZIsmfKCBoIqtf7pPenA6W+l
BNKIRzjEvt5a344yafHXWg0gg0aStokG3eJsJNpWt5pCKHcxg4SEfseBnPUBugdKTtGMhoVLKkcm
YeMQxBvkknrCUYEi7ohAe2ehrNRJzklYO6NUIQ/vwgbdrIgnUx+7LQK7K1KEm0wZbc1ykCPPtVUo
9PU1SGPYQgahXxTTdb9vfT7Pxli1rzUgS+qqkpRJ03qoRzVEjYU3yTKJoKQsUsKd4sEFzkD6PnSX
X+YeFrNTqV2iSJFJK6BHgN8ar1TnfocgwhvfraGZTg9PLhZ979Be0vxpYqyLk+WNb6xQs1g8VoSG
ld5JnubqNvxnLz/rmGXH3QHMKx/+H1NO/hj28bWBA3EDOwW4NSJvbWjyaX6ceFxqf/FBpPsWORjN
/thWpspz+fDJrN5cYo6qJAxKvtWAVCkOPC7PyQFffCd7Shait6iU+bfJ9mIz2sJltD9e2C474Ibe
kw+clVTWhCihN/1EzzRPjF/nuM5yq0lvvCRvnJK3cq9Gfa9HUAW5P1/oWo+5JjiAU3kYnx9TlbXc
elVNTAhNYjLWa+YYZPhs69N6oGGtGGRl8IaNgLdLeF3gCwnC8Du3QNtaztOsXpwwg/DYW1tCmieV
c5wZvlpSXV762mrRQM/k6pqAre+Uk3k3+1aZmnidcWl4fLywKzgQCQ8HYMKTgNy2GzmwrwiL3ST/
hcASKuVvJ4kVnahK97MKc/gCiESx9roVlr1ld9BCpl1aUmF4iOb+mSXGGSfGaxsE9ATH7To3Js5D
OGVwrXR4rBnd/cmisaWgvTzyLr1qYrLt1napRdwnVjSxxjkHsI95kMNCb+XPRYgsPCsdxJWxsdrg
ezSnqD/prFB6CgNqBK6CtqLb4gYsKjXgxfD0j/7nSzP8usiqxMIDSVbNcNI7s8PPQUU30igyJQRz
/MbTRg40uIE2Dwld95qHUl0F9iSDMkkiiClyVP1ZzzBdSnr2Z1RhrIvAC6Eecs/hUhWyYp5msePG
w5hEz31HpVe6k8+e2Vm0k6PvWadcnviH7pmavZZQB+CCxdDSJ5q2ouB46LKtXByGNDP6nHBeg8eJ
Sxbj6YxIVZsi6r3EIHM7PdE307nfoUJ+y2URFtTs0g/Qen5YVGSf2MuSNcywPmEF3nIeSyPbe3fL
VPj6DSc1npxuSMFhheRWnJFsoQGFGJnm1/FCgWLxt8NsiW+Tjb4FQXEGoL8Q9Ia0nre9ZsWupy92
mIkXkcCRXoGlTeUQ6iqppC9qycCbHWoPZM6N2TxHJboOx/fu/F7QTkttsJmUmqjfbBJY9S2YsFTS
SjFFRW6sm53hk37iKVbU7fTcagkM2AYVq7w1v8vbIB3O4zxUoHAv0uzfm9hLZ9javuaO8AGiD++u
lh/0NgiraQmGK9furRu7csqz+eYnS0zXJmAspawnPBI+bO8jrIqUQ2Z2QHiB4ShBq905VJO486n9
41DRFyL0ZwosZW30qcj6tcjKQzKt46oGjU78uerxoFaHl4IygB9M7O/px9vMoOuuU4PXXCAVOvb7
cW5EBhnt6Jg1uSsucJ56PxlfeybYi3NUY83DLS3i2yYrJqKMFINzHoyvYFuDkOqN/sZdg2YT/4P2
BLc9GYU71h+HOvqLvyoLVfQSK98SVFN+Nn7wvM5MKMyjFUA4tJY+bTx3cmd/9oBAE/oBjnLXfNAL
7EOv7leRLhpCVUqrEBQ65wAvHc2yFX4SZqno8g+J+Zx+5u/MOoseJM0+sIbsxEoiJkN4qD5ifGsL
tcOc/HHXxflM/3ayYuzZ7b1nV5sBauHPrM89dCsfma8YEvmZpvpxsZ9Mp89oB86aScUwWmk9WLe5
V3bilyq+stO73jeV16VfX/aDy48nxl5CC8UhStEjuP7p0BB7Bom/XuCFRjOaojofUxe/dQqV9bfC
M9fqUJhUp5PbGa8mvahAkoc+4udHDhkaaaUGozljT0EIHRXh2tOS/dRiZ1/yW0XVAisyvBA09aIk
cgPRp3FfW94igApbIIRP/1rybc0zCl+MPc0yUVmM110rhCmlrgpZu71Sx17rtAGYb5Qb6fWWrpz7
Z7+n/nf6ic6VnK++Mn59YJZuOOkX0ObFE4oxqn891Io7HFOuwvM+5cD45orcvr/Djsov4OobGCd+
b9KoGp1BDsCiZqAthgJCEpyFIofVl3VVUPugFMx7ZPtETYCj1KB9qFJVXKc10tIuRRRNL2Q88zCE
G69ioAFd8hW3hNRM0AH6C61O971D4VSZ9Ivhtf6fIa1MrfaTy1b0LPIbM3Ch53XwfYhSm1T9iNNQ
ybtE+CIbmGorUA436huLzaBMnbJf4CVWmx9IKgxtYXjbcQl3/Vs5ut1wGIuQJtxRmywf8BKUnsIj
4FIuI0E7lewT8aZYzcef2UjLE6T/ApsMT+x9rPo9Rk3jTAbshLuVcG10IkPczrjdmVIb/6YWUcId
fLzK9QKbPTl6JllFfwzsyoRJfDwW+pMZ+Y8DFip6dYEi0VvdE/m8EqIbHWKu1ujsmCxdkyQb5+w4
T6nEDmA8oPqwO3P3sQr1CPVTl0kNZ4G37fmFQgpLHrfO5fNeZVXlePH8NyVb/y7CDb1vhiyTxvKo
jpBiAsPMfUJOCY1fvbdt6Uu5T6MfVXzcOpmJm/3+qZNuvJ8sdCcG2P+7Z/KQq4EZ1V+ntgwAT+JI
mWwgUzyF31v3OXyuFid6XSC/04vGK3HR6SwCVaAGGBqJRO3XRBo4pmeZTWawi2TLsXYTfq4A0Cvt
k96W1AusbsYFBxqqZ23QpMXUiOyTfuMGDSXHrWYh9eRDXMtjnVpbzaRQybq6vsZSp0B5KXnR8CyA
QdArg+ZoKoMtdVA1NPL/izqVm6p3RVlVOSXYeDcR+k39V9JcEM5RVIdHyQurnkNjnTtnM0nssonr
dlCwRz5p533Npehcd8bq7ignJBNufVtfO6sKxFiCmQNNAmZN+oIoQ/nPUpOlz9HkxtZvssRu0VPX
oyJWNmJylgYw9cnWwF3o+I99tzE2wXs+fZA8DUuCC/sbiq8KT+9LMc/fznESz26VzFjOOtCjep8E
pujV0gIVqzj9TDma+31clOr9FcJ9+91y6DIyPYSlM0pjBkQTzdYFGviV5Y0Reh7Xq/oW8YCxiUK/
x/54qBtlohQ39a/3ETd1a40sQgf30SS4Ro6MyR5Oq6fDfCL134spALfb/bbgj6aSUWOu1qTrdeoo
2kYTnER2DALTD+kQ6v6Ehdrg1oQ+L0ekwLDLanFYk+tTD5ls+DVN6b13QRWzrcca2tXVJB18EZb+
WYaHI4RxPXX/uxWoLftEVTr0cEQQgZeIIRCwhrMQKRrpprNGPmd/4vibTQD9icEirYUoDu+EcxvW
v6qQ2x4NHK7AuaFMDvh5VAgcNDmlZ+Sf8x6ECdmALB1TmDAPhvNQPSrYnhyeH30zdUshMiirTMk6
ssbMQ4VTMe9XwIcEvCMI4ZKyeO3odIHrtKSjXY4p62MmIXR1NUaZ1DVUQ0yKVOt2JuCxRpBiWUba
AIzo4aFKfudbRb9qCqZ/0qVDvrOtc0PBrcauEgmE99R6uuhK8ALDPRgxaZeyi5rMmodMFM5dav46
88bTPdTaryuivTErXTxglMvuzdQvzf1JiCP9e7lK2zA/7aH9CbzF1h90upyd3jpSmj7Z1wqwcNoL
E05vacnsLFzxBDanmuhC9WeGzTHe2b40/O/UDg6mt680IVwM0dWfdc8pFgPFJgjnw1gakcSF6yAq
mPqciCLLSUnpQpM5P70Fl25KSvev5B2bC750QwyM1xtNpwf91wzmUi96xMKwJwh27L2sqUqfY+Al
+XT94rKEZYqoSGC8abIAjjLiaA0ibes7mjzPkt8Fs+EfOQ3cVjlpIPULOrk/suLGousOqr0KxoHw
P1SKnaAFQwequ9hQvJ0OO1z/pvf6PRbbjnlFqzWCuSzW5Qp4BcXJRbjlnpgj7tIhD3XdkYKg8eT5
eUa/k1GHrapZcbuBDsRffU3P87RFDMoP8pEb/2wOCTtgHz+GggHoRKzkTZ1rsdIqe6ElG/i4HzlC
foZQMI0zAoX8L69IYXNsnNNmSNthsuthCrJ+2hCiBWajR89PGxlzKCPSjAKCesx0wtLxIdcxEtlr
ALqkO9Z9MbpySJX9H0W7O4gTrWpvfeHW7CaJOA823ohnmgyeJTdkm/9QzEdOF7H7owaO88Cku3GF
Kufq9OD4KY0T+u3X4RJW8w4esYC1j7vYfB3VlRRwYYz8FTFa+B+kctx4yWj7m8B7716ysEAqfCC7
wj/VEK7S2Lhn1gesjIpKEy2XYZcPLyIF4NBYpuKFsgvPV1fXJEec2FCon4vupNtueJsltCKt566i
0d4pTX4GQLPhSk2WNRmN7sI2Fi51VFsniWik+5GnuEQT/ZguX65CiNfqMe43MpK0892leMBae54t
XAmBWvIdOY7NZjEYrNAQoKvrIAoOsxlwR03eE7v3GwWJxWeODVm0bgH0k4F40HKtFOJdGvdzjVcV
G1zGgVnsMZzhqB0FkJpGZL8Y0i986/yeCMS5SnXdHzS9pD0YOSJlO+Z5CAB3CIHXiFv3DsAbj00T
frXFGB/LlcgD+qlZscOTvrP721fWhig/uRSmrhMrvWTy9808+l/vEFYe3I5tzJHLUjc+7Hs2vPe1
rwfuuPC9hqsXtE+izgv/JEiRTZZk/RApkctIpnWWepAA/1yp+I3Q/guDMRplG4cqCQ+kMxUrAIjC
o1rwfcmyBDk28KPrsJ8MlGRFPrMIVOPyMavJn0gJVEDDyGrQRw3/vVxEzgyqFT5B5WkQEDYMGWZc
7eFwtlCS2AgJPFrfelZMLT7l51kYe8adL17r0SGIPevaziSRtmcNyKjWxWlKQ5qSwS2UuUfivHIf
mNhGhM8o84Ab1dg+PlcHXH/lk6rBNzlB6j5nJC2k3KYaG5ZHAZaoH0pyKvooOu2K7l90++y/BcMu
g9gGpijGpxj6L+zlF7YiPlGIyCrURlz9v4qZF4z+J+OqRzfHH3UxkKz5EDiUGNYj4tUXnoFklrnL
a7XYh7lu1xIMbPPG5McRUIwpI8W7iSfCx25TkbPYMhq2YsJqWtOug9VQOMJE9ltgGtUUTs7drOVu
NWtVIYMwzWNAb7X1VfGdjZJTRO8TrujYHFjsYoq/RyBvzVgwHYmd/RC2OqQUjFxSTAdItVUHSTx8
X7PGfgVyeMKVXpyQF/KaCs20kgfyVhrXBngu/VGe/rgxMe//Aps0NOzMuB2jmOT61yJu4j/4bKqU
kW4LoVFMRks+/eiB06eFtZQ6tLL22VIk6o52fuWHpx9k1S8RqMjsC4Q+Xn/vhEPxEOBedtvbr6hd
Hhi1R1lyZtvgMsys3zBEaqVaZKg0ac+tH/Hp+eZcTa1BqoWt6PZfKPQg6zOXMJGd/gvFIBoUZ+Pa
Hnxdwx2LhkupD51QklyRq1M/AQbL19aWFu7XRsWCvoXVIFc3St2ubVvNFzOz8g6/XEdFpeGgl92r
ulRrw4/vySsBh+SuE7QHPVWBVQtcDsZYpnOtME9tFFjtw0QEz1L8N1pgHkV8GtX+aPc+TyCoZ3VX
ddYqCC6xKsKcddhE3ShV1QvDaBGN/4DARuy9TKMLRXrzbhdS8f+0/kIhij/Y7YTFyb6LdD5DZOlk
Q7ICP5U27bkx84d29s54hXfMiYeknIa2dbT9gCk7NYwk5aKXGelPN/k8ou/iOicP7G7IH53cLcTX
F1nRhgDWIV1UQtPLK8oCu7yWKudtwyEgWoiH5XO9B1XeFntdK6WRyhdk0BS/ITyacpdBXJf4ZOM7
mnzmf3eOfYVMIjNTaKbjHXik5//IUH0HsvM6yx5BS1ylUUyY6aPtVyv43g+24NNjAHYkSLK3z70t
hpBr2nvNBNhRkcodpkdtM5kB0f61KYHNX87hpI7gYYWPTQ5Tz4NRIho0Y0dbxhPIdr97wRGtgctY
rgZXp4sqi+lsz5uOOwmUGGj4DSa3CX+WcKJKinqEP3c+1eLF7uW9OkFiY9FsAIyikD/6s734iKXI
Pr+ujYE2VaefyHUMhQgkUVEzHl45g48yHSbXeW+MDoKX59n72un9UfNM7d1pNDoArBEvgyeisHmz
yaYXcoN1QVBQuPZ9PonsDYoHTLfJo1LEFcQ+F2vhrueblry9+a0LaIAYHKXGWN5bfD8OGQPvpx1p
O1LjlJ57dvY9n2yasGKShbyfKvrbkuh43kgYiYv8axFaY0eKRb41IRdtOz3tTeeE+IYWe8owXaMY
EexBx2pgDjF90TiW5/43f+PwJhBcV1UYKQJ06oTS5UVuc7NnLL66+RgkjXEwtcli6eIM5+ODn8lm
tMJ3J4oDa4XLtCkRK9fbwyuTWidc7mzWWkkuR4ZvJMat0gNjo1bWmlqZU3WQlPYp7sBv8zauvajU
qGsAx8XaTOLk1s4vG5XzLuSH/ndGkCioKkBJac1I7JT6CZ6hoX46hWaGo1YRuOdcdHHQcshsVFy8
iqFkSMCUzrANrly8Ke2a/z0HrW26pXsYQxrI//8nHtWeOam5ubnFFcp80R05WRwBxe/KfZrY5Ncq
/VCvoJumjP/HKL+J5dRS0dHgfRJb8L+x7qH0UrbF8o8UaEO/SE6bPK7hKGsn1qaLDII4fRMo7o1U
RCAVoJim1KvbjYyHQXOMPuS3er4X/VkS5/E+9uRf2B3n6RPJV0c8FIJ5WYegv6AMir9HasLsLRHX
hgx6JwuGemZxgjh8+oL1ZuvUfZPqyG5s9dTjZMJ3qneh3uvSwQJ4a3JlYl8+e7wtde7gTCSVTcfl
VJmSp84/5syiRVaEaVhwU7PtSzNm4nHLgrq4BGMYpxjt1QxearWarldDOeP5ap4Ux+Aw321kDYiJ
ittSUPmjvm/ZYcn0ztvlucn5muqADFPq49fJhOYvmBY5g2NQPZlXzs/kj55qLH/mS9FI6DtkkbGX
8KIFY5rh6cl0IngOZ4TrzUkGdHah6kCdJNHUA21mipHY/F3RBUEqkBz2cZm/yBC9AcjFLtJtUZmR
YcGbIHU1DZXkaxqYilI5VQtpQePJD/TmWkJwyFStGrIp/sebV3pvVIrf8hdv6vPhTtxy3oBBwIG8
QnktCLXE+IUE6J9q2KIqjfL3xicoszEVicudQ8Cwp+RIfEqzMOQ8jre08ue9nfhQIffko+q/mCX+
TpIDaXksBNff0tHmqNA6nHVFqstOOAZndPxWMPLDwbFCOj4lYqmRkYSEm4U3TV3LeQLrjxdHw/QW
/UdawzikCdLo32cBDZSLsL4S/ZVt/iIDlHtqGgtsKyJ81f0upSpE/Jqqf2MhqFoQo+QcuHLSUw0/
8vW9A9QzIenF+uTxtIgJmPgBZggPIg2A/fTJ83hPsKKn7Hdz82Fxtex1W7dpCr7Gitwyjasl1WJz
LBrrt0gFqa3HSRtnwHdMNYajZZ/0+LOUfGDB3HO4zn8eO/myPeitIRXsoHcuMgUReia/D/97epLR
FhApaKMIVeMI8Gvac8jZh99IHYTuZIawEiazzEd28D0KcBeTPYBxurPc12H76MWFKB/3dJb6Zis3
3vSSueZ/gqjzj6xGJxTuF+qyQTJB01599lZaTO5M4eMzCmWvIrieRB4iaTHqnb0oc2lcLHpDvjWh
G+S3x4D0g3dSwvhou5Kwq02kQr+7R5/8LjWq++hMDeWRfXxfN9gOY8r48shotFWlFOSvS2PMy2Xt
GIbtyZxjwSJPxGb5cJF02sv0Zd1ObtdVx8Sqbra+R/GB8Ar4E5DgK0/+BsH3i7GQtMLX2Vz08kLA
v1qlE0AIxdG8WhtjZAyhTlp2NuIKrtAi+m3toJjFEXqHoL0zflGduj2/A2sWA2l5bL62x+fI2CQ8
fhcD3CcpR+fMXArMs+emn8J8K+6xgOVAMbbUG0ZBaJVeqDrsTL/j2KLJtv7pnGqFO2jzsosqkR6X
cdpkA0MFs2T4BR4wpcKBiy3OTpZKhmPspYTpZjwBC5YD0cuOsS1eepcObgKOa+R5bCh8s/hb+QtU
P9We59g8sKsSb2PDlGfOWkqGmgcPn6C3/2KZHIOY2aG8ZQrTH/109SzCkOvG00atnc5WXGR9jPpT
SJXNvTd+i2D0LztCOyhcKnxLYlpTg59/J4K6sWpLf1cpoGwS4bKOgWLpGha2kg5OHvdgjJ0yZS+d
LeKtCbdgGXfFLnc4D2q0GaiLOigEUZhJGIfriCsjiO8CXO8U2HH0zYGLSvokbku7+vh9byeLpw5T
zRbApM2NRh6sCmNiFltjQO21ajow6Pod23imTSs3XpDVQspanFCm1djeRTufIj1xQaD5rsK2LgAb
IC2g8oAUV3d6j2jMgSCk22WTEo8vy02qI9wa/JGmgkr44MhamqtJlbj3ijA7AIqlOpayJs4fB/KR
Sp1RERJQ4H7X431gSeAFBNoZCFsjYXO1GoBJdRz2SOV95pZXikdHW4r0Ce2BrpB+Nu8iU7TDM+/d
GYy3Iy/XmmOq3l2uAl5M8AVYjQjEDuRN2fIWowe23ORHf3nIt1LHDgCKrAxFwqa+Z6zlV9K8+JN1
cUnAouSNQwBnpSDeprvt2YQYqNEWkjjO6nfFweJJqlthUFIHVNY3Th4djJ+f2/xWLFdclv3krikV
6ZPI+epKAHvaJtgNFPck7ue87DbUEuRIhewsoKn2m/9OnWXOnjUObJzK1f6LZjW2sQel2MLF+WpH
+e3ofIBnL1oWAjvHXdcGp/aNxPIl15F+TULep57czbiaX4LxFPhwI72SbDvmdadaOdalJxd+vGGT
wGQmNL0X2eCMs7x/pAM1pVMNJ67000LP4fup2wZae/lH63a09JIX8B79lp3dX110AB8hEe+sILAO
g/GeLv8zLW1+kF9HyuBLH9d10+DAOIsLSCA+uvVwVeDeehd8pyskIDcFZpLn5LmD8Si58V0mjmzj
gAsTG7beNbSR67eWgHNWE0TCkjek1zK+hHqW+7XomEIXMwyEyZyXWTUNCrrV908oq5IfHRRtS9xD
tZzoTSVpKrqMBlE90Iz2jhPO2fJUO+G4VtWIMcNvRAWfBRzfCpWAxThkJV/JNel0vNI6bD93Zoci
c//9VvoOj84UdJrjaMT1auex0GZM5VeRjeWksBz8qXWisgPx8+/u2YjFTVwY8JZcxK1FbcHmjueJ
RdF84HAYQH2Xf7wufLS5De0MuiFK+r/sVBSGZTrJpKcead39FreQ2psF3d+si2QMzCTslW89mnqN
hJHPF8QPjaArZLye98pwmOA7Lwq/Mi5Bxpr8MmZFYG+rosW32jE3mDrmX/ljjqfiO/ouYHg6wxRF
UH90GqjDTlmf3UdBOHLnYnIJSn+I31IFT14dHUIodRavYslcxVJicpZAvu1HHsaD4Au00i611Kly
2MzzjV8SRaP6v15+oiTSq7zY8fuVaWG3UYut3AFTmYRUmHq+U4mSo/q7A2MER1iogGbWYxYZrVMm
Z7C7zyk4iWXnlCcmcc79t6djxhItgash1u5jbyZsuq/m7pVsPeNHAIn4yHaOcz4jkl5kxtaE7Y61
UpJQ6kWYeMIZbdX3GWZDAjR+Ha9LXnjzGJNMeO5KNhM//WN4+kbC2IAPAvCGLQoyw6dqAkNsoymM
NE9WI4IUJl1MJPHkqJHQErv4UMTpc0HA44TwX3k1bnSmqHFO6A6Dai/h3Nv6qMREnWxpZw8iEwR5
RK1GEoAh6x2M0S38/KyMTvy/Eyq7n9/oRyV7/MeBvAhANzthUZRoZ3Bc2eI6gwUTtR1+C/nAopTJ
OEobMw1GfPj7mzo11DTRCXOyOTKj/dyXGJiY90sJ6YMeDFjxfsYWrqqZnEyZtY7BAHFO8ZVxVKVp
dJICpqNvwLyYDblvUoyeRN/eXRF8susOhrU4IJU09sElm3l6Dw+2+ao2R4RVBolhwSrkF2PfM52m
b8DVFS2czcTA1Tvi//0TckCke5S7H/Gzxju1D7z18ZwjOg9KMCWgd2Amo8lAc5eSGRDVmuTunn4e
uRpBqJ3LzqHmVv/u87ATFiytQUqoYP7lGP8JV5kah1oRpBicospTggIOM1VCYataaAmLAwQ5Upw4
JLK3ENiuGXwBPYWs0k4gvWNz7BgMLcc2GMZNqD+GAxgM5EmmQIv14sXv4ergWncCixVqGfJeDJlc
l/QRmtu7KR5k4WpTvLCdDt4X6vo8A6wAi8XM1C/GvrEP+MGHzRA1r1r5pvfWIwrcPw6jQifJeBMY
4NoqDsi2cbJmUreXJTnndlXJLzMoDh4gqR5NYmX96kC7iI+lMD8243dr0xrnhvXOfBDMaSa/DZQb
Xh7eROfQ4BFgs2gl78agI4a8tdmJw99MA97RLhL39y1SWgBYGVa6zCFoYBLZpMcUz0ysDmP0wzG3
2eX4JB3C3KNkdNlQMUJ3BoVfQjDhhqfjdXVlouyOFfwW5wIEzCfnXsxSzde3iSAHlu5Zn4vWGABg
jkqVX5V/22xgjO0BgErWr4iU3DBnj5BKowpJaqhHS7IlpQ9+vOb5ql/a8mZHZtwA/YAjrvExA5bF
ZDdRqeQPVa6+WTZu608JVfUP2l0R9DqtSbMQI1q3h7ICCmNAVCElPrYszwbB494kfagrCfLWvlm3
lzUlQjrfad+pM2YoYBiaJLy7GN9mcZSidDzFiKUbvXJ1o/sHCGxtCfRryqs0cvWioRML8RmG5syI
uwbOdjFlq+Mgm5C86IR3arfddMO6He6IJzQbLLMPKQw4r2tTTXKQDLP+W4Dn6sLNfJgOVjpQzqFf
peSpvVjLKtgALS47K/c1uBGIrOQA4mIo47k6gc5NktkHSWO2kVI20NVkztgKxo9vmrKXzKoN1v30
pixwV3Sefg8DON7961s8EcXDQPjza3Let0D/TxpTOuV9tMGj7gKQkH3QQh5DJxOI8+PVdlo7jPEG
2HnVrAKmEhPkDWPLia5XUMIRxYPCbdonzxNKAP+h+/HgxOmaZrVpmM0YGbNy5zRRvs37DTJb63x9
fLg+Re1WdobBxEMscXmq+jPtL3gOAbx0xf+ac/PAMShKxyoCgdB9g48cw95Nk8DF1wMPFba7rn/1
YwYi1DSTWO2cm2kaN/Fw6wwUYvz6FjEXzaXwtEF44FTd73nX7IFgclCt/bvsCXhEYNT8q3faGuKv
mXm+l8ucaPdn8vnl3tvxrXNHw+urPep5EBx6L+JkCW02v+2xSfUH5bXdjqau431L9U7WTZ5w179X
/Np3vXOhEy/lyAv0H9xI3+9+PBQvDNbL0wT65sXDQqKkc1mG6xiXYcqPRXrfx1i6ITZwJILRS1r6
Jl9YCn9OVMJGHu5OWhCnovcl3MtcTsQOqiQmZwio3yYIzVDKeL39Ht2MKCO86ZH/lSByDqSlsqqP
l8az4PsrkCwzcYRfEJWT3qFS4wtFWzAqTE0lJ0P5tWtpXBYuOBUIxZMUXj6yfPJ3OZKEmtSrU1Ck
3NasAK1184aW48CwCCRAL5tru94xv7QrIJ7oxjSp+eIrI1JtoPS5wmB18lGxueGJfKAwub2Wcz6X
XfeDKJhgRWVssL6paRlY2Ks6TrthKayEOJASqlh/KoTWwMIWTLW3AsX9LXu70TDMatl03tUtXXBp
If4WwyS8ozkya5Q1DWm/rUVMxU5L+kx3vrmhkT18Bq0j6oO3p5+pMYHCazqbWbq8v8nkfPmrP6yw
OhF0EEsDtj93miT6soi3UpV4AxwR9eNyXSiU68FIgs6ChZGUypUHYT+OWl274fIXdNxcxoSmbdgC
W4lfud2A8UOMoQ8uLHZAKLKKWcgpAxGdH1tzHBFyhBHi6c8OVJTtl99H02JHnyiw27cdzsBEit9z
629X1ryeSszmmzNI6QpSiNbCg/uuL0GQXT2l4FvZTcBYquuPfVVKgCsyDJ9TSldBTJbvQ2pZrWUR
zSNDUYgLj5ZaIDrD0yq23ScSzQjuMARawLV7MCmEChxr83WYy/Prn4lPCWoELfgZ003oJ7HdF8Wu
00Y8Fn3VdjI5/qhFIr/KcKkVuSpeCGcrQz9BBQhLVP2H0FIUfMJJg+lQ9d8sZ+aixlWK/P44me6L
9CA6+Nx6u3kXXCb6H4D92uwTtzoRDGoAN0yrYvPgRuTbMjbJVyLsTtvsC2GauLsb/pKlsVZjzMam
4Wo2O7BeN1Tlxfz/Xys09ONkHh1O2KloFgJEEuzpZUJnbeEjuyz1fyqRTdsXZ9pGzNyDt6qlZwfs
NXpt28TtKPPA5qnE9oFlaua/3lCCNYPGVqcJ4bm62k7W+dzOKAZSBPXlZr5m5NKl3TWDWtJDV98Z
sEchdMwiq4TskjKXS/lBnQWexJRcVk0RB9orIbo7VYi5+T2ExpRvP6wr4XCM2L3BQWb57iV42PzN
vHH/i5iMYG9yYIWcZKDyHteB7nrunJJhTF/m8EBS3B7co1L2auUxYhaPcj/dmm1rN8ZGHiMVszhE
Zfs2prgHSK9uxjfhF7oroWcdq8bWatH1aUDFN2xBvjMUj61n/Qbqt7D2GVMzjL3fuY+tI6fkOprA
G5mxannaghjS+IzVTjChAoTE3u7fS3ryPpVEFNjKQiwDQnIXJjK+hIOXIRCL52tKV2W5JtE0W7re
hKXj8m9JJ/svNCMrZmqzt6EjYiMbprwVuLTOom+egJEfmT13m4L2XPSwIK754h+oL7NgXXPSkN0+
Zf5G9isgKcIzwXQ9hXj0RcaANJuc5/M0SwTeppu/sHVdTw2kGxZDplY7pr120HAn6u3gRtLJjBfe
AxHoVd6vtPKPs8eXcizXV4QSitFGz1pyGLRL2jYRfHyAbUwydsW9b39AUrAMPMhLgGZ4gcO9x2Qm
oTgtV6hPY5uHnW660l6Wl8XaK2rF7Qj+1KWaH/JB8g1a3ArO6p+FWt6JyR1gRuvlHZdkDBEb5h49
8rsygEFmPwYIs6Spqjww3ckW+OBNBSdFITCUJdx+5fcwjnVuoBa+CBBmxVgHu4ES0uRvozQoDZHG
cm7WFqyTMcLzkOgKwteFi1A//ANis9k9ZWboDpNFd6ZAbz6MPcmhasfwQIu6gScJmGi1LrG3Xhcd
a17YW1L2dIdMuc+EYBhBj8k12xoqiAYXcmRwcfCD0sfr7/rNchQw33XuWlWSyZC5nd+l+77MHwnI
r5WGPeWEl3OKlBRohST0qNj3fkiZsfxMlzLoUFfiCsvgswEYQPKJDcBlCeZJuwRFB2uXuD6nv998
aLo3yu323EjVYkue8OgK+1xv5YVabWnBWmwgAH0V3CvPjZb+skAqxAvG6jec7JSNpkGdNh4hZqak
fbPSfZ10kHjLnsjKM9iAUjZenhDkYhn8VtEZLwOXHTqibcTlNu40EjACuVMeAwER5oHwYvW53BPz
NLbTcuOq+1rUpDZsZqpXt2wf/xp3s1CmMoDD13YP1htC8Lg+kfBf3WSksv4HDI5bppbNRxKhT4hO
HDpzIY/Fl45WRxQET1qIdGR9MNDcvYJE9JdIuAE2CF+PdlaCMsNQbQO4Qj8aMANRou79dtQaHTHP
PqE4EQOOoKFPFIBtEJYoTZrQG15Vr2lkb2DNDY3QNSat5pKhIWOYcvmZRIoAqpeQ3pHEGVTTou3P
GQCkoDBhKXKOHZVJo9naFjXnOwkcj0S9WRHAsG8TAcviWGZStN44ta5VQpqe+Hezf/sEetjMBHXt
oZPTvp9cPbv2VIyqAdYORTMNq4Xpvn/GhowzAPQ5Kd3WyhwK1isMs79Y3O4IevW4lw2oMRtYaQU2
ng8eDxtzS4ITk4BNgrbuYNGnsDqP6XVOL/xF1eZH7W3tObbk/ms1+7LrutpIrEs3j2HmcW6nfjLA
cKxt/i4kvziAADdtGPawHs1P4CHiaDKjeFMf72nyCIm1MlWDIkJ7aA1oYOOei/uzPc1DnsHXMSr2
7u5IeADA0uFvHwce3uZHQMbzv7FAgdNNtQAH0beXiARuPjMS7Xq/xQh4K1McmY8CE8nKBEZnBrML
HUNOgUpADjSTahyePU4n21bpRcQNmVFeb6KtSZ7rxY4gi5SHlkuS66rMrl7KrfYvnhl8VucG825M
K4RCrZYi0tDEn/vImB+5MoX6wdxoQXDoY7k75C6MSWr3Kq0=
`protect end_protected
