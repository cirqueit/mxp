XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4��43n����<n�9�|~q��ֆ��������;a5�������x�S"VmU�k!�N�|f�.ytm�!�qG�P+*��m�b1`H���|(*NG�vy�����px�%,oi���m��lI������.��ʫ:pIFKJ*��t��aD1��7��/��E� �Y戍Y��?�ƭH�(�6��l+�Y�����}��8�
�wB�z�"f�*��d������M�	@n�5Y�5�,���?/J��z�wO�?��AX�Su�C�B�����~s"�L�䢆����ÐAap�}��s�Z~#݄��E[ԉX�F&�84NP�4��7�Tf��ݎ ��'lE��'!ع�x1O:j��.�^����r�����U�=3O��w٢�"�j��m��uI\�)-�'�9����,�j��hs��	�g��a���/y�D.�t�9����H��؁�c�/Y�^4�q�FMb{,jwGj�#+�Z_wDR?AZ�tw�4x��I�$-D�ʓ�Cz�O7�3Z�Ӕ+�oGi��rT{��W������+��2�9dG��u�.-��a��9�\gV�]A ����(����Tg��ǰgz˘U��2]�1?bB11[��`�.���n�^h�JĈ���U���Y��M,8�M����y2�;�e�?��L����KOYD�-R1�$Z��I�-"J�qB�3���
�o}�})�e���n3�c�-����%c�k�',�(����E'S���n]����U.XlxVHYEB     400     1d0��&K�ꉢ���c�"�ٖ��Z-�\��bm%M�/5�����3��_N+($v`����CH[�� PmUG�є�~�
�����zk��5��":�ȥ�M/�� 8Hg�	�- �&p�9��De�?b�3>��~�P���ȡ�H���k���(;c�{T('y�D~��Z*Q")��;��e��iB��z'�F0�<�_��ť����0�_�yY<①=&�Z����iy�����r�v0Ӕ `d����U�=��ii[�x��L�����E~�$����Y��E�)�N�9�LAF���vD�i�~ߙ�)� ��s� �L�3�$N��������}�R$
��e1��n��m��{_���I}��k
�,{�Q+�������b�����������f����$����".�Qj��V�ZR���oV�w����-BGWd0�X�񪜷��kXlxVHYEB     400     170��S*7�P����_������#݇҃
��t�ۮ�!/t��7V$ ��>��tPЫ0uE �E�w��i��t6������ ��q�{o�'h�tU������Sj�+�y&!4&��Ag�m"F��~�(�O)խ��PQ���V}t���[� �^*u��ၘm�N���9�>����,�UI���1F�}�X�y͚E����ᒋj����([s���\i.�D�T�Kֹ��yD�ZZ�Չl� 3*�Q���さ�A�'a��"V��]~K�!���̷ ׈����	�7���G�V�-i�K�0��k�Mu���ѝ,+x�W>���X��	����N���5���Z�ùXlxVHYEB     400     120�>$�r��L��V�Y�7 %R�I��D*~O�
�ȸ+Oc��JX��#��Z?/�s��Z@���׏��^�3���<�A�e�׶
':f ��Y(r�����V�� +��\�+ݸ�P���Q�W��'�qP���D$)���[n�\(d���;%#�0�uIh�q�gs
\����2�4G1G6I,�yE�45����#lY�?�PU}ت@��}^��	h����`U+�ÆV%H�|%kt]��X�I�z�E♦��]��1� �&�+��$H�e���X���.����X|rXlxVHYEB     400     170K3"$|=���7<A)!�����݊2�j�������t�I�a�6�~զ����/����񎑞X��V�DlT�ZY��U��\ק���C���Nm�"?
e��~=%PWr8SL�)\��'�?��|#)z<&e��}��ƬY��S�Kc��.vW�BLX���8���R±�<5�`��:0�tjŪ(`v�bd:|�S���w�p�c�����;������� Yv�t��=��,������G�q��>h�{��m���Dh-P��N.��_�w�Y�o��c�M�6�|�����EEv#ٗ�߁n5o�z!��t��_^�E� �LMտH!4s��yw��lL�(e�*A�;	���f��][e1XAXlxVHYEB     400     170>J:8}��;vB���[ű����fO���Xe�o��6�t�S��>̶Ċ�>?!�&+%�<o���l�N܍�i����v�Ga�?��}�3�Ɖ�� ���}_T��D��4%��5ά��M߭& ���E�X�m`�d�	2�n�x󏙈�����}t��@%%mΊ������;�آ܍tG�Ul�%�\�BG}c/��k?�'t�v�l�Gf�Xy3~q�ӊRj���J��z�m�� ��`�����2Q<V#$g�Ċ�\����*�*B	ʐ�����Y���O�&9XI�� Dp���>xo\Q2`���]OMN&�ݠ��2�k�6E)lx����ǹh�C$R�F���[�_ �"Co�XlxVHYEB     400     140b�(�p� ����(�������+�*U����C�f��U�Cu����/���Ly�M̖)��F�G��us�D/�(%.�E�tee�ף���Y�j�z��\N��c��>�k��z��Qd��ǯUyu��Ra�N��Z��;r�a�y	��'A&hMG��ޑ�J�b^L�(*�f��Z��6{,���Ey�o/&/��f`fz֯�=p䒁�G������l7�.w|�r�[X����Tx���C��a��%k�ީ.�m+�j'yw�..w�� �1'�K[�j�G͡!9n��O�	p����Ӛoy<b�\GL�
�e
WXlxVHYEB     400     100`��K�*J܎Nw�+ƭ~cf�^ZJ� s�ɳц���'H��
,���	�r���Q��|��b!U��O��� �*H(Y��#�G%��+Q9�W��tP�1$33H��\�B���~d�{�Y���cl���G|K<�KpAtn���M�4ܩ����Ƭid^x��W�R�㍍�"���QN�#,dCq額�����@�6�,%�����Q��z
x�~�/�E�l ��)�u*Ab�<�ex��:�)�>��yXlxVHYEB     400     170aV����Dڌ�l5
�u봮�a�F�+�3�������D]L*zT=Ff��h}�ʬ#�7��I���*_@վa�׆�l�% ���]90�xc@61��r�|��w�&���5HC��#���z[.2o�|�Iݕ�p�qܴ\d`v�?J��dC��v�HR$]��|��G��X>9�N�L-�C�
wm��}5�fq5ִz�������T�&�I��]�f�A��{�"-,�Z܇5kz�S�Ѻ�����׃VQ $>��D�*����zj#�w��X�!�m�0��a���?*j�����m����PB;I��F��֔dSZ�Bm�U���ι�,�3���smײ/���Z	P,�y���ǳ�;T�XlxVHYEB     400     1b0��UhM�"r���N\��G�%G�GA�{�q��t/�6?=a������(z9@�K����i�AJ� �EZ��i6�T��<����=?�,�l�C_��?�#�Dy˵�JM��y�
Rab�%����s8�k��.^K*(l62,L�lT1�c\K/��I�O�yi}Ȣ+��.��0�ʯ�{�{^������<�E~�4�Q�!"ź�u]5��
�J�t��$N�3��hB �S��[<��i(�8���c� ��ֻ����+e;/Ј�����_i�l9��XA�V1=�xZ��vx>�M0��U+��{�'�y��4�'�-Վ3(���oY��NFX��ʍ��Z~�%'ϸ �/,���.�k��0�/j�i��v����$�c*@o��X.���#Ve��%�Dcm@2��k'��E���ߥ����>�m�XlxVHYEB     400     160�W�$5}̹�S:��PbAk��@^��<W���Y� ��e���#!��N�e+�<^�/��Z��
��u��9W�P�h�,�����c;��芃��I�r��+������+�b;���T�+�O�	z\C� wC����]�XG��B��]���477A���c��DO�cWo�:#�"J3��	l�;=$<�3��a����v�G���u��К@��{��/�O��RD�
&B�u��t����7��N.��Ϸ�.��v�Tyg�V���o)��ǃ(	s����	����Iŉ_�#�ÃL�Δ��y�L���;YL�2ѴsY��_��o]�& U-�K+��QXlxVHYEB     400     1d0�& ���@�h�2�$5����x�+�X�&��-����#�NDNg?��R��j�-�$)��'��A18�C��ƿ0��=c���w�J�K��>H? >�jHW�*˘?a���6����Y�	��nDw�a�3�!��U�p��wG':��0�l�Rg-���>5=�>n��:��cje0R�oω*�\ǖ�0�7�w���*��~��|�Y�F+?9=�o��7����x�3v�������"~�u���ٽ�E�⤈��e��2;�U��:�z� V]t\f��mm9�Xm�@������<�r�$�!�G�@�{*t���2@�5��٣~b���̭֣upX1��d@��Eg��[^��#���J�����i�	jA���rhC�K���4�y+�W+Mr�,G(#��bF&<��[^"s����(L(8�yR{i���ev�S�R�,|[#\�p]!�
��XlxVHYEB     400     170�l:P��2�P�&��L_i����f��E��MmK_T=��ZUs��S��Q�d��͖i��>�����־kV�W���\/[4É~�Zܪ�A�u�NCK��D��y2�vq:!/?˸�&5t����q��@H\Q�]�	9#؉��(�ĹcJ|9o��G�߇��g��R�%��&h8j��MC��|�O�8�}���\��A@V�Z8�ob�L��,CB.6�mJI����Dz%��x���x��s��!��w!��ˆ8�=�1K;1U�N�,��/���W��������	�0�PD�k��F��y�.ם��],��1�����AOAr�l����ӏ����F��O ���`�n����Fz�'Z�z4XlxVHYEB     400     1604�����MT�|zXR�4�[u[�:J��Y r��9ؔ�na(k��$y�qf�p1
A��"����ďX�ݠ��3T��ͭ�AF�1���[B\B����;X�~.x4 [�X��w�z��ҍ�WAkb�Nz0�5��5?�н�?�_�k�Xzָ{
�M�o��,�a�O����7�>��wn�O*�}~�kw��F���2iH�od��x�x�S��鍣��R:��O�����й������!�����j�A�#���xM侚ڿl�+/�@��^�.��~ r->��czV,�SBQ���KK6$�܏!��G�)p�r���y�(Ÿ�LR�?��V�KG U�b̠���uXlxVHYEB     400     180M���gs*�Teu 8�W}3q[��_�B���rF1"�nȫBa�����tA�ި$w����g�&�� ���K+E:�ӥ�`&�����b�������n��Y����E����i݋s�j���|kq*�׃PG� �n�Y~�>�C�@�4�%���r�.AD	�*-�����H:�֋h�=��D��Q�2�%����(G��Pc쪂T~w�礅��3\�$ (b�m�����n��H�p���T��z�B?��MH��N����E�q��o0Gh���Y¢�=��뙕�2lf�.�(B�!aYۣ�� ���~
�L|�Ǎ�_D�Ӣ�C"e<�M�`�u�l�P�{Ⱥ�#b�|f�߫�Yq���]�L��q��e;K'XlxVHYEB     400     130(&������o����� R��y�������<WF�=;��@�AE,g�x-B�<ơrj-:�%���B	vR�����ӎiE�����:`���x{\��V8��ۀ+���T���e��B_�
��m��`���0�9�dl�e�H�{�5���ll�0e%�2b)���O
��x��� 8����)�'@mo��e�0f$U��w���rz�w�g5�c,h
[��u���b6Q�z-��4{*e�
�^�7%z���b���k���q88N���������@��-W>Ǔf�C��}N����(���i�~��XlxVHYEB     400     1609/������cPk���mQ:��p&`����w��8�ͬFk5.u"����t+7���.�I@sJ�Q��4f���®2��zaxs�VZ��ʌZ|l�}� �����J�SW�v\�U���JF}��ǸTf� uTR����yѧDE� [D(��:�8&�N�ɒ����!k�
��:ivL.�cI,�|h	S@���	�R�R����� �"�^$C��	P9�*���e�M�t���L��I(�NJ����_s��b!N�A%j�A{���h���6Y� ���Qi4&��8��4�r�4d���������
V�ڋ5�te��E��l��0�k���?w~��uR{a�:)XlxVHYEB     287     130^Q�Muo]Œ^���1=%S�����\׀���j�d���E��(����^��*�~r����*e���̦����!D�I��J���v�	�YAx"���:ڋ�W�?ӄ$���B����V-�Q�7���h�X�	t�N��d��C�^���&T��SW�,yܦ��cQ"�~bDLٛ��.��*���9�d6"�~�bf��@".���x�F����*C��v6�)�,^5��_�}�
��>#�w��t$.J<iͱ��U���/���>�G�P�3�g#��f�/Q�~m�F����d��HGi.