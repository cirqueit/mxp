XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%Q֯�K�u����I��M	�ύY�8���{%���仧�{(���9FO28-�~�χ��'��a�T���豣-;��&��F��N��b����k���(*�O�S��>Jd��
�C8�
RO�Ȅ8���e)�C�7<T:0{ڠZV��TֽKg7���UXr"qgߙ�4}J�I�t_7C6�����tm0෩��c���M�!í)G;���'H�XE?79"�pv��'��߯*���c�Q��_�;^��C�<A1�jͿ��w>o��niD+��\Q݊;�x�a���(pn���
�L�4�r`b����?L� �&����y�tB�=p}�;����N�����g3��'g�՜��bu�?��������H��Et���6�D�� ��Th�o
�8��M��t}8����]�D=˷���T�B�\z�-&Z�o�Q#��-��s���/�������� ��{8I�W��� |��9����*NDw`�|��7�um�ޯ�w��~�fA��l��Q�5F������ţ�.2��/����{k��D�4�͛2�ee6�ֆ�H�oc�Uw� #���
DSkU��������l*����#�-�O"�ߣ���TyV�=�(XW�@	]�GF�s}s�2�y��@�jўר�ID>ϳ��@	��0F�\�)���b�%���hH��(x�)���	8r�g�`b�u���j%0�c��0�b��h-׸z�J����D�CXH���`D�Y�/M#�u���I�nc�eX^XlxVHYEB     400     150����6��"zl?�I1����E1K�7k��I/���05���W�H9Û�v.K:��Q�A�} ����@&���S��R��x�`U�4M�8�����}�pQ�����mԿ	���V����ʟ*<Ҧ���Ǘ��0��˗c��Y$��j��F�A�2�8�49�pC3k}����ҵK�2���2���"[��)���E�8�V'�	B��U�ZC�-�6�#T��+>����u0�u�0�[#�<�~�7��4D��y��%���9���"B������/�U��n9;����;	���9���O b�T�g���]KF�FʊYz���xg�]XlxVHYEB     400     1705B?�ԛ���9iR��q�R�q�osAqF��A������<�*j`[}��/�r'���#X�Hŏ/������h�C�ѳ��$�tvӟ!t�7��U������-O/�Wa�� ���0��6(Z63r9��n %ј������>�`���+�Qs��� d�cfҜ֮7ơ�p�x5us�	W�KL�<vK��~q0Q��U�N�\�*�
P���#��7�?Xu�'��ڞ���NVj*�gF-쬜�W�#Z����b��O˃�Ý+�?�QWě;����-��������숖Β�b+�K�3���`M��
��)�Gl;s�������Ҁ&�ϴ�}��cR�Z?U����XlxVHYEB     400     1305�o���{�`�Q�=pe�K�9N�v[4H!��r��4�`U����0&��y�<��++V����T7��s�Q���6�;�D�N�Ӑm�j�������� gzz-��3��"�!"7�\N*��
�R�]�{�7E�u��`SgUV&T����V[�}�%ɵ������f}���e���k�C�M�n[�zi2|C��q���#�q��W�\�ž���!���'��|�_�749ALA�� Q���Z��#�G{m���\�1����j|d��XT�����S��[Cy��*�\XlxVHYEB     400     100v7'3t�g�&�����&4��Q�<�'u�b��I_�tib0�,n�ȋ��
[��Xu�P��+�ԍ=(����ԁI�����漟Y�1}D������CBv��b�a9�v��N����X_[A����Jx�~�[a��mp�=u�uZ	ş��[��[�-� e\�,/#h�}D��@7��>Anj������*F)F�PH���j��PofL�݈l���eQ,Z�oE�	�=�2�7�%uX��O�T��	XlxVHYEB     400      e0�nd.�����pT�������Ņ�p|�'��_��\6�`d�ߔ;`?"/�����������O�9��┐<h�9�#�]�jd�/ b�=�4sn�9'��J+z�|kA)-����.�9���3)�~������s#��c�8���N]��G�W7�`�A��R����'�=��^N�RSPvO���@�s
��#aB�M~�3��	�;�#�,�A�XlxVHYEB     400      d0�rPe� pi���R�Q���=V�t�������?%�U�����:�j=&��1��N}ZIe�Պ�R&���� ��؂��o<�@�jv�P�j�=Ol�&J�(�3	���u��������\�<�������}����1*`p���x��w�W�;��6ћ#s����ɺ���2��\O������ȣBM�ʑB�$�R;�Dj�o�8�`XlxVHYEB     400     120B��Wa�s@�uFqdM7�7ņX�~�	���ڨ��?��Fb��p_�k	�R��h3r���Q���=���Q���&��\�,��}�0W(���;Y�R5"�����r"Fg*o�19	��B!���j�A����~�08$ �^��_4�y�ӕW;�c�U���hV����=�>�٥�e�K��&�~�r$�>�φ2�.��i��X~��K<��* �-�Ӟ����G]��Fޭo;ղ��?,?�ǣ�!yת+�Z@���Uc<�T\c��d�sO�aV�=��n�XlxVHYEB     400     180�P��B����i�<�����X�,�sb�	߹5�Av���v\���Ȏe%�a[+��1M��֔��O�a檠u��P��� �P�m���U�U%�r��ԴO��_�w�޿9$�:7����`֗[M���O�6�g+P��
����seo�11Q���T=��=/~�N�K����:��6x��z�(ț�]j	y!l Z�c��ͪ�`��Q'����xXʴ�~*h�KsV�w��G7��"th��iu#��8L���M�Zzd^��6C�<f41ՌL�ƅ�O�u����q������0[�"�W�him�-�1���+�$g�F\��ȸ舢��hV��e��@ 5���A�c4�K(�	�$XlxVHYEB     400     140I"���Ѣ�D�js�Iz����:b��=��d0^�I��:�	&iXk������ڰ~6�YG��4��&��"�kfw�EV���{_bu�N�ufȳ�UY�۸� �]j����S{��TK����_�:��k�h5�r�sRP�?a�ɔ|e6���/�h�T��h�"�|Ѳ�*��^�A��f�+L�+����xHOj��$ۜ�U)@�k^<�h��>��F��ٲ�(�ʚ�	�����Xc����|�AEs,8�@�JA��r��*�6�a��'�'K�h3��'~��ǀ��0��B��v�L�v"�P�M�-XlxVHYEB     400     170`a��yz�C�	8���g����,��bJ�*��k��]��ګ"@��
+����|�~�� _�c��e��炏#��U�(���&:)���s��O�ar�;kx)J�uR�"|����p��'��ښ��������{B�c�M��>u������r, H�v���7L%۩'�����D�J:$�U�+4��Z��&$B��{@�]5���d��� JE��:�L��]<}�o�\�Ռ�V_��b�E�e� �0�X)Vs�ٍ�$;������,��>�5����� w�\b�FV�ϰ�?'�w����CrzH�y$U@�`�����<cZ�R��mfb���feA�����-5DG�C���/���hLix�&JXlxVHYEB     170      d0sa-N����h�.~^Ԙ�.���J-H�k�|t�<��L#�t�9��������h�4a���Vz��e�'���/<������q�do�`�2�w���%����Yg�?�W���5#fݯ�<w�5<t�r�f�;�<O+�7�iO1>X]���zL�UΣ�����A�UbsQ}
̴ek�@#?7'X����	���VG�WO1�σm"�