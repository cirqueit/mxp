`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4176)
`protect data_block
xX7nPnoite0fUOxyondXIUtYC8/QpjgBsQ1965navbzLUmei53KXbZbtyklMArNITCmMnwuXlTl6
G2Is/K4kwt35fdkO+0QMRI6rhECo2Fvgc4ckFTfjSGN8w3NbakL3oPPrXct7y4lgCIPmsFpZlwNA
129kp2EbnIEI/VzIFXPJWC+B3SyhX8QwU+g88R0IeH/TSpjkfU4Us1PoSjfhSsB0GqtHRn2InDne
3TgoCp9iCiY7+9d7GAu/icnzR9LXS8oDDPK+vtWHtbo9R4ZRCreUkmX4OXrdYJSUv5/nRqafQGJp
KVRbHSi79mjlSZFiIi1y6OANJPuLS39ZRLMe+iRiEm/ij7QF5yPY/YEtMEBAZjsn0te9Xy69MP8Q
CjFUuU/ls2dbUGP0h2kB+Y0qIVKf7OWgE6oI/sLKKgYCgIigNwvIioTnAvvY0LNPoFhut7IBy086
ErB5JyWTLutBSAUyBriGCqp219Kyqx7EVqL+KlnkFFcun1zuv96ywdkHcpVrsawSck4TOBmEYlZA
KaXIq2yzqJ62KgpM7xTXA796xkRlSGYFdl6xE55YnTqst/5lS/09MrepwP1vSW4XN1yREu4JjH9i
0mA6Mwn27Js0jSVHNfMDmODJqU+f8XRKLChddQQXdg5sHO9BO0N9bn6go+RHe2ObFZCL4Hn+UgA7
SSGUe+oOPkGlBS1vi2SHlrcJMbyAxqIpSGbviaTnyC+8XGBQB6iDPY38jTUQdO2eVn6m2kNJAu8B
c1w/nnY6zqvxV8FdTVqIJu0g0HRHkoQJWT01TB0QurUVjx5y3AUoWamnwQHCTMNTdf5I27V3aiNK
T/QnFq1rJlM5B5pMuqhrqVFw2hrx04KTsv1cIQ2t06IgvvgafcEtECF8dQGwhvJaJE9BhbSh9DzX
n9pZuAXE3a5trQK4ddpceyPLkzRJnvM81vU/aKODzL3GhCNmRsZIV9K76XkMFuw6Rb7pEUlbgep1
zy+7EjU0X/IOoOeBvRMfYlPYeKRLddxvGFwKM5Dx8uhy7sEExiQAeIpEqpGVq4xKuuCjwd5NTq4l
ubE5JbE9ywEIfkp6pRinPaBRPUNVjnM3OY6aSeqxWD71M+NG5LAONeSQ8/XJHR0e5SdRD8+YMVm8
Uornb2C4GBZxHyPil7LVvWqdSJSQSwuGZlKdYvUr9r9HRvtaW7fzn2HFTssVGhRzsLs9+sTeyKI6
KCrV0StKbOwM0/itcxAIZO4axdoR4wCcvJExYMGg+7aBSvtnIUO04zpys/0eWphwA8TnPdPCTs2k
oOxECCtyjtFIaZ9JxfWrfrQiTcjnm6p9xXq5rVNsJdDXFUbDNagrz+oPXZyxf9Z0PVCM/UXI8c+S
t0RkKjnOT2jgZb+kCI1/p2gYOKW0TCpZpKdmm9LpIaHfXg1T2l6MlZeje5MthXC2fi/W6GXASKdM
rXyiWPeJM9+6kFH9pnwKFFMwqhK8MDpTzYsQhBMvFHMPIYjEf1womfzKyq7ByT3jUH5CXzgZ7Ghw
cyyS4LZSWaTxML/AjxCuXlaZ+weAQyz6Xiv7Zk2BShl2bC5SZVHFINFJA1V6hCUR2qvGMjU64+o/
1v5hXeFuw4JiTfisLl2BjalfsGSeLHgTYdHlVwvu/ZKPRWR0DwW2Sw7Ivtm5v5ZdHh+kg6Z9M9Ez
FMcuay0Fs+zw8zQmQtxj9WGsi/BmXqPBnzboTRND5G4LMNo5lEckmuoovF3nIY8Tx5Sfxndb8Qcz
RxIdkJKaAntr9QlMlYrQR5Y1Jnl1LZI3/s4vLw47Zg2Mdwj4rOsaJnvMkdw3te599FDP0RdpUiLd
Gwuqls5x82ZyGsNYOE9ygJR+sB1OIYZnDV12SB7gerOxMb+7RF3IMzNO9BN3L/pD07eBzvcT6gQ4
4Ej2uXcwTHaATEAxvUcBc8ZNc0yofTYBHPU5tHHrCGxprf15HWjAluwGErMXhs6zJkgZcsukoUw2
it6Pg4Kq8eZ0YwZxNsetUs1QL0hJfos13h9JPtQp/tp7iOdpfIq8Frt+3ebB0x19gZYAeddZTCVK
7AWWbfSbL4VNBhNV5hmJNTUl6/jU1RgZkQH0iP869aSnFiCftelTS30ZuvcPm+xFz6NL0ljV+g4G
1sdSRSqCKOyQlnA36cpoP4SrPjhEvFHWMdxo7fvsarpAealR5AiPAgSugBeG8wGoPKjxQGGjOCVn
aBw+p2VKu0KdrcAFq9lKx1xNCl/A/Ys7b71TiXFxNIcZUL/xfO/zEpFMrScXArcALdvxS5A0boqN
S7f2P50LkeED8IGYYLtd0FfldMMLUX18SPD1uA0LTDpWCUqGIImx21cKJR/Hm4vnNtHYQZzKm1gc
Qe7fMw8sAgyo3XUODDnfJx8ncAPwXO76miLIgf4pV5ZuNZd/WvYMxB679DXqCGpU5VMYBbZ5d9fZ
NjEAFtvcXXq8Aqh3huf0uqWN0hS9bNQzM+5FgsBKkcpf6Q+K3BgMxcajP7FZN4TZP+00WcYuac+k
mvWExJ5bu4XNiD7g0pfbr2t+AFxPyT+RdFwETX1BX8DB6ZI/oUN0EQUygLcSHo1ZpBZfi4HYdSfo
vNSWfb6HrwHkOxv5pWsojqr8opUp4TFwsLV1rNrgWqq3hTG4enFfDrPJaONR0I+bUAZbuSUsNWg/
hcPM4Nien0M/4j5aHL03SMbIKQJV+QAc9xFtXu0qt/YsI4LLl8PWAKs0mL6ddblIgdJq72nwaCEo
rsVMrsBatvvLAZXF+29mE2ahIDZFWSMOBw8fiM8RJ1ZnubLzTL3zvdFhRMMkW0p40TUF7tawrx84
o6BzwKpM13vmzOIR/AO1dnS3wJR0vctbEY2Im6f83wQ4xlyKTeqI36RIi5QAaoRDJxodXZfngIL7
aLl9BY4Dy18LP4xeVPcpHueWFhbIe5EOu4cNo0xDiR+CCjY0zr7FPHS7h41IlqKG508ew+rhbjJs
p8qhEVG7brrngXgkJTWQnXbLSofJ3bQh5e1dPFukyCa/kWJoNsepzVdaSsdCnLveNHGQsAICadRO
l4AKOpg6LCa1zXs7ZukT8AzKv1nCK9eD21aOB//7dRiVU/ZUOZ8/AOu+8lCj3W9wblfTxFB0/U9k
2dAQU32OgAcaqKz6X690/reCENZJSQh8i7+Bhf3sZ97tQTqmpIixKsjMtHQXuSrMNL/MYBsGdUXw
o48simAq1oz+ZpRQ+OSGLJoZy9r0f3zH4u4e9fDsebK3CCpN3GWv4KkdT6cpDVIUbe2Xt0NbWWqu
PLPaal/H1vB62ndCuN1xjHRmUbSInKYginFRGWpJ13KmhNDrXB7fIMozIzs9kSnjCqd79e3HGgv/
OROhJsCXnGPXc6AXv6ss80yv8CdEJdQaImaQCy4IZzi5qpQsAMDEQ3zUrOSJGTrpKNiJOIbuCZSa
A3s1GnANDBErqT6rnaz6RAC5hy/bJFIqfuP85vT4Epg0Qa3DY0kIjhoelJJK5Ra9hzitlVejXoQh
KZv+BUp7o7fP3Jn/Bl5CCTk54LxHvX0w0W+aZEgHSODo5oFb8P3VVn8GOx9KCzsgXL21n5kSuGKE
XkUJn+M5VtpVtx71FLDOrxt68B+EUGJcXOucX97SOgprcFNHuwS0CafWKAMbEwpB1XPQYREjDtlT
/OskrefRneCIPz6aRAIU5g6/p1/suwPLTBshRtCHtVHOnMbbO/lX4lf9rie6XYKAFK9m7cdmorod
uUb0O0AG/xtHp6GfpQgDKrRXzgWnb3SxNUtydPzxnQCGzTKQvJj11BXdI5owvrfMW8oSubx/X94x
mhmEl7pzZ8gYl6vMI+VHVd0k8j8ZAd2oJEIpmjV4m0j6o+ue14tM5XHWOW6IH8cE6G30rgWKQxbt
ibcwKqZcdz7JmYT1IP84Yoi10yOSrsgP55u7HUhtppcXaaKqVBFW38iN8ftKA3MY1GIF/wCK193P
BQBDbea60kAOm5Hp0huiv4aVKfSOYql3YYHHjbXSLTIk7yJ3rNhJ3csIGOdklr1O6F3Zr4mLxdoX
bdMUGM59BEQ+jX7yA6yf3rdJ8m3PygCLWdtSNhQ+gLl0RfSWpsMY6uL+aGbz2RdvGPc5GW2ABG+E
rRrn1IQeR/jeBL6DEHwevMTjpQZvseVj9vwQlOBDXE6wcvP8pUyzBTRoF0MDXmnrKM1b+F0RgyXP
DV1GyR7p9QxYZ4xM6Sz2eOF0NCh7Gw7mqFxdb+VHwaXSkFaVXhGeqMSH9fZEV8oFCDwm0MLYm70r
vInygZh85P7eL5KGFmFqAdHpOWr2U6F9Ym4TdZIdXxh8RZp6q9rI5bt8gqhxBiDg0F4+yzIvYxDX
SveBqZeOH+9wQdrYfh5l0Dv+EzwHVBx/BBmwkFj0w5N7P+js74D5w/DZPBa4Az7Qg2+kVRivU/DA
56FOzK5bMu2PiyQv645m+9HJYq4koY/eWIFWlAhtfcO+d4QpzmcQBhYegMXaBQh9uH3WAOILtJZF
qiTAx9e8TsH0ylJls+jEUopQ3SMPLE63k+ke7famAcSnLeGYe5nBCjdiX1dFrQFB5ElIaJynJ0vL
ilmmwQ6IbKofPwZTjYrS7tt0MFm2bjR2CQ7fJ2Yl8Y9XaFqqK+uMT45u11k833dykbsYqg6gC2y8
FxNIJfGkU5qEFxxJrBijuHk/CpmGvPEkuG/lfRIN42CW+FUVDHVyUzM7KkuECuSeOQbzzGdZkXyB
fG3o8uPgN7KPtIFP8o8XjHdDKKTT5blpu31apUClRYqRPZ1CNb8zg8OQATP1KYfqFgPdiusu0u9n
HkdiGpq0POL4IBWrZzXM6mck/GaDG3MHJ9ImuocKnCVgadf3cP9m5cP6U7nq1GTb8Cr1x6+1woou
K6nO5bXVo2uka2x9LQWWEcfg3HJxRgiA9cnr3y4l0eXALzwtTruhX6rhYqgl396gGJoGtdB2e3qe
ky7jWb1wre0M+xJDoTsnNoWC1cT631RUnYnwLxU5LTG9pjbzjySKSBwDtvlpSdFA5EOe3kQxMNIu
+gd1ZAR6q+7152snjE9R+lSluG5drsrt3jeNn/mld0fXp1eICHXWZdHFrIp8Jfo4LyI44R1kJP7h
0TEzpBKnDkoHN7DxYuqSW1kxBMM1mgfZiXOTaHIlFXvxkgq9JCBABy3hS39LLTZmycpVN/oAuLGD
aND2EWXJuaLOwOQSo37Hg5AhLTUrjv+nRWaWYIJhCcFsDMeM+o/CMcptluHxG6O7SbIud5xpjmE3
CglZ7XmYnBwfmFUYHEKJLuYXt5rZnmj4t1L3a0yJfR8ICJvrr6Ao276tEUMrTW/MXHoTDgjp1r/A
2GUTPwTY/qNvV/UwgX3CQiryc1SI07pTDyM+ef0HQS96cfrGQ5c5XrG9a93anMrFwKdGLX6TTNV9
QPi0xWKMnftKNeZlJukwrSbr1Lz81isH6909WGRFCjSzWLgIUGf/bvIZ/KYaht6numboQT4HCFGf
236p9kyuDOlc+ryGegVAYetdcVqmYqTnuc1mtPRZvTe9Nv1R4Z1qzl8mdxjk2KkXeoT/0dCbUQex
Vk5rDKLClRlQE2KcEorz
`protect end_protected
