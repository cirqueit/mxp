XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��dB9�6Wg��#�2uyd>��B��yv�do�	�W0�����F�ղ�����E���z`d�XF+p��$���+����r��^!^�6BJ��wmq�0S�\Bq(�6��Pw����T3N^pu�p�#�~�����F���<���/"ja44�Q�t�2��F�\&��v�:� ��g���Z�}����Xf��M����m�e�='	j<̮�ԝ_�j��a�:K�H{v�(�H�(!�����dy7|5~� ]
+�֙��14D�9/�0G4�Uh������]�q,�j�i"���V��aU&�i�ߍ��IG�
�T]�����������6��dI}M{�"��2�_����<g��f٧�͈�mi?������H��o�� B�k���MtU�#x����S��,:;A}�����5r�-e@��	��e�#V�b`�k��t(�ՙԖ��R�70$�$n-��e�0�(Y�ƞ���{����4Q��.�M�w�z�T	|3D��0B�sq���`D��v�i���"����ǁI�H��Is�w��7��k`֎���՚�t�O:��)�0��K�>']|L
h& �?�.��MV.lܻ��c���I4g���]iJG(�%$�~���N�f�
���zx�p�ҽX��Q�e~�u.��|WE��׿��İ7̗/��C�ժ� +Ģ�$�-��+%�����̑c�����b��c�ݰ�v�sP���^�X�R��5!��Ӎn��>O[DJ��*4
��XlxVHYEB     400     230�X�ڗ1+sv'@|�|�c1u��C��R���p�Ś'D��[=},��.���4x��k7_�9��6�݅�n,��W͜��B���5�`}Z��Z��g�)&�1{�i�~�������9:,�T�Pv��p[
��9�@����Β�Ѫ����^,�S��k_E�6�t���E���]</��6:L��:�I�k���٧��L��/F����C*~��������X`��,19�t��8�HT�.���E��X��T\N���4�Y��>���u���}r!'�d�Z��`�L�P-@~O���[`78"��a�aT�j�=f���3s�5.��Ά��^�V���ä��o����wC��t�q�`
����9��I�����Z8�R>���7oUzI�5�L�����L�F��X+ʚbiyd�Z�񄈥*-��i�J��r�p=g\&��g䍓�B�~��q9�"`�l`�Ā�J�q뗶�(�?��Rs�,��_SkG�.2gBK���&��͑�^1g%�i�w���&_M����J��O惙��C� 3TXlxVHYEB     400     1f0�>?�����D!fgꍘ>`ZWB!/�C
��P^���էjxep��/��\FM��r&�WO�*|E;C�s�}I�JJ�20}RU	�����ܛ��C���T��&��i�d�`�T��h��t�*"�O��&�y+�2{N��j�DY��x�i7-����h�	�aB�;�?h��;�]S�i�����߯@�h�-@ҧ@���$���BI:<l`z���d/�(���xS��HSq���ľ�uu����EMv1����Z@��i�H������		#u-�͚!o\�?�o��+�l�u���C��iT(�k�
ԣn;�]�R�Txzz#���
[�BR�v�E{۽;ِ"�t�j� ��;d�'��kҖ~T��&R(����`Dv���_p�)�ԙ���|1����4��K��֠;�p�jd�蠻w2;K�/*m벹�^��ƞh��jE��8q�J!�E1Ǌ��];*�8б����P��$a'�j.�XlxVHYEB     400     1b0A�����$f �Xɐtp���A(�<�c�0U����Bo����v�q�W���Q4/>�b���:��� ���l�7)x���}�M��<��oW�3)}0ܟ=�k[a�2��eHD�^��p�\����O�D$�qd��Qz�)+d[����wa|��Q�uI��&|8$yG�|��5H%9���+^��iY+n�э�g�H'��O�!�N���x��a|���f`^Ug�Ѕ�񒸒��Ŧ�W��6�� ��I�D6��4ICP! df~S�^:�8%m>�zy�Ņn�/x�cT� ������Eě��勩j�f�^q�J��-d��ک]�o����9�PQ�F��?f_G�9eΥ�V��[<��'F�ܖ{�Ʈ]>_�X.�#�W�����L�_`$���\lv�A$UG��~XlxVHYEB     186      b00,���c�4_�-@��|ٞ%��0���	&q��0�A�3�7N��U�oi�p�ö�uc�B��с6-�T��Yvv�6��H�XK��Za�O=�_u����b�E
�i$�-C��J����`���#,G�g�2��#_�إ��Le�r�����~ew�ﲨ�.��̜���!k�pmhBFn�cKLZ�