��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���v�d���G�d/3��a��3�^0�U���薆2�Lm�a��Q#O�Zc��Uw�_�?��u
�����v��j��IaT�*��i���չ��O
�G��x�O�N���|!����j�)��,�d	�����c����Ds��dR�}�*ln<�L���p���EQ5�d�V�uY��+��dI��j;X3h�5�R9]gw��~�]�|J���b=�V}�;fo<*�����&��r�*PU�y��J��"ΣZ�Ǥ�_��0�N���ЯB��B��r�w�)Uߤ���:Mx��T��g�L��{����%��!-b���.����C[.�Pm�<WF���š��{�;�r��xT=v�����fюh�t��e�)���t8c`�M��=b	s�N���d��o���y=��en/5.Ae4ǐA�ТK�Yv{�Z@#��.�t�T�z�u��,�*�P��%�$�T�bI_7r��W��C�3*��,��1���]�_�n�~����v�4O�xڼ�ך�b�Y�w���}�9 [����������֘�6/8,�`:�7XJ�~<
`��	��&ɑ�H�Z���(L	N��^�PQHcjrk�E�z�ʿn&�T���3t��6-
5�KƱ���ܽhڸ}�a��|!�Y�ƵP��#3�=�Mr��<K_�x����K{Y6�o�y�ݴ|/�V��ٌ��9`�Uҷ���!��2�T����O~�@����U�����\hp 7������M��Ϊ�E>����DE�4t^�Kך���k^��+��TE)b,�0�|��^5
>p�a�u���x��#Ļ��#��FԴn��
2�����?|�8�zGp�k�`��Nk8�1��?�!F�c������ca���A���橊��!�Cd�I��x��f�:�n�ǀ��0�T��I�,D���Ց��8ݒ�_d��Y�J�'4aߝ�q�.�/g!��I$�� +����ƒ_"�Yr��K����9T��t[7�r�z����w��u�9p~�b�ߴv����^��I��x�O��>}�gE�;��G�*f��qՈ2Nt�SSxY%<Ӳ����%dZk[X[�oC�dS�?��u��(�_��y��4ā�N��
s�r���q��p��G�/��d(L�[��KV5�sĮ8�2�~J�׿�>�KJX���g�i�yD�_��8�z9ף�̓��c����3��F-'ҟ�PU�*dS4�*G��?`_�2~Կ.80�w��h^E��y����g��F����/�$!�D"��u��E�)��C�G*J���'��Q"o����;�2��u�6��2��w��ę/��z��<���p#���l�є�r"��Uv���Q펆q��M���^y�\J4�B��"'9��<h_3d!�~�p��V� �{�L��
�E'�)�Wۜw� e����s����+�+��N��v?��G���rY��Ӗ�E��)��N���:�����xP�b|�Dr�������P�"�f	t�>�KlS/���v��;V���%f�̋6�\XCө�JUk��	��1I�#&��\�U�a8�����Ʉ3��7�o�H:��汧{��vWw�K�M��^�V�����ۭ�s_��(E������k����_��"O)Mľ:��_����<y堾����=io��z8ep� -p�����e�֏9T�&U�*z@����l����Eu��uu�)F2�������N#d�8�H�Y��o��*�Ҡ�Q0 $e,�'\s��S#�#|�F�����Z_̎�v�s��"�W�TV)��jX���(��B��:e�:�2)\����2��N3��˯�P%�D���wb���?O��OZ?��+���fʸ};���!(Tv|i*k�}.�<x��+���@ܳ&�[eg|h[�V�e ��C���4���y����5�*lȓ"W�ⓢW:�����?��U�S|'R��a�Ftm(,��;�ы�)�6� �|/�Z�rrZ�B���#qB ?�\j~�g�a{��Gۏ=<��w�M��}�4��L�x�ȏi!����/�7�j B����a�F1�o��B�^$��Qpzgݤ ��ft/.�+u-�W�ۉ̏PU�̥�r5���Z�,J,����c��T��<���Hm�����������8O	��S��(=�V>�%7�&��.�F3�!Ϧ�ؿ쫱��2���zJ�/ހi���Qbqz���%mj��ȇ~�m� {�وG��5�vk7��:O�V���k��Z	���}�&����؅�c~�� �1wd&�1Q=W�~=���s�.��I8�m�Y�� ��{�Э�����J!����(�bݨ�5�+���*<�_"Oߑ)/���W�����de��0�Ѽ�P�x��ڦ�L\D�#Z_R
�����&��d=���r\�{Y@������D:�%�{��YJDA ��{m�,ҒN@W	6ef�y�)Ϻ3M�1e��s0}��$�(����xW�H:YS�h�*I��$~�SÂ�6���* ����M-4L{mg����'��E�A�jq� 8��_M��Gs�Ɋ��!��!��,΀�rl5q**�g����5@�f�;��,p��y���w2�X�`�6b{���r�j�l�.p�~�S�F�L>v��21��Qti�u�������38آ�0���ڀ�ɓz���}�i0
�ϼ�p�*ƀ��`TH�eM*�[J�]�n�B�������G�[���E?4��b��̀�R�b���)�|�4���X��
*�^��e݋��l�ߦ����>��2��|��U���޲Z� �O�LP�0��eƭ��}��%�*e�+���@�:�ǡ�3$9��L�I��)h��]<����=��n�7��U�U����/w2T�+<����H�����^��Q�W���h����� @�����a#r��u�Ln��%� }g�~mQ��8^��hBe���ˆ�	�ʏ5��/���]˟Xfr�C��ܑv�l6�5�֪�Q_gY�/%� $Kػ�5syN�N4_�ˑf���c��o�WM��&�G������'V!�JS�f)1�]�_�%�kV�P?�5?Ji���
�j�)|��\�\�z%<s����*�vFQG�G�/X���޴.한4%?��Z�f���L>x�A�L�G��w�k�5��X��\fBU��8d̨�G�%X�C�g|k�$���]`s^`^^�� �pz�4��� *yI6
�
�v�)��_��*|��SB��؈�D����3��d��E�����V�S��yrMK5<t���?��B�m�b��odl��4YfL`��M�l���1����{�h�S}�f۝!�Wz0��S�*Ӡ��;`�r�o5v�qtg��A�z���T&�m�1�P����GGr/���2P�컖��댊�[�k8'��5�Ѡ��ʆ�;U6�D��'s��(@eKq�$��ů��k�vQC��y��o��,�l@�nv��S�9��ccڂ~e�%?W;�
"U�M���y��4R����r�[
�g/l-���A�T�*P����Ɨu��;�U�],bd�	t0�jCV$ȋ��P�U����~�ߦ�{^1�i]�+�-9^3�n�Q٘�o����"� 1ͅ�L@�ߐ�[m��`ө���Y"Z:,H����?k���j��n�m��)wF��雈�V��q
B-���v	�Tߎ�<LDL�	�e��t9�s�O&�8h?!g*�\[��р�q����%g�+�E$�����|>�v0s��{����(�rS� �蠠%[�wҭ7s��*&��q>ث�O� �~z�?M��y'P�ڶs���^��3q�����XDD�$󧼹Ӕx�`(�~�m��g�hl��_�I|����lYg�]̮�ʚ:�{��ɻ4��_�觺�˸/�(ϼ0SQ	$?7e��_8K�O�{�`�]_�y�G�!a��p �
@7��3C�4l�EJ��PK&���N=H.��28�>�m��5�:#�4utVd0Q��������)����p�,�Ƴ��G
iI��F�ꀃH�'p�iq�5�B���3�B<��6� '6��Vy��ݱ��.��`1��|:�K�U��z�4��pw����+�Zx%/o�e�~Y��i��Q�ШV䖮@&3���#cI���l�� �\��b�p<v����)q5�����������ZҦo�u�wk��{��ȷb��nb�a:�����*w���}H*G5�s��W
=�㎨q�2��s�)es{��}�Ϙ"4JՍ@j ~iA)F����*�)��pk�q��d�}W���\:�.�p����;�����yU�'c���Z�z�dP�e�鍪v�e���ٹ]�\ÖF��l"@�M��a���P1Z�{?F��6ڝh���Be�K>�t0����0�4?���0p��w�s��y㧼�Z�)h���׬�G��{�@���<�����m�v����u��e?���l _�W6TP��o6��;fW�J'�@�q峞]C�T����rt>�;�>X���l60~m`���HM;�l��{:\'j�[���#���v�F�a��"�|�j,N^r�Xb3��J�&�@㧾�z)3I�i�Ⱦ^�~����gx�ϮJ"���+��D�"�*�>�;gˉv�S��aꓵ�q��Ss8��!�����-���9*�"��3a�����!�'��yab鋋���i_ q��xz:ē=0Ȑ�/dY����w͟Y�|�x�a�R�c�n��Z A�V��2]d�}h��~��	��[".�Z>��|��[�Ru���+Ы��	�^�|u����V�o�)T�f���qvu��8�9L�}�چ>y=+��@�[�+H���Տ��%��٣v�h4A>4��Wb��d�_Cp�f�"��ԙ��7g�^���'pm�A�2z\�;��7���=q3�����^
6=ͩ������2���[_�58!ܼ/+D����m��Wﬅ�U��G[��dF-�)�xYPHԞ2�y�ت��Ӂ|i�adA�ɘW���Ƣ�/��8W`�n�l��(��%��w:�A��X��i�=���梂|)��]�p�n�&Y�`f��8�!�����sg�{�&#D��/�xgϝ�Zэ��b��W����o\񃸢�ӳ ��򧲱*�EQ�����/��� �Ao��/�SO�-#�1�b�
�OMQ���\��̋A?&�HP�w`��"�I�N͔;k��j���b�w�.4��k�ʗ�b���#>�o9V9�^�N�K��̼��[�5n��V��+����H���Q0�{�z������KE<�.���a����p�Զ d��mÁ(���:E/k�q7:�YjN�.3B�+�-l��|�4����21q��Q�����	�(VC[����s
��G�p��=ȷ���t���n<���{}��'S�'ᄼm�dR`5�+]n���"�._N|�z 7�ͩ1&�����y|�4��X�<���.�!�S,�Cz��/��,���J)܌���y�WM�.!ʡ�u�?�K6E�@�iC��P�	HTz��{�ù���JV4&�@(�V��W���Y���� eX��fZX'Gp�<�0�����2�縄�h%�xP2�$��l�7���X��������	9@4����o|���=N�%�����m>X����:V�B7��)A_��b�kJ�]�����ݏ���s-�$�O��{�M��{�xK���Ŀ�5�x���OY��+7���sD�f�}^�a(±�$��0�D:�����+��.�Y��ʶ/����xJ1�'(Y���
�l���~]�`[7w�,R
U�E0�;��W= �}b��Ց��w�7k������a~��*��x������bbᦡ
0�J
_0y���Pϗr�*e��C�j[noK�ȷ�;���n*��}�������mJ�Ϭ���[O���t��x�����H�VD����@��7�@��)L�?��!P�n��]�C�3=�Y���^m(�i�F���e&��j
�",�]B��޹������(�B���b�����`|VIU�A)�r�'u�h�i '���J65�<��#��m =Z6�6
�ulXʾ���z��!J|i�-���Y=pn����g�ٹ��R����_��7��/��za�����!�RQ_sZ���D��#	��(4!���j�9�6׼��{�9�����*%�V�7S�������UM#"�v(�A̓�����[
֚��P�ѵOj�Ps+�g/��,��z��c��UGh�BN`@��}�WR ?�s0�qZm�M �\#\��a�����]��E�K����v�ƛ5�S]�x�N^�6g�� AZ!~W� �%C��"�č�5��&l<Ҿsə�������s</R9N�Gŝ�S>�T���y�&�TZ˰8��`�r!��8 F�!إ�7y@��N���P_�fUQ�],_�{���U�fR�*6'.p�|���Ԙ>.��{�~m����u�&�b�l��2̅��։�08مSϔ�B���+k�"�����mu�z���h9�:�%!���9Y�8�۳�k#�Rff�^�ꑓ�m�jM��*���d��6�l?�h�^�R�a�f��Y�tE����悌z���M9��?FAà}��������g�k��R�xf��v�׃�����Cr�^t�	{�v��|�pm�'0�-���.�[��������'`��K�#�0��ʂn�y��K��\�x1�rY8�x�mU=�{.3{r��5o����Y���KU!�mIXp�lG+��j�;6�}ql�
�4���*O߽�[��PϜZ\����şcDK!���]�l�R����xn$��+}E�sF���O��ŵ� ���|]BBQ?@qi��}��M���A�g]�=�0%f�;*�O��ڙ&�Z�i˪`f)>D)�pq_�)�0�Tǫ]��T4�#R��N|CgYR<$F��T*�J����@�G�BhP�G(^��,��t��t��k.ʍ�IY�2T8x�IY!c,!';k�ː�f�L�!�n+p����ϻ�LQ_K��L���kQY�q̥�'21��� �p�5J�I_񠄦u����W�� ǝ�{e+A�R�m��~~V��+D��/$w�J7�e����.~"ux�cu�ly.6��;:3�qL����Bj�*`��#Σk�`�c@����ӹ	c]�Yy��y�\���~������A���6��C	��P�� U5rᬂS��ݙ�q5 v��,�t���$�DsD��v�:Ir"���U&�a���)�\�6���ۂ��/3�5�-ZC�sN�����U�JȎ�2�k�,�<�.��
��b�l�'��ARd����'��Hr�Bn�A+
ܠ��mH��� d���-)��d��s,��E� �����[I܊J��3p�h���R����}��r�f�i\��7��e"*�@sRt���b�,su���-B6`����IS��j8	�4puO@ �T�	�i��?�u�nj=p��
[Zu���G ]������@qd*m0��va���R;�	�
�����NE�G�5���D�����}���S��yV��v��lߥ��#�Tw�j;h�L��ŀP��7٠*lSo��, �H�}ϥ����U6�RCc.�r�O g��b�h��A;����C��d׀�+5�=�˷�Fh�W�1~^�R\y�X.p�I�N������<<��1 �5���d�,��XkXH- �����9N��2RG�.C�2'��CJ�o�k�1GH�؏�ɝ\���W�#N��T5��qXף@ǥ�Q�"o�̆{oП��g?$���©�*(�2L��(P�,f�HQ��bƞDz�0P�ry�;�g����Q�6�Ϥ ���.�qp3��/�0E-g\͝���FH�}�-�����(�7N��!;�@�~��1�;W��ri���v=���aS!�7�[�b91J�p]�.�5>����QoZ�\v�տ��eFHj�rЈ�y�f�O�������v�>�J��;�9�v���������9~F�C��w���-�T���AG��\�>�A<��m�'�/�3l_C�#��X?d�������7|������rA�)��}c�p�yi�[�@��1*7��WG�=�<��[]- ���nL�{d7:;�7�!�~Jt����-�a������!����A�����E��p�Қ�_�� z�i,�t��~]�D�Z�E.�eG��3\)R^�(w9+<iⳛ��e +o�vZ*��A�iv�ɥ��m��Qt�a@��Z�~t��~����qSq��{�>�M�a��?�-""�(���^�����XΟ~xg����!Ā��%M�I?���`�+2��FQ���R]ֆ�i�ԩ!�V_`K�3����X{�ԋ�����0W�kNZ�Af�)yg)j�P��v�{F�yhݾ~�F0+/N7�%��'�N���-�n�.p�
�^G�1/6��`��Fq����^�u�_ɫ�c҉3cA�풔T���u9KE�k��r$�	��5<���^&���R�
���1��>�NbF�8���E�H.O���g�ԝ�M��z}��0�|q^��!�@e~f���jt��u�n�1:v�6S��$�)�������܏>5�����q��0�\�@R�WT ���
�(0�eBZ��)Q'9��L���ɐ�0Ԗ�J� O����(�R"�ip����Y� Qڿ�½@�=�6�i�;�6)� V�j�b|�q���Qf4��A�ˈ���T���,�1�S�Ks ^ �e9q�p�����Z���H�mQ�9X���ǯM�P+�h�¯��+���:��w,d��ih_�LR���iԋ����D��\����z0�7���s�%\�	a��9Τ5p3��_G%�սcCu�$��f�i����r.��=oq|5�	�I�����M�E�9��!BGe�~���=�o�>Yf������h7���4U�[�2�i����VQŁs�>���룯l��f�+��*��0.����t{̥]���C`dI�a����ޠ����<\��F�8<��h��&c	�[��I:L��
�'f��#x�v�i�s�(OB{ �*�/7G�ʿ�o�#�ޟX�Q[
��o��;DyP���cє{M����N��<5��n5`����rB�-,�tms�v4%И����¯O���t	�����;��=�.`e���Q��vf��C��JLP�C6 ��c|n�kh#?��C"�J>��֘�F�V [�7��7�� +�5��e^�Z�WZ�á�Y�>�r�Gt=��e�,��lA�p���zL���3+�w�7Ӓ�鳳5��l����r�":3Ƣ�!,�F�� ��KF%I�`�T��:9.�Ɯ@~�d����`�/���?./7D���<�Њ��2��B!wdHn�����BT��>�x�[]������U�-;0�0:v����sny�%�	C�]7��������'DX���	|8�#�|?��{���+K�C��6�\c�S��2L]P47�ԧ�)��Є�Ƨ�x���� l: ��E��M��jK��^"���h�c�C�b�|�[k#�b�w�s��GȆf[e�^gX�%(5���۟\��݄����#@n�o-��C�����r����7�~V�H�:m��T�H#��n�~�<�}دF��y�������n$��t���jtV�]X��,��w���?9���+}Poج��47%o�A�]H�X��	w�E�#��M�`�LFZ�{������/�L��:PC�l������,/M�42N6C��WO"
��ډ�J�����c��YuǠG^��+�3��S�{Lp/p!��E���#h���x�YG�>��%�h�I�-�@���d�C"��de�o�[��ڥ%*�;x��`�����Q[?�t#��e`4��#��&�����,��;��W/��o2�$x�Zp�����K����.�/�)�F�Q#z�f�Q�[p�6O� �Y���^\C@l��)3;Kb��7��;�]�}Q
7�=��o�!�-�S�p��u���O��d��0�C�	k��&�1��&[Q��� y��MedK",�f���x��m������D�_Z�9��f�͒}�=�����PS�ǥ9@L����\��J��NH�DִV�3�^7:�bd�Q����PZ�#M
������y vț�.����ۣ+���r*��ſ��������6C�(.������|X`��O�d���i�Kv�45�!�	p�L��<iv�f#�ibܭ�z�����L�B�6|�;� ��?(�[�Tq����I��moYi &�T8}V�=�C�Q�'rcVL��UɎ�X�Ɋm��Q:�H����D�:������ͩ�e�X�`����W�6uӗjk���Y]J�چ�m
"��x���9�5r4�k�X֦�+(�@~5�♪�dÏ1�b�KM��a�Ԩ�6@���'���V��U|���Q�� W\������D�[����L�������i��J�>���^/
����-]',�U�r��j\�\����F��w��x�&�������1�|�N�e~;�u1�
�n�CW,�������k<������t
�%��hm�gl�][3y�m�ʙ��~��E�����4A�p4��$,XN�,�U����j1�u�56u�L�Vz�h
�C^ �p� ~�f��8�1,ʺ[��M�GH9�B>����Md�~�y�z̚�\�ʦU^�b�Mtf�������Q�(�M,����]����3�`V��\���`0�>a����Yu��j$�F _�߀�b�-�fv�jٌ���:�qik�Uz��]�i�{qaQ4�
QW����Xy*R�?)R߇��D�Sw.N#��V�_?�)k��V�-�l��gh��/���zm�0WB�A����lf5\�
6<g-�Eh����&� �6��'�a������o"=��o���K��Y�4,_�ޡ%�`\"#��-�)vo��Io�<�^Xa�b�2�@v�c���30>��يU�;͏�}��\=t����,��<W��R��л4���Ϲ�t��k�1����/���4��@I�>P��1"�A���I�&Q}$Ǘ��7/�� ]�M4s��ݽ�njv��<`�����U�;�*_'��9����A-�U�hRo�E`�0��RI
�a����1ˠ�%��E��G������c����6��dJ���n3}��W�b�2�}�V]�����OIJ�w���`��e{L3�J����r�	�'#���$�eo�v�6R��tK�A�zJ(_�fwxj*VM�'ǔu�
wm�����+�a�F�H�_X�e�b27�ҟv
��3-h�	ͳ�Lzn���x=]�#�|c�G����eU5�tMYɔk�%�s��|ZS�pA00p+�x�xi�9F>/�����Z���1�w�κ�n�v��a[rg5��Ro����m��v��$/@odyRS�A����F�	Fa��(6��.��]����zL�����KZ�jA�d�a�!a����e2�������Qq'YAK�zb���'�I9���V�A��
o���Q{l)b��"�R��tև""���������ψD{�9s�{����@n���D8��p�׫���׮g�[f��-�*�PAm_q�҉Ʊ���G���(�Řjj�L8����� S\B�y �ǹ �����N�/�aDkf��Cz��#P�1�n�!�$��� ��((��`�C���T�k� �S����-�"�쪐�&��k!���ҋ�:'�ړ��Q/�v*���M�{���(�aB*�/����F�������m��j�qG���Eؾ&Oe_��Ҷ�V�H���1DW�(S+��}izb�E��m+7��{�Ҿ)zM����,�f���H��]��0.�L�E��.�O�~^ ҥ��N�al�O!���D|7X�1����^����s�=9x�X<X�^4�y6>�2��խ��ݫ*el�!7���D4��v���K7.CN?g���ZQ��$��E͸����'�A��t��&`��?3=:7v��47��j��v�V�~e*���1NnE��$m4�\E3{w�A���O�#B5o}�����D��%]��tnQl7	��v&�x�g�DhF���%�R�1��ɤ�Ε���>���Dٷ0_s���j��x���TLľ��ݚL���!;��_x�����WRY#���}���@��0�{XH1��Ag$'wu�U(.��3tt��/��p�ft�)lذ�*5�aA#/�	�m�?�#�ӛʰ�5���ME�ܫҞ�y `�����)#�p<�0\W�
}(|��o8���<5٫��!@>u!.��Z%15b5��q�}�B�Krijx,M��>Jv��8�����o��t?P؈G�Pș�Z��;�)� ���h˺�pLL�p�W�$��5^���-�F�J=�Y��P����F�"������� ^����wqq=p%��_K�5nw������zҐr�#bXH8�n]	M1���eaR���Y���D/�x7lD��ܞ"]P~+�&P�w[�A5�g���C)r����ܧ]����a��M]8���C���2���)��>�5a�2%~�%c;N��ݺ*�����-��Cn�z��t!�!I�v�"�0�m��c��.�\NA~��=R�6uݶ����IR8:fW��e�ܺ۱�C�w���{�9?���܉��S��u�{(|7�L��tkɕ�M�p����,�#׵�d�Ƃ�(B�b�����u;|��w �a؞o���)\sH��AX�]8%�ԪY�&�f3鏷O���� �v�c#e�X{V��pd�#��g��/q������u����d�[�ȴ,��3�l���t􅘫��;�%�����R�;����H^�,��%*�_��M���^��V�*���v{�Z<a�n��j�Q^NJ�mDh#$r�DH�ys��¨J��h
�,j��d3���w��o�����5�[-�B��)vS����b���>"�gݬ�#�����4���Se�� er�H�hgS��V�ʑ&ڔ�6)_-�`P%��~��eCw���8Q������nU�jʂ"r�N�^Ӈ_��b��OP�K��5Kq5�c@�=�qڱ�s��?�S9�@
��d��Cb�Q�	�/�u��	Lu|(ib���2ki��ʄ���n���s��C��5��<Fk��eֆxK>��=���N ���T8���,������d��&���4
��o���i����=B�׵�!�H!�snc�1�o����a�!pOC9����yh�|�Ӱ�������a�\�����oPm����#��E����=�F���~��UG��V/�v�U��ܢ�u	_���%2�m���k>�':>J�؉qߕ��զ�$W(���0-�@3�h��~/��q�k��� h��fU�*�Gͷ۶�XLigt�[�f�ڋŪ�N%4��g%��$�������ɔ�D�F�}����Իf�ѣ�'�KV�5�õ'Ín,F�ل���hY���0���
Z|R-�����2�g�M�	�<�*�6$�N�����Ƥs(��k��4w��/��d������_�ፑ����}�e#N`{�B� A� ׹��Z� �s�	�P�� c��9:�Di�V���*z��Ķ:|�x]��s��S�U�ۖ�<E�5:��!�<����89�?߾�`�ZP�E����J{��+e��42۾d�����[m��p��j�ބ�>�${~ ����ȡ�ȳ�a�4�����?s*L<%��P>�Gf$艉��-7�%ab����
�:�)Qb5@���掑˨((f�̅/JgUvh.�����ub�(�;�X�]�s�U�:��3���s_��F!�L|��-��K�r��)	���,@*i�TAX�2Z�zJT�����Ȑ�I�S��T�BG|�u�^f&����<�M4FfY/Q迺 Ν���2xw¿lO�F���O����)`��:��jE�|X!o{�O��
�����X�@r��M��Sde>���rm����}x@��r���	Ǩȍ�Ɠ$��2n���>�U����Is�K;�i� ,�~���������B�'� !�Z�$�7n�����46�t��W�GʒoٍH�.��~��d�B@���X����*�+��#�h�kM�d�h\h���S֥��Y֞?z����6���ey�M�E�:}-h	�̢�t'�~R�#���}��\fH�o=�v��<��++죊j���������B�N�^�y'Ձ��/��=�Ҫ����<���Wx������+C����s��(��J`�|�GW6���GH��u�V��)O+���=ͪɦ��G�y���e 	9�o�햎F�OeӍ��$s�s��Sv�\�bZS�PV�{q�n7���Ѝj�7�T���b���B�4�4�,S.�8,�)e� ��L��x4͈��c���x�jI�l��Q/U�B��q���vb�Ca5������IN�y���\w��9^�'����n�Ր/D7A��S1�05d 4���2LJfpʯ�@(C..���K����&h?��p�M�k KG�������b`��9���`S�#BO��=��ϥJ��C�b�v��D��aN����T�Ռ���}��T�����3 ��1�����W�X9�\��nN��\,�6{�������g�27��]K��~�7�pF(�e���k��kp%��i�q
�THh�gvY�S����8dk �Ġ��Xā��C�oJõ\LP~8ڔ�ۇ=����C�ɜ]���B����C�"�m�0��`��hu%9�$G�g�w�����b}[�|d$"��Q\N��^	n[u#��A�8L7W�12��%I�<NV7A�<�N�l`�s��U��fu�Q�/�	�ߤL��3�o��ݛ+/h"�Õ���;{HW�|5���K[Sx�v�=�.�v�����d4��0�2�(�j�I"��?E�]��ȁ>J�pE%�Lj������s���d�U=U鴉����Y9Z}UM��ep�I�Y���3�@Ë�=rt����+�9��8�ӧsF�����^S�f~��~U%+J ���L{,�<f��ح�+r���D����I0�`u���g��ԙGL�u��旼�U$P�:���^�z���uQ�R����ZS\<D����
c �
X�@Ґu�w��"{Һ��{1unW��33��z�Ъ��cJ�Ae�4�*&�snk�P���j��1ɿ�yޫ�	������R"h{�#Rr2yh�Y�+��&�g�`]v��Τ��ب�&��d5�v� 6&�g]Lu��YWx���\�1g�E��V�j���K℈'M�#�.��H�M�����!�drN��S��g�!R����;u!S
���vX��γ�͏n�pۙ ��|C�YP�@����Y���yK[��H��@��HK�����`��$�{��N��tV۷�=�'v�wB�)�cI�z�,d�Ä���{1��Z�W	��Pc�px*P�uX�2=��q*������$�7��Y��m0�����4�cjE1﷌G���.6F�Bo�ԫ`W�9�5]���!͌��j.�zܸ��7�L�#;�g���L��MO@���R��3�g��BV��6 ������r�����j�ElZ8�16"I�~.��P'5�W���/��}�=;c��X�� ߻ۢ����x��s��{੽�@���"Ӓ�Ǳ1��9���d	�&��j�l��-�=N�~�.{��p����ãm)n���X"
�l���(g�uQ�+ <�CSy~л=L?`q@���>�W�)�@�&�,L֭���E��&��4$����>�O9�Qk�Y�X2�{6�{��Z�f��'T�s���z$�� �=�dZ����	>-�~�׬�%��-q'�9����Ӓ��!H<WG'Z��~2<�ᇾ�猳of`�
����*�ܵ�6��_M�$sOtD0bw��|>]s�Nj��i&�� ��ɓoqu��@!+�%?En�w,��v�ɞ�:8rS��DL�3\�f���l+�~z[m���W*{�,��K.�s��W&�������[^��y�i��?����뻮`�[1���펦� @̝m�ï�-�r��b5���s�!�}..16�=����2�;&�fE�p��x��aqYrk�κ�֧�{rB�b���%+�q ��=�������9A���î-t1����k�:T+�2�|T�Pҍ��3%tM!㜹���Wdk�����E�@��!<����M��n��n@�[*hg-�ºMx%�.���!?Cx]�{G2�,=X]x^l%����%��ZmqT?of�"��6A�ت=nyc$]��f�������~c�2u_�da΄�o<BL�#^�E�:'�I2p�2Ћ����m9�HP˱��@�؜�3�95n2�vPg�Hy45u�َ�P����p���b[��,��	0�u�������IG�����t�:I�z�ͩ��p������*�})���p87 �7>���@ {� ��tt.jî�)�`rӯ��:1+��NRq�i���Va�<�V�-���������h
@;�_�F7�Hz)hH� N`cKR�%?{"|%v�"%�܎()4����$�=	��j^_����,R6����^��}�ԙ9}q\�%y�!�6qL�(`����e�s�[�벢*�</��h��#k����7<NF���mm%=�P���ާo>~w	
�MD=1���3W/���-3�a.��-O׾ef��̓�%�	! ���o ����8Q�L(y�]kD�E�]ռ_1��1/�����IXZg�yO:�dmp ��