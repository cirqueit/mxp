XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��* ���R�[R�9�HHe�>,5��O�9v��#-�jy󐻁�ePR�o5��E��2��v�j�Z�
�ɼ��!����f����pK���r8�ào\_��t&^g�+eY���y@~�,��cNoIA�:����is��fr n���c��t#_`Wws+5ӿ;��Ѥ�C�;�D~!f����{�Kň���`�6�&����nݼ(�?ݡ�W����o�X��Y�٦��-u����5����'<�.%@j�ό1�m9t�"/fZ���733J���@�T�C^��#C�h��1k���Cӻ����V!8/����]� p���G@��UA�S��=������^J��6��Y�7�Ņ�C�6��¡�8qV=���m�O�%��d���u8�Po���n���f�Y�~ɥM�^�R�����z1Rz�W�{�;2`�S�=�Z>cV,A�+�W���HD�r�<��t�R�k� �~}�j#~�U8�Ҭ>�6&�_��H�HAD�08�I��w]���}���0�	�����oS"hMȭ��wݏ�޵]w�t�[��� a�ߡutC�	y�-t|b�mɟ�s�&�Kb���|� ��H�rT���aE�U����鍷s7��)�X}�U�'�O'��Љ����1iR|AK���S>���z�K��6����ήE���tU�M�a��R&9�=~a���L����#�	/yg'��_�B:������D��t�c�8y)X�Ü�>b����J����4�˞� �o��tW6D���O���XlxVHYEB     400     1c02�7)��N^��:�zS��u��l��w���L�?��/���)^��:��T�`�6�/!�t-�y�V��G���2ѭR=�#���J��[�
a����uA.K�ɑ��s����>$�ί2K͂�9�#QSy�t�)��j�A�G��PC��U���N?b��>�r�N�l�	ؕZ����PӰ�.R�={bqH��A� ���h~��������$$��ndrue��P�1ip�O�P+m�ߌ�b$ߨ�3��Q����=P��Y�0�6�}����VC~��{]pa}q��R]^%�m_��!�*�_�%~���yuVe퍷�wzU�}�K_}����M%>P�l'l�\qՋ���Jz�_�O��~��"�<w����w�Œ��pΧ_ú��Sc�k����'3����Tr'��xJ�#���m��ae�k��hI�G(�)��j�jXlxVHYEB     400     150�j�Ö4�P�������Z�X^��h���ɜ��V�2:>:�o�>/O��gb*m2�Cp��ANZ�{�햳��f������	��>@���u���PȑD�[S�{��q@m�|���nHmKom�ܘ�377��щ�)
Ш��re��>h��7o$:~.P��0��иAX��K~Ͻ䋤m<�Lن�ǡ~̘���I��ٶ+\��Ꙭ$��]�5��� _�4��*Z�F�v�u��ƨ��Rm'�L�4k�JE��6<�x�Σ��=�w��[�>W���S�P��b,���TL>�Y�ڈ��ju�zCMc���Ӝ&Y�iAL�)���
��9XlxVHYEB     400     130�ى�2z����"\�$P�q�z��T��+k��&xL���
� ە[��UK\{F���Am��ക=�Ws��Q��Ӊ�~���ͩ�[�y-�-{`�ͻE�/J��x�f6V��7��{��F��}���:�I�1J#m8�d����!��w�7/�%w7#��x�R��nT�_`Tǔ��+�b�'�I�}Rq�J^���0���㩚��N�o���'���;��$c]mj�:�e����Q+�R�$|x�Qp���a]�����Fc6���e��`x�@kc`��iтrz<Y����k�����XlxVHYEB     400     160I$�~HF}�����}�-G��n�V�)�)�S��=��B���H6���-a�y�&S\!aΎ�hG�KzH+�G\�\t䘪�ql�!�\���;Uk��p>Q��/��Ԓ�'�]�_��i�P<#M�߈7BN�,z�w3��WP��'�.q��w�U��jPP�/X�mT����eQA�/�Z(�N�*y��*�i8�]���[,�)�@e�_j�̿�#cǀ�;|Z�a�y������2�9��(L��[��L=+�ȳ����z�^�Ǻ퓻�������ٲ��˟�U�mT���7�Zh�B���0�wf�bx���0�=O&3p��y�i�A�d���$����3���XlxVHYEB     400     1e0�I~#���<�φ��e��v���g\Gp��A^������ |ϔ���1g>�O�@��'�5b�`�Ó[ʚDKV�*���M����+�e�DH����0��L����5N�.|��)C�;�1k�B���ٛwr.�����ɴ�z�h�"O��݄�@b�dx>�	����M��eu,	���Wtr�⵰�$(�a~iw���F<#H�E��%.#��7�G]��w%��,-3a���r_��B�/	p�Ɔ�µ'?��ME���_%�oP��L.�{7����_�ր��٤�_d�ȇ6�fE9Ϝ�m��udj�G.�[���2�&�z�K��e:����Sp�[}���|�z~�2�J������>�X��V�i]���y��6>+F|��Y��xYG�K`^��R	������_<u|P�-LI��P�n}/�fe�v|tB�Ĭ>���,�,BE$Y	)�QQ �B��׶;() �NXlxVHYEB     400      f0Ӧ}9|��y�/�Vz�e�f�9�l��+��`�v���-_��.�Y����I���{�0�ѡn/��)?3��2Dm-8�}tB�,q[bf���������C�6%�%��8�s�,�j�(HB�(ߟ��#Ͽ�Dg�R8�Q0'��;4���X� �U��Xo��b=\'��[�5��`�� ��:Vk���)yP��Im������PdD�J}�]���z Fz!�6�)vS*XlxVHYEB     400     150\z�%��3y�`w�ʟ�������^
x�t����-6%M`���dP!ss#%����*"���8���͹7���lը���m�J�$y*]�(^��YC�p�F��t ��OϤG��=��r�ۖ�EE�2��Y\sa�Y7#����8K�g G.�⭌���i�~Mw�E�1�?�B6'k����V��v�2>���
�,��N�0�u@��c6L��J		XƫN���}�&�2�no��_�Se(C������a�i�6��"Ln��+Pë�?
]8Z鮿��b@�# ��܏�|��Û/�fK�2���SCs�m�_B�j�XlxVHYEB     400     170JWB� ŭ��ƌTJl3��1C�:��u��N2[l>K���?�q�CQWG�	\P�9����r��P	YN#0�����L$�m��~e�B�6 Ħ΀��8 (z9�<�(���m ��_d;�٣1V�Vb��4�"N��5��&�|����A˯X�@�,�66w���|���}�j�jՐ�����}8	RT)}]z��nf0~�a�E�Y���AXq@Q���N�
�P��1������� �Í����R}B`q� ���6;��J8f��E�U+f`<^�Tσ�ʭ�����[�/�0�%���p�)�ynG�֘Ue�i@�n��ػ�(�ݧ�����1�3��bk������^`���fJXlxVHYEB     400     160l���?�Vّn2IvŒ����A���Z�����˹Af�ej�� �O>��a>U8�@�7�49~�c���g�B�<_��9��T�Z>,��0x4��sV �����bj�щ�u�նE)����քp���α�յO���'���u��MN-R'�y�>.iVw����S�XO��yz"����Y�<��{���Qב1I��~�;��3� Y;���4G!I�6��"ӛ��S�W�
�������?�񾜗�W^J���>`�Q�eK�(o�o7��G
�)���da�+jH����eq�D ��.?jo��fѻ&Ø�C		��c��`�η���|m`$������h�XlxVHYEB     400     180�(���^�v�"P��`���k$ʋ��'���Ĉ(�e#�o<[�8��������Ed�pn_i�'�l���qbI�����I��m�yN�XV�O}�`�ٻ��J-Hﶳ@SFj�_ ���HSs�X|uH�� # j��!�� |?D;�k� \�F�m��x�|�a<C0�x�&����{\:n�=���0���Txt�ǒ���e�+y y?rf�e�?e��UhE 	�aŝMƸ��,�0<k���V��E*^y���H�9����/�������ޖc�7ͤǋ�"`D�2[�n�����/X�[i��T	o�H�&����ʾ�ѷ�;S��$��,�Ɠ���J����ӎo}��x�Q�
�`v�
sXlxVHYEB     369     180r��]*[Yo�$�n�[�Q#���_�+;e,F(L��o���$�[�2�\�`�[S0�8]7�/��
w#�Q���SƄꝋK7�ŝ[����.m�T-6=�_�>�\�X)bX^�\���C�SV�u����0f�ll�� � CPX�~��K61j��Yf�+��R��"�	3و�����������Dr����������{���\�1�1/~���B�1a��I��=��)���Jgv�8���Η��v8���uN���q�kS��~���)e�
NM|�ϝ9�d8��ƹ&��Ϙ����ҏ���en�K�YJN�G	�L=�Q㬲���i}������eG?+Tzo�I��'o~һ�?S�6��Y`3�	��@�%`