XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Q.GT���p�%����� �͋�w�5����i�����(Cá��CۓI_U�Q�G%7��E'�NQ�Z�I���]u�!!b]�B�{���8�PjZ}�U�W�J�M�H�<����ڶ�m�>�n��5��������sHˣ�^%3ӌ�.Hzfv�̬��C����X� F�]�#?{�r7�%5�ErL�@�`	��.=��R_>��� O:�a�T�ҳݮ7�<񨑚>�������e�hl�m�P7�u:q��D:�-��{��}�6Y��3SX�2]������@C�1 ��b_֘ �B/�?�2��߲2���6^�D*|��S�wI�>{!nŜ -1bGx��% ��^��B���@�ˤ�Ol�D,��Ѐ�r�zc�mS�(���^#�ds���+r����4���ttss M����j��k?e*������L��@�D ���tNp���SQ�����S�n�}�8`��[)J�T�q!���W?V�΂�yz�r���<�_d�8I���Fry-k��{�@y��>�5ޅ�����y�o3��:N���qYs���!h_�����睋Eu��8o��y8�j���ܖ�qI��h(��e	����;m�X���, Z�*�`���oq�!
�~M��[M�_+�(m���,�'{�e���M�0Vu�,̋ڥZǤ�M��4��$�Y�T䘆W(�u}�F�h�l��#�* ��pՃ
¶�F�Q��sߏ��")�n�pDXlxVHYEB     400     1e0�9Ma	�O��ߖ��Q5Q�X[q�Q��*F#E��W���!g䁺�l;���"�����nU���tDNzg��^�?t9��b5��M�M���ƤG��nhm����<�����B}6-�U�pK4��R��T��<W�nX��1�ѯl.͎�	�^��$�I7�i�>cx}]�
��ut6x����
���S'���g�� 1rȻ�:��b�o���w"[T"qj=<ك���&�u�b�D�<s=�]�[��IOx�_����5����`B�"A���J�Lp�@�ܗNN�cg�P�\��Y">�-��#3M4��[��+3�(�~]���HfA�34�>�H���.��D>߀�;�;���W=5�.�q�`�+mS~�����|x	��t��3�O�uL<��OglA8j�)n��3�	��O���ғ�3�L4�g1�='��g���Z�_��ބꝋ���q����F�$2.myXlxVHYEB     400     140�.L�F�'�<���t� �թ 8kșjĞ�e������쒭� L]�$WL��-v�&h����r(� d�ȗ���s$�^��H�e����.�r輚�*gP	��B�~���_6�V�U"������l��j{�|O��\�\`���K�UX��b���|��d��%�ۼZ�22�<: a]+>t����	SսQp�B��!p��)%eCx�F���+7�P��}B]~}��:��Q0�[��6�$�`:�M�$�,�\�}��q�q!�'��/�ǛW���])�.~�v������
�)��w�r��0�ҷT��ɚBXlxVHYEB     400     140�b�L�8`����)5�?��[�A�!�ō��F�i�D�E�D�[v�A(a�Ta��p���7T��5ǅĵ"T���ˆ��Gd��P�v�a���[�tR*5��e�bVq��
�R�lK���`�ݯ�;u!�6�ѝ�'J������C��޲����O6PR�Մ�0����(FX <��Pg��z�b� �[2G>p���cf�>&�ʾ,��ZV��wzՅϡ�����S�ן�p�""E|��V�OU�g���l��y�5����V��Y��c�$đ}���U;ŜU��E7m>.��N=���	�竈��\�=��{�XlxVHYEB     400     1a0�% 	0�|B����g%��|��^NOD��P�x,	 ���G=�0#ד�s�R�v]7�^��2�?_Äd�
���d��}�7e^Pk�>�UK'� ���{�G���n���e!~�t&���T�4y(�O�����z�{���;����晦(�AIͳ{��Lʁx��Y�@�7�n�d]���E�,��fNB�Pd�PL������b1yyP�ǆ]�L�i��+��Y�u�%T8G�qѰBf+�� ~�Z;�O���I�$���n�|W5�ޞ{�8������M�ד��V�c\�j�]aB���J���F��۽���U�fD������&���)�k1���w� ��uCI;X��>u���dC~o�҈���qY� O�ȑ�	1f��8���x{�7K���t��.�sue�\��%�A 1XlxVHYEB     400     1301d�K�.�o(�f��*�&�a�,���e�"�_���j�3�%�:繇�ˮM݁T��T[ʹ��9����LR0���=�Z���!���x�����+�Cm'���Ǻp���!�e� ������v�׭����WiS� �ѯ�
�%^ �(S��I���������^�Y�N�j��3%Uv8�;�,�F�6���� F0+AP�%%m����$��.��?�����aۍ�%�2�j�C�}���#���v@Ԟ.l�.4�ZF$\
�	��:��9#φ��O�62�~��>XlxVHYEB     400     190D ��&#�{�ݘ|B���Lq�p��W9� ���(�.��p�4�����)�c�;����%��6��_*9��n,e`�V`t�fZ���XXc��2`��V����|�;{�y��%fMׅ���?O����v/ԋ����E�ߘs��O!�����r,�ws�ލf>O#�������F}���/�SJ`��� ��s�и��%0)2ڙ%���d�f��0Ӷ��/���#$3<����e������X�[�܋��Qe`��s�n�������#5���EIY.cIX
��3�|�0�[�'�� %��5��^ԻIn�/1�h��3�H �8�R�b�P�����Ji�]��:�b���� E�Q5ղ��=X3�`�&��3(���U9�L�3XlxVHYEB     400     160G�_�^�y���:������@!�,�3��a�����AS����Y.��	Y�)�WH��l#�<J{yw0�16D����_S��Ѻk��{l��\m,�,�?ns����K�2�k�?[� �~��u�wU!?� yPe��k}8s&�y���
�x��xr�T�&�bˏ9]!@��5,��":��뵥��Y�b��^x<b���6�q �`���1��d�sOY2����i���b>lQZ��g��
��ҪZ�ЇN%jޙ-��DW��LժX�i����R����_��'V�:z�n7�ȹ������"É��2�pI8��H�$(y`B�j�[�
�K�4���XlxVHYEB     400     150�nS؄���k����4�����zv�w��3��hs�l���Io�g���}�2k�q�'�O����_�/
[#.�,^9�$D#V^�`Ih���EBD+a�-�+�[w�^��tE�]�ն���X�*j1����Fv�[P��$�9S˛�	=���[��l����1a� �t��sW8(��� N !9R�Q/U�f�(�%�//#����=���җ���G�?g-�>�(�h�͋�l��'D�&ƪ����!V*V�b�7�δ��kH24���-Ku��5�z# B_���%��n*���	[�le)��?�E=�,�A��:��aXlxVHYEB     400     1b0��`~?R-x�����֘T��S�s]����:/&E�����O��$$h���/�K2�.'�O�M��Q6F���Vt	�����2�N��0���d��U.��r-�;���Y�35t���"t��2˅�}#:[_Z�w�2��^�C^ :�h@��P
S�S�ވ�$�I�_����H2~��.2i��O���z(�xK��`�?B�4���R�UD~����: �j�����\�KV��-W�t0{��/K<{K>�{@7�c(ԍG��V�q�A�6�TU��J3�%22�v
*s$��l��%�Z�RU���j���Ip|5�J��>��X�*>l+���`�n�swF� �})�ıo�+bFOtMZye�!d���g�C3�:��D��(��u��.l'ʒ����f��%N�zi�N��E�XlxVHYEB     400     1d0��I�-l���IHSJ�z����*m=�C��D�ɠ��@mQ�k���7+=�� ���%��	?_�G�S+�>��r�"i����k!B��L7��!ƕƃ���Ӡ�+FjMb4��9_���'b����*��9�Ou\��{0���^��I�A�}�x�m�k���uN��?����nx�?C�_��l�ór�	t���	���I3�k��׉��㎅]��r����x#\)�m�V����&��*��0��g3����!��_�,�T@C��;`]��{��DB��*����"��� ޞQEU�/¾����xU�F<���ZH���?ز��>CӁ�:�j�����4�����q���;P��E�> �Wc��򁭶+��vgy���|.4�O��S�a�M?|���72sX�W��ǰ�|4c���U�wy��"	5�{t7���c�����)� ���XlxVHYEB     400     160��S�#^�x;�Yۍ?9*y�M^/�-^�鼗�b�mv�K�����:�l O,rk_˗g��\�7�B_8�2d����/��n�����e�q�x��!w�4���sx��vཊY;A��v��Z͕�z.~=�kO��7�ֻ݊�6� xbD��`ݩ�(.��з�*�c^���{�㵐s��<	�.O��,\�W�	���^L��b�kK�R�QW~z�q�����d�i��!�V:�6	<�Q�qں��Nl@vr�F�"d��3��Ec�	m-|�g,�x"���3 C�s�����T/�&� K�1��d��0�γ��1�-�H�lE
��h#�c1�[�_�XlxVHYEB     400     130�����Z�ob�Lid��O£�SON��	o6x�Sp�L�����L#����L.��Y����=�Q�x4?Ɋ�;�&��6'��(�#�u�\[~yq� ͚�t���Q��n��9�5��~"���A((&{7$�ńSi&~hh��Rp��'B��;5�=i�!Ds��yg�~Ig_9:���́��0+�;|�7o#��f 8����5눀�jd���BWѧ�X#k���?��l"�kj�8�H��(�H�{��@��m��gb�p����3��i�z<H�E�i��Gc��^��XlxVHYEB     400     180��!�;@;R�k K�]�&�S��_�ɱ�
���&@Ya�e-"Lg���6c�c��Yx��q��z�� �Ä�k�|+D3ᅡC5�:��
vf~B�/pW0������?�QZ�#�,�+��*�9��Z�y.�6���*����d��h.*n���42��*��[��A7{fͧc�_��?��y��?���lW��? ����[��}=�D��]�}�{
�G�q�=+m�����H�\�d���jj�� ��/XF�j��9�tn��.�W,!�f�+��f�� ��<�&�Mû��Z��ꖺX|[�k�ľn"��1,��,z%�`��Ip�<P݅�-4k	�,{��H��-<Y{�����;�>����,F٫��s?���XlxVHYEB     400     150W����o~"��36N�2_�!$�w�j3�$ ߪ����������[�j��ꍾ�?���Y��ԌP�=���&	���>85-�؞!��p�ݴWRT\��!���J��Le&$a���'lE(�ÜDNZ"T�z08g�m��EP�$ ���@?����B��+�AY��n*�@;m��B�'*o���zdZ�����a�����>p VVz>��1C������_	��6����y��� e����ꊎ��T�L"@�'���X_<dC&7�@$%A2F������d�y����k|���˼�"�'���9Dzl�[�)�&��B顒B���Gm�?����z�=XlxVHYEB     400     120�,Q���M/�S�Mm�k���0�$x�9�T�'�G���	/<�5�&�{���UO;~�s�-���

��vYB �iA��2s w�M��ju�EG�,��<&ئ*����A�3@����^b��ͮ�C3)@���/�n���ʁ�\��}4�G��!�8�Wk���I�h��>��r��x����X,�����#\�F&*�hΉ���o�	D�gR����������ܖ�cZ���z�q$��e�0��)Zj ��%6��1�o&w�=���Nn_�������5��G�:��l�XlxVHYEB     400     100��������s�)�<��;�?.U1_�gn���bb��ץ�a�pNN�Y3�i��7�6�g�W2g�-��@�X�����[� u'�)~L2tFs��ct����E��)�j�Eq����&k�Zm����G�揢O�R%x�$#�c���/���蝅�ʄ�an�xW�������K���4C�U]�}�k�%D��>����n^��HW��7�꣮8s������v���Xnet)'��b�*�XlxVHYEB     400     1a0�B�$�:o`�'�qVi��0'���gTQ�k��si��<����)r��}�T+��4w;��/}�L���.�X���N����-ZvSO�-$��z$�XK~cc���,n��#L�G��\+26�hd������n��A	ב���J�>U��18}�"v2��uW�Mƞ(���nys��어�B�,ť�%hI�C�W֝~w�*�#��W\�x�KR=$�u*����[?by,�/��I%d�tmp���,2�7�צH��eZ�r|�F����j�U�~_ B�=�1,�ֵSJے��{md@���l�=��a��LYt<#��dZ�9	<Cx��'��s���%J�<L@U�&��̇�#K�\+��~!�8���͵dnFd8g�ݗ��(�*x�ѱ��u�k�I�XlxVHYEB      27      30��њ��6}�1rJ?��ލ�k�0K�p������n���T5�ɦ�