`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
1nKbjIgs6wYZinSBYz7nAgZrWOkjkvwO0IBAg3u5sDxPwYEPSCVTQFLhIhQuobHEkwPMdzksg0PY
YQvpljpenZRVE84RHUlL9fsIW6qD91InWn0/w/ENR6NG6uFx7MpG+M8wnYrnsccbwfih0dqar9Yy
RSQbgcMhd471TKrOz3qtR+X/UQJh9ZU29HpghC8fdKrr2rVdCS4mStOl7WknuISuVTSZvRarn+FF
Y1IF1FysDrwo9DzCWpOccmBDImnDQXzw8ANiKQmkGDN/ub1NqF76CUAwLTcZUKeT7NH9cPwp/bDY
j8guN4B3vsZBzPyTBMpmyyJp7JFLVz0yYGkFpZDw/0BmECO2b5dnt8kmipK+O1oWjeAf2LT4Re1Q
4CrbxCpHjWDBQbi0vlEFlIOws2Q5sNFKeIYF1tC1cVkW4wB6NaanN4uSMWeBImTNpggw1grEQ/4+
YK+ZkpGzBmkJPTI8agt49uplsiYqQwWExC6SBluQlg+wWKFKQNhTGBAe7IWBjW8ZI8lWaCC32aQa
zJkyLyphJCl0trRLKZFBQVS9XQFB5JS20G5lUt/yrpVg0iKgXiBdVVzU8gdN+LgsQJ25ZiRZQ2/x
r7Os7NXbuAJ6QOgzd6uyBP9dxn+qYKt+qmkt3RMnoQ/hXzQcniCuUzQb50MaaguccxAUqhWvZQVN
4PzAJ1diLQxUOTvcESSfvUqEi/iWSxXY0T8JGx4UJKUlA+ocUjwmv3uyEgtG2ocbtaR3e4qWYO5j
5scWQ0/fCe/URjh1Rb4CoBednd6OpDUcYNnL681hhm36087wKwZbHVOPXzApqcmsLyWMEEcJJNVj
yy4q/3k3zz36hNb3vRbC5WQ+oeq4+gD+vIYCXN7NQgSqe3hVlq6/1U/glhSaiJzuYreiq7iTbtCk
XYdIoIMG2031An0gV218vdAmuzG3lOuiu0ayYZvK8lEUl9rV9H7R5Mct1pTEyYTwv2QrYjbkdvHX
YoPwpxH7jbpiG4pdzpeT1cjbqYVwq7G7btavPRMTPgrSZfS/B3F+lrAc1ItYNZADPQh6DphHPArB
AZAexrOt/Vw/5SE5DelzqQdyXi5R6YpcVi1TqeMwMU8lxJ+2qYk4O+MhVJ5xGwy/oVElesPRZdpB
l1AwyV7NuyZNxJqT3DE/pkJ21qdZdljwx+gmjDn28Z0v8GtfbqazRGwrGHU2zNY7mv6c6wGIAly3
hb+U+S+kEfnvrmeEadYSev19J4oPRFkL4DKPJA7nbMeHRqvLlh8zGetUVAvA55gFFTTjDj+PeHTx
SI60laxSfWEsq+wkU7dSQP5Rq4k4/+EMBA7u/J1fTmoryKkvUAHG6VT5t4h74WU15ZWfXHACm+SX
OsGB/U9gXpTQb5mKW6qIbXiZkIK0u5wYuo5pUQbPI9UFyTbYBWjsyTfPyfArMAbNDq+jiJyCpW3W
HV10JwFShXsBadea5O7ne54sJt4426zpbFkYp83PG/sGZgz7ZQ==
`protect end_protected
