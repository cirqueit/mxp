`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12016)
`protect data_block
o1aQI+nw6LpnqPxIUnuewrk4CBLgBp1N9YanimWm/rluqz6Zd5YLa+6ldc73HIM6fgjfBYfG5Wuj
KPv+hsMwc/vvVkqMgt8/xkFpT3kL5mgl784Grac4wJi0eNITlz96Q9w0E3u9Ss4wjrXRdz4FHnma
VyKt4qGrXWOxowXyMz0bLccb7iThltmWm3B7xURhXGXCoj+S8p6F1Tait+fXtJYdIbjcgIbbsnxJ
61diqnd29LdNZ6Prh8sOQGBCqnzRGJebWmEtYmidPxr35OgQAiFfJhDfWwle8Y3MapX/fDFxTO1Q
GUA935BJG53vf+6Ktqg5IvWWQ9d6x4ZiAhr98/23ewkY9jK3gf2oAoRHg0Bzf6i5lhV80AUBwRqq
LX8TrfAod3jSZuw3AZkUhOwrq7m/IGcZRJeRfj3edO0JDd4r0zz4Iz2chtHyhZQJEXQ7+SRWIql/
tHVFGCN4Tltg2sqmzGuqmsRiKD18yTYE7VuSbxz3peBh0MixQYTzIj1wMaMP5FbujSNgUuKXgTWR
1W4DEUDrljVGdqvsndXuAI2s+JaRAEemPzELFD+KIpnOQWvWpoxTU6IYYQD55/SGRglH7lN1SOsm
6EDBHuNvXU9em25drYcFsfwlo5SAPUhy4fHCf0zfDoeP1Dohy5AGm+1U1qS4fZxy8Cfrtj7f8+t1
XBn7TF40nqYoQ2Dk9qixzVVNtmWWlRwm1b913EexjLvuLVJr26nEYCI/4LWXzvJRyqx0rwnQmxSo
RCLCwwViPJ9nnXTvR4Ls0d879SUHHrU44XwnMoqbEc4zdX0X6ISE3FqYSP+6XKf+a7Sh0TB0VcPP
76K45Wo5FJZOqsrtlc1+C0C3hqFMwQDBbnaPKXnc7qAynemwSkIjpSpPWz7WIGA/36WS9t1b3fw6
88n5ODkUEZh6qfLsaxYLc10TiMY/2v5aXZoS9OZ11ZIUUJVU+cXntTiVsoj6pS6wPp9+R3Bj8ewJ
wUr2CWl9kukXOHOO6Tlfz0ysMSTBhPGvd7bM1hgFFSM1aPU+8yrYOvRZaazqECp8aitNX8av8Rx3
UK/sCDodGxvKB7/zeO4pzUjjD8EYny8xmdXD83/o3PPJn51Ijek4KimuaxECYTxz0NrhdQQ+tNp3
220LMmbG9GcIwfbDJMZOQ/7p1II94GZcJNoHgExJ8LP+tfbw8mN6aFUziaKYH7sE8AZpjaW5lAHR
F9TiByP1LGodDuqMkM9JTaNkNR8wbqp2h6rYNXlRXUkTGGmEGIdEpQHUf2lLnn0oTbH7XeNVPLvv
KPYr1BXxjHJDb+DeOcERI3E+djO8wNNfJlgF6oek38eXH2dfjhQn9Dfoq48deUoXVIVzJyHGLhNh
TfzLbp0vMGBOlEnqcq27NbNk1bKr1y0NR+/kMw87RkN4r8DxlSSFQi3vnpEFd4yXAlqt5aFjJmip
Q5lWX5FzqAhCjagD+eC/Nn/Z006EHMzqlL7HFkWp93E6Y/DUtCc521fjXpHlKjHf0+cU5KfQaABw
wtq+uOY7tL6y97ttRiv8SOcv5VDuvaEB7RKale2htCqA12gTp9ST0Ojjrefrbr1vUVdwRah/cyJb
v026p388imhaIVEfCMODItvdUsXRVotFwmziGoXcisIOajUot5XPozZzGSQK2ovNS/n4t2mnT5mv
X7g0+sqKuiRyyQYLeWMBwCcPWTzKtxokUdW5QeF3pqzCPP9KJ4FbiuiuVHoRUbffHC0x91I0TJJT
KRJj8thdswZ4b8y+ywD8qDP3IKanEdHhd4IaYijVguui5agFo5HE/RlzmoAV6YMzeH5UkNL2NiUC
yMAyCld6PEqt0IQ1ozbKtmppfx8Xp/jM6WUlhsqs1ylMpcAc+uSRILJ6JpSnmu1sQoo5QFIvGRwD
vWFcjfr5myMIRxiE8qeZ5ir/QSSG48kPbndmHH5WRWTmyhUqoQA10BlUdc1zIXRg6LzjW/aB09Fh
UQEjJ108+UXE/im6/gZah7pMtsThK1xVOrlBTts2HmWGYor1cEZVLuZUUcK6zDDWgu2TwxAMr2FJ
odZrXN0ApdcNz90zUN5jMPseYl1xPtu3CjePp7EIhp2ItCCaMJpaJKQmgVWT525BSPECsOsZH7s8
kzk/50fojvSWIFsTyxts8iNnBTtCuEBwynb0vmqIGBiIUZcO9lwk/c84VqEWG7PnLccs9OhZDESz
y1U2TetCMvfraBYtQn2A5bEweNl2oA3P0z1E+BdN1lITm6Ar9tHN/K+4BXwT+HW0M26r2i70XNmn
D6dr/wLE5R8D2rMhKVFLvHpWNIFsL+JypM8JKow+kmM1cau9wJ7KAZoMbnS6GwxdlMDpmByiv2m8
2WOCsfB8En9Pwqf2ljqHWiqjh3oAHx+ooOUkAHmBfsUB00pnwjL1o5uylcUpbh6eWe8k7A7ECDUQ
CnYWtXKag7sB+9xpisHktujvngiw+49CxYvur48ShxRwUtoO5XhEjwoBypTB7Yr04T39BrNDFr7w
1wwZqxjx/796kfaUQUr2BMgaFc9n23VupQXGSP3otGMc7brdLMP0m/hYPH2WWeKDaDYLK8mvNae7
2+lH721a+iRaBsGkTggX8XncPktVx7kW7r9TqjaDvDcbkarAEbhMe/JeAfy6ry7Ir2qkth7/G8G2
a9T/9P9Vx+0X/IzYoaUXGpdxgv0SaC6wsZVSFhoC67T4ualZX3o7MX/QNQSQTj9hgpEq4FpKmN5U
dbSHYM8xbqCsS382K03GafyJJjvo+oR91fe7mb3jlYJvqVbemKPioFa/Ng2sgXEdIpe8SLx9UDxF
+cBWZGcxlUyqnTRblH/f05yeFvn9WzZaVIbb9TJB/OjHQkDUyecasizovATvltJ1jLpfUEhM3Hf7
w8SJerS2MDHuZwEAIw9JOigK0GnJShrPeiM+/F/ckXgAtw+qAiCEQ9pBvt0YJzCS1I/STlV9+FPk
RmCsRLFvnNCpxoxuqECgEIw3zevckwuBLcbJ+sWrFpa+JPgmvU48yrWg70Jiv93RksU/E+uH3DsH
X7tmMMXGRFFcHanF0W+Va73mLpwt+TrClm8aOdgTC9qE8DRpCsF4DVty4RtdcktGszom+09hcXh1
5ez6XzVw3g6Rrz9B3e1flykK1dimXvRn3ifOlF+V6Iw/6Bt3wn0DJvQsE3XAvk80csi7VlZl0x86
+ezwp+HcBmbG5OYH07KgZvhb3iLcjFuUmLRA6jl3fl4TeH7WUNi/JlRV8otbc9RtvamcF16wPQ/H
E7PK8Wfb6ITX4BjkwHruynLJVmiuehJxMhKIxBa/2g9KTNFL1BPmvTr5SzNKBvf0oTUrU4D8Olss
b96nXKURC2JhBf+vPUEvP5jPgK24vwR+r7YkPj9oQiOuE4Usqo3uxyZ59iFjBahd6TXqx0+QYn1k
X7VJuXpFvOK6faV1pwt7zAnYi//OMvqavKXzqZ5yCmdnHHwyKAgPMbkcqgm1pSdMjM9wAVFut8LJ
0c0K8XEUbdos2orTpVbjhpSTsniUMk8CSZbJTEnQFdAdY+h9/DqH8CJlBei9crpbRWsq1JRy4xis
HvBTASpJTy0m0TTCLFOb3/y88H8W1vPk8AbGIJ/enjwFCsFzMy1haZ+MSzB0kWli9iFbDwoy2xyt
GzQd6G+l6EIyudPAMYLIE65F2eAi+c+2KLvRREbIxvtWm4pefSD5gMKuCS6VWRT/9Bn7j5KfkMSM
IVhYNqFPBEgbg5M2cqHkyDbsXUaCMgoi3D0RTJL75dbkwZiVOS6+Pp0GfistRK2vHQMh4YA7eOOL
5dbkGwBJcXC3Gch/gtdGu4Q1nl6mgzQ7H49f8lQQ2YfV3veQ9XTfHavCxBTRHsddu+xG09sn3F+Z
8OwLD7BaU9oJ7ghTK8TLwqj70IxVjNt0A3EbRNCMRDMsCTmxZqcliqMjaHdPDQyh3Gc4IzpsA3pc
H1MU+9Bh+PdtDAsjUXofZSq9istRcPUcEwmVSKh63aLWjLZ5n5pEjQ9JqCjHhyKlJaIkQiawT4VC
9OjTKilrPNOWrx/WM8QVpQ75OfjjNE1SvtojApvcda4x4/5D4PD2/S3axn3Fclof/48QB9f/ZidB
+qevXiqp5YxH8rdfpt8EKewAhzC32ZgwRGudv+UIU9IOKR9xNsnt24E0SMHnK/vkzx5rFybW5rZq
rOEUHgGn9gLSzGWXfRItf2b7Cf8MCz3tolWUOs3swDv1LwcLkjK5DzuxGglvZqDSQzWvIhyEHVxr
927XpFA8iY6ZLLBSLPHe7jCM29VFgQIlCOHP00NYNxB2DYcUBKnGtYVqE/W1QkdHGTWeIQN3jfiF
1bnkZ5+8kCrJeiROcItQGxo8swRfyO0G8cXCokQgVfJUGDtowNALT9bFDBCElPODtV4VFUIoS9+A
kGMCh4Qc4HmjhzzDF9p2XRGPSM5knegtKR67MexacInbksbNmKq3xDAKUpkI1S4zMDolV2KExddb
iQIFLJL9OAuUfR2f6LfH/7pImC/CE2AvDVX3Cxn+7N91YDz1Q/WbyNu0VCa//Be3n1DCi/pZnrqw
koQehlvuDM2Ki1xPFpJBRZ1SFWswFgkIaj2i0f4eyuZ0XfoVVdoPKAvwNITlc6At7r9N7+TOxNJz
tc9nW+pKdiaoe7AavswZTLp8+Xjw2hsQB9hQXgfsZ1aS/mVUoxxjC8kiIS/6+Zuql/iFvBgzqUxw
jHCZsSH/xztwyBwfJgo0T2fFrx2g+TPe8Aa3lGSzCcd+Y2PSOtT/mbyA8cJqdn3KCBkV9UW6bu/k
gfYx8qLSHT15ef+xKbD1/7i91Ys+gOnPNU++YmaBm9wWjGHsdYzkd3Z+sDjbpSfjqDW4OM4TZQnd
A4OKhomS3wx0Y41ApYfuTE4clJ7GaBzjR0fTLijwdtkOHTqZVxe3Gs5R2RSWohMij1kHYNOb5GSG
gt5m0TJGJj7evf51X2+um5cqN+76EQ86Ag6OVY3GY2foe/yc6WtaNoo08UxcSCBxTQGtGzTwTsVQ
da4hPn4sQ1hxztt5tQnh2+nZ4wGlfes7Q5o4Uzibnkp9k809LDo314FbAARFLZLJUah9r5F4rP/F
NM0Bg67SHUdcOYRIAdOXlzncnRPVGYsNIPqlphZmUeN5Gi2P20W7jjc/tNxfn6Wni3PbEBDMVy+s
RDRBwgtK13quoAuynDEL6BCTgVLl12kQ/J/DsDYcl1cGckC/6jvZdfWBmS4UQLbME+V+ASXNu5oP
DbD0mDZ2ZXOB+pU+mzqHFPwEiPUkzNi6xz92iD/v/apVj8cqq5zvpYjr5obRB8cdykdfQqiYKqmP
tMZVvo1vji+ovV7rQaLmHzh391htnv2i1r/CeMduW9+vRZMrTfXs41JCwuri/JRZG+p5MSHCTBiU
FjXGfyVfBjHciPREVIfFbB+v0jIZhg8mp2qTirIgbaVex0/DA40QuQeyc5hswajfJu6dyxbgJRE1
3BoT4cpRIdH5SKJ0buTVJMsXWyVr5h54NI8XG6pYyLK5s/FGGwtiFDwgjKwQrJiBtvVGB053YgYi
30ANjw32w7HL6GMuwhQAeHQWvqhEzTp18YgIJ/PnS6kxDx8qgNZONEDHNohcDpPcs8n5Qk8SyY66
Zr+p9vcwP2Kc5WWX5iSPpFR/6Mx4tc33nhSyJaPcddnogDj6uVw599AtFXECpdKTP41LJValX62c
nynaQF5bVOdEkKOeS+Yat4LEzSTRbmLTdHTjNIGBaytl1xUW3LJB1UadqgEdfh4jsGUfkoaDkyMl
C/xfwvXL1GXcHKNZ6vQUJv0h0gDJiQ0xkZWTINvC4I+3nVUUdGJnCEnQUq7EaiX1mPyNk6OEJT+X
7qDgL/aEcmN64KEpq3XCBZLsfv5F1GlyDwK90mUg8YmAh8qZEZKFXpBa3yRnnWpHfcygeyuQ2+Sp
fhbW6f1guiwUhSInWDHk7rERkHK8Pj8Ib/5Z/G9UGxkb+KwR9kQfljDtEaw9RjlJXuFg0s59lBmy
y+MRlM9+yhznxcL+ubg9Ajhqm4WHJtOOJx2Mxm3a0+hWsD998j7gUXG16Sd6Kw/RovTXJDaWjaaU
N5qkymHEsKlP+0d4a0JVd6r/hzabx9nf5dHSM45JUDA+egCCWJlyJ0F4ZBsJCSD9abEdriBUSwqK
ZvStA49fm1Yv5J3F5gOmz8WmiRiZdOVWwWdTIfBW5uftNB6cJeB8IbGj8y4Kd0nhhVPi5uKS4GGb
hwsZW3BoWpPM5AXS0g8wrmdtLxIjRF1N1ljjo6H/8yGD5km27x0NcgaZGBqRlCPMRYfXqy9ZXHYj
IvdVUvKvFhx/l3HvKLAzn46sFWfCS3aZ1EdTBfLMRrBz8LhwF9YiJ+lnPc48XLXrRdCcL1BNi+av
/rNYz08gKoo4pkRvxDDhSzLgYKTdPLTNOf73WeYvLk8pwowb+4S7+1b2iPseaiFkHSlIh6nOKD7K
nkbK/lFw4rrwHW8207gat22yfXLQfLLGatw7JDtcm6rAD3bIvS0X2lXG60Ep3CMdB5MlKwWoj7Xj
qOxyztzjdI1+SlWmtEGfH4Mpp6nBwLDEW+TiWRjtu3otmV3f8NlWiT3x8+uwQH5iKT2Px417XlGz
f1/9j2MmP6jT0xtiMe1MkCNnPv5D2Im9dK7N4U6c7fBinaSklmDQMFikhqvIvbzqPGUSvh7x6n0W
Byo14wCgi8pfyux4iRJY3DeY3TAWYevYJdmySWInm/9x1SwO/B/3uGRf8PtKHK9n8LlWQnIiqRk5
xQNuosJga7dkOfuRDrvPdwV9ZAvQTcZrTV/e60uiuceMv1XfHjDw069en+6WeH5J0uMo4UMdgiMX
7jZDVtseuSy820ZTqLBibVaWUjim5d8KdCekVbRsrPbOsmpk6dBsV5gQOsaHDVPcP3XrwEY//IdL
N0IDlc1UgYFDbF0RyVJ2N+bCOUTO1aQ9bG4Y9CxUPoXejJGZU181FpTuxSUJpa8Ha62yLmXVj+jB
+NU9qDh3w+9dnlyB4QeNjM96SsXneBOHjezk3yvG28rBM/K/ZlnnDAuCLN2okp4qBrLn6TGKZtvh
cUJeETE6O8f8dmaArRxZZR+D9Uo/BESjND7MOLjEEMPAyNZ76UcfVLW4MAapyJHO2sVbf2/QLg/k
hMQTPVZv8NoW5TjAK9IdvgkQs3bo20QP7OKJn/Cs/Mf+h/xSNE8aawBqO3kZUuttiSR0gdIQtnNn
jiYwIVeoemSBFkYvgcmFUZ8gziUVskzrSiXzTWLoumvBYm8so1wxxRxpDMaA54ZgYlIa2x5J3LXF
LPgqJgytvVuvt8fGnHd8+kmHq3g2YCRQW0nPvN3V8QMtJas7xAH1nUf6LHlddLoXnPz4HCTCkDTw
8yZHoVOJjOvJpvtsH2e7g5PvCIYmmbjBjbOFqvwo2tH+YQ0J8Lpl3xRBazYQYccDO9cQbE9DM/oP
7CNRH7QvISLmfeChbYwHy3AwCNSJEyq2vKUljX7dHBPjI2CHvCbad2SxgLhYubDK4WXSxAhAB3jX
Bul8t6q0aTQIgrDWvcBfsi/2joPac2YrzEMoqCTHUWos/S2hRgdRgwvP4zlQS04uyfoLVVJuEo+E
MeRLAzGJffut7yKgLR8FU564XeyrY8t+nIWhFCje99Uxeb2Zpmz1rxbwjwp1Qc8K6d0ugoiYlgc4
j43xkNVUqReJXG/tAAENB8VgJz874bsBb7rIhK/rbIz0XYhIdvHoxLsDEKi9epSBxyWxLgjVw1e9
Bj3lut05981Yxt3aQBdCNQc2sZ7zkZ2PRk85t4kjdK3l1vvnPrFmmnmA2GZbXC0WgzDUA6/gYZ/D
Jfh8U+joX6/A7CfGFUSSNQNOEIotD9Rv8ARnYiD+hKRUo957c8wLnQgnZsDGfnL8CXf/VRsKcbUj
cjmnSHcKsCS6O5NjQVGqd4hYJvhqyRCvyzkZlnR7vesRpf6sNjE0AkCitNUSrFtdfkw1CQpYq+cZ
xpvpJqmHtc3HCPZJNjyM2LLZ9Z3PgvuulvC9gsIaqmlt7215Yl8pcUknaXncvrEX+F4maNWbQnov
YbFLfJ5jHVuxYsJVXbLWzgN+ZeG7EcOpNEygUXeJkes+1unA/SVDSpYgKJXR1gWeQyf5Nfg8f6Rg
0hufYblpxp9cXvjBCvTr58a766Dfjdvbxj8/XzKTO/ioO3xlOoq45gLKWHKPrwZgrfg5GTNrOCCm
rpkDJPcUZxKbzrrz8E8OF5PxJSvTeyEE9xak+QNvAQ+ciRVnzhuJiKkqLJp9KxPsxQHbhBZ0VJHp
Q7YEWGeQQVgNOHfA+j4oAQ1+5pxk9YLvizIaWS5F41DuxuGz1MR09XZZI2v7Y2jN5YS6ZKABoLeP
JnuqjUWSe/S6K+KzVeHiEBw9wqMqTI4EnZibis7FlXjKiH6+f15g+T6VBzSBK2vfjg5VPaG+Kd8q
40QWNLPBuA8BTSpp3ooQouKA0rLRTfqlBnEJ54xjLj8MGO5XQvSn2UKDKZXCtT22hMVkA19SIyL+
ZAwPofuyMYFxbhezGdhd9c6aKAtYe67H3g+QT0I+lPEtKfqIiUL7kHkigQUE4JkRQDOHElz0LEfN
GGxKQpAwOdEt4/I6b2WTCuShEXztaDVCZ7bMbtjRfUnWgdUmL4JWEacCVkiGDgA18XpJAoSVa2Oc
wV0kRIGQ9VJeh9JedRTDNiIpBX7KFGAB7SLuuQQ23ibgMXPjieZfWfxqMt28Lac/u0dbkrN78qiA
ERnMrHzktnrWTLkfpwje1Dj+2BrKkhW9jmAwPlHLtDfYBm+dUhVJby+Pqpn3bsT4lBkH/eXlP5pT
d91vdgnLi9C4fLlGdmRtoxyBXkVQcG5oa+DyNSK99KSTLO52aDJi+yAS/KLXDYg7hO+wP81eGSPx
9cU0lySVr25twgV6c482lF+19acjqYdz+6k8PVg7s/Lqk2Y3lykuBUjT4LTV0kJqY0/S81e+KJ+H
OvROOT31mImjdh5DJof8BCDKLLgpHJT9vOd4FmqAR7CHJ9RJDcfE5kIgpgDX43rMKpaWkF0R6Pus
10dc5dr1yQW1fE7dkmZK6lFDMCo8sQ/40Bl7MMfWajW0vsnS8cmJxzKhMHtgN2u2zqYoiSsmcy7M
3F9kNHBjN8qkyu36n0YcKMQeE6C3jH7RpqTZ93tpj7GEISeOcVpnqCuKB1N509kvkb40PFOYwzZP
NiN7emefN6HZRmXcUV/WZrNCtT9rl9Gwo8HeO9ldhm7jf8OqKARz4UCisn7UlGLkIU8lWLtnqmiG
MAT5xeUDkj+ysqj0+d4aGNIyAxDcumy7lgUFscoUaNG+YrDcyABfd2fv7nsTyWYfgniF4CRzBHfI
QcPQljbj3AVPt8hBQl+sYY4Bgt+xD082xeYsmiYsI+VThda95C5WyovAoP73K1DYyQfirEbAdIUs
r4TDBzhvWTCwxawlFj4Cg/ShRNbdZOVS0b2swnAovdstSGfvjkSIDSSzUfRNLH5wYJLdanwTPfaL
chLpzDlOrZcG1wF3RsDtSS2ZNSNGQMC1tue+S+rWQzp0yAKs2eWPloY/kk2ZsuC5C1RB23K50Ow1
BZ0NESUZnQFozUtVUZc97lCMWJzgftg0/AE1JD1N4NAEMOq3abpIOHSmQUg6oEhJ5RZ28yq3HB9A
oeg48bE/17fhopqBQC91ocWbYwlWGpN4XPMjvswqr3PTWP7v6EW0auf0b4VTaMG/Sn6u0uYqdW2E
HMhluMHh4bxo4SgMSHZBZOLoS4Rs8b/8gfsmJez/kGt1EFDq8aaAsNOX1m7yU1FNqFAxANbdqpXA
0fLNus5Z7NxXE8z1xb0EBuAsoMSOYVzmK2hbE9dSlKbbcI0KqP7FhO4hHby4c7MbSHubVJRjvxEC
4U4g9z3cVi9Y2KQDWMrHdCybXXyRSePQaBz7dtYdfOADlnxbk8LUMQwgNcutiEc6mo7AVcfPTO9c
7HHYl+sPViDjh04lYxaFCm7KI8ECwow+VcGRLn9vh1C3WQjD3pkwRHZ3ati1nEBanjBpHTa6SIwk
Vzc3+tbU0IC1qe6h24ZpnPTzUg+tt51RDnFGEUrazLMjz9FPHwZz36KjZevLXqhXQ6fkkezffnvF
EZNGW34c6sTCkdqrjJLscwno26JRUejfox80kuFIqmvpTrJlu5mSika7LXO1m3BSy0HwtmRcRFHM
TrepwK8x4aWYWRT10Xw+CVp4UD6lSp6Po8cs0dvHRV739HbX+x7oQIRXUtJUeaUExfFqPrpLiNKg
4BhoaF6TcaSqjPNYaV2QUKOEGlTVVuO4dDpkUiSoXGpMICIux8lzmLcTtyXOFNLrVZaseVgVkZ+a
u65j9ssGSU7nALgnRMWwYsejbnQDiio/kQdAD/2p3zMKiawGpUMH/cwxmBd0ssfClbcQCCMHmeEa
OSCGmMsbHsGPz1WN4chDFOEW02kHV20T+DLWiIJ2jnkE3g86zmEKXqF0VEK9a0f9umGWRb1o+PJU
qJQIRkwe2oGtFJ+i90R+9BgS7tIcccCjtUboFouQ/xWlyxdlO/ad3gCD+qmob7mrV7ROGLGNaCRp
pH7nNJxG53nRc9isgFnwTrJMr3zKBAJtJUzXgJ9a9uPvMaPbTZGwutqiZQggtv2a7bZCWWFS/kLr
rAPj+Cba2WfSnurnxjm4/VoF9KOmkmVdFZfdyYKwOKnMobL4SLuioSRTf7Kvk8trsi4V3bxYfHBJ
PafI9YHXJWbWlbBxkNxw+NDb42tcBXBwYfwe3vAZdgKN3tWptAG9FPXm9GvUqHNW5C8RMmmYhMeG
fg3jThHu+Wvn6nK7aZk6BL9fuUTZWBqA1eIRTBLxNJr7I2ZDQ3Efoq9P0kYGru/UQwBXAkErf4IK
oefDLClyFuizRjv8fyjKPTUc0YgdkinUM4mXfwxj1CHI0oRH2qrXZAvQrtqAx2c18gnLbSQd1FPj
yieU9o+3Vvxqd0XQw2SAnsxAfSAoECnuAgoGEuid6wZRJLZKOGhFoxuxgF4USERLYl1uyX5/ds2P
PEaSLp2D+4FKlXYaN8rM/wkQ8dQawNTW/VfAq9zE71yXXoL+lj80JDLQH62EJgZZDcrlEwvvTISf
w8ZKbAQf3/InTTZsOhYiUVhb/iuohECnCAfxdL4x8xMvUZdkLOpZZ5cvd4PlBWY8ZVz5d5yr6ebI
3eybZ89EgCu/vsRVb9JgfGQEDaMKx9k9kyJtFwzJ+7ZoGrKpjhxGQVMNSojzLe0dokr6hweAlc2x
EyaEJTuu8W0hipJ3ITmNEY/JjB0U1deffBUY5oPYU0Twnl4iWtGSqlsxlJ+Hms45Knj7F0u4uSdz
ISoAluu0g6lm1ksd408GV5KD1O+o6fr1BzcefKodUJhcxFrYcLX4iFpiKnM24pMAZHh4YYUtyMPg
/X94OvlLaJQ3OlLgsA1ruer5KN1SwH8+YX5ABLDkyIlTX8YF5y6vXy48iGPXsc6l/onG2vQi3KX6
EmBUgIRTtwrRRBd2hQkMzl/VOLziJhtXhdGorYoct1FPIqjhBsg/ESyFADNMeiLX7IG98ZuGeaLx
rcAUGa90q3VqPSkyJa5KJ8cUm34DGVx39Xr67Ns3MumRyHlAJo5NEWYoqGk3brSyzchSbp2uNr2b
1XbMj5wlapDPrR6Rk/4iZVACFH3Kpw5uo2PCVX9XB0gcrtyWSagDWfqIZM+tkD8YP/1DmR9iNYIv
Z30eRPMccpl4/ZE3eAePV37VfWkAFmAlgQUMgS4EPeErnJrQuZJFTk6GXHwJZCXfJ/CkC/0qZbzy
YfMyBrs8cw2PZqddcbDlBTZDVk9+L2G9rXnldm2hDXn7oiWE+tF8k93KtwH7hpYcY3NzhEmfEdIE
yYq4CyRD5SsDQ7/0lgHA/I6j7EnJzGprtTO6Uv7ryDW5VkvB9LVV6zsNnTGu54EWn+ji3ESfg6eG
o+yafePWtCrJjp13+7iLIuLxdIue4mUeZz9MKsgoMiGU6/gPyK3yItPnKh6O5jWGmoRz/QrJwfBQ
TadhSZ5RQOJp521ySss4F3b3nK7TaCw2Wpi/rjSfBGNn9VextcLgj2cq34Lii4qs3zU0iy/BcbtM
M1xJbo8WSNqeCEjvjsgGJQTQdFeXBLxEw1H+bOPtLLrLQ1FfHuBMQZISjOXNIXBpwUXbivxG70BL
sYKJ2RboisPcGhcdwxVVSXRNgPjJXa16vVsOl/Mq37IEXW2E1nd8gPVDrmtI/oHbr3FZJcmsYu4C
bNW6H+FLvQy7FcKUG1uXqCONhZJUVUZXYYys/7+VhEACWcd6XrB07djB7Ndq029hCQMdSozYu6iR
7rOq6T4zL3ol3sfYzXbmuJWNcHYYcNNl1PRLYKaImz1is9U0BJtwlDaXKGohhTMukaxuyzZ5U1g4
4NtAdTHot/NXd9IRPtANnOCuD66xO2qHy8xlsNYPXRLeFBABGjJu2C5jQynHjZUeyHuBIzQL5A2t
LcSA4UzqKct7qO9vrw+HMeBTqMrfocrtkbjrcqTb0mElJ+VklMuIu+BfqE9Yrx4m5j/ZF/eMRO20
xF8QA+1+/ojfvi0gcGnc3TqrYwhS+BPr8deWS3NvjiccWaG1cFrJiv9wB1k3r8+CfqIUIEISl42h
8jIuao81U4g1XYUNbqW6TM/UHoEhLGt1mrVLf3CE8qBf2eXnpZPSwUKcuzSYqpU6BwlkLsAX9wNM
MnwQWOB91F1tK6YXV39LqQi3SX8yh3nCidcFx0eJ5PKf+7/grIr548Ig/AE5z3TWPqwTNZ7/2uKg
nGI+z7JYnPQdAySctduDoupvzes2vtY7hGOUr7Ga4Ca4W2G1cHo8AvQjKMCRBNkgSbzBniSVEvHs
4Yjof/tng7TBPZRIc3tbA/3awYL+JGX4sFmP/gSdomdNhpce4BDDHM2Kfm5UIYUX39tGpwXdQnQ6
iM919GUPYSgnuzLxbNk3Jqdw2hiIK06yKUB2hh9THZd+0/wHmQWrWFlhPrSh9kpIRXTmhgQpWDDA
0P1C2T0nW1pIw/OOLPiD7wblsvPJrD/j9ZDjCSauF0hsqio5+fLmOzoE4mH1uuV7EXOQsDY/8YCl
uFNaQHtqgNYz10UBRw5ykHyHGAKtq6KlfSi3RPZcZ+Iu8dRVSjYAmmHLNSeJ2q6jLw9lc2hOshBB
hijRTAXcBLnhgMASgAewiy2BkPILLtSYFs3YW7jSBkDUnRnNXcWVPg+myJEhhie58scgUzsSn8lW
/CX1bqqF5XdhRi+Q5NS7jquPNZSyg10lo7/cTazXb9N9xqlaxgyV3P1yYY5EWwdY3shBDKEjc3sg
wbjvm0WVgFTEDwvUDdGULuSBdTiz05FGgBdvmQceDCseqLB0ncPyHYMhsNwCW0I1YDuAIOhtWJ49
7tulUgv7XjPKv+8qW7PlpqJ3uWXIZNVErk+plNP71mW+VmT65bipfyPZfPo2REQbb913vWUxvK/7
rd8UIHpHrR9mLiCrAa8teYbFQxhpE9D7bgyQtmZRSGE1y4NQ0YwAGYom73lbTjshQIqFVUHSOlST
DwWeLUnOMpV6W5QYLvCvpnIcsuRtn3KXhp8n25vD7uMT5QerFj5qFUFf6qHm5T5phLiOPzRZEfwV
7YlWNkdoDiq+9QAw08iK+2yR1mnHoOpfCzlA3r063VQ9Vfye6AeBMzkDhkXw7SrGj4exn83/CpVZ
fcLmx2m21cvFZncwI3bhQmYT7XOMGnTwumJRn4J9Q2YZkJ3fGohrIO4/yDzEiXhXMr1gF78QLJPZ
lnxZNDrMzsjJKJfbODB7RrgZW1rFOFoZo4EksM50zlep9ndIHio6d4/U4ebDiOUU+ajC26XaIDIg
TvGiFu6xPYXzzlWDl6SjJUYnpRkc2O60Tq/IGxXIsM4LkXPPMnoOlNUBUXiE/JwgWnXf5S62sDXu
51IYrsoByPL9mZQi7xs76x85G+CsW/mhdiP2fR58Xh6zWxOhelo1QnS2w0IcuwZzAbhmRiRPfB0b
qvcdMlFaUxB8AI3+zX4JfFuqQdXz/wsieTvIY2ebj9jLQ/TQ2feMXJluka6eoxAgGKAsK5BOAhr+
7//TMSwysANdR6DCtODG0IOq5VjbQ1M4UhCXtt4oRSA2tqwyQGxrclF/NPN0GqJAbA58TdnLM0vH
KFL7kqsEq+uG9eqetRP15Zf5QGCtgUDzZHKqCMGlOc41ZvJvSmjB5cz+FAQkiTr3VuUilkEVIOir
MsNvOcPV0FvCt9kak9+q/mZdkjGswHnHIAUARPrteq/4HrfGf4idQ0bbmxgbfsKdB3aMawXKYeV5
+0gUYoMgc6DJ88Zd8e7AqjKda1zExDzgxdogBWCWs2HvgSZqKwZ7aznDcYrsbD30pJ0dJh1eAeVf
GCe1F72XHiNUaR55E2jdm0Y6rx6Y4cLSJ1AyJls/9R7BgpSc40gsgJNvqYqxHQm0wGLMQjkuKkch
MBWWLqA3pnxRxtQgw5DVrVkC5Cr4MNLU5Iz2kByopVmtZNslZsYDqz4muUrPSZw3UfXYzpgjAJMZ
SZYRO5mGwdr8ldhi3HAkiDQ3GGNMDVmbbhbr2mMaGyN2uNuY++FDT+1p0SeP+lFNt5AF2sNzpOFI
7EM04psioXfZwtQz9op+4ejdOTYmr5J1EvvxpIvr3y0zFbb+UWcHag+j9CUIsz18f2RVQZMm/UiV
GymNvvvO4MITVlxXakEoS3oje9bZGclptSl+sMD1c4OOb6keWfpbabGnrwAK0S0E47RyEcPeIGGn
bdRZOgLLzYOHwr5G9LoLtbxC95vIiqSrqa0VFQWidxhOtsz9Tlzj0s6pjg7CMVC/SfonRClVHFyV
607N/wI8eowr8rjq7jO96muzdxQy32abB/g/QCzpWVI7R3q6pszAX9qGjOUj0Rv/wDfNZdF5272U
6ztW6S47zP0PXQY5zcMvvnZ921QgUSbisaxSfPa8AsX+wUegmPHnsB/G+151vZFiu3U7q8M6xCTn
f3tI4xYro0rlbHSwTAThOumWE5ci/HDrrxWdUn2+5Ax6qiJpD2kH9ez9xRTuHaejqPghSjs6HUWK
4qmDig3mMIsvQy0DjKd/n87BdskH7fMtZMYCFeC/bmnvQCuSokTtdyyL66KeUc5LsAHUNodiIB+a
1K7kMH6IgjWYLknbKcRt9eDPpbuDo5bfpXZJFPPnWVNhygw4xGq45xMRwMzbfTl/BE8WBM+vtsph
90d2AeasOEgODYWz3CCuezoIy039wQUYDwilcKNn+xtIHTvOk4JaoT1WaUmoJvjiicSygrdecTxt
SAZ7Z8Kj+GWICDQOBX98yEngu/ziCdAyUlJKUVZTcc0o7hN/r4kikNpABVNkcGhJb8727xAK167W
TYtPzNTwOfmNeFP/MYfl1c8w80hYz/6N03Th8AX99jvDucngpdb/spf/LoDS/ptzAli01xmwd6ir
sah8vHXZGYWwxPZHdEso0th4cPgmEwwmdAkYbQQjaH6hvwGwBykmpi4r/k69AIbDA6AchAq9CTiH
+y2tplGPgIAOieUvMWKOpIG38iyV7r2gyTIaF6hy5M4Ha06j+bjeLTJuAvZi5lRIQCxO+hlCxAvw
tE2m1R9GvdhagriDTJ4cH0ufWBOVwXIgn5UZk0ef5TotKJmKHc6wQ933TUpOu1dX0LxJwoONfEA+
074ye5HVsaHsomDmKocgmzjH46grJnIouSbwZE2tLzSvkgZr9ZfH62EREMZL9lHWWLAl7p00Odx1
tgz8wWxKPjxp/TJRSjk2WYazRTM8TVIpGnIDlxsYCTOHPz6iWBPOtF+qOCKLnKnUy0NTNsPILw+r
Vt6zLyFFAjJnInLBK6431P7tZggN2LxbFGbSrElkDOTL65u3SB951ieTWpegt2gfcyhYVuBa1b+R
bufyGU74kBarM7dfnz5berwr+qWXG3MdwkfQsFNALm0YQIIHCyL0vWfr6esBZnIi2vR9tkTQDz0I
CPoEQY3z7GriSGGqjNOhaVgTouHWFZsS77H7g0qlqoiGX9PghTdXsLSv0peqkg==
`protect end_protected
