XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���{.q���eI����1A��པ������E�3���~��i�kWŌhդ�azca���E� ��Q�90�?���~�Լ$c(��[(H-�fN�_2�W�r���d�5^d/�`�ry�_^Ǯӧ�>1�9I�� ��� #�/�4t������Z-o�x8o�x��ڨ�'/��Qz�dL1��Ѯ�^�d�ddʹk�.���ĺ��p�	 ٚ���4k���㕀4[Cx�=��t�{kᴅ���a?����n�K��i�ZU"��l"	����o�{]��B�N[(.���RՓ\���qn�q�^�IGq\���vB�Z�^"��ـ�Ƣ�ä��,t��0�����?K#3,�*����2�����{�$�i��������HLb�eA� 쇧�f	E#�,�γm����z�Ҕ;�*/V�������e�5π_�d{!��|ѡ��q�U~��@�|�It:5�ł�~imed��R�������H�c�n�I��ƭA����û��x�~��PFj�И�
�Ur�Ĝ�
M��k'b���ýM`g@��|<�g=�����t��#��G�@?ʓ��Y	�5��bX���Z=���m7��ඡ"� ũ�5-vt��H���A���QY����6�·i�9_�@���2�bRѬ���i衩��ʗ��I��"��U��]�W>G(c;���_�;����@M�e��&�r�6[��
g[��h���cAS����[�26' ���XlxVHYEB     400     1b0Zo�O���/|_�K���Μϥ�,��r��ve���dw�������Ar>m��9���W�"�ʢ��(���k�+C���JUJ�.S�I��NP����6����cy_	�N]���1Ƿj�m���~��E���1�ֲs6��OI����6���Ob�#F��@��}9�߷k���a4;�ߏ7q��&w�p�T����ћ�"ʽSc(�:���59���t�lK(���Z09�z:nf�GƔ8`�K�B�'Kra~~�. C� ���	�HB�HH��,c��;�q��@ydX~���[<����}s_#y��K��U1�:�+i:���Ce��qx��Wx߂~OC!���6,6����2Pv�<�cZ!� BG�t��섲kX��a�(G���a�IZ��7�?F<$�O�2�/0!��XlxVHYEB     400     170��-\�IW?r�oܟ�W�2�������h$���P�t$���_��wl�`�'8l�b��D���4��o����n^�>�9�ۀ����\�2u�O#���
�p)�э��y��8խ��]�n�� dc<�~�Pt>�$O�V��+��d�Ї�Ɍt�fm632�8������-����3�Ǝ4�P&@���NDU�E�#�����_먗GHK>��,[=D7�D��ͻz��xap�,��Z��3!I�i�����;w�1��PMU���+���Mq����1¦����4�ºnq36idz���F-o��0�?	���h1��84��8�]�b�G;�gc�_�JO3�o{fS/h1L�CN�z�V-XlxVHYEB     17b      f0����Q��[�}5:����!���ay3I�]<Ð�5�[�4 -F��F�un+�
��/P���j&3X��` ��@��
�Q�;�ҿ��h��~�݇I�B��:e�u�n*C����L�:oܖ^�+������@��C�d�H~�}|i�c�tQ��G�O���kP�`k�tK�Y-�R��t<:�7;��
^�&�!'���U��Y�AiT�S�p �,�U��T��6����$G�uQ��L{