`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14912)
`protect data_block
TiL+Qi13P85uc/NbHa7E8SorsVwVNgULpftrO9F7u0gchfF/DUCWjKL4UpaRe+1R0Vpp105LMyg/
tX6ZrhYINTxFAP5ocDpYMcYPJFkYP1bQS4qVJ8rvocuv4hN7UHCuN41YrUQK8y0ISWYRghtBSn6t
JUgfF/mvzIgTkLJ8MU49Fld9Lluee+xFTJhMeAxzDuJjiK2h3xlo0DdEN8dD2FzTvWl4MV6Fg+rI
FVQcQXUXIBLL8Ao75qB5c/KUbYoK0yPodo+bsrWK8H7XxtwVzSE9uzwzBA1Jhoe6NMN2joTYK+MG
uxz6EV3f7u+485getlCWqlswvguHfMnpjgNJqlw0VBaeTsjfvuyLkyoVi1wIlHwY7/LAoUMSTgHc
J6pI5vrRoSp3qb3G/MFKtuUEnomIHMXxWEWdzXjGdp5BXgXJPaaQS5TmJWNVy5Z0xorfelfojQac
nJnDmswuGCRPk+z+Fn4UqlHPKZB/aNIOGFX+KNtWhao2yOvqXj3Nv73oWKz0+zdJyKsVeFqDg/Oo
jGJtdfXTUMhMgIoJpMWtyaVdyi7yszD26fkpmUjs+wzSl+46nLuKov+y6xsc64xuSG07anKc616l
zd/Va1CQ1CGBYHiQ63r+mSdF2x3TYhkxZAFUX7NT02LiGc5KlB8jJgHee1sKzukgl8G5EMagTcvF
FHHl4BlLnUoxltQA0GGqhI3hxc8ldgTVJhN5uY/Jzsl+qXJPDuy1q3+YMSx7UP2j8VDO/gAFca3q
6MFKZHFK7fzSPX7bgdVV3EOydBajVsbh6bqAto2g/1NzPANbgJiOh1jHFcMHRKMI7I4nJ2+XaqxP
jd4oElOl97Yv+HDTagI5zMkN7VoyrYqW/hHFiLRqpUcBaxOXMz/AWlyRNNeLGjsOVC53e+Y9x8Lh
6EawXk6My1f+w36DT7OGmeaF1h2o97qOsSsCa+eqwZmP7irKTVQ2/aJUTTPYbOQ+tIQeRGzygRet
K0X6CsLmNCJ5l7ie5fHUxY5suy9vpz2PUVTP8OqM2Q/1PTIVTQvxBsYnT7GJDWYDgNJJHJU/WLBV
tB7hcMiBJWa1xiqNoIIBL79xTtHoaVe1Ij8pGxnUF3R/QBD6VBIy6cH141yA0tWvGcEPPuuwhdaI
xUTS1lA/NlvB7otn53F2ny5pWAiM9uZ++LdnQuXV03Tjz+o+CSaNOZCZFDuRKzxtMCl/Fv8zjOCy
pKW4hFJdnPGPwWpO+CnFjF/5+SJMGBF9PnJhFJOh3L5jylIdMzkURQKEApf40u5OI9ezLprctbuQ
FzHGFDUoPlwB7kSPy7QL1Q1gxXW9zSEyDI0UpCLlzj4VsCj/tP8o0GbXGtL0Eu/ce9oremCMidg6
ffYAW9kJdZyupOYqHjgW/O1lz8rB7Fkh9EIlXRsIMK6uHmL1lHaUVCgXSipoWgnVL4uFfLNUnJyk
38HFgrpUGyJFer9zXb+BgYpkhyyrP7ieduWrsp+ac/W9pawfovOk/OE8pSrXyXNLI3t5Mi1wykcX
d7EJcgfPIQ7m4gL5JCe/njHY5A4q4wTQFsQVe9G7yBQA9h+AKJO9UVpWpJWcBmlbH7KX0Chbp6jO
K3YX8v/RUQmOZRqaPTV+MBeGhyHOqhpVgwmHy6xddBUFgobSUrUWiQ3iv7ODxiZPetdn1SCWjm5Y
NkYDtDjPdf4ooG//wCEIHaHeA+kf0kMKu36qV9FtjJWZR+xzgR9YJHRUcrqGR+pjJbUm/WdvJE56
hhxnwVzJycQfINk1dhwPhPO1CVKUYk4rB4ByLhH8IgWbI82SI+IwWmOQ5EmRriMM2wfX0Wc4Um/+
fc5YfS6hiYFJynVdfvUYRtlXntv9Gm+u8ZZN+KeW2jwIRQoZfjGOpUTf4nlaA0IJYntskf69tEwe
KIWk1nq0d2CHh3hU2Xwvpp1QdugIVRUkm+7kMLyJZzJYTmbJH/tGTOz5jrcC7dVNHGpaCnApz79Z
xh1St9BPYV4H/HU5OC2RxR5MoUTThhfLgO3DTdM74190K+bGQp3HdcFzuhIx8CozP9eoLXIZ1di+
tfeyMfIVcjUu7A2gABSndWNJriU2/HfcxpB/Vt9sci99wIBZjE13S4stXCz18VoK6eshiCH0FPwQ
hYTsaD23gFQz+BhsdttNQZxm/scvty/HQKt1XBOooDkxGP+GuFE06SOg4kn1N96305ZL2/5PkB+k
kpooy2sApACt8SVYVoV4LHBpocfaOVBqaywUQX8JeudEovon710Pm7Dqjpr4J6iFMe/wU+ot7Xhb
cm+5CaAOah1Zke6QeJVNIDqSvpWHE+HwxK9a5vrtiLmm71otb1udI+dOSJxuLZfLv81Q++t3aDa4
IZCS//dR2NaAYWbtAtIGGsjBCJWDlknx1CkZrLMmOo2CaFr52eI/MtCpeK2PdMsDtCFWOvS745mM
YBVEs0wOwEszuZFmSmZUS+mJ97hxtoPjyGEnWU+TC/FwKceccKpPwZ3lc8tQ9Ry0s9ViGkV8tIci
fBW3uz5p0oxy91iue9QU5aCIJKWoX2vI30hCzrLpbn+xpc98QAZqWKUpUzqzRnok6uNcqPJfWB9L
3gvu8EvwGf9OM750ZT+cX7B6vlsPTAKZGW7hLxVQZ+GYnsgN8GOG2esGaneC4wttjq3M3CHOHq7G
wqs9S58o1t0pw5EhY2HbVWBiTUGts4+VlzW9/fq6Z4Q/tubIOBq1ts3eXWw8BEPklcJnfSiHqqPW
z/PRDrZ8GEJ+NvnSKipwZGbah/zO3mDW7lisQvt09hgIZuLk+ngTSIYmbINIFNHqNDMg66qB2ysw
68VWIhqN4mLTgh4WyhGxkS7K7jKmYwEjmFgUk6nfXHZQOpB0d+XY8oLu45u5uH9M8WTnVC5fbXpE
pltrq0K6h8z+yLhZ/Y1ZqM2PsX+QuC0Z81h5/V4W+cJCq9BI8p7DyskNLPCwge+CREKzoKI4Cym/
siPyXe26RMvbxvpeRGpq3KYwjiTstY4yT6iRxsWYkNti5ccHwuSd9c3QqNhnQKyV5TUIC8Er/IQP
+b1SgM80LP0pUsUTGwQgFXIvkiPdJDAKPglWccCWi75UclnUBWB230EemK/+2aAOtpHdADa2zu6g
1sEOyIkZ0mC73B7zmiQzIZodndyUEzeCCbjR84Xj8a6cx2tdPByEywgDFgx1YPHfNoaOqzMVQnZH
ZwRlFUdW0xktu3B5sFsK3pXYm//pCSM8tZK7j55tN3Byul0O9Yq9EQ69080o8KgL3lFWvTIztvQQ
1hR/z8CzQjHDrG8pqxu0LfRLdKGpAHJr5ZP9E1FSKD0BaNBEbhCAOt0mYI+sL2Gzb/BCTSVixcSU
cD9BSwRkikKucEiTqN9iCQxArAJSYEqondzZVU4Mhie10BuUzp1tw8VMm6dLgAz8uJMhoVgnf8Pb
g3B+Meq0nt3r618nt5hvgOi+bZmVxRa1bX/BVcyf7CoSStC/myvNL2ylrZU6TsCPA3xug/Pz+3XH
4ivQwXfyZu+rkpVqPwqWzTZYom6NC4Ab1mEmKrr+8ORLVe1oudREKXnw6CZNBriakN8oVfHTPi4h
79UvGUwm7t3ApMy9vZ08SjAtiQ1yb+uRa3kgoBdiMHMnVSo3VV+ERwVj+MSEqSI6PiOAiQmjYpbw
1ovqeqUmuy9BiJ3QW81HZ/PWm/zzlwkeUl2bn2LiOkExpblWxxbLwGfY0KnR8HNoFwMRFtDY9Nhd
KF+KRxNGaK4ldXXch+HzuhyjkdUacSh+KlU3mwZ0NBkmeb9zkrPukJSXbQBp+AoqWq6UqIKsB0CV
uhNn4LhLE3rrF1OiMrOXp0p0jT59JHqJ651EqIh8IvQ9ym7iGkC46fYCRTDxXasHBLZNTcrNmiio
JngK5t6BatRQWbnRtHuaV2PrzpTnt4zP+6NHi4Vv4fRrh3C6m9GwN6tEcHz/kTOCS8sz+edSyopG
LX69DbWQxKtZ2TemunKYVXCN2okceyGzpwBW+coDNAl/VNl7uLLTuIm855NEHO85A9luX2Rm/x2c
sB+G37AQ9g2wb3HzqQbwRoiumsKx0aS2dX9ERuYDSgIxQat+0KeLq/11+ozoB4+BkRJ1AzXXMsh9
+uEorHhIuOxGRe3GSKbOMBXl8YRnJ/gCBCRwcO+zKWtPSNP54h8No45P8RlDd0Lx4X/WLF6K2bst
28RUb+pgD7SWJgx12ydu/0d9l9siPDUvl8iL/6UZDN1ZjSBUzFm2a2QSclDX6vMPnINUGKTcnkmb
mvjAkyBORf8o0Ls4sbvem8CauAXyeEipOsgt4Xz65uvpHxUEa7GpyFSpWH7x1oId4tKeyvJGeIV+
gleChNbJ13KEj1vQCgPPH1aieSvvKIy+YIrUJBRwy1v/cqp0BkrVZrbLTADV8/EisuqiM8qnxnZK
9HGpubMEDKApSp3Ed7ntDFvgPXHgimPZ2wtL1PqmESwFEn4DNqgj3OGK2GGJQ/F6TSr8E48bjDAv
o5o9W+f65whKocrtLnxpeNP9khV+m5cF16PuzgblxYQUoBSNwJKzsB+/2phyGA2KNZ4AacUzysGw
w1lfYNdSpkgxcfLRwvfopEL97ZgIw+Wn7Nx3ag6SZctgxPxrVgfSC5J1PD3VO5PCh43546i7OnR0
J4axUOLiBXBkAQoHnTKyvaaPEi88EKcigQ8cW92erjL2iLZPHfyz0SUDqL5BQZXxq8JVz4X2tO1b
bkMhzeESAYoLzVimTz7nkaKbsf2ukRVLJlrHkeD99b5P/+MgSFXQliSO4EJBa15ItoKtBG8ChIlw
/bhJca4x8TD7RjL/OwOxPA/z1B1chiaqPf3xkGMoxJx4P97TubmCcPWopYPa6UUC2xdXQRurggLM
VXIC6QyxTo5SyEE9Pf03eNQEQreGfUBKGCN+yuaVNK+ox8C3v9Q7S3qZqgs7L94oYBA5iazCcmEZ
eum5E5GInLv1kT5QU2bOkl3OWUEkLmyBy4NpQ3iIlhEz0tEoTRyEVoYCqBxIDBiI+tIshVL2l6KE
3fizSiC+bUcGnHWmK8K8aWY4QH/47GjP57Ofik9S6P4AsduahYZ/V/pixoAgsqUgiB/TI6pUO5GV
0ImIt2dhOBEcRc9JSsHnuR0t6ho4qyiMhVUmaNumQkefGqAIhSZU9ZinHkA2ctg0Kvey6CXM6fSQ
Q3nrTGgOYJXqU9u4/vcGSZUkGPz/NTA86oqH/ebmkq4YwY4abUKHNMreXJqR0tab1oxTZ1LZfpHi
TDPnzeQzQFk82YI+3/Z7r7WPaqoeXU2X8ejAV66H3GxcoR6oZTZKpEN1RSY664xjpH6nPbtWe/8P
0sbFoxuqSEly71iGCjivzW4RoGRjLnLXor6s/eDgfnfeRT5lHt7yw6Ee+z79TnZcJzecLMjAuBJu
omwPw9TxmcP7pVP2TJfyE2DkwtUWJ/AFaO4b+tjAFtlCd/9zlEb19S6JDEXQ763k3sRgDPcU5jCz
Y6zKGqabkzSI8v9sQT8ffkbaye64Cm12iebJa7IzcGXKv3Xu6+ZAyT0zdVeuIz9YEFAP1SMwh5KX
tT2lfvrAbEoqKuESwH/VGSNL5KTLBGHL9v+rzp+0oxtpe8yDJStDAGYRCDJLGEnpWHlnRaZrs6m0
9CDUjo5ShtzkKgw4TVgcJcf4jJC753FnmmCQEs9rOcjW5Hj9GLwoPjoY5xJ+kjj3xFt4cavnxFit
H2ouRQig/vRoFgI52zHPDlqBDFZgpM+Xb8C6sZ2SfYwOzqPBUO9DAM9EtjCYxcwG/zPCQZz9AJJi
1MiJy95YQ+0km0GOwHALfVyzlRrNblBJP965p4Hmcr2XOKgP/bqX8cGNhUFW37hfWsDFGcUJ6IZ9
sCXCFppkT9kl1gYmkfpkja9GZkvcnDNCp5AmFpGUl9mMeXbeQH+s6t/3x3mL6ATLYE9XtB3xkC6Z
BLhWG/ntl8AxuaNwUxf0FOLDsm10v6Q9S0AD0dnty9a3ENwCNh35MMrkNRYLwhvTGX4c05lgwzja
UHgBxu0TlfxZpUBG1p4mK/19deUTK0ZdL8O3P4Fj5muQuxIgBwnVu1xnVEUck8W0DO/ICliW3g5Y
gO3xeeO1snvzVGj+s7BfANcg0M9iGWTH7eKF0nY9BwXdG+P0A12y94M43GWwZyPoP704rgdXK1IO
N9woVVSj7+QJb8MyD4BGsL6fi4gICBrPFsP2Bz0njjkmM53ulYyz5nenqc632/G59QDzznv166Vm
dsYEClFrsLNQQwdpxekzJfeqwq0rXKROHzTkKM3XERwjs26CZaRGPD8qzJn8+BoRQOe5tYBMsokx
btyKZqKRFCxDJvleunR17mGRLZ064IvOSABNGc1hUNkVGK5fPyXkezmMG/6fFGMgYIzPF8ZXRfXI
wQlBgfLGTIbrZCPp7jQn/lJKH8Yy3JPDt/pgenJezfPJIBueOZaZa3FgZ6sHJ2/KlILE30zX+xPK
ut2NFYQ6lkisg4cyjWiifoN0EQhWFHDj/HLEFkpksu/P1cw2g4MHm1emBpt0G/8qLSobOmvKHnrV
btVXHI45ryB488eXK/V20bFDqlbEwUxGwEn07hmvbppLp0bXX/mWcw9I2vEoDgW7NsUx/yuWzue5
E5LW+y22eANq/vqn2weJ3u17b28XVphQag9n6BgeAvErplUf5yjrY7d5BzuuLFThmtS5PDc+LvYu
RbghfHvXNBcsdNsSHQgnera3s5LQyqANvN7f819ulVyL/DN0BUcaRys1FZZaC2ATE/xWaC4qTWsY
nX3h3xASM64k958kMTIRe3oxfvUML19TbTBJFcfsyTlucPO+0OexlFp3O367IYn1xtMxNBYfJ78E
cO9ywX02LCSaGswXxP5v608TkaYP/ucZbkZC3TzmJBbgwgMZaZo8rp+eI/xxhBemU86Y0S8cXUXy
+qPS3RFEmu0n3GJKYCnt9bRXYcts5tFCo6ks+U517P03e69sEAiXk+xBB8G6/3o+IhlxXEctwxvj
kmYYsBJy6QloJwiaccMU0gBHfyAS6k5+lKW8u1pOcKyr1MBiAgOPPFibKIFwnJ/bdIIXbFvMRcpX
NLkxpHW8+ZgKrduSulvH7t6farvefPRUJdLNV2vFdf7pdzYQHh9XIVAtTmvjwhD8sln+pNR+ZRCB
SIVVjXC8uYRGYFR3ATzupdIDjahAFURuywPGHzPEUYooldbhn39J/QPyu6Fp8R4LPmZIjzYearAd
OQEuMYOtCRkQsOjFSWET0WLAHzRPAPwwc632+hbRCztDSs4Wsoh+uAdiHZEp6mlp8tMFG0gxJCOv
H2QdqQxTzwgg3oHY+nLFHnVKmtSqByQ3wXIIipddtnFeaQMw60KZk6JvTGykdFZ0yoCZDXbbd3lV
jOekCzmheLiX64uPoo1b9juLujnvhEuB2P4JnmynCIO7wtnN3aaXpv5W6Qz5r5BxS905mkhPvgCC
ZiFjGT0oZC7eUwbXCk8yiM2t5sbDNFBt4IU2j6VrbaDkNCewDXB7OmQ0XRY9I02ZBLUvRK2T8JYy
HcSXAG+e3pxBPDTudTfNsbywh3W2/W+g+eweCtlFFSxRemnilPS8uIwHrAdyc4pkFzGnHeoeb+Zg
qu/SIoFPPNaA1UZOcioL+sLkUQhRB18Y1cyGzUC3Z+JZoZ0vB1Vguo8iUPDe/5KXK2sLAZgKA7mC
befG3pSELCHL4q0pzu13BxVzfdsaiaCRXafDUuA6lnYClfwMsP5wnZK9wFnSqjtqWZnidQdvs0CC
gjcYkPQAhDgi1pW2X45wo2bZqp3ljJoiMIkZJYLPE2fx/UbTPIXODBrvHE6FfRAuoqipopoCY6Sd
8Rn5sbgY9G9TIhI1t+2c6dWWhiB4j5/jwSM0lTlcSYQsRGjp1SoU8++1eKtGHd4tIA7NU3qMlFUc
n1hS8AL/AloIrd7ge0G5A52K7Vx5S81p72CjRnoYiZDy+4kBSWv0hFHv7Vv2jqfDh5Xwt/HY4p7w
NyN5yjPZzhOM5vO3GzTWAg9ybIIOqcTcPTFzta9PiCLPr/Z1KGqdTsinxwIpHkM8RHRj734CxlsQ
e3uKHpJ6gvQoCfSKzZc5ZgYtp9vyQn6kX1TRVOiZfQLfI9ez4po1TSU4X4Rq+pbkGgRHbl6inH/K
3zZ5sfkTbBq/ArLdfyqQD39G4T4T9GwZTt5ahDcLHA4toOOpje2yesL7u6n3N/lnwS7i4BPlH7Hk
DV/DJ7cg9G86Bho+hGEeR1T9TTI0YbagA79eBlvrO8CZ6v/E1Nq05VbMkdHGdGoNBoHIlaka+0uk
SmW0JUsFj7txAN4QXnDAxemnyd04Gbui5y/s75sdOCxuHHVic170y+iU+v6sFvtpNhnW+DR6RnAp
/IhMbpGpqWpbXKUEqoR9EX1BkevPBKbw0Y0cZbl47oSB5nVQOrlmfL8HKha+USOgHKuvRLQCsxV2
w9mrzX1FpFkjz9ui2m82mHmGlMDTJi7LyvzNy67AAbnyClsu1Nsl/ixz025WjsHoB8vDvSd1JI2j
JBI0a99hiNZZil+7tS1919JLjEvT+wNW18fDgtAR58TP2qvdD/LBCckph6+31yq0EzAKr/ns+t8q
7wdMGcoidiscDCh2EWuY53TaxzRh7wGJ7zdzguOfbyoon2j/RswF/sESxFVHFIzSGrK74Uk1RSTK
04nOXL0oTs2szF4Q/J8Bii0ypRW6O5mOhPtP3Z7v7NF7bz2n0ZEQPxUOzs4pOsIZhbkvfY1E9JPp
e2odQtNZOyoV4jk4j+Enu5ml///pKPhF4LdmZvp2wfFnT0j1e1iSLKRA0pe59Sed0TgXAlQcwDdZ
bKYW1Si9OMwtwRYzm5/+4SsZkDTjh+oJBv0gE/yqb7SNfQUBtoe0sNTwecJp/SlmWx2jcnoJuRLi
D4dJ3DiBKaw7OX+LpB2xpjXh8cZnGxYjUhG15+ZfPyBZhPOWgG7WOiLbVoRWJas+ZxIhi0qpUqfY
lNqqt/HRqUGI+FSotizgqeJUU1ApuTeOo3M25Z0dGXJ7vFmhKJk1Kb/HXtj+uR7cGQYfndTLIbA7
s0qLmeiTVnXPzNrBOWy3ejKqPR4CbXkGQR0Mm/PZqP7pa3jI2sbpPDgWfKOoYhwP2rW6TnmMnULq
+QTLt4nSInxmdo7TkizCWGkdmFErRfIsvfCz/xvbsw5KY4JFk9yN294gNp5oEjOciMZEOmQOLitN
T8Qs9wXxBQ7eD4VBmCIAmu0r7bZGKU0EJcfEaJ6bmMkBo5B553He3XaKq2Wzx1w4JmDGG+aqHo4x
mqvwTZsJm8Cj5fuYd/OmDCjicvIkSkIO9T3bnvFKcUed+TXKIC6rOYq+dqP63TEmq/TVkmRTviHy
zAwlz5oJ9d/WGAYEwXLlqEadU05xkZ3CSC+RURv9Wdb6gybdDOkft3CRP6PUI5j11+i16qc2OHY5
bwS7ngTtD+gAkK3KCWOm7xcNhrIu1ZDIzIx9H050y3MNpjX2EFChzQmssmiAL94CVnmtza13wR0w
TnHZ4/SLDcE1GmvwpgvRrxW3LeNejG1l5iVkE90w7yoFAy2KKNl/GvG5G3ztbDSM9pqjYWwHS7T7
F7Vf6ojiSTOsKGD46EfL65MYmrvhbBwtvE4c1LzIbx3xZHdICri1JLGfiepOI4++vmlIOKTKG+dE
IlkA5Ppx3o1mALaKIOfOBojaRJ4FLx4vhPq8/AzhYPpLADqwjd5Unj9HlFl4fR8mhDEhVKAnOiHZ
6lPBmfV3fEFet3J8lGd6yS7T/E1S+h/HG4VUde/R1G9glWZZsY2n6/s/nRZmjX5O7Vs+SE14vIIl
nZIUb8AMpvldOQVD0r5WZIDRycdTG3aOAvG+b7yOl6zBxHHuovTdscdpi94u6hRiVsviAu//PlI3
xfH7VTJ7DceMrTV0CBxbFG/yTqslNGcFmPT67K0w6nWLL0Pokw2ARDwnYF3iBYgFNWgsRzBfh54c
awrYU0urt4ib6u/jduPCKMDC4o7mC0gwl6zDiDZSCUpAE581wqJMi/pevAXOGOJ0xWkCS78oi5kQ
ua25wzVfXBOotAKRm2IV0H1+slHyT9+LpmwknQfwOjjCnBAbQICjR5J4mjYKZjUwmvR3X3GZr4tV
VFwTkPWyeo1jNKCsAoHqyEsVTShs2x+c+3cIyGecfIW8cH72WLfXBF2gF4M3cfrsK35f6TBV9W1s
3k304I6QXHsHxsayXZuTVDN1dwohNEgFQeZZtJIlfTr7TAgNZ8gp4+ywCRz+KkIHYTV4R4tkj+YU
zqjvFB3Q8M5E4jeDJqUkPUEpEv7Vj6c5pQnlyZPypO1T9tnjFTxdSPpG0RvKWMEWa3tbZtmImTvD
VQ0h4LJXckk95xZOvEA8Ys+Us4kKpFEjXSv3KZfhTM1vCCWGLJALfWwtYIid+53O/OtwraJp10m8
aYXrbubwIKs+B8UUEh/xfa9TO0b8avWdkoLwaRgMutDhHU9wXRkjBjNKQyZwYcR8eZ2vXj3M05Tr
7PHWW/z9OETJasQxHCFipSf3jywAFUgBV7slAbYUF0sR6ZWwPuqp9tNTW48Mx+6zsvBTazFNs83B
jhXBOMjHjYmeg3s3ItKd4yh8iMOXBqw0tiKDV6YjqnYzf/2vmI4yy6YhJFfaPHvDw+L8V4VYEMfj
OScWsraYPZabbD78vQ7Hfx/H64+2WnWNjvYDtQoVRgT1VOmN7HMHHMpdkliUeeObiYDRjGSgz/Ei
uHh456kC/b2JpnjHR1TF63hVXeT51dKCqb1v4VZ2JxWWHK0DoP0b5kix5iy981xM+hG9kyP3aSJr
+u+RvgYPf1tIbiMYnYWVabuAJX0BVGUEn32WkSbKNmA3xF5qf19uiIHzg7618cF0DKAZc229vg7E
1rk0J+rcFwh2Xq3bum2YNajazOMiBh4mqLPB5+YVKLxTdVJwUzljXV2s672pnXVCu09zE6zBKgdE
quuR6mgN5u9fiSqeEl/7pomC0X3rt3ERFyQDTbgIu2TEpLQK8AE/8jlc6CuTRo/fz2WM5v6T0MLU
HWklwfTzbxVNmq+F6dNmWpmFzkVoIViXtL6Y9LOdMPsXDtcxw4TXibrZv/cQDBjW2oIgSL6dyosv
qnLfVGTIIUBvdTvD7SFK/iIgyTGZTlxjxsjzLOfQCUc4Hr228F+eYeBhm8UPqM0bF8my37nQhzxN
KVEKrL7OK+oAqhPSQBihud7CkrIN7Q9sVSKnfd6muY4GbPT1lEJ5dOJ0O5Z4giGbzBpelRXbw4Sq
JIGBeMySIYbI2LvetX3E+CvLXl9gziw5rgQ4n/QfSvBzqN+fOX55+OS6gvyQ8cM3k8Z64RwrgZBy
nR7GArCq3OGByhCFtDVpMkH9QkC+svVcnzBqvk0AQl07lyYVnoAGlgZON08UiGSklnoP4VJ7lOAy
cxZpC1hth+nQngeAW6WYIUfeswm/4AQ2IThQDgmkK6zpu7xOx7CX4El40abL4a299DB25tbfbgN4
+TtOoUyFzf+TQS8l1JD+AYOWgENZppjlVL5pNV9/qE8TvzC7uvSXhjZ/ZqZIVfEKY+VqXONWs5k4
HbIKnGJspJ4zaPWmVPkQFgqDp/BrUa1MZPcB4VpqfpN3vcNOgCVz3vSQCN6IWCbr6ONE45Dqjlyt
P5VLsEsf0dQ0F59MbqxY5CW/YAoxLXScBhMVe/9j/Q7NQYCgc0xKyknMZmIgIFhHfx0ix2iyG2zc
CCJS3uJWn8T3yQgo035m9BcGArwzQlsv9IKDgZYe3FZdDQTakeQp8tAzEbw78tbjct+QgxR/NwFO
5CdX+fq4GCvOz1l/48tBTDsCBbAfaawXy1jcT/4hcncH23vLcEf0C/ydvVROTXetmiuQTK+Io1Px
5zAjCXNMCrDJ2+HlqKu1GVOqZlSbMyQN1FcdEQiNLYzt5PUslTYjRewD0tWqJ85+get4hW+X0ytx
bUuFaG2dwTffyxWE5FHZjK8Ifz3Wppeo4+Owu8t2JZv9/EjjHnGL14DsSBJ1NcyW2WYmwv5VEoxs
bZQVoZwS3+j12OuB22laQTimwOHMmPs9xRh7xXNmDZRb5QNWDe4DKFALFA5fICcDKMvDtctbJsFp
jzQGrHSsH5r/cCmGbtAsACEtzdUSl9dJD3FY4/5BFTQD7P2Mwt2YCDTe63N4Igxw2ch6Z3PG+Sk7
Gh/gfB0Deh3DoC8OLNh9GQLdozSyyTFNM9Q25vObzAfj88WMG6UbaOpKTwcEbVBEx12RN7SI0ziD
v9dbmAum/RihZfAf8B9CsrpwJ4BGGqFfd9Eg3nsAUE+uYNm7Epts8JmVP6o/6a3G/3PF0L0gXlct
NBe3lZO0Y4laLjPlwz0fghYFEUgNZzwhsRyOwHr1VRm5GPBqyyz3aqOGU1lgXGeICdhLDcW6MceA
67VroGoDTwRCQZkQ59fgIFDjwQnu/BmutVhmqas1jVfNQo7J+TmZYBU/PTJOBqCGokZHHt752X/w
4ErT5mbnFI2qsv9P9kcP7+RqzfIis49YUuFOzCvrZvVYnn2NB4at5ylezEKZ7ex09kE3bGD5V1OY
fl8KDYHTg2DSaEqBJBUIBputFnd7gZUb5wRVWLanE7gegA6Q3i7p6XyfN9/14oHofZ++XI/q2IqG
h6/6UxpWwO9PoZLB6/lwzbX48H6QO+OrHNA6g6SlJfOD/h0aJJCNWZEVfS/MWRBVF+DOHj/nhUcU
QLrfQZLIdqaMkCUaeuWYtdbpOM00ju8EyqOBPoT/sym6LrCJsHLbMWIxAhfYT6yUqTPvkABmjy9K
b3Yl1hYh8kSg3xPN0Bl6M/FKSMPzxR0HV6NfBMC6zBQ4sRzIxUVu6r1fN94DbwM/M7VTXp6V2mcy
3aGraI5qfJjp1equBcGFCvRAVZZGnMfG8d7qagtk7l+3ZTLMuO9wlasubm1iZUfnMmIzAKKW+Jf7
RFhSdyra7Fhv/FbNBlKZh8x7ppkBjplnCDo83cIpF2Ec+NYwia2NIwYD7tbW8V7beqnHJK1sV+Z3
IdiXzgnYM8TPOnez64BB67/ufeKCXbtz/o2Qdx768GAvVb2qt1jxik1rAQNzuGrEGpIqJ6hbC4dx
+ZhKDkeQ2yK/bQi0kvP/Vh6h/UeleYKKfxNjoLK3jMYFAIQtMg1VVYyrylVC4jMyrkC0aVJ8896i
kyX+HsGdPLwHflzjUGhptbAZ+hfbOL9Z8LpgKpj7HRO5vkOp6nfKxjl+P0yl3gLSMYVWcioTU+i1
rA5EBFYxQSHPMYkfCCJVTLEHUOAJjTGTb803nBZ7I3a4vyFeubBJdSGsC852wKsHZ2A1y6NREO8L
WvVLPUb1M5lvExO+zxb0fOXU/7PjJwEkTh/GuFpRm/8+xBFaLZQ0BGskUCr1eX5FN0EK2kQuoAFP
D2eySPKbzAuHbv9g2+2R6Hr/6dzX8ly5d+xJ37uVP3VfbcF7NlW20WonU6of7ydHGYpA3NWv/H13
9QlMbTJEepSOjeW78o0Ks8Y0Sm+tBBuBDEQ6fLKXK9W+KStEpOMVvCs/jNelWe0CSTNEmb4BB3ER
m+yDUhIFLcHjj1QiiaXk9CjwKqinX0gPOYiMhULSQR0cUrfqiTevg9whZf60+mI8b77mDAbCgaUX
XNqOFDQxAXCo1KS/yC+S2ST8ZDFPQrN2KwaTh+OeIk5lkzqQUSITLf/PBKz4c4yEM/bMk4Hqi/bk
u55BwPm+3hhhzlx1LYkBrZzTnXWj0BYyHgwKDliLHCMc24kl8i3WvHrZ95J380dw981kbJKo2mZv
qqUbBY2X2sJ32C8bGwoVNsStFk0TXcfRF8hJinwIv47k3JWXw7tTC/jnDEidoAzPdVPQcOSrf64+
4TQXe7Ufdf5kHmVYzIgE+CYw7uGCQ+6twteLSr4XlYT4gTioxVv5KzxEWi4G8WXY+jWMoUM07ujX
3/0vYbAU8L6oYbeL4wjqv9A39thrKiuR5IManQeMio8icbGTPhb5Ugqc8BoOufqzpC0OMwKDBRQW
QMX6hWLEtkIX1PmK3A84HHHNhQTnkRl0u3q7qOOCMbujARtq4J8r/kRQgIWuYKLRyrJSngzp4gxu
W4iG/cE3sYNu8gQ5sdBG9rLGE1Z8eRXXGgRfQIe5dB4O4kEPUzcPpXzuORe6KkNB5f//pOdCUvA/
kw0TxskrgVwA/+RVC1HnrCgEOIKgkv3BhTAM2sZGHXedbwQuVPvjcbrhGkcklBbT7sGz3ehoLR0O
HqA6cWZZKqM+03hEl9B3+IIw3ukwDEqoJ0+raQ8IJEEYyEKQTTW9EVwfrwUUufDqM02QIpLrZ206
SCny3CCgrnz4ZMzLIz5c9mP2hKI8NIGlVQn4AIUpyLZdKFtbgqCuLaXlGg+hcbklAlB+nkmVCy54
hufqWWPQHubdTiojeeGqUeV5q9LBAL1BFCZ6RLI9BVx8T/gL0k/RDMNxBKOJAAgCUyifcKcLtrdp
yDpgIGKp4DXEH4d679T2sWrjR69iT/6NS0F9Z73FzlvlVpfNtgIZgh0ks+thwdhkixADi6LDwmEU
zvbasX0cr1PbEhfZRiEGcV31GjaqAtlziB4o9QDiVL0ipfHgz4u8wkQqJyIto6b6N8W19CvEH284
Wk3kjsbVWEQbp3Sd/U3oEk5HmnaVfw6Xm2Esh5IuLCRNFAUMinEAI6ym0lFqmjzbny68N+Sk/LOA
a/C/bNozC9V7faeQLFku304wrv3kdwjOoZScRV1xc32K+M2BJ00sBiFAiD2C5OXbHU7/bPXJzHBm
S5y/OijO7F7c/vIf01Z++rPz0vw/DVyo0y/30U4t/nWnInZ3WHgpXVaFaD+OwXpewegICMZPsBOb
jmJ48xvYwdhaj0KslyNk6u95Zq1pO9ygmHqZzhRUKCgl8LvAvq3qyDkL5Dj9Gc9o02u+kCGgopwG
TpBRIMm7fQm98TgO3TTTj1Pp4PRumgaQVWeatxIYOBgVMkD3iJ/VT/aXllAMuco8KS7RH808/YFD
U4I+hYMUi+c/Xjujt3qfusMQnlW3k68t0EHHoynuILzGTZNO4ueM8r8uYQGzPOOKAU0wHSMBnFcJ
nLbktIax/b8Yt8mE2DCcGk4Bwx+d8LiJl1QB5xapWsjUQEj2jMfiRWtbw1EanJgbxV6sa5gWQt77
E0FR7CJ/EhQj2Jp6rlTTjf72/R0+WlhawDyuHCaZGcuLjVHOAQ0BX/M2lalZwCGwuMGiYX3HL4H3
UG3LO/oFIsDrmh9VqpudyHWx8+yMBdGkj3YKgdUNoYu0pN1T1FdKiEtD8mR8Ns2Hb3BZ7UktHBgW
HeIJe8XOnTfp4euhPIQcJHwPIdaCedtws0nByGMYCp/tWR5OI23RDtGE6h7qZOt9A5+P4XhS0ip7
p3saCSWTxBzorPnFAD3Ae9Ik5DKAHotjFMNSxIgpCdX8BnWAaleR8UsZ2Mn95UK6Yh8Y7tTpisBA
4J2nGh0NpQ/oNVtRpZgLf830/kU+9+6Wjhyl3hqXJ0YRIhxqXdyM8ar8u0vKVKVBQg1qAwkyCOtz
BtvX+nEUZsaTJ8vdkt7BqA3S6SLBSmfAWshPpgUer1x9HrDWsrPxowKgUcTmwB4rdGOAnzHw2fVf
7YbzpJx6uF7H+EGgimVfqtF7JZWfQJpbsgXS/iYl/k8uWfDNwM+mDF3MD/jv1B1iK9thLDGNPWS2
HAJgd4tPyYiyOV1I2Y71IgwhO1m9hj88YkdSgFvMA5NQRJbHfjH6vFui33BL3P+Ix16GhLg+eX/z
q/AXV5Eyygi5ZbJG9SjPHoZHJYZwhDUYVn3b0pQG6V/QOYr+nKQ5ECwpgndmQcw/LZMKRFFxsVgQ
RBy8Aeu+pwKTkwtARDMi/svN/JJpmpv+wP8RN45opy6EzDZa9zyUPFqwepXefF51A+jz0UERga/5
BqJOKB3ehhXngoSXqIRVQLZi96t5eYQddx1/vYFK7ymJSTU8GNGdtHOP3jilDWUFt1S4DO4hv1XS
FYEKsuHFH9C8xoOzFGuV9beZLeYzNsjM9wyjq8brHZsCLJYH0Kou5v7Gd2Gy+Csvvl16JYg+aSz9
7vbdNx/zrbLx8kTJHFdK8qPMQr3HQkEpqPJ91V7C24CdNDumUkUaKw/x+8MhyXnhz3utqjgJbW4w
rAVcUm9AfVK9iLowK00lFMlkwEW1ifIsYUkY8wQglDcQHQ+nSZWNQht/Q1kcbGqw75efclzJfvBp
df8YRbj31V+WCc1JxezpaJTFXX9yrB/I3013eSCm7A2o8vI+lJ0yoXFDntR14TgBUNLyS91J4lJ3
N5slu1hjThqD4p9ZWDy8eDfDcYTknYdnaS3WhWZZ0sdh/Yo6xmNlISbBr5KksMN7DgvSKZywcc1Z
a1FfSpw2OJe6bbw11FJKiQ9lCXCHFEOMZD3J8Bx75VFrhErL3Hace0BoKOpcudB1Hgx1kKp9A19r
fA9uB3V9UPiH9qb9BepRDCCqE6TknLNIyOnMfdUwkaWFzdVj1IVu8HIT/9niM/yiTY2I56ToPbTJ
+H5JDKrc5Gh9aCbNgGI3ORBIEQ3kZ+PVCJXQ1pGiH5ZbBL9KDO2aVM4G9LPZ5/XPoXcb6mKaxYFq
SvrnKinWhvpkUzKO4O9Is9E3Db30+WicVCQGlGctPD1wPb+S0yX2JjYZvHmH3PDeGdkert3jNMMu
hWsE+/n8/k8MjoXexU2v0om4td/GJf0DMGLIu5ABqfS+RPdh2i6kftIFzltgvGkATSYQrNftnG9G
gARiY9EMxWeRnFFL5KalsJOKXMtnVbXMYeChKtENSsaxyz+vdW4vb6wmifvQ2GuY/BphW9zMQRsi
zHrsXP+i959LGqgDhTf0vJZ2qwtiYT5hI5MuZjOI7RiaG5GchRmpZwIrA7uygcs1Pcrsr07V94R5
Cy4NKRinSHfccfEGFWwewmQ+rvs0k6ps9JmPc54t471ckj7jVoR33mr2ItdSko7c637RwRcra/v5
oYWva8ZkRceE/qXkfHZvGVX1e7pCfWw3cSbAlX/I3C2j9OzJGWRzabPviRshCXPDeqJgtRQRi0cp
yA9xBBhYogaFA7UAzdtq/3evrLdAyHIidq0Nm+wflYGnEml3OoBZFcxqaZVWqo1qPqOty38LYw7W
Dym5ZmErsFrAGWs4UNBiWi2bXOjopCEEnf+A44JX+P5H1hdh+7B19yF9oeY+BX41S60Qfc8gAnA8
bVwcGVfFVmKCcJgYlD70Trs5fdw27418D4pZWWMb2+OW35wOvMcktPdBwafAQ0hLAI0r9dIvBitX
iQXVCFmrqbRZLMkyA8pFXhJ65axXBYJjmJStVXo58vIBDk5MX4G0iHXVhEh+veICt63btT3Yidrr
iIPyuA+/SToXQE9xwOIVi1sMhEzvUl4Y8cPD5c7E3YxEkjdX43E2cw7K52J9QVZVvGLUS/pohNlc
Xy2ERtcu8K0JLxsJpwd6NYl6VvPEZmKNWnPPbqdYPMdQ8wat8qVLKGblwRX8AxqJNRG644G8ErxB
OWCj/2kYhr+uN0w09HcdnjURX2HEPvAcY+aXF3DM3LbhI9ZIwv4vGn76FfUcTkVLCymMFO+W0VBC
Q5Lj+V3TsHhkFXj1InqRJu+B+uqBThTLDAWgIFiRp4EHNepHmA+e5cBIRwtCy/gmhNEnMzyaLEfM
t/g7KbeSJzb2v0orES7k67LAS4Ng7hMxHoOcXNQTnQx14RAUz6FAo5uU6NwXaio4z3bjh4AlKUO6
vOTQU8ShFC4mgULBXRQhlc/oLjEOFd36RdvG0tzvt5DfOtQ5t43SA9C6/FWXeAcix7XOhfiyds5u
OGMi/1RWkm9wF+cLS6Lgmdi2GRUpkTChAhJVHZR69244JEeE4P3ywQE8Sk8rkV/YAXLkk6+wKco3
fX4Fy0qo2C5uB8OoP8Aq+RDRey7KZZ45j60WMqh7uCvhRVdVUr59vTOQJqe8zns9KcISYexU3edk
sfi3ATWiLwBIwXH5OxdQNsQoYb/bxA5OWAgaX/ZnJQULqjOhcyldemO83JwtoXsIoOdW79jTZtIq
ivzkwjxrc58IdTedcrEPcKGlhrnAete07SulieNxWW3Z2dkkUR4XjexcHY50cHq4ynd37ka8yVjV
OnHVvsDlCa9giuGU570Y+IRW0eik/6rbIOlrHQWhHkiI7EZVNXiABeyIjaC+TboqHEOrDeyFHhJC
B3qNXoZNXgik/ONu7KB8OgKmACKA90ObjsEV87uzJACr4oWbt1cqCQv08/gc/+VLHCmtpWBIpS6Z
6QUZA1p6Jdeu9D7IedpYKoGpxqPmRfSc8xm+h/3DYPqoCSaZXjl6o5YYJ3KhT1P1a3Xa82huIC0B
eNiD1MRLdNIbBBM8Wfm/M4Kh+CcTEWjAef6vWHlThnqAx8J/0jzEKDtpdjHXlj3ljNYvgwKz4iX+
eAfi9RV0tflU2C1JSI4AMuYHjTQ42XORfZz+0bPX+s1CBa7V36VHVjC8IXERbJfQ9bIXfSZmjYtZ
7uRSaMZ0rhd+0drtkzUZrG/HQFRdWITADSGWChfRo2lfZBZDWyioTLwUPyll6JtSlnAi2+OEdKCt
pm8W9rsNO/CZuhVL/wvIpk3Y2wPowGB0g/0NVVr5Bs79y0efwhO0NY39lBzNT4RVQbgnPUDVPepw
/Fh5/Dqrld97qHavMcCgP0OEoZQULiVSvPCS2WDXnwtTcxTaADs+Gjy4JLYmmu917rK4pz6xpGMh
l6jj5hnUl5O0H+YRT9WUgi1CZLUm/+HQE+FR/1SvFX0ZUg5MR7Q0IeUwsEiCIMeqUlRxEhrIngUP
f/Z8lWE1ebCGzB3VP4z5KabbzK9QBoRLFYqFV0AmhKN2Q7fiCcbqhQSgL3tCbOdde0L1hqWmrZw/
DGoD3Z8dNofMJlays5fMT+x+NC53+MAD4pvreTOXurVraFO9Hn0RHIRkyxkpsP1JkYh7ixpmdqZU
9k1ceGITSo6bjW40shSx+hbd+E5ah/ser5FvWnYT7rSfKMqMZOasJdZi1EMEr1izPGQYgnhTZr1H
n7SWyrFUteH1yYKDEWInYfhHwWXGOfeDNnf4P0MtT2bjknvWNQtj5wyBQ2/dTut86ICbgRnfSRd0
rbTi9PNbpjRqTyxSstHkxViKEIkf+iY/Us7pscY7gBFWc6HB0cLb5LhtwaAhZu5z0rdMaH1P098t
fMw60Zfgq/2PbNIdr5XDbhJfxwSkdxYDe9uAwtAvLBMulAg4dhdsb407+log9RfnIoppLbdLO4DH
fztoFfcrlP7uRDrbBb43AZxnRSGDWfN8CEEtNhOJ564jJjdzYuVGiWw8VjFC1YZiTsfdommDHwo4
7XEn8IVY3hGamZM+awZf7D6g/65Hjpj/lS3SuzlGlWipNMOi0lrnoaoSrvCVdUjCBSQF/f9JsDKS
UcIxKjFXjT2Np376MJf0n6c7MdxsYOM1EaDm+MTgxjsezNyWjfFNq0AvlLwVKCUn7uOthTDteovm
b/9g10+aaxsDlKy7tgIn8uEmLzdFpTnOf1CIPKwfPSy4Z9A5MTtINYTMsFl69I9M9GSo5ehC532I
ncqnwBZSLQWMNItIrGZXG/h5/9pqXTPQUY4blKaKpI4t7gFSwyrimxZCc8JyncFkVdyhEeS+5utR
KY62AaFoB8rCScxmfSjVhHj6dGMnzSY3MGc7Kuygmg41K1oEJ7R2A94dFB2eNiSSbLWuOKIJ2+WM
yM9LQR8J1nNSEiqaFXf60Z/FQhWqjKDIZPIrtixPcSvRDiAvGdKqZXVWkYaX8uL4NynWlNkyOkrc
pmDbCFatFj7W0qiylsd7zLAcd2VfhjeWBbbJksx/EFjThUh9CrK3/Q51FsD5S6/pAJ2IMlCHS4GO
1lg7yin1defmlO88x4jsL4gPrZ2YuBXkXGzADfzB5b9O4ro=
`protect end_protected
