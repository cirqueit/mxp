`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
1rhrly/JiWdZF0abEWQ9+6v5vFCxmAq1CuPJF1kGpLMpZAQa6ENN8c0BdNcRYbilom1sCozLvKE1
fmQNOz6tLuDgmkiCGIMuxO4hIY5g2UQHlHMLNUsY+Y4lQlqUcGbrDav0G0dHVXl0WjYRXzBUnLFz
fS6I923f9b8qsij+zYiXkl4SchzBY5GDd2YefSvU3MQ70YjI+zUJrz+RKlJ4PVJbu2u02Joed6G1
+Oq8rlW1Zd7T45hb3HHOgGBhYizTYjLxRA6L+H8aQvUkxiikSNB7FLfywCWcclb+pL3nAFveiSTD
6jTVPIw6HM5BjqZKA9/l/8X9ogZm7Q7rbK+MbOB97eVd22hQrNf9ln0sHJyq7UydrYjV8nhJ5q/e
0CfmXM0zg5fEF3iUzDwzeVI4dxKzL94dGCw+KWExUFIfh1zKP4/vxKcc6B2KyGr5qskkNGAu/AwK
HrKGsUXnJfSr1UAVASbkJXy658o1q64Od1dWRWED48TafTNLsaGK1cVKsW2hJe/qBXQgvcvBVQLE
c2Jnfrk9wDLVLizj3fQpkYWCqV3su2K5nM8/EItQkKwvcK45Xaju6/o8jHjTkuFEPGwWLlTnclhZ
rLMuR1GiG8nmuuaqkjriuwG1uko/KIJlBxdRp5q6OZBJCCEEvv7QZ9knLXoVeJkhP4pXrhptD3xu
VchVMznrPpqUtZGSKyrP6sIx9SWEyjBtHmUlcZ5FJDAzWhvlVemGdhLOTQSx7BsNBDy1rlPOq5T8
ZnHuMYqiiRJ0QwJbaVgZMbydiHAC5tB6+9JFoi/w7MC99069aIBJf2/IGLJDzIcWptZaN4RNLbu4
bp6QLhf+/FUPID3NM9goibvI2lgavu0K9Wq+wnqyzpaw4CLWEgZl1YtOOgiaCwN7R39XOVhS2qn/
PqSPGGvQIoMYoHdFtHBqirOfz/5KQWOAXkDDjKRDwkUtzqhNgExZwRxxk3Rf/bGdJPbhM2Bs1Dkd
hZc2J9bVHUZmGJ1QfzXiSJFAVvp9CZUTODmaMKuWmpjkdE5RFZb58RY2YT/sBX7ga53BOxfqfJ3Y
1hgq7wIXtnTv2Hg8V6RR7IZMmL8eETiByZ2doU9+Trw37f37q7ouNTyuvzmh3qh70yUKSTZi8tNe
tug/ZXRXyLHxnKFCrYD14oQbLpfkfWHy11Trid6mse4Q/BVU3NBNiicWuhRQWNl9PHJ23Xml6fND
v+9PT0zA3MYz9ZiF2EDJTJ9SHR9jsIloiL18jZfpmKMsEZD/npgejzj8Z/I5dFEKzgoZX/BERazz
zTZQLct6g+Vnbupsu6CzwPymPU+5ppDIFw9K4j4OB3q7dp5GID/eM8qenXKrDPO9E9OD5hQBMRfX
OkMJUlfC8cU1L3YdXp/sICZJ86nF44SxLjaBjCuCsj9mZp9AuxLRv/aKXyHY3xBc6tGl9/d1EKD1
5SyRgw+ohpgt52Sr/YWTgx5LZZqS9eZMZR7JlQJ0hL4VpV/5uw==
`protect end_protected
