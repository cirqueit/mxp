XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,5�K�q�`U��%k�1B���8� ��I�.uuU�Z�l�
g�WD���>gm�v���H;J��K����6r�l��V�M���CVC�V��G�xv��h�)� ���}�;1Bl����{xjt��w�e��Aꋫ�d;b�^�k`'�ާ��;x=�(t,Ξk��|�ٯ	���u�̒��ǳ2��s���A�R���qI`��m�+�,w������7v�>��T��b��Gބ�e��E$_+��k�j)�G��a8�#ӿ#�9*;U�~M�eE��9��X �}#p7�� ��Cfp�1~�  ��"�Srn�d.+:�_�	Xm�ǘ^j���'���/����`2J�rKf��l'NB�J��=Z�^T֯������4�L.V��IӢP`��~�l�ʛO���!.�����Q�y�sΝX,F�xX�4iu]X�%�|�0Y��=�V�y��}��r�/M��F�X�q��La�/���4��ni\.Xy6��+C��8���l�G����~7��b3P�.�3a�i��>�!��8���rؗ�7�{��\�RF��ؽ2y�Dn���SLq�
���u2k��'���M̷��^jH��Դ����%L?!���o��89YҰ�j���$z�B|j��`N׀�gLKRa���[��a�S׿���8�����z�U���+��v�5~P0���)ш؇��ݽُP��u�����e��B��x
�N�Y� �Z�~�(��n.-������3�ٝ�XlxVHYEB     400     240�G�D��f2��U������P�	�1�p�W��d'�Z�K�xN���(���Cx)]�)t����%%NO-C]�������y�w��4K��+����܋atl�ج�;t
�!��V��-(�<�������	�C�.��'	��*{�D84�}^��HZ��u9	��ɴB����ȅ����,�!g�:��HJEh�:v����)��2� ���v��;�T�����x_�|��PL<oٴXo<>��׃r�����TN����cRL��C"���<#�	Y�Mcu��l!ϻU8�5U�������q0����)�]�Q2��X����Q �eA?j?�Qf����L���Q���m8�r����ȁ���Ui�=�ݼ0)���_��u���v�DTu��Z��{�%�����~��g�N�gEx�Y ��XKh�hx��BU�6�RB�vx*��j�W�CO"+&�FB��ɬ�I�/;�t�P^ӣ��!���+����.M�X���ۀ?�z�x��^�Z��l��a����7�FZ}��A|b�"��}U�
�e[Q��u<j��I,H��w�dXlxVHYEB     400     210�0��-G��ï��ۚ�fI���c��(2H�P#��H��j�����)Ksf66���k��9Q<��1=_�A���[�îj�گ�:�3o9f�>\�C���qQv<�:��n�����VJ�E۶���g$:������˱B^�Jni�u���`����
�+O�aF�$�>$����y<���0*����9C7�|M�"���6��7�O��3�e��Xi���Y��m��27�w�1���R�GFOi:�w�;P�_�A�%9X�~�jRpf?H?�, ���2�ˈ<��K�7<�g�D�.����˲��I����'�v�N铟�j\��������L<�3ތ-3��p��!\��s�ԉ^��0�;o~a��{�4��D�܅桏����Նj�h��X�#��
���*�x������*T�8�р���#3lf||�쒵�b1�'*a�"A5����8-�
e_OęJA#��(�	q(�$+C9!�6�n���$�[v0��xtXlxVHYEB     400     1f0��ҥ�1�To�SA�'Y�azܷ����_�yX^PJ���2�T�$F������dY`��g�z���k:ZP@q��wV���7�4ȹ��NX�,>hj�l�pCDL�H����7KB��­� �E&6���-?�(+	ʀjG�|��	��4)��i&`�i#�Q�Q�S�K��D��	c�?�km?��x{���+��z���3�Te6\�Z���̃���~�#��>B��%\.�7f�1�V6}p��􃚺�z���s�v��Ѹ�`�գ>QLà#��a�#mq��d��X�}z��?LhV�*���br��VÛ�l�y�\��ͫ�-�~�Fc)�9k�F���6�,��# c�}�b�]��Ț}�D���G=�,b!��E}�C�A��U'�+�	�-y��f/�.�C6mx�3��3%n�2E��ae�+���P��h�!���e�q�x�t�(�i�k�HQ�/w�jm Q=� ���aXlxVHYEB     400     1c0�t&��.>���-��a؄��2%\�x>|��#��<�':- �_�+��8lY��%�z��hE%.�d54�x,H�#���笀ZcQxK���/WD�e������kbX�"�����C4n��Ǘ~[����&�F%��Ĕ�M��w灸?AE�8�H�%�3�x��o�2�̋��)�y�g��Մ����v��R����/����Y\E�ڵ�ZA���SM�ك�u��+��m۴� ��=� �
���5G�#ĝo<��<r��'�^B��C��Kۤc�}��0����
p@�;��ܲ����d���у� PM�v -r���N�ΗP��%\P�W�yP�����v����G.~*S��hK
l�C���>���yy<˸'s�°ȋ+��Y �K����
�*�P���4��2�u�'/ZJ�PŐ�d�p�XlxVHYEB     400     2005���,�TqkNދZ1�ˋJak���2�-��cWk+DH�`�k8N=����⺻WX�8����Ic�̽���9�^�Q6Bl���q�6�kO��PQa��k�@1Oc�o�:�$��=Q@S�����\�`��8�)��6��5l�p�c�B[���2 <KN5��{.�]`����i\|X��C�#@��0�嗳�xkO�$�Ľ?�k��4�ƻ�(��\ǉ��@��y��!�=�VYC�.�sK������8uڵI���z�/��������&�}]ŝ�1�uDH^4?�z{�O�|�_�i�Z9@&+1�.��,�7�͙�a����ǉMP]���{}����m��E��&�wOᝃl�L>ts�S�w�D)���]`���V�� �[;��oF���������;��"%Ab7��!���XI��d�%�i߸�](P��ͽ�z�=����>p7�Q�陊��F���t��Z@͸?�"���:�>j5��L+%�%kB5�A5XlxVHYEB     400     1207�V	�׶��`|���D�O*��� �x_3�ވ�
Oƈ�zぞ� ǁ�f`��ҁ��"�툒�OY�Y�f�A��姟��������#n*o��^�@��)VTJzqS��s�T�?�F̧!�
nn�ĳ6m�3ZJ����$M�V��_|cY��G�Nw�)���^K	���<F�T�M^���ȵ���wd���4��M����᧨�'�U��}�6���������í�Y ��fj`sZ&*�D&�BT3�l3J�7�ݨp>$CMXlxVHYEB     400     1a0
�p�"k���hDn�"k��/cBF	ů�sU$��?����~��g�R�֐����I�LzUg������jO�l��Kr�顴S2�4�E�#��7-�/~���k�IG{��ڕ���7w�р�oAᲽ������ײַ�[ĳ��7�(��l�s�+��B��͠�y��s��^��)ǆ�x�#���k2M�_͗�B�	��pF�V����N�Fūj�����&���@��bO����l2�ö������v�����ԓ���c�Ӵ�p�٤RL&�3���?�*�ur�_V�~����.;7���SFx�C]>�r4R�p��3n�%d_���=�h��|P)X�\R�nd��*��n�v?�Rn�V�S;,�=��	F�q��e��j�u�ȶT+�S�����XlxVHYEB     400     110�u;Z��-�K� 倬�߲�k$�"��}oӄ��-9�dk���qv���L��\<翇X}�W����1�m��k����~��4�Jr��x��!�EΓ+Lȍ.�xǑŵ��^~����J��^���w��Rc�����sFړ15e�����V���r!�{���Z�f ���Ҟ/��X}�n32��}:����r_h�3Ƈ�J_���H'�AR��i����a��5׾���aڥْ�!��|8�)�_փ�ݟc�����XlxVHYEB     400      f0��/�F�Q@GZsZ��;���� "���D�[��q^Wg@�zͬ�����j;k��ɹ�/�_o�`��=�m��ǝ���J��iQ�l{n�E�N �/\�F�ܶ�P�����h)����3HR�ߴ�=I�~�Rw�f6��&ݘ�c���pH�鄂�j]Ĕ�P���X��w��<�1�:p명�3O���ԯQ�v��3n�k���,����c�F��]����b��[�:XlxVHYEB     400     130l]2��z�f�/�p<e�|=����zAl�V�pi�*Mb�pG,b]{O��bn{�M�N���__�.T6�B�����i)S�Ri,HJˀ����qE��~�ƨ3k��5�/oQ�<��|6f�Ē#���$��y��/6[J��%-�B�j3r�`�����,�Z>��5�s{J�1�o��tm|�܁g�7+څ����զS������I�a{#V8��?�9@�T��e�S���#�s�rp�ق���"��ݣ�.�Gv�W5���@�td&:`ԓ�/ԫQi�4�BO�ucǽm�c�ZXlxVHYEB     400     130	lng�h"P�ڥ��јޞ��z��0��jֻ��ە��WnC*�Ϊ�1Eg�z.+4\�e[7Ɗ7­�u�*[iC�@�n�(p_��aP�Q]�����vZ�lb�����Z;��Om$�>�'��Q��a4�?�ϸ³�[ĸ��r�(M	����A�k����Ux�щf*o��[v}�� P�3��P�2sH!��O�:� 降�)PF&Qr��*G`�O�	\��\�KL�X��G��V�1�a�(k�N�SoV+�ij0�۝gҪĦ�7Ss4E&�x�0�����)XlxVHYEB     400     130�X/��2���(;He����c��7����E�'�r�<�4C�k�����	����W����������Qh�e���|1���v�H̟���\���}��"�'Y�0�{ܽ3��=/�� �.�G�@Hun��=�nއ��.D�v������%��rT|r	�����m(�4�p|���S�&�z��I�����O��8���ۭ>��1ws�Y;c#<Vg0;�Bw+C�ȓcl��%K�	v����1&
�x�c�Of��J���O\�Ol+J�Sq��a"S�XlxVHYEB     400     190�]M�3Ma"����:ا�9����!unB�o�*�wy�9�[xPY4��t�G�EW�j�z��N\�Kgjg�O���.�P���u��K?4����m�06CC��6"e&� �y���� 9�ڡ�zY���gkJ �R�W꠪DA�;7TiRK�ְ4��?&G�F�g�G=F�O���9�,���Y\]ݪ5� �fmR�E�:���aIA�O�#G����4C�T��b¢�#$ɑJ��"��P�3,�D��C��t��2����2K�����.n���MIh�}��D���K�x�����(�pH"�Sg#�.q�a�R�ʔ�`J��c�(�݄�l��!v����y�s�'����P�������
��|<��,XlxVHYEB     400     110�fQ�h�y+f;�d�0��@����>ˊ��%I<-��)�W��'�D�D�1j�j�[f�E��*��~��l7�:m�9��X�M�@�6���Nni�!~�
�3K�q�7|�ԥC�!��P�c����n�1�>�ܬ���E�)2������P�E�h'�(iN��T�k�
�Zt��UqD]�\�l��]{6H* w�Һ��FЍ���ڜ8�)h�u$tQ�.�f���9�~,|�I��%��	�����
*���p�䲿r~G�5�n�aY��'B|j�	wXlxVHYEB     400     1b0����9b�3gN�ʎ�D��dpKN9c�M��65��'��:�ix��t����_}	M���3�8���b@��9\���z/&��j��!�7��U��h��y5;�j L��	�&tՅ�G��1;F)�$�q|�� �X�}���Ԣ-�|J��>��;��JyJ�̏��2q��׃:M޴D1��	�ߣ�N�t�ݎ�g���#ҝ[����U�	d�T1f�@��s<���t��ja��V��f}=(~K����	�1��`0Pzc�S���.��'��q� �t]��I�@�ڐr�_]�	��o;��K�<�$ �ʰ�ϐ� �'�FH[4����]�.Q��u�*��*��Fk����_��n�������nA�-ox=�퉃?����,���
�W�&�d��R�}��a:�XZ�,��X�� OXlxVHYEB     400     190*�VG��k��C4��9����ާ����/\����:�T�]lN�P���0&����@�dv3M�8I#����(Ԛ�;����Q\�J*-�w"[ :r���a�IA.���~t��)�gl~��r�� ��%�	��*��k��ӴӺ��y����T�f�C�{q*�?���~NⰠ��"B�T��?Q8���z)VIp5V�����4��X����4r�Ż,���'h渰tѼ,���rwia�ʁ{�X��'?\ ��`�c-|�� 7����*����O6�_�4s�P\�I�ؙ���<.�N�v)Zot1�.���mRb�[��^�E��2濩L#w%w ��h?��&���@*�ܚj�4�*s󧣳�)$���N�uݦ�L������Z���XlxVHYEB     400     120��h�"{�C=Nk~,vԶ�Ŗ���|qS�}�'.��g�ս����!�n
E�,a1�������K��nx�GO�Q�����逿��鈪��:���`��H�hjG�ʪؙ�Gm�di=�������Ҵ����6��lv>�~����;}� ���Mq]�`���>���	�qv�E�l�ԯ�|����RB���7~��]�7Yэ>�ЃȶկĪg S��N��4�J;,�62G�T)�JĦEq�
���a.�4���̦� :�Y�G�l~	Lb�XlxVHYEB     400     120�rڰ��NL3�?֮7ғ��O�����$r(�  ZhIe 6�ͪQ����<K���$��[)�\ҷ>G爥c�u�8)"����Q`2@:������z��[�O��lt/���9q�*�R@7=DA0�o��W�䓾�x�)�X{��O���S�M��L4W�g<���<��'!��o~�{f���&�e��M���B�o�h���t��U����Io��ٯ<&2y�h��D�~��v��ޙ�n�����Z�F�Ei���k-� .	���$��ˏ �XlxVHYEB     400     160#��S�ݱx��+�/�۽���1��j7��8��2���`���M=����o��T�c�'�,��E��z�p��!��Ϋ+�,��d#��z��%Y�\R��h��m�]<��>Q�	�]�f"�6���r������t�I�C
��}Ԋ��2\��rTo%���sE����ʄ輪 �����({���2^�_�h(	��/tuN� �*�l��x�k���J�]����ȿ�	�d�������uD���_��d�E��ѼN1?��1Z�(0F2
�#9��0�,e��z�K�x>SB�]c4��"l�2����'�f���l2�D�����f� -��J����I�"n�1�	�Phs�XlxVHYEB     400     150x�Ų��bԩ-Ã��O!��A��������Cnj_�T�ɩ�ž��We ���1��7!%Aq��&�[ƨ�P^�m�Ζ#��T�'O�Xzj��ڳQ��ѱ-����ɦ�Jf�f�$F%�����ɺ����$���k!��������(l��P''Qv�P��Ke�9�!в�w�1҄�de��P��t�0�7�{�"���xh�M�YIvKfw�q[e��� q�V:����1n�ݼ�}�����&�ݵ��۲��Y��;�(��O/+���T�*�[����53?wmfC��3*�$�v>��ʹοá���O��qz��aS7XlxVHYEB     400      e0GR���qх��e u!{9�٥SO�JC��;��\h	�O�D��5�cJV�+�����[�(	,���Ia��;�YE�3w@������\�/��2+��Ps:n���ܚF��̩qc�ilɲ;��H�\����9f�<�����ieUL�M�*�!���f��I��+k�L	\��p��oҘ�`ޅ�t@���H=�<y�P��ZM����^s�֙N�uXlxVHYEB     400     130��h�4������a�U׷B�����V���a���d6]�O�������{�ו�B��7���K^J7AG�[J��)OsB1>c��r���=;p�P��ڎ���7��d�	?;����閑Hg��@���{�eT��9�h^�����,�:��Q2��n>�� _QO��+;�/��ϖY/35�C�x/�Oj��hӵ!�e�ʱ�-�O��R�0�Eh/��Y:	�&����/��6J�8D5ۮa.�S��9���T�m1M�։9�u�g���?�5=X�7��;!�I8�Fr�D7�(��XlxVHYEB     400     140���3�df�p�	7���9���Ü(�L�R��'�	���RX�Q�^>U*��y��,Nc�딲}lbo��ԏ������4s�a�E�Ͼ"�Bq,Z�=�R=�Z9�jTv�g�,�v�պR��B��n��1�E�d�0�3�՛�R.���뙣B�m ]= ��X~O��{}�-�N�d�|��C-�\��݀F�e�}5/���5փ?�U�Œ���C@��G	�
�t�rW	j0&l��Z��
�-����U
�G�p�6o�c	b�`n=�+3��D;���y�]0r�<K뿾�7g0�I!.��u�2;XlxVHYEB     400     150�jC+�ii�ʰ�H]�ڊX�h{��;b������㪛N�z�S�e�P/%��U���������/Ņ����&s/<e�Ȱ��^���hщڍrŉ��5���@߯����W��j/������tP�#�.#�ɒ�v%��CrR�,���X4c+��uP�(�QT�ϲ��H�@]��l0R�R�p������ٗ�j�Xb�їK�	6EN����U�:��8��F�_�����o����pHFU��Q�$Z�]����<0�����/�a޸����7�{�`�|�Cw#�=�=�T��n��� ���@q�ttY����<�PS������1XlxVHYEB     400     150~�a`x�� Si`�YN3�%�Di�%q�Ք:2�Ո�<�V˫j�M9�Dhtw.�f�E�s�")���m��x�pfX����^�5��(�mcɣx%����#��l<����C����-�z�@�&su���AQ91EB�KqW�8"�a(j�ή׽��Q��&S��u�#���3�^Y��9��R9��o��d8dCR"�c��;�X  Mp�w�/e�J�����%QjڈP̂�R�uS�`�ݕR7�sO�+0j��н�	�KK�<ˠ�0C-�[��n(�~k=�n`���H����(���
�y�5���MEw��.!
���	���XlxVHYEB     400     120o�ơ���k�i\L�A�Kw�mS}e)�ɘ
�έ��̎����N��÷[��"0�f� `�.�EJ	�fm�YDų"ʎ�n�%�LE<�#���J�<�^�*J�,�y�C8 _\���Z�`,:eo��>�)�V�mi��ێ�M�1	>�db?`
��#Q����m�W���@�� ���R̽J�H2��,QI�T�Jw�{�� @5v�d�_a�j9�.��W�]n\hzsc�f6�駍�g�ݬ|�g��1�5����~E�
5�Ҭ��R�e��Odʢv�[�̠�XlxVHYEB     400     130}��%��C�����l�i�~A�*uP${Ȁ@��a~�\�#��o���˗��tQ)b�n,������y���e��-��p���)z�AO�� ���ehAy�Ӈ�+s�l���bϿ��� v��+�0�Pٲs)���p�C]Տ.�ؿR�H{��jh9����_u.��6�����������F������kZm�<j���	�H$��V�Y�Z{N�g|��ll����ת��ǡ����8@�4��4������cXC<�� �I��3y�My'6��^ )n��"ۃ��XlxVHYEB     400     140u�#���È� uV�M������H�����_���C3-�X����� �鐻t�=��Qǿ��%�MR�i[L���o�xB�Je�,���P\�]������옣®�ߢ䂑��v�,Pi��Ϟ���:���l��+n�i�M�>����\��.	!B�w�LNc����2'5��B�`�T2ǘ��Xۚ��Ԛhh�a�!אr��Le��� ������Pk��AL��Ϳ�!V1{��0��>��{��\1)���|y�ۯ��<o��}ڗ*Z�ivh�{j@�*-q�+ym'bPF-;�<p�3�M*%֙i�	�����_��y�hXlxVHYEB     400     120��>k��Y�,���9�{�a��Zl��a[R�`�#|���&����⪝t4�kC.���*�"�
� q֋�0��-����F�f|�+�X7�!���c�<$ױp��:O��)��Po�o����
G�`�0
���N��	_���v�ݩ��jfX�|tm�3"*�кw6	/���tm˺�\u���,S3y����dL^yT�t��ʆp�'*!�
w��eCS�BM=24i"����+�efFԼ!z�
zѰJ�1�:��Y����H�n&�s��(2��E���^�XlxVHYEB     400     150��U���-koG�J�3���YKB�ΆO��G5!�� '����5�f�A�0��i"������]�xh�P�z�_�_W�Z;=y�{��'(�)�QR��U�}HӈX�<?��iX،'5N��ﺪ^��@�T�ҏ��ћa�a��ЛN����k<nF�n8BY�:�>vt</�B�}1_��F%g�djP��?�:�w�u�:ǖ�8G$l�E3��T�4~����|���T�q��8� ���)�T�-Hۯ,�n���Cj"�3��!���(UH�Y�r�pc�A��M�Ry���s��b!�P���l+�-�"n}��XO�t��l��dbXlxVHYEB     400     150����ĝ�f�'��v�싳H�S���*�bIM�3�a�>p��Ӷ��t�L������gOj��QBsNV��F������bBޥ�E���P]`U܂�;d����,��EЙ��'�;���ș���Q܆����J��b��S�+F��.��;��8Ԑ�s��z���o��`�
�=����ۮ�6�U���4:�n$EN���XW"�p}�i�i��t&�N�~8�ڀGѤ;���5�9���m�{���S�N�%e��#O��!x�@�&�����ޟ67�٦��ͽ(����&16����!�P��dB�\Ԩ�HIz�n�����"��XlxVHYEB     400      c0n�I�L�H��2��r|��O���M���&�ӀB��P���b�>�<�����#��2#|bə�#���%��̊��>�iG
)C(r5y�y�~}�X�;3�!�ϑXfK5uꂞ��ʻf�<��F1���&�x���S{�k�(%�ѱ;����vw�f��;�)~|�\��Qn�d�M^�g��x���ɸ�XlxVHYEB     400      c0+o�N����#��LJ�$�ȼ�[�d��n�a&K����Rޭ�E��8A�����ĺ��^^&���{����X*/��� �v"':Y@�������q����1���D��Xb!J1�!xN��T��kB\���������.�Y:�ᶎQ�4,Ŕ�½��`΂<����#
�&6�Qfⵁ2��2\���(�m��~x�XlxVHYEB     400     130r��>��2�ZʷFc��T�jDh�h]�� �Q�����<)3���W'7ML!�����@�şQ��n��N��~f#�+�P�xu�qn������4�?Oz����+�J.�0+Rf�7�n��9v����\��܁�jZ��T~6�
��Ф��2Zk�&[�@�����/����V{�'��<�f} ��s�!�*,'�E��4��4�f|�ę࠺��i��B
�53�L�юE����bJ���v&&rXbc�)[s&�Ƚ�p�'�'Xʥ�	���MWql
��IA
�zY
��`kXlxVHYEB     400     120W�}>����D1l�>$���-9����|�2�"���D�jm����G�߶o}��ʩ���U���G��6�������h6 E!ʼ�� 5�ϛ39F]�۰�_�$���<r�e͗8J�p�������s��1$��h�\ڎ3�(M�+��bf�I��r;
ARA���O��}�ō��1�Kٱ��C�9���h(_wK�B��2K\�6ՎR	��A����ݯ,1�������B:����3�Wʒ�0���M��f�2a��L� Lz�G1���f�b=XlxVHYEB     400     100'��<!h�lR��@z))Dj�_\��E�/:�\e�Bm'����k�Q4+�6YB�)��I�2�����b!�߁8���5���Sh�I���7�ۅ`���-Ok�R�j���I�Ϟ ��e���vT޺���/��`b�6�NZ��Ƙ�.�*��h
I?�"��P�k�`����#����T��o���B���R�b��fb��j!���ֱi�j�s�@����`�;�މv�*�m�WnADJ$�(��h7�XlxVHYEB     400     1609r�}
(qUvө�ӓ[	�D�f�� 2&��+�N��{cQ.B�&�lf)i��M�_��5���*/6��EaCl�j��j[�:-0����Y@��
�����݈}�Cs� �7�ە�6��'���4�DUe���m���̑��m��+]Q���u�S�$`Eҋ1��2�	��aB���#}"g�f�qB��5:O�zfx�����
d;յ�i}0��-}��$��*����HQ���V�WD���xf1S�UO�X6�#�$�;����?q���x\S���׊ڑQU����V��oif٨�+���<� �ۇ؝;3ih/��p	�$�ア~�9|1o�=M�2��XlxVHYEB     400     1c0�@��ˎ̬��&~����阮~�%X�X>�����V�Hct�Ĭ:���%N�cs��U�^�L@���O�'v��S���1D��'��,n�k&8�%��@X�2W�Z����	��2x$QH"����F�ZEʛ<�5Y���K�q�Sc���4)},���:|H��D����)}Aز�����[���6�dH�~v�c���-�kX�6ٙ�]���S�e�)�� q�y1�)�XGH,Q��^��rk�5�>��ꞺOn{y֟s��T
l��|���+�F�?-e�u����M���u��ϓ��OK������7�cX1�rvh�C�z:�Gx�/�nkD8��a��[S����4W��O����6ǵ�ۦ�x@ �c�V�d��i�N|zТ�bxJ2pRY5�����:5�
��l�N�߯��؉d>�j�Zq�ZFt�ps:�XlxVHYEB     400     1d0��`�õ����0Q�eD�9�>i�9���1�ĭ��VG%�D�3gɱ)�G��������1���o�����7!�����o|3�Kc��z��u���{N��.�ݱ�`ٶ�]U����M2dxn	!<ZKEFEu�e
����8�+z�Є��c�=0q]#�/	\�� j��^p���랍��b}!+�&ݻP��0��g[d�H�h슕/��MO�0�*�tҔ�v��{�wH�#8���65�J�����\�nȒw�S��́ux���	�Z0
�1߶tȻ/ԶZ���W�����7]6�v$��mp�c�	ˁ���xT��u 2*��v�;߱w����P�&��>5i�*�� :xTs"kǈt�����U��4���S��Ӄ,���#f�f���0��2��}�&3�_#c;�aOOd�D���"�ҏ���~}@[����Ð�x��yVN��XlxVHYEB     400     1b0�A>s�67K��"")��r�YJ�_�h&��z�'�g7�*s�D4�=����>����D�-Z²ٛw��;ӈ���ix:��P�0��g�� ՜Hϖ/j�ɏ�AS���Ps�����/�$C�������Ox�C;J1�T�*(a�ޞS����^V2�x/Ę����$?aQ�|a,�f�5��K�nƳ�!��#^�B�PB,��u�w+��D�<�F�x���j���d�<�<)���{ijJ�B�hkwo��͡��A�]����������{�'2#�	����U6��׃�T{�?�����<Z]?��K�w�DYV���F�ofXZ�4sB�(_$B�O��\�6>�b?_���kI2�<��>�i��@(��K2�U�B'��!<�	�l��|�k�%���Y�H;���$�b�j͠�Ԑ�XlxVHYEB     400     1a0MX�?�!��긻�R�:�J����!�����wC�%�������U�C���;�}���ګ��V�i᭘*=��y�B��/��W������zI��/\|���c���헹y��'D)�L�YA�8�v&,hA}f*�W��b�ϫ- ��=�"�0��-
]k���G�7\��
���Tf�/���h��&:�F��Q{Dc�=�
C�U�J#&�6�P?p�nh�y浳��0�V@+W�����Ðp��c�"fS�w�O�!+�h!��U|��B�ؗ�i�a#Ů��Χ�0�% �a�}<ׇϞ�f���H�V%�I�D� �ds#��DL�j���z��dO#ؚ���oT�>"�1%̻D��6���C\�Z�D���_c��љ�n	B��=�0&g�\Y����(:X���XlxVHYEB     400     160��H�;�lR�Cx�V��َ� z?���#%�O�cT����,&ǉmA1e-[��v*BVɐ
!�M쎼������?�Xi�yʸut�b,`�;���8,${��{ijJžc1{[�O	k�J�ǣK��K6ժ����ߓǈ��u'��/�Nz��c�Y_EkJO�U�����G!6O�H���G�H��Z���'���a�\�����bxt�
���� ����y M����%!.,`�9 ]�R�_�~}%��l%6i
!�S%��KXV> Q3�hF�C簶�h�jr�P��6�z�5-B����j���ಗ�~�@K�V1rZ*'w�� �%��=�%��XlxVHYEB     400     160���V	R^0%+8ih����6����^+�T��||)�KN��(��Y
�qP:=��fU$��J�K��X|-�f�9z���R��`J�����H󹢼�k���œ	ؚ�5I�I9sf�Ҳ���)��eY�i����ӻ��?�P+�S��B����kG皞=^&�Z��<EB�ɷK��k4=p�σ23��"����IƨX.���*�M�J2-�s���~��1��$�W�L���"{yAK�q{3\'֒�y��L�� EH
�J;
1l�����1`i���N@� �tY���b�'����Y�� �M�H~���)2�<֡��d�dRh�h�n/^>��7��]{'Z�XlxVHYEB     400     180���%��Tr�S0H�ޚ��CK �G��q���v|�gB= KE�RG|G��ϝ�{.�m��?�hؤD�uʱ��Y!W�"��JS "y����۹�>�3^kM�m��,�U
�[��q����|�H�-���ns��́|��u'JɎ�X)n�����:�{(��	C-dM��<ڐ�Œ0��D]�V|���(ʔt, �,�<^��@ʵ��L�ι�*�p��.�|��0�~*��F�[�����>~K���.0^��o�}�{��Tڨ���a�-I��(3k�����4�^�S�m$���}𚋱w��#�Et�X���&�ip�^r_�Ȼ��9͝۰;X6���E� ꩚��]á����Gi��T�/+^6�d��:A�XlxVHYEB     2ed     130~�3�֢�އ&�w�ؑ�U���я�x�쳧���^c`A�~�ӈ5�<-���R/7�"u�U���{��P<+~�동7�Q��`��8>#�p��	��(�`M��	}�11k�\�ˮ�Fْ�B`���Fd�Cʷ���;�6�� �6}��G���6t��w�`Q���]&'?;J[O����V��NqF�HX�l��8�AU���2
iM}�^� ��t~��+����&�3�㵬yBS=�T<�8�v�O��A��LQ\�L�b���va�����\/��1��]	̸�i�E��r