XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~g�8��8���8�M�IX��{\N�|!e��;r���A�\�BWB 742�<Iz�$pN�>��O�b���A�����Z���@P�)�z<'h-�0�g�%'!̿�q����.�ɫnc�Q?� �r�|�oj{�|	�Ly���+���;:�i�~~(��ǖV�с �cj2?��:�D_zI��b�98��1�ψ�h�~�i��[d�m�2�J_{�M+U�	�	�3.zw	+�Z"���8��c4J���o�`�ތ�O3n��փ����RثM�3�I*�o��B�����VXҡdU�Ar��")�ٽ��=��K-�N ���;�!	1g��9�XP��]�s����B���%�ÂE�M�����`,)�ـ��C�_��7w2�%?��ی}ך�r�(���e�=�`!��102�Xmi��3.���@�X��Z����r��R���ǌ나�\,�hD�%�z�fZ��g�jQJm�,� �N�ܹ��������w��c_�L�@�<V_U�a�`䵂���'�����S[C�лB��V]h }%3��z�G��x[���å${�h�Dj��i��o6�y׬1�덈�;:w����Ǿ����J�D�ף�����u�� ]�5X�*pAx��' #�������>X#�R��\vJkC~��n8�
�Y����C���\�#.�#42�܁Z�0�ƶ�9M���)J�e�I����}�'@��enm���׊m�(&,$�T6^`�i5ރXlxVHYEB     400     1f0%�F�N�a�
��a�$��u��~�7�p68��(WM��2h���|	X����A�=̌G`��3#���۫��d"�R�X�%��]��]e�;�Q�9�[��*_b�v��AS�nA=���֋����R���ۇ�N���;�&:�a�qRX�W[D�N��=yɆ:�A��*{[��`d|�E��HH�6+@�Вܼ�~��=���M/�3ᶋ��7_�#oz��*�%:XɸT�l�)�hr� ��8�j��̫�
�i�9�?Fw��U��������q��آa��*�xFi�� ^����������'�}��a��E��g
�D�s��޼�X*?��E���/$�ĊQ< ������R�L��T%���Sk%�D<��º�?@Fv�����9��&pCLG�E��lϯ:QJ}����Mz�\���
�~�7���0�*itJV����z���{��E�d�졝t%�6��,�������;=p�_�XlxVHYEB     400     130GŊ��v@� =a5�E�jtub���x��7JM��Iɐ�cݍ9p���E* 
	����P|���≛��NE�v�$ӈ{H�k"��4F��:���u�#����}�(̿ �j���熔�W!M�	ŝvJ[�-��[nʔ=~��^TJ�Y�ܞ���`�0��@���ycZdZ6����?��4RjѪm[yh���.&���|P}=QϤ֞����؈�g�%0��Q�8V��bOq��eE��&Ա�x���މZ�6��r�m�=��ʦ���߳��7�3\C�|;Z�˺vG��eXlxVHYEB     400     120� �Q{,��B�*&�΄%���5��ۆ��F�7����U$�rR�'J��=�W��u)�1��
a��(aN�5I��*r��]�5�i�]�����|������'����Oej��KA
�ݳ�e+�� �8���I��&|�L�tW
�������[�nD0��V���J�
Y��H1�͉�I��P���\�[9��XH���M�Iy�Y�Ā)8iuX^��c�o��te�Z|��N}H����i©�V4�y�#�X`F��u;����#��)F�R�/p���h�XlxVHYEB     400     130�%�Wޕ��>I"c\�BVS�G�d!������ ������Ar���ؿ�nbz�\���@���QK_o�� 7X.T�K)2�d��P�&����Wг�)�w;��n�w�_�����\�4I�*��[�Eݬ)��l���8��sM|px�m�N���y��b�6����d����,�w��[��hH3�c;<jΠ��^,Ug�"ھ���k�~_mԵȻ1Gצ��.e�tV��_u��Ea6�>���^�L�zp�W���S�[Gws�g��h���Uy����,c�G�1}A�,��aXlxVHYEB     400     140k�3�����	WE|�w�SQ�3u�uj�@��hv��(�G�?3Q5+B��mQ��Ƿ`]�vZK�MGH�d]�S���5���/�(���e\qO �3�Y����M��Pw�@��6%�?I��Xmq�$%������y�6��o�"|	;��&@?6�by(�N3E�]����z̪�0e�%Ѽ��~��GuˍX�й:���a��T��;��(� �'S��5���3S�ިX���T~��݇T�g{�}[�*ƴ�6*�����}�+/��oI[��K���߼&`�k��(���y�4�������Ŏͭ�5XlxVHYEB     400     1807ǧdɲ�զW��^PA���2/�k��T'*��9o�àn$a�CZB#T�����-,��ԬU��N��
���(kD�z��s��'�/#�h�)2�]�(���p�L�U��p�>����k;!�Br��ggR��PD޾�����N��7I\��J��ϝ��y�ud�PrP�{K&��sQ�_��ά�.cP'ک}b����=�+Zښ�~��Lv�s1���f�>��1L��{v>?*-o6�ר%1�1e]�W��D��i�]��������%9��JR�%ʈ*��?�K�1Mq�Sٛ$Dy�j<A�(vn%A�ʥ���W�+ok�x�G̑��?���5����N|�O��-roe��Y������}��[ ���H�d1��!��C=�w
�XlxVHYEB     400      f0)�)(yp�D�b!뱻���tV�~���O���]ئ	lܚ���t-f��L3�(��7?��s�˪������,�qhh7!���9�DC���jTo�2���D��x��'*����D�v�E,���aȰ�0A!�OT�t�Q5��u�Ax�������Š�hJ0j�6@$�ױ0U��)}�N�-s05��f"w��2���yO�b����dc�O:-&�/MѭqCx�^X7�~�P >	�a�4MAXlxVHYEB     400     150;��ee+PG��TE�$����R�R��Q�S��`�
����0��!�����
�9�G��a�,] �����C���4�FM��sT��bo�ݧ�va���a�ʪr�An2�W�G���;���|B���NOE�qeXWZ�%Nz��UD�(	���j���
�6�d�g_��E�L:��O�Қ[KmVd�gƴ,<��E>P�x�
*=ᦜ�C(ɴ��l~ifex�A����e�3=Kq�;χ,Ѻ}yT��R�
Z(���,[T	&]뺫�t�
4���C:� �֋�ϳ4XG�j�70��zn$�ʼn֡�K�Q�Y�� ��8����XlxVHYEB      b5      700VJmV��K�fCeK<"�m���HG~.�4��h��&Nf+�e�g��2�70ښ�t����v-q��Іk-� Љt=��`�W��xF�e�dBi�4^��V�ѳ�օ1��K