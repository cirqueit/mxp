��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����2r����[�̜/��ć���t�9"2?N��qr\�5U����b�yD^O|�)���H���t1H��@({w�?�:G��T�>�c�nǪ��	���N�DZL���
_u���,�5�u�P����ր#�A�� �*>Nkg-���]щ;g�xJ�"6�Cx�Q�l��;��JG87N��^��ֳ�ta���5�s����������6�=���/��=(u@ػa8��N�Qp�F@c�"V^>\���ʫymE!�	���Q���п��\�Ҋ�h�Hդ���F��<�ci4����ru˞u�o����/��f��-s�x=��S�?7༗�-9*�A0�?�\�C�ꎒ��+�kVj�D���\^M�)6�8������PG��惃z��6��w��cԁơ��ȅ���=\��	�h�58�P~��E��-疄0Y�.���y���d>��t��4�8������f�B�`��ܻ}��|k1�ː�#�5F���Y�����'�!x�DK�2��$>Xcb��ӗQ����L�s� ����u0���b��-�e�pJp��'�_o�?���wJ�B�}���v0k�7��ěC���)�]���0�#$���@8��>��ҍ���'���U����&c)��t��2O�E��"���;�<�KƯD=�ƶ��X�I���BEm˙�Y����\��kK�8�'a(%�aĮK������2|(����qG��z��a�9?A�`�8�SMUsX7@���<�?Ivk�g� ��dM��K(7%����,�Λ]&���fB��Y��m#Q�*�_3�?�!��>'��ao���������<`b�#%���P応Q��h)��~��DFoQ	�q��eoCY7��2g̘O�(�J�}+�R��f���3�2�t�d5��=w�.�)C��҆���83�h�c�5>����%``�[��@y1;5� +bHճ<l��K����Ӳ�'v�=_(:��#7������'U�4{a��gt1ƚ?V ��n]�7�s
�.�X�߅�5_��r����#n�p����]uH�w���t:���/�^�� �sZt?����իl�*�]��yχfc����t�������EⓁ�@���6"�]�
�8v5�J�])�~�dl�T	U�LѲ��>d�R��"�\S�v.mo~o�~���bݔNLb	0��Sl&�^��}[�U5�ڶj���\i���� b�����,4(��]���@��/:t�L�z��l�pevJ3_!t���j�]�ٍ�B��͡Zk�o��W�^�a��{�ڷ��� ��.�VLp�m�(t`���/��O���C�����ڪ�2�(ʝ��QZ�f��DBrQ@u��-μiqbW��S��t��Y<�֔�qJ+a_͞	���e�r$�Vи���R�Ƣ��!���w�/�@�ܲ_$���[)>����g�$H�j���h�
������R����;��p�>�����B��"�ʅ(�]��l#qM�	�[N ����d�*��k)<��9R����@*0+ĸg/q��Y9��p?8Ӥ��ȳ������O8qĻ@M�R ����p�-���ͩ�$U�z�n�װJ/�.�Y�J�}�\^x�y*9��3���-i��L�wi�Bc���*����'�m��Iz�h5���Z}�������O
�%t�K�B����23��#�įس���^����C	ف/I9'���g�(�׀4����=<�?j�:�"av�\Q6*�/�`ô0͙��tpԢ
�Ps ���\�M�����H�a�	w!����c�_Kn|e�h�Ki�v!�{�Kck}���r�כ;�4���P5$�'�����������y�c�t�ux���H:qY97��NV�O@~+�����Qia�����ݮ��#s=O_�z�A/:(˭@#�2�5\��:"��A��1�����1�a'2趫���Yu����V�,�x��������{�����n�����Ņʆ�E�����5��^T�T*��$��t�d��IY�����%� �s�G�A��8.���l&p@�Fb9����G��R�t�̡dz	�����Dm愸�&�7z�L] 3Z�(jU�����p�(c�'l����&��HXBf�G��b�1l�7�g��~7T��{u)��Ww�/q\����΂S�I��!��1�ݫ;��Cڶ���Ì�u�?/�F�@ީ*?7���gY�h���(���D�s�P|�!�Z!�k�w�Zg*�Ӵ��S�.�Aefڈ���Zi�����)Bg�m�(���J�Ǧ548��a���b�&_R�-bz��܋B��A����;d�|ߢ9w�1WP�~��ih�`�Z�G�8��C�"�rf-���=�3�S\�i�S20ӷ5���t�8.A��R��t��N%�0p��na}��8(Ǐy�:��Кd,����"�Rَt~RT���  ,C�~�d�"i�~�� ��`	��Lߞ��r��� ���=�����!��}W.+Z�vv�:�X[�/7e�Ey��_�T�o��v �^]iy�i7g��˄�?Os�{/�ۑ;,c5ĩ�[�hYS����~�[�����uxjh�1�F���b�g��]��zz����1�sS>��}�Gn���M)	�8������X�]@?�ND�u��S�!y�|�Uބ��2�Ki�%8J���iV���-���.�xWv��\����4@��A]���o���e�a�����g�/g0����<V\�6�Y��fy�ͣ��>��kƁς�>� k"%���Ƀ�DU-l���J1�l�Es�2�̣���W�gjd�uq�@��!Lw'Z�K�6+/4b���ú�T��1X��f�����_�@ү��w���Ar[��Ů}B�}�%��ϥSB���*�J�7�YyF��Gv���7k�9�r{��7���A����e���} �	n�<=�����r 
̙~w䀁��3�y��H[bV:�G`�{�<�1�K6L}�������8�&����@j��!�4�|4����n�hiyol!E�`]�Zd�x����.�n"#a����}�D+��g��*h�w�3Y�WxV��?`5���M��&GF֌ditz�\85^[�[B6Z՗'{�����0������a~|!wl����e`|
 �}� N�����͇��*W%���d)��0_�\�v�R^�j���b��T�z����}a��	�e�_���RD��� ��JӋd�b�
���m݀D�]��SLx�7r]��i���k�ʣ�����h �ΒFt�it��LY�G�E7l��O
����Mq��|��E���"��΢����y��Cn��NK� �������Gj%�yC�1�q���%����}0��®y������A�v&���l.���h�2�M��Yh�{	���$!�~����~R�݃R�Ws�(��>OI_d/�� ��v.4/>8�6�~��?�*,�6G8�cj^�b��fM^�o�������1(��ۨb۳�O· r6,V�u`���Rƙ]N��b�%x�����FԊ_e9C'���,\�W/H�w�+�h�zŧ,[y��/@C_ђyV��0����I�s�x��8X�Ir��8���!Ŕ����Qؖ��'��h42#�:��H��O�b~�L5,�e���)W�ڻ��`�ۑ3m�:���>\����b6�t�	�H8z��ϡ�Sv�FS �b�������1�y�!�����s��Yc^��d�U���@㧘��F]#��a3i]��A�y����k��u���lۚ��y��SMjny�'� �\�73�%J�5�O�F��Z�{/F��.���:�&����mt� [wT��!�+rQ�h}��3p��/����}�Tzx�0+҅r����ټ�ڃ'z^�Ծw ��/�>UcIvS"��ȡVo8m,��}�Q�~�@2�4Xıl�1L��wk�jN
kZ���mݸK`ƛ+BR ���J�����u*�,&��L�Jr�'J��_s�H���AͩjB�m�C>�aT�d��g������/�c�Ꞔ�~��sѳ������>�N:0Z%�����?~3��2����tΨ�7U^TӐx����xj���בW�,�"t~k~fnv{,]L�p���f�
�n4)±7iO�Am.=��j��u����*Z�e���2W�Q�Z��!�#Ȇ�R���6��e����s/+�I9�Wʴ�F��3����J0��S�ǀ��X��[z;�u�[���9��z�A�<��s2�ٍx�d�>*�&_�7# ��͊7R��wNZ���b�F�����bيX͏H��~X�RM�a���1��v�vո�m�e���ҨA~삝��){��Ws)C�4�ӹr!�c+�@a%a����ER�g�V��y�[mϖ�Ou�W�NHM̝��m2j�}?d��qݦ��~]�f������������'������r��c_����Sh�ْ�G���C�7������j5`#zk;�6LC�S��W7z��ɪt�Xm5��g��;�mL][��s�*o�u�co
Z��⡽;������� ��4��-T�Q=���?<Fߑo�����oj�C�]�������tcr���7\w� )��g�~(�� �\��z�X�L�����]�0c��6�B� PG�E���h$�1�a_�� q���>?S�����u<V����֡AQ�}S��E��v��2��G�~/�g���h*t�<�������u��e�꣠�'V�Yd��Nm�iӘ���H@a�?*��#I�uj�RxzL��a����v@��o�MͰ,;Z���=�v��
ğ��d�4���i�BG+�jl,^y�T�և��D�壙[�/�5±a����m��~��_�?zv\Đ��)�_V �&��Ӭ�x̘��<Fj�J@e@�uJGs����Q���l�e���>�:KE�K�n�3F�m'���*�a~ƿq)���/[�Oဃ��m8g�f"��n}�=������7j(42aHrTB����!���A�n'��F�<§/�`��sp�NвV���b�6�SFp���F�4�(�*q��Za) =Է���G�pW2X��T'�����e6��y�˸�81������u�ç��ü��k(-s�AB�����<C��M��Op���D�ek�ڽ�Л�����W婬/?r��'X�-#JH�W�,��g�Xj�4�Z��i�Ɔ����?/���e��g2i����P��Q�&A˻��{.��KT�
xd^�V^�%+FZ���`;�LW�ЯԠ�z��k� �~P���5B��ZT�q����@����sUeH�<+�6���1g��F�L0��\}}G�
|s����5���g��Y��o��6xt r��W�T���P�x!+c-᫡��:4�JS��������C�=����[@��"����.�?����.^��:\�n=���ٶ�wN��̎[����?����4ڞ����Գ�
�K�f�K0��ap��׼~�H���1�nύ4|e�����PR{V)q�'�Z�7�=ñ�pMUD�:�$�ɱ�lu���N��pm{$��5>J�Gf_���^�%�AH�x�pv��{��2��2�j�)�ob%#(_�M��ԡ���i}����\^ST��T�u���qZ
ų�,㎨I���7rL�]ϱ�l��M�h��nzN��������J�i*�mk�W�8�zmI��q%g����T⊼<۳���@��ͅ,0�c>~���s�A��`���o���X��Q��p��#;���9Z�Nq]:�����Cc��z�C�O���l_d��9[�36���Q��a������q1��G9�m�v�	U?�6�&)�E	!-UL�L��`���e�bR��7{9ܢp�F|�~���ԭ��\�1���
]W�jch-o���ĝ�K<�j�˶���q��:g�-ő4&�I��\�Ay���o4	���y
���'���T��36r���D�<'�>O��p]�uXY�b�T��L�<�lW<�z^=��z�쒪3�b���z/�ܶh3������e��OB� rj�����f�0���ݑ���[�˃�$cݜ�����I9����`��m�
5=��SC��	,�cn��G�>;݉|���/^�!�)�l��M�\��O�x����=-z���gڣ���D�5�m5S5l�i�/�u�M�{�W^.�TQ_�E{�p��i+����:!���!�ٶ#�Pr#�L���eު%��BKx��=���ނ��
 �,��D��3%|�֓� �

`y,�&A�U
Zso�)Ru�n�9Z���s��[�Z�»�U�;�mU�fՆ��K40Ȱz�O4�� /k�i0���g�UrOPTq1��/ �ɣԝ����yl �&���g�<��������ǥ"1��\w��9r=8#3�e�ⶎ��!GbH���@W��t���\�}�@o��%� �;x��r�p�ҕ�\�~S�����ѝ�I��x�5�9����p�O���~�S%����hD��&e�`/kaY1��FL��Uİ�R�c.L�����<$��j]��c�\�+K�"�� A�h��CF��USy��T�ö\�#ng��P3���k�u�����456"���dKBW��ԋ�\,v$!$:,�8��Z������u��Vy��I��Rh�^E�y;#]<n*'O�/\r�]�k.P��G֟��pm�Dɣzh
�D�6�Y��U��NG�1�ͦ���K�k�YbNDL�j���:Q
*�
9�%р8�^s��+# 7T��m�0�b�'��ϗİ�>p�`�zՐ�n��#s@Ѫ�`��#�m���Z��h��p��V,2�S/�Wf�[�:E���qM
~w�ʏ���(W��FC��џ��br���8�P�����vrT3��.E�H�G��fOjj�p*��� �ֽhF �pw��N7i=�����d�z������� >ܣ�N@�k��l��;�x���8�\Ȑ�[���B��qY#}����%@�����X�W�bT�^��R�rs=�F��_L�p��ݴ��׽̤���b*p��"�T=Q���ɬ$�*q��7���i><MQ��~#�fy�5@y�oV(�y��M��7H��v3�BZ%�[×kT-C����:��в�~g�A�#jW-����Ks+&�r��|{-�J�m��� �z;F6v�0���2Oak�*O^`�^(>�t������o.�`���Vk˟�l}����?@!�w)��|��G~���8����H+���^��bӯ*;-&(��8�!�e9���x��{n�&�W LԜ�x|������I�f���w��~�m��w�M1��E�9�u6�`�v�SK�9��4��$~^sPX�qJ���8v�ĩGc� n��X��iUv�S�Ã�a�?���jv"D�?s�@>��v.��"���KI�`=֐�
,$"���2@�5cW���N�'��(UkbH��W�	j��s����v=��R�T���=G��:^A�a8��F�R���'�2������c ��W��*�$7/��Cv��<����7	��qz���.����f跕IuѺ�3v�]k�A�?�"�{��m|(��e"$<��W�1_�������0��R�%�̍��R\��󴹜<Z��Q��<�#�luT釦ӘS]��1щ�΀9f)μX����$�0�>8��3���f�0�R�%�_>��*��ҩ���_�(��<��u)d�z�0�;W�H @d�Jb=X�S\��6ڮ/��S1/�����ڱ���k��8�}5���ޖ/��A/�~YZ�I�����ksG��I]�K���fY=�ٟ#�O(����.��%t�a-�0�/xx�u��>�ϠH�<{��'v�p�>�-��	tb�N�w	p-�!�4=������>�d��;HюR�y���e�*���.;���M���4�Ca�ѓ0O���#�? �(�70��
�	�������"�o�8���R�"�����]]p��K���l+��bM+��Ɖ�������i/>#�I��<�$5U�7Sjrm�r-1!�����M�6���h��u�㤗�"N>Ym+�<�R��QN���f�W [��-����X�δ��F�aĉ���v/YX��1qR�2�qi�`��W�����3�����_9�#�&#BG�]����C&ER]�L��B�1�l�.1����D�_�_t�G ꙍ6	��n��f(�A�¶�Y	WA�N4-�f��kg�Y�Ϻ��nT}R~9o�� ľ>�D���',G`����)��!��/�.<��js��u���!h'���n��^�1d��3�R�����yb�m*�0���5i�\����C�#H��M�.�
���I	��:zl�c.E(*4i:׎M���P��ʕ�.�+7BF����5w�bL���L\u*\n��8b��+�U9R�}�Sq�)f��V�כ@���-�����&`�P_�<?���<�1��r�4��R�T��0��琽�P�.ȑ -[&J������ c�r�i����N o��Ű��I���w��z�G8T/n����6V��tv�K�e��"w����$c�,T�ԼP:P�iP��q�(�כ�r
�Z��	�@�;��V���e���,Q�-���::�W}2VW��w6���4k���M�7'���k9Z�E�/qz�B�@ǝ�ۣ'N
�be�V��I�t�����fd�$��h~ �`�#0i\�Tg����?��������q�_�Au�捉쫉="��Y;�ev wX �q&
%YE�w� M�%D%輺��&H��x3��|)�zx&�:/|Z�I�d���ز94#{*��	v.{�U"u��E�ь��n,�2f:���k��]�����h3
ҥ43��A�������d'�鿜���1/��矸�3�ULwn��v߂G%�N��l�� ��cnsr��#��L��x��(���n�O���ӛ ����������*��0���ױ)�3�<��C����,ʥ$�y���ʣNՉ��s���u1�� &yC���>�vn�� U�~�����
�32��� m+,�
��:הN��biw=!DR�� ������;�&
Q�_1V�b�h�L���'�
'*��)�dXC��F��	�> R�/�^x���1�f[)��~yZʗ)� e3x�	�P�XÁ����/[��b���	�=�C:��� ��5�,��mܘE�e��݃X���P�OV�����+Р\A(�n׋n��L�+~���wUHK��g-�I~3��*R�c�D?ND*e"G]!!1%�K�qd�-�guX�P�Y�`�~�?�}Љ���2��t��'Nt��b�]}�]����I���/w���h���t�	q��r���<z�_���?*5W�.J�v��S�ô�^|^�+t ���=1����Cl#�Dm5����w��=d\q��+���?����̓+�Q��>�W���mud�8ɏ�7q�6��W,��|���_�U6�q��,b�	-�{Q�J�D}��C]��,o�-�7ێ�x�������X�� r9��8��_6�$�c �M�	F˧=Y�!P��T�NtǮM��.�׷z�=px�2��=6EN�����>	8s��ڄxŊ��X�XM,SbH�#[-~�̾"��F�Gu+�J:W��b�X��i�����-�Xá�	m!��l:��s�H�m���HD�L��	v٫+>�]Ϣ
�X�9�K/�=OH�� *���oh%>��A~���~�	��Ƃ����#�d!��^\H?Jd6���r x&�c��p�&gv�k�D!gH�g�v���AkI�C��W�^Cԧ���Rf*?Eb�+���[�,n���#����"��?3�4�6tC���c6G���(���0F��q�D���V�>��q����qtY�$������8��h.T�����Xt-�0�9��0�.p�m�PBͻ�^E!���3z��;=B#
bhG+�Js��h;(�o�Hs��0Z��'�dH��j�۱����8��K&���q�"�yqp�� l6���|��HN�3i�U �u��B%V�F^�LN_��LM����������9��c�V�y�4E��n���Ƞyk߭�ԮJp���ek�svY_,��I�v��n���Qm��i�U��\��<�No�����0kZ{c؋�W���}�,Ѹi�.�Tx��������[��V���~6F��.VT��^��S_�^Ib��W�7�,�k��1�y�p��@�L��9T�.��B�)N�)�H��-&Q�>�E�%B���H�*2��J��r��[