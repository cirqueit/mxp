`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69072)
`protect data_block
8jRazD6Sf07+i7hpdshP2xEH7mqUyN6ABH6uECFEKrBdfg3bhyn4cpFTP0qOqg9QfJkngIcypbEF
183geAq5rHAvJ4uxgy+U6ZmhtuHwzMDWVslJajw/PThsJrgpHHGWfRO16MJz8rCzjf8hlVW5qeVh
MSlsrYc/IVhjAHEYVnjYe6cXmx1dRZ77XolVnazo7HQinOZXZu7Qh3rae8dcqsOBjN/iGh1uCwYm
s9IPt23AXAvSch76uPxhvWoUuheadpos++mCZmZJ5mHST3xFWRGFQI9/EUYScb5rVE+hXwbdYC8C
A0ixm7rt/eXMhRuaFNebHDHYhAh+8CwdUYD69qO6W4o7dUQZ2dczywR9lfeygbLUFa3CzcM8+JsE
Q2cZcI/yqasnNXFHrEBx65zCH235eiPRIeHyYwIM7DNjYeQsmNK5aFz/ubpSMKEKNE/+Dcl/gpa9
IBU6OaYg1wsyAI+FOBM1jBeHK5lkaUGf2Uu3BjCYoPyQ33DLTG4lvYXdZqfFtCe8F3J8NJSKb1L9
pO/QlhovPIztI26Nif5rbtdc1QE4xMlnvURVQjF4SZ+Crru9p4QNe+fd2xLdy6tbRXvGxFttAdsA
ZG9kqkSMlbE/ZdG7/R1qZU84ydTwTLmTJ7TP2aGVx71YHMtQYLrfudMv2begoJVUaFIkZ8qxajK2
bpaYt68hJjnMZfpzwRAf4aB3O4ZjHCgcjOarXwtDITLFXcz/TY9M4CMGd4tVzth+ro6KaRFJwbMH
UoRuZCkI50/upotv0tDoZCsY4Cm3lNvp1LBDArc6wO2+KEx5RIHb17lMaydTpewZtymGQKQFfB/v
iQld57XnLf+sT0WgqscnemFkgc1rLwqnNvB304V+apLJm1iYHHGSQdM22nLPP4BfDNhnmzSrvrJz
OH91SGB88pHMvI+4sYiX/UCGOIbIBujAph4iZTKCPO8Vf6Rh0y9Vspx8wCJ9h/9eUCt0a0srt8wk
YUMg4TjFucTEIPxm/RA8OM4lJ++FS6u6+SkLd8JpsoWz9Glxl+CsmmAwmC2rrEPkXpWlaDyyKqZu
tifza4nYi2ChcuZ6u3izH7CSNI/otv/+qSI65U+L9UkJBEXTxBgFToe0vCTvlDqg4VNpwRk1Smpg
s8bS2DO8Vf0gBVyy8kO8NEassOpwnm31+7rK1F5N1/yXfLIIuW9BzpKmdM7OV9O3e5gmvpD5wfPc
qntMGMSVfh4H94D5a6Pxg4PabqGPFy9TiWJi8GzBtRuJeRmKMBToSh/k6hWKmnRHZSuC8dU+ARfH
0NvTMxpempwqB7zPsd7ciLAjvhOgD1JdbVz48xFDFJvre/OcEBDY42YMVreEXtGWAHsOPpASAd3s
qsXzR9qQb9Dk2T3q4ZXEehX/mefcQgTxc5WmHAjA8HyPU2SLBdo5DQM4YTBiZZdCp9j9ocBnO0Sz
8hwQXcP/scJMsQUnKk+LWa+BSqPyOQTM38EGFeESO8b5l2uoW4IENs0OIjOs/85H66sJP47tZs1w
u1MF045SQQpwLejw10eQhVGQASYa4050L4/MJtLkRIpaP8iJyl4eq5AIKn9wjaeeYD37bVCSQfdT
kbjtO7N94vAJCAtVvF4/Yljd0i1noCR6VhM3s8f0+AUPDEvTxq2SNViRhtpPZjWmLfcL8mnR/aNR
ocmFma9EUc5MW32IhqoKyQGL4rT4It+QuwFjy2lDemifsiKcxK+xGmPPYvH2GNCLJp2uFJStX9gt
IbrkNcVJXXayXbALzw5i17prckwW55NWdZ/ReZuD45vmyAHYJXTU59WGM9F7k0xIeMUq/jxa80My
OhSsJC2w4qosbMHk5Fh0NlJugtyAkXO+eImG8La2a0cfCnOmHcCWaBLXFL9WK+WwcIn0rnMWy/we
lkO1pKzLPkA9uuU4yZMcWn9jF5qr9vf421mO9SYgu464KL7Fq+OTEFD9JTCj8ocM3rs5FvvO3oBi
OANKLLCPNXgE5iKHOnlFGckfpNGyd9gDNZzr4JoyWAMQGheGcyzJTwfc5+BBf+80yi+VaZNCOsjx
WTajziMOWROdSkls8ILXdgZqi3YtyfOqgPSkxHHhPuGlul7eiWU/h1fvH7s9JjdNrvVezGtJKdGb
/sk6f9fjXbaJ6jNkUPa7RM3TfQqcRoCLhFrjZNSeB8NBBWe51JPiBaXq4rfsiHpfi5GRGysUFl2+
ICYOhBbMokpCd4tXjbmcQFK9nFk9HFf9Ch4JDTCF1VuyYQTaed0DMXXxHRdzQB1cIe0gGr9nFhX1
zncD7TMuhihBwtVVXfDzr5swdLqnLU4yX0hnMTmtBFr29lX/VeQFd1Oz4yTEFGQPmQjp4drQvemn
VTRh5U9+5FGtFYcCtZmGCazllg8vTG3P+Viy8rqevvxr5VzRm6P0AnLAWRRmUJZOQQtdnMNMd+vT
LQ+iqDp2ZJBRd8ivD6Z8UMy179js7CPa2x7ZRo/A0zHiseR40P2jBqrCwt2Sw8i8rf03LmYCPtlr
jyN2u7z7OSKtH1mF46I1EhpNaopIrjNaze53NyMdmD27IFOsl4Zal+brYwg2rSbcetzko5ilDvAu
uS3fYkvSnHxx95frRM3ZnDWXWrmC/+RDlLmrN7KYFK09TrL994ZJrKQTz+5hmGF6CLJxrjBDpYvE
NrjBOT/XhlUQbz5Sxri8DGSITKJQcCwWJD19sHd4xE5miI1zz7RLxLSh0fBNMkIzui+tsKmUrfaq
tGk2CXe0r5+OEpJlXJBnA/YnT6As3paQ/WX+ywGKbpaU/uTRguL386NjP95jO1ASaAXPBtz0L5PF
j0TqWzAOick88OAuMu46O1nPilx4/2Z0wDLk4k9PQcYMOvb9YwnP1u4alwGsCLRbjduo1MBMfzHJ
C801wYbJtbZnrfQh3ra/4nffbyLXfjA1Je2m17wWztGdue4D1Hs9GvJsecUrpFeyFa6ejwqf0HJA
uJbq/KYJtUN92YKHG4U2h3g11QYXmpxmu5B8ackF85IVxNUBq+vLrrRF+Pyq8fmY4b38buXAPZ3b
6AVt6IRyZySi+EpKPfA0oM6K8Up61wfZfPyG2m+er68wBDxs8lkSBIdQcYuKfk2SswQlkYhxAXkz
SOPl8I4Y4cq+ol04IInW5KB7WC39Po7r0qGNNpNIC+qUjyljWSG+CSEVlq6by+5l60uyUTkyu1w8
a/wIgRG1/UZS2mE3acNzUGVPMfc5KLdQN361vxe4F2Zpn3yvE7Qqp9XB2MoJQSqmGYG1avYlsnYl
vu/JQRJonBRVQAOTc5U5wseim/LdW3I3bgePH79tNahOlcsp6Y/SDnREYorKnU5IEN/ZNjMGhATB
UwtXL4uhVsvUDAKR8KVG/xOwd36vz6T4WCZvzHnlyTmtZLHC49QvGjbw3NKybfzH1MK0nUPP8eoV
cUNbNHiEgygvKdIYM/9iZQqpPD9VhXMyMnZ81fH5b5XS10qXotkHRZHWv7AFfcIjKzlOzW1B7FIU
XQmAFIR+jU6kNn6jjNeB3Nw76LwTuP6sdQnOlndRo8cTr8D6lDBUGhZMJBC2MfVtmaDrjLACI1bJ
B24J91cj8FGthfu1EaxqGoxVpwXgm4U4e771QWbAJkyUJ95uxtLlcepjyQ1OmxImLmsJ6/142wJs
HPQ0IYVc5PtZRrVOqIfxC1nLEkhgYih9MThvpsGVHozzDVJgJsRZghJoFevDm35z5wyqQwJIR6eJ
3C7VgHX/dyThQ4FRTyLA6tX79AyFjN1KHsSRD4gk/Deu+2j0RpWaMg1gGzvV9POMk7sJYM1zmUrU
On9Vbhn4H0hb0QCGAL1GF3ujxiDKMh38/IFO57KYC5ge2ih+SDXGTA+TjxGVmqHT/lzH5sQzR6Ov
KsRNeKoq+IyakjkxTpYR/H+YUTJW/eTTmW3wvZU7Pt3FeY3MuW4BaFjxc2EhXWd7WmfoO4aIaeo8
nQ7/8HjiLMNVaRu3UirCP0ct4/dESplMv7pRTXSn7zOIo3cex96QwmxfLl2RBlkwA6LBvxP/lkbg
x4B+V/mFCAcQaFVHUwhT/mk3mDhiLlhqHFOvutH91EONuyzaIDwZcKLuHATStZ54na1E0fQ8EFyw
DZx4mjNVlCXZwl+QP/v9uWV3e7vFBmkPAJF3aQbldmXea0RRI5L0add8nq6BPW0YhStvKOEIOKzb
vpToGLE/hqhqb7sVsPpl2BO79zI9xgavPOx7bTp0fTKg4sy2llKSmKSJg/Pbxna7JBac+KMdzFGp
FZ2SakmjRxX4clB1TlpfkLurU1rzoOIPNheygqh2spQWlGjqHlY60OlMi9gaDax4VCQTO3u09B9b
U4A9B6lvoicQVzfiarw1iuFcbiWEok+vYpBrjVpqZ18w3xNw0Bl8VV+5Tk8duskUps2fxXl8/IsM
eWaSB2XeMxAKq2gx8ysbcDPP7dn57s+M7avZVVrUkINr91vOzozU3/9tjCA7pobbkTQ6G3nW1s6R
oseMJqvsQu6VeXcSc39frUfM6XyMeSrbTBW2+Gg8ggLHrNS9us2ne5l/T3CS2XxlgWmxctTvD+ZK
wGPtsb0oxgculKZJMNQc7ArSUXnbxgker6NKkRhpWh8vLz0cUqcV8AxROb4OFVLHiLVg7iBl9HYs
Vcv90uQV5TfT2SgeghbFUuL2clJ8J1aUPygC/TRoPrZvIyQlNF4TVLdnKTeA4/l696ILfFGtN/B2
vJDgRrnZiN+BY4mnmIDRMLGLqPQgZAsWWjTJG/gnZJaBDg53RXlQ6AjMVMH90BYgDK/qEczEyPE6
oii9c7B+GaMhmQvhFdxNZgbHFrLAe/8VtF7PJWfNO5Q+h2gePw3LyrKViwr1lCmr8Q3x7Ks4ROYP
p1RMUTz3UXMCy0t0IxIiyJEH2oX4kwjtzNePNK8IJ2i1YeJs93Slgg8Yd740QlcM7A5UqTN8yxU+
zR0HNJyJX7OCy4o2bThtSy8g+Q5nAu+xJzp99ufJSFRFXiBzCMxgdG1Mxe2YVlYJ+harMF4VI25v
WSFIBGXLiHxjiXoX9N6OIynuHYQfhZwgTKOK4jEotr/p9Ud4l7QYkL3LqYpv8fxNP29iYUmYPT5p
zOPx/Cu4noUg0g96cui7FRnoJTxlYEdq91qYVSr2asy/4YUiaVsyjhRo/E1pNxvs+C6kDnkDS3J5
PFnipFcaESFJBT2amFGswBDxBAWm6rTsDTS4xIGEP5m/xJL8bjLfCRlsQtGuPKmtidb0lRlch6kL
1uahWOb63lT6/0JVP8oQNEeMG/u9ce5/NBh7/7ivZM5ppoLw7BwkGk6BThjNlzCGT+SR6fkDyHkZ
q+/S3WfPyxQdNtaZqN0BjxCjD3+Mn35nb0C/h8WPJKohE6dP2ONZyfH7s054ts21Pml6eOpHTvbd
SP7Aaf61Wo7yT6gEu3aV4wlbE5kIyVoJxd8jdLRPpxwlrkp14m8vPDnUIUjr5/CXO7PkFvlMFwrK
YhFiLqP567hRTb0k000Ha5Uq3VeiYMye1E4Z7Ns8RyExVO30YWdIFeWnwenSXrY7PKjjzHaVoVCH
BF7djj7zJ+5d//7HzotPkEYrR6m9xeXd4CSgxlhsl8TLQAI7vVRWrxLSepbi/rDEL0ZAtjfaB9SO
dxOX87maiZTnuvUzXFdVKrEgjpJUd0A8DzH0CtHCYSxDb/63oOWpMQdV2TlmAGKeGt+M09VvTEgL
5pwO+6vQAkHWK6sqXDfm0c1WXvJRzVoek+wadWBU4pqxTw2YXk7Qyt6pvjBpAV0U1PBBnoXSvhI8
iSs88xsBT6K7PCUm2RJAR+DizfiPMRJtS8/1Iw7NHozxvO4j2MJnfP7Cuxg61j73A0BsxOHTCXJd
HQGQP/rdHFzWoTuAzLoUFGwfirDC1lPZVJieGIYFX8WybhQzYHmH+W1KHQY/QBbrV+tNJWsLolAz
NusDuW31P4U+X5L7uCJN9hgOsEQPIs5pxMa/SCbMdKKWsk6VRszTdKw4K/NVW16KBK+ot+KE+sho
S/L6foCwABimZ82zUdT2bWjLf9ciz5lU28NiEy3684s5spotBFdxTuxkadCnN7OGhnYSAowNBpWc
hDvmSg/LBNOh3tMx2lL6ZTUWBlv9psz+ZjGeXV3fZEvwrIxTO8JCTigocEBUFJCmHo8n9UUHZZo1
ueNx64P/FvOk4yd1iulbGkrnixMRciDcqKonXQ5fXX9yPsvLXQ6RsFc4YAQW+v9obHqPTJNHER+V
JreM6VEXAjL8TnM4eCmuZZ7PVNzYQMGOgnCY9dFoIwrfC0AeGu4q3nm3qK8RD7lDUQOVjc4AGdth
/KEJmh7SdqGq/ud4Z1JtJnlxXYNwa0T8WpbM4+U9nViKCeoVZYK+EZujQUdJHzoaTnluvtwqmD7i
Qq+5e7DzaQiR8WuDuXfJftDT3hiqgy6aA/5989MhMwyAYdxV+ug0eVpZBQnUxdWktYE5FDqnhh7x
s1jmYrOBbzDOoSKGK9D8OAROXAJcwOMvSRdGo0+ZxqIG+hZ30tJstzxBtQYNFkOByDG5J0Evasp3
KkcR3gS0lftT1UMXj+/3CVvnlwZQsHFSj2ko1bzGa+QZuY8juFlEAK+EBTnSkA20GFpZ5leNLtbJ
33zK+nRuEhZH7VtKBh2mHtdUAPRunbJoQm4QVSQe7m/qbxyw19UChiq6aeVK3Gwc8+BP2G8Uvxzk
GEta2i4gxzRKV/eRLLexiC6OoMc9uebfCnib6/XylOoKjz48F7sSEcDXkmqChf+MMsinI5MkWrmQ
5uxPAQn54evg0u5zPdGXjH/f7VnLIKCz0l05bL34O12hS0W/u5EKstuGR+WlzoCaYQFF5tIkKZYa
Pw3wM+QP2dkgCSqGNYuJ6+7PpPFhobvAR3BjTGqJ4NQIOdYTjNDjFs8UcbZigEPV+D/HuR1/JJtj
7cZLpveorNM+Cr2fIdfOHk2Zt7HVRYLI1hFHZ2zHLZn4x4+MP8M3gJXd9k8apRkSjCO6TxrPEC8M
QIHW/MoCsENRgEge+F0ByhDjt7Suk9GeFD6tB9eFi5+VPm+wfp9IudhiXUA/cwDRVCoW9EfHAqLp
rHm+NGcdijWyPW0+CBJS2ypEY/Ew8O9+OMjXKVInMy670c12N3yFGopjZ4Lfm5E3/y5hm9OlnB42
4zrMOY5ygDgPQu5iO+4AvSStPnt3StTORilSng1xMm1DqUeB+n/wjgT4ilpXwjbPZvtLMOzYckwd
3FIEBRoeZYEka33AtwpFaR+fsb0rSSn+ze5BrsBDj7LtvdICt+aAUxxs50iQ5ecGLdfWSiQWq0mX
MmVMfZEqozjf3ik3SvnrBGZdF1EOo4lfcVeRSYEscpopVnTQM9Ox1V3iao/VGkmD0TzS7Cwva2c2
NHJXYpKylzLokFy+edHO9D38K0wB8i0A+GLIZzpZyNywamho3BOyGZCrF/J7cKrX3Kl470jzYjX6
XNKwXQp0bmbMUwCh4KBAIFkuMcWU8ReFrbkLn+jGCvckBp/4itq57ZcQ5m9p8tYfGtNPfv6OLrbm
jqupaECtErp9ZVmHt4WzHEhsRSLg0N3owKTf/qOPMqr68/eEsrZo2/DOnCK9jBZTAPRgoKoAnRgi
mhU/FlAw1iaxnVAlzUBJU0Vi5q2fCGjJmyVRsGpTJp7QcJqU3diOermFmy9vZKRM8NZVd2oDk2+C
i5RGvhh5CEbk2BCBWHJe3FoMyDrHBVeKyszF24XBtjC+QdLzaBKgsLO8Me728s6omEUDb2XiiGBM
7+/0csZ/1r5ExH5ama6qIDX8cxAAbPE0y8SatQhwWVGX964/GQQ5ovOwXrZTAIdgpC00EPY2gym5
1i9sWiMTM41gUnJ8UlPwo5J0EIu16HHZNg2NrJaPquMxTQG13zOa0Gr/WkPB5kUQNsXhHjtZyG5T
+psjxrSze+//fZv+PuiG/iHWprUKRQvfZ4acDk5m0/BPm1q99GejGnL8i6OuEmnQwCR4eSaB4CWU
BH3WjauZsP4cZ9TZnOwA6l7L6tSeFO2QRFo2hzcy3f5kfwqBgtJMnSaU/5KMRZbR0N9Tvpe6eFI/
3oG4Wr/Q1zGujBMgH5lmJrTR37r+rH3NSpEM0q2gPkzvbWcDeHD9uBTpMv5242Ocuy23uJgRDWTs
vM8TqtYmem4ugoyqOsq/tZA68vzy3/tnXvzIBv60wL1SCzqKhiCQdf/vx1WPEaWCvdQfslPCjDfZ
asSjPofwdj80DAss+EjNyYu9+XNEmW8zm5Jsa3sTLVb8dIxVfMDc2n4vKw8mk+eJuVd9Cy5jZgSS
WeFXfPEcMIq4m6kXmXcDk9YZ1BvyyIAKArXqbnq21ENvEGAD8+D6Ulo52RatR7YFRF8c7ihdvQQf
mnJ0Qy4lYNgRliv83ApQsqXqiIXGnSKE1rIIBC5lOz8WzP9vvsXfL7Ff4qoimHeM00KzD9iDIR1n
ufab+CbjUv8mDIsZhNn5FrmJzVbOoUmYLOQjgf5wE+yUBRb03Us8DwJtiZTm7RULvPdH5FjskQ8Q
d1R7Wxde5/1jZgmrGt0OuD9mu80P0fq9qCdS9akAArHKjYsShGLwnqpJqDSm8uJeooN1jIq0RE/4
puvz+t/6mEVEj7GjA6d2itmPJ3IpvEZ16s40qh/VpQ6/olt/a69GDUcJ4eosR3fusrjZZVfIDWBa
heq4nEu1YpbcQKBbURWT6VL2yp4A5mdB3zVvnPd0Gal0l8L9MBziNq3r51SPw7EFpURddhRE+eAF
fZYi7zilHHQc4DL4fXTfUpuPwo0f6Xi9jOQym71RlZf4/R5wpqg2scArBFJeFPt7VGEClYiwcm86
OINKil0rXPqRfE2FBgAfE6mS0FVcw2HEH8pOZR04htAX/awAyJs7E1b01OUl90Ivz+LiUXiR+TC2
rrbgt1CC77+XBuuR9FW1+e/DBWE9jiIEwlVgAZhpLcwTzTMOP191Rn+0WOetLBVmzb8tKjvinyJb
TswpqI7Z++ZNoZJc0s3eFoqmVvCNdqoykLnKhq7b7k+SQjEpP7AcdqaT+W3TWBavQuokD3xbPYQ3
cTxCbP9szBDSjGOfoxO71yogf9Ym4C0Bsd2Ew0xcykcSMJvAF3GXZ6WfLN8v8/wB6uLL7ZGv9rJI
6T0aWSGlYPQ3wmaOWUgcb0W1kmG8L1Me2FE+Urm2vpQk1HUtgz7h6qtzRdzaSfpVkCSusYizSV77
j0BvFWiKkh7QPaHMQGXiBveRPxSvMPrPQx7wCwPzLJyNbqrfwZ0s/+j1z2R+xHtcvmCZZX5cutaw
MG3fHle5x+urltGYI8TMI/Hcnqfu7evvJdiSIissiNPL9REs+Ozf0C5cwUxDRMiMtASBoGs0oSV3
BPbOGL/qIyldE3d4Tq0xcbX98Wb0UlLGo/EatQnuh8vDdZ0Ofb+vvtBQkcM+7Mj7vVCypac1mm8J
CGg59PFaK28YwXG7XvBlg43c2urrN3d+FUSejOProtYAr8JkNHALarICJszgKqmjs2on8XigT8kc
qfoV35g7ANP8zJRAM8rTOO65bwt26uQbNrSfPTAHBoKfPO8wngFAV/MQPdeBTcgMEgoxjhK7O8wP
05TouzmfvorlaPJDXFI5L11BuZbi0G6xZidTOXkcMyI2EqMZoZjM/u0FGuVeDPqVzOJsqjXPtUFL
0PFGTf8UNoiajN4Lkq1Bu/pv8B/qLqb4Y4PCF4y83+omL4xvlvjBg6A6uyFDBeFDYDio+ypCK6Cq
2dc34YgsA0ovLRK5M7/iVa8DKoMPVrRdidjTC+uOefSw5Xu/CT6Vx/ISoMD+AxCUMjv78iIOXlFJ
cs3FS9zPC3HGnaJWirbXQE/HpvHC3c2zvSj/FBLduTrCVlLdznMdCo3E7zQR7NV5KlwcNUQHViXW
dwVpFaeBLRpq1pVXjUbyudw03hiroy78vyUAIOO5ud0pE0kIKdzMIyi1ivAAv20akM1N7ikScUXH
Q8W1pYJ55ZUUMbc80kd4/m2f1iya9h3fSogvUmKNnOZFpohWesRd/hmwhDQxH01oBiFxQJvGkMHI
M810Y+gNSbjvlhJifpqfE8fgIgJkMfD0a4gqEeBacFo02oKYnA+X++NTs0TTe5209V5j9gGqs0Oy
MPfp/ybasfaVpu8ts3B+Obwt45McqerdStbeRJyjXZtZOHFd599odr9ddGu2auxtsunJCMjuzwuO
l5PLDaHrGc5YcYowekjPIU7HhclCS8RR0Sw2pKV9XxIpBhYbkzwtnoLrZYFZ2SxplG0JCeM6W7u0
sMGNeV7KjJh5Coq5P2/2h5hHC9YKjhtCA3X6YJhuTRCHt21uWk76Z3vR6+cx+h1VLhxH0ftwPsGf
7BwDSr5tDh1JqDZtf9ZLsKrzZ7hq8RpAfM1z7awQOIQsXW4KFbnbKCBVQad0YWJW5tUWwnDYx2Bh
htlT34Ko8Hjt8lPoqFpBQFrxN758AymYOXCiZfX2YGLZ/Rq/q5I/PP/jk83n73VH4YPRgX9cZ6yt
9d7OpTEI83ZdDr60+XiFWBWI4zEQZIxul2CXgZNjm36eLlxXJ9lKHbyQPPM3DjK79dfeLTqQeZQ9
4uqWX6LLt6dPWHZsDsV7eMMp1pIakzCCm6oNdIyPDWDpSHQfDZL7eeDy6ZMBt0kLCkoBvkb8aUPi
IjSKogPE/U4Mac7SX8MK3jvGyG5VjhdrJskxZZnOoIobZfMGSzBRqqEk8uBlhIsh7VKQoU3ap9b3
CjneP4e4RthDSX2sSSe+uD4trhTUN8a3UD6fddExdRKkivNSkrz1v/DNNYhr0AReFO/5LuepgLb9
rLZi64Ep+bvxFlCLQTp0kRCn6VVDgXvW9cIu12Zlsj5toHC6aj6OjIINkW6lJKl1I2VxllG7Lqqw
yAbrJiklf/NLhq98lbuy288OppfaDkJBo2iOT3rr6TKnWZBYbGcZ6JXeyXMGw3JoeQIe84lIW97l
KW8gdzr7+OvqVnXobccTf+XUFYjfFfuFXb01F1ripGkmrPexSsbdOiMkpcc25B29FRcOpT1aYjYv
gWq8TkI7fllX+IX+DC0tG8hkuVvcaq977ykva2N+nWiDMsMgNQXqm6OGfisT3s6+U/GpCYwYPKea
4yAQexCfDL3+yhZjrNdyyHkk+a1bGT8L+2wQ2dNWaO9rKYJ27lI+PiUUfoM7nHE8x1OG5IadnXjR
W8aW14yzzK1gr1p6RDw+jq5wHVGecuOgfGinKJSsPcWzC62OBJJxzLZv87hrqcKy/yPMEEEe7PZR
HH+GGWCwlqmc8rzQxItr9sgLW/12EWrQCRiEocnjq/etXag9mdEI76N1FS3P/08NeG8915yRKXwQ
vajLDOFLCGG4ZTCIF7oOgWf5xLPAQ06H+6KwC3cYjRYvkGuutc0xXNuJppz55HbxkMhn8yqaszqp
LxsM8QNrsLSlzpEZQZdmDT0R78+Os+b99lRxVqvt1maBVBljRy6XGvSvstEiM49XJntyVIdshzpg
nCHZ0USOaeqzh/aoyF8bTwkvRZL6eF8LRM0ZAbWJZjcbILylkYtfpyAUxwF9XWuc1EX5CAegdkjU
B6VE0/oNiIBCzBBR+fEfyfCBNBkBMRiS2L/OgTOhJJ/JXND1laBI22Rhe/XjsagKuKotbZuUe4KP
R/gHnn4Xta11GqkmJlAT4o+QQZZdWpv5FJ6TqoeM2KJz1Cct/ejpMi4I9vPKk8JNzgy2D0ccAOPp
SF00zY8im3uMdq95pQ3WqBB+9cQM0dnR+q99nfZO6dUbu4zGILDxz9Lq8q4DZhgy4f+8mtvKE0FM
7kGpnUNxoe5h3TynISVpvvnqkTBwv8pY9R6zP0hccBciy0zAiriTQ3ZpA60nDc2B5WPReblE/Icb
VLTZluTrTkOnHHqwwEsk/z87g2OywY2RVprFnj/6Xb4rdaZi/OfuEwQWzdCbA7EiUO/XixhRNCvN
jktaYo8G0qDLk+S5F3+IxMjSquYLVZtoMY89CU8o3KcxNJyU9Fko5OlBKQHxdJ4pjY9Bw0ftsOcu
MvyupNwisHnlQVIFlYZRHFbomrUh2ABXDjKO0AhQXIuJtGJJ2rvekRsK9BybErqMlOvspsyaB7Cu
gxvJn/cfPCLuKBqMWJPo+Sfc+fUAySD51zfBMgXdvQVZbS58LXxtav/JPIgT7Jp09UmGXGlPy0zA
7iGbGOBV39HV0bQrWTSPB8Rhl06kkHKG1Icg6loGuFuziHnF8JIjxyAddFPkfiE0bS+zBdx19w0T
ZMPak9BKjes7s8w2CCyzrVF2QzwvW9Muft4DuwunukpOEX2tj/85TNIHv7Jf5+GSTZH4uLM0Wey5
4joBFtB/97XlFd4ZZc9NUgm9TYbSX3uCPYFTB8Zr4YhpQi4KcFJwOf/4HqdkuxoPCLW2BCa6qGeU
q4n+8dLDdYoHWE0EwHqWMhv/KdVJuLUksbJXFnSDCYvEi7MKfX2yMK6QFxOqCjh/Ky2aqUqDNI8A
HU63RvKlbtktS6qoH+k1u7zRvdtwrsuP6qFjDL8HiiysarDyfVWMYPpzIIpBk6JKD2itQbKunnHD
TbDbBE5Q5nkk9xJUVvn+6pP5FcwuG0KihErvhfuBhDvUwh49HUVO8pAme23lJp7cMkMzF5JecP7U
eK2KUkEQfPLEz8erRSgOgNIGcEnaTMR+vzl8cMbDcvvWZSHe8LkrIwAmIedimZ44KJzOlCFR1778
Q+wyQJb65Qd6Z+zrkhyeLcHgZz798QMGFNCpMYEjlUaWj+0MRxdTIodKtJvCFGfm21l/AONOVoPD
xmuidiWKFbo+egVRHUZlKXwH3tyV9HnPA8NKyP6lW32zYvNu2UNYCWyXIpNpvLwvuuY9jmTaKXjY
UexqlwFzutEg39kbyd712Ur5KCpLafTftWbbjR/TBjnAX94YHS6kqqhTbnazqJxrsCXA1Ubxh+m9
+PfXOp9/bYU2SKLdktoeB2NKNqGC1NVKTqymbqQ6r2VRqLLG6KDKzQl/vHnC1GLEXzmFtKYmlPKp
mz/fuesY2LWomR9knt9y5DwOn5KbAUcG4b+YKtVmhg+YxGln73LHdZpSsd1NunuB+Bnu2hu9dV+z
9EFNMHB4hRsOSTuI6rnKjJuByP0HwB7gGYRFThuB7C2V2t101x+LcDAtZq6cGEcdr9DzPaadWcB4
yX8Zsd5QA1Vhu25QUcZvHqE/Fjb6cT2wef2CALMs+OyXmA7U09crafcvsbFXbfQyf58P+yMpzrUF
IxypL5pEM2s4dbYsfOQu8dBxe0z7PsXraH/HuRS+j0yhXW5dIrvu7i7CYApYp3g/iuIOSr4jmtYZ
NVm/xl1EGUDQxh6e7kNIlBjn3S/Ulr1bQhXodiYzQ1MqMtxJ9MlYFNrdspcSs8sa5KQ+3eoNUmNH
C3NNBjliG3qpKle/2dtNJzSvrrlUwL/1lqY4xJxQfOkoouBJxesLe/lPvjHKf9OPbbstFE9ST/hm
dNmtPSLbmsA3t1KRLIQOgUx/GHvy9iKVIz9Qv9SwpMB/EAUAw0LgpOWYpZNbyEw9QRCUVmvZaul8
JoKfjywCd1FYFrvVdJRnRg1v1psElOVflCTD6Y0zFj8TlaP8bw2uThzpgepqaZfCTOZlfF5LOuqw
uLUrBxQaFc3czFPIAYLpGg+c6WcA70DbDp9q0hLVK7o6A3Oc5LFG2cAdagUyAC/Sw2IymWx6kae5
hQLmnZsabLaVSWbRE+gaIdzTfIKUGA2s6pJK6wLwXbCrfelWZAHmjw44borkoaoz5U3rZHJ1Q5Pe
kDUmigXcjyIKZjfvmA/HUpkTIsN4K+HQ4p1Y7LYEwZKiKLLDavmAQvNSqP6zHk8gmyF/x/tymXxq
jFS/+psuTZSSEddNvas80soQl4KEyjFSDC6oiDQl+Jq38q9dBClxnEiFZmRjHzGQkC/tjwH4lOd2
7RNrvoOt0cFbvdd0OOVtgZqMu/PaCDKwkkTMlPMHNuFv99pEYA84gmUWNSx2a3OEA+B6tTH+9Gqr
fUbgwPYHkiYj82MpccU0HTmCHdqZm2AP5HlW8mcmS3mErNIgNZclM/a/NjyEJtpcec+5lYIoWjiq
ld5HQLEXwOc/XvOO8IODclnv/ozn82HHLWgTxZwQPn1Caed2AeSTqZdb2dRmrH9XsLa36T5SeHIJ
N/mlLIxK8SduU1B8eul+3eVI9qHRXlcuK/hmptDycuHk2/IYl14V2SUm7bBooYzthvgH9q7AoeJ6
QJgJaJOi6XIojzTHkCjbJ/giHxvTI3/4UQ5mObEagpdCXYqzlRt3VGV7hA4oylbqkCBgGhm3tOcs
/rdseBIU+AO39dFOssID2OFuAylO1+iNd0SfrGfKYqtR/uoPtVWlB5tNzxfST7999pltnyzsgrJD
vwkkcliEtrrZqTHJSLVBGDhoOTL++VDZg5zMocC/K2WCoVbE/Bw/hubO2evnOWiUUNLSyj3YpaBi
aVCQfg0cucSkKsFOkKCqCUBwRBasp698SYWrQAKNDPXf9xjITxpcGzndgVdzZWvfvq9et02hC5Sv
TOF/yvYnoIuPcQvjvu9HDL87AbBes9nP800FAKXP+ner+6vE/6pzxPVY03wLDCwt49KmvZETRVkk
Oua8TQmK56loHlZ0l+u37ZQC1v4Oo63NF67ka4IYttdLy9yb8TbpgCFvEeN4gvnLwRBwDBzTPTuu
6B8O6W2JsBti0fvtnCEjbxC0Jr7///66hqe4BCc2R55U3CF0/9ZPmsOhfF49oVNmkM6IND7rNcik
UQAcI7E1Rxo4uNF3+lKX9MPszwUMX72Y9Wzh1jk2uhA3b9l3T88WDgy0tED8pcTl7wAev+sXa/ym
hhyFkA+mCqZiHeJb6UV/jFu/5m0PpcvlEqLGpjnCkBpzicmhijjaI9mSK0WNhKbIL5g5FGdapgdP
Jrt3UhipZLz0ZpyEPUN5jqX+/IOKu944kYC8pQ+Nqii3Ffam4jekm/XcvMp/vEV8gEJQcNDU9iXS
q3Epaa5nprNHXOFx1fbv4wY1R4mnuamzXMmWwLSgu7cOFprMpUCljVEpMvaFYCLg9+s7FJ9Xv/PS
2vRF+3QKA02t9IsJzmJE512AR302VWPjwopW11VY6sgHYAB/oGdchLY/zUmp7/gFau+f3QVJSikj
Vle6fxoqDmkUeNgYFJgANSnHOfTn761v5zIlcBTMvgbZixD3UhEIR/FGLdncpvKCOrmWhgJrOWoF
RxFeQyklh7eZolkzhmPNS0wbEIZVVgRd4picgdksnsmIslAMkSMruyYgmvgt1Z/g+ZSh+aA2pTnU
DjwmmlnxwrOQn3XccsxWM16NC8O4c4zYcXPEA1Kg11Nd+ZnMfVLP5vNz10pbp47KYLPU7k1tKQL6
wF597Sswr5hyc6xYhv2bzeuNMIrGqyIduXL/+8ywTo7GY0SYvF6C5gu1jamj5z36FiFxvDQdxppr
OA7YzW73xxKZVyRc0uz7LkZr0mhuPGDxEWE2teLyrtdcRiZ87ZGR0L8Qx23FdakwrC8PvfpCHXvX
Et+36Tq+5kIQPl7BNB6DsYLeXsIEuriWYeq5lkTwJv5fLsI3UfLfwAGKKy7KSItum7qrMZ9VpT29
hE4B8ui0WQVpQqh488kIzztByoMSTtB85Oxm1UlqKL3so6KoJ+zZjTII8yjrlFw/x4RYEMncxIgO
o2ZABBnRAC88APxUCokXNt/MWeYReHG/4AcIXAfjWqD6TLOsGySymkM426p4icpSHycGvLNhZHwv
buixglXYWqfS9ZiQDfxS/G5XdFEPP/oGPtnOs3hhe43G2PHmF01xIbgQPeGFMCu42cFkJTuVao5T
Ag/prxtqMv9yS6BGL6kayqWlMnZN3rROf1nbg0Wmk5zVutnoGxV7pqjJV9h5EpnMuVNwNV22WD6T
+hbLuLlhyQAYlhO+h63/1gtySwlswXIUBFALCccHjRB+VV8hygLl1eg7qf++Wx44Dn4DqJW/2EnU
V3L4cIHN+h6XgmI7n9Qu/Lp62PvIJEWqpyUZILxDvuWSMphr8X7kTlNjXvxxIBiUbsZwlqKs+jiC
zezN9FCKVMA0iWgUKWFMePcA0Pu0FewFMKN6ql1EhmvUiPSI37WNoFi13TUfJpbD4Y8nOARKmbmz
0LhxY7sRL5kXcQEzsgHZXmRN3xhIJ7/vX5Ma4xgpOCjY68MNJHAARLybE2RK2ipTU1h2BQkySQI0
italU3Lg4n10ArRZc1Ho+Uzw5qkdqxKaNyNjp/rv3HYhwuiofa+rzoWtVS6EG2LGP1xUNDa4Z9PL
KCvHc69UgYMdC1SxDcGYY/ibr/Vfve32E3BV9+8Y43AIGkMrAC/3vjffNVYqXUGFQIPVuYE7q6Kq
ZALh4RGf3z6BjRk9SPWblke4bs0clX3JUNSc2zjW6HvpSk3zMW5MCX87w0BJ6i3Pe/T9hllUjrKX
p1+8ZjbZp7zp9lim0qWwBJaQjOGeKeyzm1cCXl2nExfWeCjSWLUKmARIT8gU+njr9JreatcEtsVO
Ryjk5Qz1jVWoNm//aCxzEnUvzcMjX7V8tlq9snp1yb7eQr153TFTJgPQlOspy9y/krGa4xXRbyYs
iyOm55kiJDI5TdQqahQaU4lFUQOdgYh2XOYPBFe2FPelByQh4+aLtdMeU7eLlokso56PKrGxMhm+
9vd139/l22swdB2OY+2wRDk8a+z1BKcIqT+4NernBfoBzlZyCJoo/pKcB4T1HPbkLJ/IIDKeer8n
wpFrBN64gTbmXzwLD+/u30eTbAVjGt6wAjVGu3v5xJswUT92bAmvT1NUA2Fy/HqZRzsYJKEP6UCk
2fZj1fSdNWMjTBdVmk05jHikOoWBxp1K1b2TCTb9wMBom7mtkJDsNfvCR7zAZm+sNUWb/5xVKVTi
s8wOJi0HRWI6cIUIles5JB7Ygzc7zps+i/QyaYx6iQ4R9au20el0xmNqDCQuAdo6VXdO89KKuWol
WSR7kyuEHeE5RhERsE5JPIdX+81Ry+nKvq3wBDZotRfK1Eo9loXeyj2nXkYtncAxW+IrxnaVYvgP
lY8qrXppGubd+xY4Z6b0wfaIEAPCQWIa+4tOCmOOacXWO8wqazu7IAAfsbquoc99VV7yXjR3Ouwg
mavh5+WVsIAUiZNUnBwm2so06wS3J36wzEqcAyCz+OTpquKeqL649RA5IQp8hXNVvgc6l6M/6nr/
RuGxJ30nHn30KytBXs3E4QMWhkqHFQCOjbLJCp4NKnD6K7kiwAAXOfqjOHIPK/c/TJBRCGER+zsh
q9z0qQPXkNYE54mvh3g9VtB+qmic44Y568Yiw2w0NxQcuzPEUQk9IiaI0OoZzWJlXLD7+++8sxGy
05A+OO1OzUQyNUqsC/aKfkRI9p6hTjRop6il1P6xOoPGZh7PpcIzWwu1raNiR5UcocnMP20F3eYz
lqlDOyQNctxz6N3Nxcj78au90tLeES2QYd76+lIRZ7RbjgRU4CfOK9hSmWa2In690qb+7PnsMohE
xVwLWj2WOzNR+ONX9QT+7H63NR0OfezuLVyc5Y7KDDVjMpfj7WVcXbINOrpBJ+wWNrqzHnyY4LSC
cXQ2bpaKLlikL8wjd2uJMUt5eduXSMTazhPR5+siyGiOGUTdHg7iiAhuaJdWITmK7h7abt/b4Yzn
ATpHXp6WXny6ydyT5OIZzLFyjp/22xnQ3LswBndZV8aETq+rFt4NP1B758Q4MvBpi/1TNJunbFYP
8AH3yaUBkfwUPAQt9W2n8SOxVobkeZvCG2hSuz5OrKIgz4XjZ3eAgSlOg52+BWZrXRTdw450aqdq
M1HCPkYCxRY7huK0ugFGRYqXZ9bCqMQcXktmbGjJ2RimLRelyMlqjVf4MOLp6s1sMQir5BQ7THjN
wJ/4v5VvfffysZ+V2AqMO31Tzhhta11MbpDuOT9nHDsnpVVeJaRyOaWrU/8JPbT1ICNvVHqSN6oV
W3xvkPeuwd0Y77F/Ohvm3Dapc+9RErMIxogq4qXVn2OU+xXOnqFCSNLpgRHk0UEi0Pu5ZbqChiDN
HX6PJyVYZow7Ho0ObT+cd9QyyglHOg01dMBOoiKVgzF7MhZlIIIqc2C7g0nPThnQdFipsBo+lRb4
ZnsFh8AvLWNnUFy6VwZbmw/ly4RgvBdO1YRGbrs8NgmCmkVa3iih18Zql8R9AMym1byjWDQ5DPAQ
FauTiPzAF+uEFU9CJFvSA6OGbZejD49izGjs3YmYvawQ25cG6/jhjeIogvnrMO6TV/8/uRM6Zlab
eJkQnSHr6C1ttPwb/4qLt3FbMkV7xEIUVWApNrrOXomLNXC18d1JbdEpCtwVWWrGVcsGrKgBbilX
cDYMEu9nQlLzO1IaliE3n8fVhq9qKvDQ2BUeEbQDnjZ/Si4ycuWytW4GKM9L/0MYGeRapYQA5rI1
qFbzJqjK+tonnIT71dxGt1KLBXbkVg9HPiJ4cQdnWgnAM+hDI3Po1RE2mF8u2eymSg40JOctwhXZ
3ALFjrokSWrzjAeopuQ9ZF/vZgCj7cmb5wXrHLg9/sozM6CrnUsV3xjH8Rmcxxbd+jgX/BMBD+4H
nnX1Kzg3+evDVQ3Qtumqx7PW6HsvxEXgXw3M5PQHiH6JxgWXn6O4Yj4DkzNWZeC0RWCw9H/FEJuf
M4mnEKVWly0PR00lsqqnQONDKxY5DYTIA3yOGMu1b4tYWvZD3CRpWKaEvYGqSf1xMkjKdxDYgLx/
ZicobqQ6+pOfoXhE1TGC9Ct3QvfdPrmtrmx21LLT5WVkAfRYK57M094eN4CzfcECmd6Kl8E5VdO6
siBpmMct9x9YT99T6fTzRvOLwNeCI9RbMaHtwAuXEZNKo4ECwq1KXSlsdfe72fOBRekegz6zzzTo
qwr0wiE6b5yAk4bOVJ0YeD3k5bov6dkwZlE5VqtlDEJU81qOQj5pXsB2r/T0DCVkhyYVaQUtQlYW
WvNbbhK0Hk4wI4cw4wO3cPdnEs+sJbvUTbbJkj8uTAcrm+brxurUol31c246756C8waAST3jG+iu
fy+Fl+heBaRkJwPLVhjzziR07rKPtmCDZhB3HfG4HlBA+xsYCbgQ3cjAAMFmcgTG/t+rhGMhs3Jt
l81GCHE5vw/FSTY8dC7S7iqlBVmP7CGMvnHlmltrm6uNlNPF4Q3Q6eNfZX6KPdiEuz/rbsyITh/1
ZqEdjHLX5ieyZGYxtFopQAqgDZM3Gbqm7itqwVZivtLsy8QUFd3w9WaILRBNdB3+qUothQ70Bm9/
myaLxBBHvIeLxh8yyqe/b0VCw4FqQLoVoKDGAcWUaLZzSFfGSmYfsoFSokmcJpFbf1AkfQ1DekEC
VsKthsb203D0DhO0Eizdf/sbS92BJBTUTJOPcApfnJxPXe6sSZLX01QQFFLK6o4ulbkbfIvq9CwS
wcsBrZmHlmQVktwysB303XCdhF5p1jouUUo32Kun9geTH8poRF7n74VqcFJkjrWpCm2hYsxBMhoL
2Q6cOPFTNzwrJXrp2Rf1rpsgPUkY7/NjgIead2Y17WdFtp6dZxUS6iOXnffONjxBGS8X5ON4FXsT
AplA5Pz0f7BEYnBfb7Hpr5zOtLr95S/UO7gUNwYt8C1qqTrmFm2V/Bx9Wt7GD5grDAFZtZDKRK+0
o9x3vWsg6sqRl/keJolbej9d4F640iPnTU2msB8DXZMweiB5ZruPoumC306z9g/lfspFt/9P/OV3
Eoas4ixf/cv0icsEVJMRhx1aNjNytv2xBhtYMuUp+xZfIAnX2PCSackHjf91pS1BijGAfRQL53Na
hYJkttf7jCfmmqkTu0DHhfNC7HTEXFR+yedrJeV54A4DiSvp7YF9QA25IMZkR1C+a6RYJKBqvlUy
VEO/94R7biAObmtwS1SP72JBqQJRZXLqsYMsJmgwN8HFOOVzTbXTPQz2k3eGBpEVr/TuSG8h8AR7
3VG9Q3/4o26N3EGfF5rKl2cWXZd1eCrgClpcZrvKwsDapk0ArOwJ51bLzcaJdJc1IlFY2lZKQ24a
zBg5sX0rOAJb/Kl8akLJlGtZb1sv5JJwovfSHKbL6jjqMRVvXEDFugETExW4tV87+PfaGxIxN4zF
UxbnwGFImXj+uiuWZ4xsdo6/4jHQtaEEe9bAmS7k3QJjL8TsARsUpYJFBba75iX25lu2EbF2XItM
oIk+cj5/avwBSYYcfiJFEGnh+B6aDqVwT0wCpkrN2XecMz1rjTdR9wLrvVOSXCSbFP+lkdLUOsk9
Wam/aCLTpjU9gL4hSdArkX9UdbZryHDVQyfDUaBp3bl+WrJc6SUkUxQmLX5h3vFPWTFDkw+XKnsx
jSNZdX65fWmwbR+OssvRojVlGhGRdEBP1mnwfWdUfrcLfz+QTWxk/CJgbLLGq5s8z9c3bjoZbnrH
vwehq1ZpkuUAajVkiiamXOxGqH5wKRHhEkkyqgYoPgxZXCRN0Gnt2v6VTwF+UWS+oV1pUxGGceJL
pmt9F4Xg6rzFtBul2tepVarDAseEyDdK8xrBvxzrOH5hZG8K/yCWxYevRUSXqyBeJsoM9heJdqtX
+giMXhTpcA3bY7qjSASHOIub4MDiPq4VsVeIwkP/1lIOv9cRh3i1LzdnKdAhjiNxUU8867p+SNC/
2gIyONprClPZxKKTmZN4DLk+lsEQsoWn4T9IkYr0VnlC6XWRPlwHGJcyLE91ZMOPO6KvZbO0I7+Z
C+PS0CgOcV5NJZtRQCz8F0XmWcbVv+TF3Zpfj47av7ToqREfvLYiIWioGUWvxfnt5NAforiGMaHx
Pamrkpt+kITNxRq4F48Gb1/1xQTOoLCozPfBfzULuYPcVVyqNbLC+RRboqUABpx92PCyx+Z9NKod
iUKGmGKYed8QXfsmuu4D10Y/uiCA9+dF1iSE3R4Iu9QXkDUj5V7XL8YnxF2QpunHyAlnt4eTLIj9
k4kGPJQ51WRRvVQa4W+SeOS0ncKIG8F6q9RSgciOj5mHWvl4N+4YFZSpKSayWn/CR0aLWGJfnZ8g
HWj+IyvwU8VxM4i9K4CvFjaJFVbN6cPy9dc+GLYYx4kNlNPvldts8m7QKp0fy7PofcxHQg+rykxQ
IoiymtZaTSD73HOYhdWZuzFppSPKn0dmEBxeKcg0+4dc3wAqEB002QUzbIvSxyk6k5lJUqHTeHuu
SFwoqc4e4cp/WeP3YEsfESssFgy9boU3MSnyroqnmzxcQXOyVDOfxzvifidymH7ugyGla1ONtWGC
mocbzgVXw7MmeV7DHmwATMGJpsO5B1AdpytRLmeMtQIe3WnhjRB2rJ1Ay9K0FeQv92hc1Gz/MNP7
JDwoc4MPMXvjVDRxQynfSKaNejGf3+lm7YbqEow3QZ7cEIMUzQYz5KhIvctF9b0SeQbZ+89hUazi
YCzs4odToOKkAsMNAVMUeK8fjqVL5cMh9gGrEtpJ2rzvmBaXuIjV6nUVYak3TSCw9Z3+okSx2orP
HO05BvCE2rsrEMRcZy08qBh79Roj0vPrDMMYO4Imj260iad3TJinAkiYXKRUreK89lJyZ1uvgrHM
MYRxvdhhktXJ6BBEe7t+pKIIfj+d+sU2sRUo/wl0Y4UtHM4Ci4SgH5TpfYOhKtrmTmihoR+qIWo7
k4nAWg9L7gYCVr90bAgxDIsW879zPSaEOZi6Y4v4SQArgmJwNAa54sOPplqYer9f3XESCd33mnTU
MtGuEgl+z8P9VeYYiZR8OrCIPzvNvuqLbWQJfxE76eFLH4jgDDm0lStUN7fep3VNHCQOsILhc+Fa
1b31amTXXic1eRPTih+jGf7eu2UZxzj/vmwsxfhwLyZJYtir0usS4ZX4896EvEttCk4w2gEHzpuK
2jY0Er24wV91Nxe4ND1vijpeeLpH3gZQdZB6fSzpOBXjfT6skinP5FbiNjjHyH9YryTlPFT28I98
tyWj1NlJqIV1i6+2lsfrlUnyQ2ic8A+cqshDhVAAR+5pLM29n3nwf0Y1fG/rH/Ec1lon9ouBkQNA
tWuU6HAEQYCmgP8YeLn612a8JwqufFmwJMA3dPpAIqH0DXZCibpIxnHRHA0rMHbt0f9ypV7q36U2
wVlMJZoyLc8l/Bh1IonY0km5yZSdf9g6TLrSGP1BwQTnoF49Gyr2yYQnqjaKY15lPHMhG6LCC6QN
YkN9La9SkF46A+kDM96eHU9fr/TdmyE04Z7NNTYTdPdc7u29wD02Q5xUbQp6GPHg2ibIEKmc9YfQ
WYaEpv9W0MN+IzvlV8bOhlzU1QfdnclyH7O0Yeopsc5yATKCqiODrZxBZ86RIivQiQnDlVJctara
1p12DwV7uSgJGkzQO0N51UHbrAWpJWVYVMdMnzuy7RipdgMAEcHmz+fPfrMdunpGUvN0PuaQt7X8
m7ZOAiw7Rn4mRlo/HqoyeyBuE1XAlIFNN+fRwyyvbjIL61HrIrWUi9rUXGynKm/GEaRIzPrIoJnF
fTuLur3QNHRCH21DmKT1+89xlsqUzktDMPE4Dqgwb2S2OUr4JRqTvgv8CWdO0mHKl3OFrT7i6Xhm
tDDYeXezGsqeOmqz9ogCpQ2l1zNx86kbwDt/0nN95JG4yx5Aq1EWlW/dhFcMZA39i9+Upuc40oXz
uazFjDxn7q9EERyxmbGHH3q4oSS3IwAYZfHdRtS/F7VtbLe7bpry3j+xDHeLMJP67i8bUxSaliv7
FTTwszmwyPlf5FEmLW9GRo5ab58119n7R/aemelyv5dpE+NIwOdnDJqUertAF9Pt6K6hM2AGCXHY
dP022138s0vIvGINIXLfQqeD5JfNxEUGPULX4gCuTBgdpKca5UsvrZSIPqXmsMJw54cNKiR+Im31
J0DjiWkBThC+d6JA2BZTp6++torKimCWZsfOmFBlpmuXhba/LB7ixPJJ9FFGF9cIvq5S+kqp7LYy
iASuLsrYp+wcXltOfLewGidmsQRbhMPg1lBdZWpWEi9DFooBfKzdMJzBzgBZXU9vacbGjr4POVgo
/bHeRIE9OS8R2+7Is1/dzHgGlsTbKKA8qHhpF2Q1rv9fHQ+oo0g4shUyfMIb+3LyJJ6Y+tgGd3XV
BFvfg/fpA9u4pMohUpEF0nC+J1JT5WrXLcwTa30N8xT9pSxi2NxI2yPxaX15kk5g8w+UpJhWbNU4
A2JVLTc4b3vHd5gueZPL7l1Th5T/WtgtOk1+w8nlkjmjD0qSIMs/2Twk67A93PH2HFOKRlTcoSg3
noBUOVivQKBPCZWufOlGgT0PFKBlBODFJEck9WBnp9IfWcApt5B89iF8MTIg16tPv0oEkTrZGNpv
PUVVyKUEqivtLAh6cFNCiF17oHOCZva4bDemYzPv/EUVToGi6uFhVRvE1r0Ve3IRY10q6B4U8IAf
3xYmJz6GnxlRqh8HwGhz54c8bAh6PWE+ZS7ZfEenBfJeZdVQFMsiggjs5CE4Z7M9AsHUJBYC6Rye
5nvxMGb0vs7tNrx2G3AvyMGApqsmwHJL3ZvVdc5tSvj2MnRKAo84c0W+mBc33Hq2XUjaNHOAEvRy
8FXnrNHMGLxqD6XS7wPiHM5z9p86+/KNgK3ulGh4luIW466O1ynuqbWvrLDiWnZ88KGRyUUBYjYx
9qNJdlPygZJgCki8MTAlM1zTetufrop/YPGw3zTmWIEpSpZNK6u7ZCKKixCf9ui56uE6Flbsx922
L0b9OhjkoKQHPCf7CjrgiJVCp+CuhK61aGs3FD3bRBsrG3UP6ZCGbMOWSm7wsWSJQbeYU22calDa
ZvUQfvRDSw+F3eKVKvJIUZ/HdrcYS9QyTXEne2GAWm/AGDOLacheIjjh3swDsIJ5oR8XLeIGznKa
Iv/Wr1qAoPLqk4WiCE5D4C5sw3C1SN1qiIXgGc8loLeMs7W1050vZt8h8WZDC+mmQUPrLnmuI7Y3
iULrWj+tQBqt8hKJ8KkrLw+U5uRiNVPwUQRIRhcONIs4KC4P4zUhARFyJVQOkcnA57akmjzaCh7g
nGLjBvzdFO3DY8VQu0nB5KsCIPd29I9Qsnm643D9N93rR+VaZ16hSzQ3AiTVPCZ501LK3kylWdmF
PBboip1Gins5lkUsLcRq5HhW5/OAiKx9hUHPCiRVxoX/Igv0+aerkyicNb4KDTYjL3zBzFaJQnWv
+5BiCEPMZo4qc2TjV7PAjL0T2e8dEe2WE0UFLfra+CmtzeI6UVdj0DXOgUBiZp8EljpWeLjohxPs
3/+tLzQ5OZE58MkkX5Vv0jN0zRxwDM3mBk+PnPGjQl6hf2Ci9IGWf/exuDpz9osc2h5XghrNthUs
uu7x26g3BS+VAw/tOp517rp3eDugPAFp8HLPeOyMmLFwQFPBT8E6HguHfd9DPTddFWOQ2RPkz5qt
ZPNzuptEDZUjHjBEqYP/Y/xX3Jf1ZmeWN58SRZ3B/Lj/A1lY1Zrtk3INpQ3jTRnlH/9i0lIbIv4J
5UGrN5cdj6gCnkxpT4CYqCWtXIIhim3zmiKIoe1j2+cDZCrObEEEheSpPnQW1lf6nl3lMPIWbxVq
xLgGTDojXIdWONdNIYfIzx8jDgNaXjyifP6lVDOC1bnNnDM/g2IOmVKfBsLvZstOu9IjT9MqnZja
AYU5gswGwxzWoFlzEyd2vsN2oJ3JmHNfZKtBCqJGahhirYPpU0iDwj4Tidc+dmZL/kwJ0y6JpK5B
RQ4TioWOxPYbEcMrNSzeYtrITvdODtUilhdaOMZWNluQbfoqItoG/TGEJId9fYGUbqLJwum6bTB8
K/NFYx2bbBwuow3auqeG/PoTyDzmQQ0Z7ivu6cEg4tiFRB5Dlxe0iXw9eMlJU3WKmeQyzfPCTjk9
CeaJVHQmLg4kjNSqH8cUAc/pDFCZAlSwtnY3pkhDRYiucWrV+owWv34iguIPUqqy3CTJrVf/4aK9
G9tVL9+xf+QySIOv/3T01hvNIHa8aiBa2zabJ2D1YI91rTPR8gFFxY+IqgU/GekDb2LQ78+mwyiv
3l+V/wirCaMOeFRGyJzplWkhj5NahM0OF9WEmkgbkzzQo4jxaDVHDLFnn554ABNqgtcEymY1cgeF
jnrKmNH5tn8LuyoQ+x/JAGQv4f4JIO0GAyKiiT8n+06uZvebaZ84ZvyvKAkQ5VG99lOFGOBPf3oJ
nub9ZWEFtR2RPyhQfbNbV9Mdx9MrrD2oS/AKZY7hHfUL/VcswnuGfniAF8F02Ir2M9D8NWtcVjxF
SzZm/NLuqMVoDtjvZbpLNReqXUEj8LwPUltoD8FBzlGv1UuRN6AvmPLFP1+RN1uJv2jolWGKv28+
8ETwzj13AvFAgl8OoMgQTtF7Eg5yJJhY7KgIFLcwUvfXgPQ8kmtx+NGJUo6DCu/h1KE0NgzyMu+6
kPGgm/nWuvo0ceqesJJiBqfhkxfdoBMeAeTO1NYcLWS+6VlrhDAQ7/8wIw1dORNkNS7n6rY9oD13
ZEzAxGrbpnAP8QFKHmsQ3vNkCtuptE3kV54dtt6GeywTja9fFBdg50G7BEgiZgelQlN38jitrbk1
QWAXSIsfdrR5BIWiB+n09Hcehy+kg2BNvqE4uUTkQvsNtFDm/jATpg66I6K+RGKlOhOS1AOo7w2P
cT5ZiMTnDqVEZaddRni1BJKLxxDgkXlkzjkACkcBIrqKM5bl77xEEwqGr9BzTF5pDcr2PKtiqwJF
elWzJSwWwsnCvPrtQDg9xbbBYmdwr981gwe/lUJ/0WuD59nZV2eDoWqTghqkSL+eK/BHbfxEXzd9
DaNncSZjXAfDrsq7x+mnCQMaBPhGFY2aKLI9tLqwUEhMtBTPWnmPx4hjUkxCo9mda3QqM/3so1sX
h7uG2+7nqSYMDCf5gAunPWTaFhtFpMq5YHnFghmro1uXxPiY+T0H+v0xgnSKANFHP4svRdjHRkOP
wg/bs28jtHxB8K6vxqj5/8/dh0auR2P2fsmAWQfRBXjDy8DFhZtxho8pi9TA1zIRvaN6Gi+vqREH
aCxTff+4IHLK01/l6mS9gMqnDo1lEZbpEql1naGLbGoVdg4p1UpU56tPxdw4eNoGXek+dcc+k3UQ
v/2drE2vOUC1Z5l9nzWxe6ERwebsxNLPm4OQLO0nydJl+HxLISLGyUnsdoeI6T63MYa2uahQQuMK
EtuD9ou0zcfQciF5CIXju9LZipo6bdLkM2t/lLGNYnsM8HuoV2gQ6mKu0NLNUGP+AHWzFvFhSifV
UhLzXLQjX9rHiOghNNxC+31jDBMsCQiwXIfpMhoO5/PIS1wjVybTMvwYAaDn2QrFbcTB+KyjdvuO
xJZzTNLqHtlFpmIity7O+x4tKr8H68mqK8JmjG6LrzAOy0oDFMYDpbHeebKycY4u3HbEG0XxM26S
L/H4Yltto/vfBnesUHIA+xFuMJaqBIYH+gHF6Q/hS2R5znc60fVMOELuQWShBe1Q9x7og9rA66vy
DY20iNU3KwaJf9N/d7NEEp77oLpLg7QqPha2BFsEF1v2UX6kUcdnWBrbkWLwGQTxK8Sol1ZsvMLS
4HFMbiV4RkcXP0FEP09yeSYp473eK6JA5D0Rio+nQsTmYfoROm//EHXr9TwiUpWORJCBtLLk9d93
lyG0dp4U7I9VxfgAN8q9tW7TgxWwmHlahgJQUwwQoikwxv7CU6eH9K1xpPwtbxQrXu7IS18O3sel
lHlTGcsNQQHR22BnAx0Aw762gn0lEreGOOTyja307gk4OXb7AIqkXUVpkEQygwNr060b+MS+jF3T
Nf81hLmEorPYxCpSGGqnwKYaXbNL77t65swx9qfLIJ49/xQ4Qcrap/oBrXNnXr+Jv5eJghP+Fpwf
PrlPvg9o1VH5gkbYfMdtMy5MHImInTgEtARilsIy54WhJiCXdbYFELOkIyTWhpFeInvmLVnXOsfc
6IaW5OvBoK+D/XbAIorYGp8tn/fzn+GM9POgM6LxVUX58pIPP10iwEUncYCLjrWW+03jAT0mDSk7
05bhICPHm9DyHM0Xm+XPNZ2xQV7/EVnqX0iGBq33UEnLhcjfGG2zXhLjFHI4+NLTHyNVjAIjWJiZ
RCk1a4TN1gvidM8c8ekGqCcCbARqHk4HMfpWWDghxHwJIljQ5aMv5V/8UdRBMHKXgUaxfPqtRaIV
MOEit/EcWtEfzpSXpNGhmaT0C4g1GCtsDwodOZ1ql7wSA2ywC/vrHQ5H1XKBKGlZY8ivFDcyLaGF
cyFBnj/BVFVaKzJ5EiAEJ2AQ1XAkZ4aiJgiXyrDimZu9oHMSqka8jxG1QU9eBTSVCSWX7ctWyqoI
AGa2+JxhL2akjANGbemKlslxgR1SFbzwyMfuR4UGlJaLKkJAL5Wsj0gxIBPNHXsvnBsbWp+2D0An
PYj+1XQB45M0lnc7a/Zuc8uSrc9KrPk3PVCJq7rrdoznlPKUpBT63ChA0x+0l7J/kti/ejVaUTwQ
bGAFPVe0N8SrIEB9XFcgmtpX57W+iS2xrjLyY6SBgY8qpYSG8iC63O1yhn3+kjGx7AR0hvVLVZ2C
COQROqs2YMQkqzvigQdFxPMUufUOzBO9cmArP+5Tim7oCfXHo6T3V9S0ODCupX1MDkUlvujI3oLw
fhACBBwU6CTa3ybvPC1T4qf207AXpiuqAhUx4NFN+RkSiSJ1RC2G+T6rx6I2wfGmkTgIiBmd0vDn
yBY/cfhsRQkahvOvEZpB6kkqK92cpUtoGLTOhNKx6ptiOay/eJcEoIEguB/pXtVh9C9GombOOVS6
IqBsLWGpOv1FLEWjj1dQoSW/An9BuoNjFd0eqOp+bnHqCjjm0arF8KItisGKNtwXigpq4VbtHX99
TOI+ls/+bylB85cFjs4qdXd30xS3eJ/enVZ/J2U3hOg5CnhAaoDyf9EBQ47gMkMof/2uuciuuFeZ
5Vyqc8q5jFbVSyPoIeXa0xq7C0K+gewycPvx5vk5gtWZAzOoGUyTAzghL6AE6zAAbJqgDPOFRTP0
YrrlMf8Tz+mplIo70uNrRCYMsCBaFRKlLcFJWYtGF83z1j9ACtvRnQieJrH2L9SEwMxonXVQKJUR
j3RXpifHFj6CbptY+jG0FWpJotysxaMlxWPts1OVsnpRl71OWZTptltk+3+rIWxmeffRrpluaKKP
2AWaRajh0sDqvri9NkNmXgxZBJSTKRInZdc+g4Yh899ZI5zlPvkHiarCCsfi1SEz6De71EmgnNsb
dk7OR0x5Zp7t5HzfFixGVgS0lEF/OltkDrac/bqf6RvPzkzlLHOzmA94e0gdiFv/e2POKouWBYNr
qv9egYNYzDyn8/hvMnHDZlf7wlvgyBrqsmLXr6IxcMdc5CqowvM/FF+qCcCt7MWTYrIcFNTo3lQh
AMO4D1Wzrr63gnKr3wzxtUh017ratPcAPRJllKtCgUB/7AJKo9RllPbt0ulaVDyCbY5ExT7gTue9
rCgEsIISZRrXSND8ZdEfSxBOr1N7isReK8zh3fKPisMtRf2sjHbDP0Y+q1+Wrwp86auV4yWgzh83
dyZhfRuIEkwdByiXuO6/02Cj7pf6iRdTCnjZ9iLpjBxp7jOkIHp87FbhIBG1+czEKZPg5S0KVCt5
0uuZm0xxeTwhfzGjcQDI/t5ZcOKRZPoJg47psaomWEUhT5S4s4aT8y6XI+nsGIGEGNsjny6ixt89
R6LsIzFSkuLSye5GHWDRmtzkvDOuzwShNT4SBp6YSEiAOVTWEmdAi0mkkV83OYqKTHM1pz5YOzBR
xNzjMr90WqehILRXq0qTClEfb4DSGcuePPUjGG3ogdMpfTg1r5SO4B4mzF3n602SvY9cBK+6izQj
9S7AIlDkIqotck5wExvtq+7IOOAknkDGgjTl2WUf6RGJinCu2i7oo0/ErnGWBabB8+KG1iQox03v
HtQys8F7hN0tvrVytIQZkDYpo3rUZSMGL5g8BuIhN/1a5tKDMvgg30ER1KssHVE7RpiP4ChNZRlv
2bdbJ+LyKBl50l7amnpp8aryksBdgMOyk+bPauLbEceTxkm/1IPrzEU0vtaqHFPVU/BwIOCKADKz
tTB0wdlVqOc5HGzLNcunmgwRSvvkTJS6HjewIRIUIs1MUylbShz5qaOD6MhFl0AOgaVl58vy1bTg
QVl+BDcCU2ps3pJ2ZSmBCnBbEu+STLhEziMMtvQTnYVRFgNFtUoWFnkpTrQJyMREsVC873suS5sF
cRhF2widLcFXRuD7SoBEOyV+EE8EIK69QfJoQ6VzyQZSjM+qfL1l0UL1QGcXKcXF53qJUVZ6qcXe
FuiseGXQ8zbP7fKUqexmv1s8SGWcwxr7HvHGllH6OqcwIEjH16de7NAoe5Wtqyp+6MRaPwi+ExnT
MWl9HM5o9y6DJQs4y+xSJTqS+nzQ1qAs6+l5juPraMsPprFArakDhwqxA2qhSIsaZ5TGJWFuhUNA
0y+C9lFPhOJw1qrdAGQ3tvexif+vUDhhwIbwAHfJyVx9MpZhEMw+uRsTEtRkki2UavDiJbuxiR2Z
EEtvAuja5cb/TtOo7C13+dFfAReFhAW8ZwiAYx4YS+KnOL/WC4a7uDNjK5DC+tgzOvhQsjC2TiZH
vzxDpmmpfCEs18dAJShAkBXkPiX/xLd6IrxERbQ/pZeA1Q8ZFM0OvFjiK1u6QMlyBtY/X+s7GmTr
eJGfLkIU86tMDgxOXqedUQMbzkgNyRC1v0EdlJ21ukkI8PlpdMTHE10r3wKnZCOYuiZtZG9Dd0bR
RIThA7bAh1CVevf68eyBDd/0LBoDIl7FrXZM1cP3/xr8la+6wbtCLrsmzo1pt1DiTxOPDXXc4KKY
B/RgzChhLbCdna8w4Yy27MKtMN1aAJm9Y06bQmoH1yq5PxVqKQyTNmwT4kXr6jybOPPxVRdrBoOE
HwpNrg++Ypx64gdS6/fOX/lVDri7UICoOaMRMcTqV0I5HPxhQICyEosiBcfgZVeChLBIlHmrp5L4
QvV2UQWhy0GulZxBLz2SDlvGxoA0Uod9B8/qjhOCtYG80U3eK9T5j8st5zUfCBPdukaCGQ5NAWkI
aZhGVLQ+VVRQRv4pD2imjwsz0M0XNmscxhe6miUESxFmC3TbvI2JwXsOWOqaElENNyyau5xkHJYG
7TUpHEfIGmBwoSSWBBnj0wLJPkg4IDymrybwuUTIH4DsQxWRlp6oYdAYkZ1M2OVLb/PnArkG+Fc7
kZnR2CZYMMMNGnW6/clo/MQpYuyH7Ds6Y6hTUBEISto9qbv4X6yB1BwW8seu0sePXJj295Fl/ZkK
2KPHRqVXBJVLv0divsYQkpZ1ssW/ghpAZN6+dDRskfduV3okNTPkJyCaGqGfGXZFd7YhxS/VD+gH
yTT5TScpNWpGBg/2W+xZpbCrL8tRQNacNnt4SXp4jKGYV4mAoW4AARZK1Ddt4pZLY3pLebMTU/Kh
OK0xdoS6mCuQch5tuIFvOi8f0e8Jen8FSnYLz2kTpbK6n3Fm9zLn6lg9OqL77PiPwT+BGSA00Eej
5S0Ck8+hKo0urJ22RIubsWLDjxjzpLmiCt3Hrqyr9SKDe5s7PXmB2mqgmTDaDQX77KVnEx3RRpEn
W34Un+og6nyrQ/OLM2OKGUl5rALcJV2Fx+UB0aECpqYWyGnrkW2l9gdEvuTOL5hmueLjznSvBp+i
wnJ3dYT3nNBvzS04rU88SRY+PtWTR6bkAhLh9eRvmABp4yb5bRv7+lIbiO88v/jlMcIdoQTFwEBT
Ps6CJyLC03CWLvAKeLaltrEAW75uONVbEcPXV/LvqZfH1l3t2MuKGF81LLbsnNQhTrpnw+9g+i07
d6RHTaHFTAjocdlm143MWutC9/7wJjWV27WVL4EcGrl+grC1LWe1PvBnY4mNXErOaR/YcO4g8W/r
KKf9vw3PI7RzNPjU1wjMdCEM6Q0oNCApRLF1HmMSnWD5qyN/mY+i6uroD+9f8sLQrlmtY9GOeJNK
eeNJjCHa75rlcfh+YqP9R7gdt68mFBnlE16I30fTLxbUTx65JBmUZ2C6i4touDk9/Q8oP7UpiWz3
twsc0bbGX9k0nzm+ZlbuCl6Rm9YkWyk+pK1mIKNWSwy0RArFuW30U+G6heGH3MdfpMYE/lFXNR4i
UBkttJoLfxwDkr2AR1w3PsW2uy5Tafc76ktBsrJu8LyuadqLxoSks+IlDtTFyePl5m6w2gZaBOxz
1icyyt+cLeb3FtsJ/nAdW8lfjR2CAFlCvEVNHm5GqZlZEf3rUvQipm7m9Hggi10641cE+bUnPl2v
5/dsFA0KNqrUIPN8yiZs9eRUl1456NgAzQIgaxkaNIWenapDjpqPF0XbIsHLfAVN6GLLQpa8fFsF
2FWJVg+XVyBgpWmYbCKiaiaaMXsVfOW+YTtU/fUQBmnxKPihvUZLk8VezfxfEcd7iCMzlymui8Td
8LqncBvR6rc5jbeNgeSzbWjKQi5ZX9HSz5ohqjU1tMnSAlUgZnrl7GdYXc46d4RN3j28ci5v0rRC
WpyKnc22v0KCIdkU0bR2JT1U4WKnJLOgyFwF7Mf1btD+RC9oJLzTFXFQ94shckMjrR1dkFlHut1+
5FS86rlcFYbjl2dokY16mOIpvlCJLBQXNGV9a+xOUKgpvqM1o6GsgQv1gZZoJYpmDk4ZrN4SQLk8
MBmK03dYwCDs8e7QyAflo2clVsOZyiQhKuUaJgl69is4LMZX7++5MxidQdTxgts5i3pBA0ogWNDi
W21tHYfTM7HMho9m49Ohpd7jbeHwd3OtpmhmsmEt74Xfd4W0+d70Nkunz7s7erQ9wRLjeFtRB5x/
sQ+0rRIalJxrb2vYo06UrTp9K/hYYDRn2BEIXczV3sIyyxDCh9E81Ma20TJFEdNLll6u6KYLza9D
m0LqsuXRisXRL41YA0NmggfTf9z7VRqItUIt215dAiiVq+6ltxiJ6sCL7T5o/pNorD3Hy27Q/4J3
kzaP9SZlrAC19t7p+t80zITkIHgNWvq1soHPoiG7Q7QSpdBGIk6+gcXn3CeZAFc5k0oRlTEO8tAn
ojWY43M4lN+sVOv+1iMHJlH4MmGuoycKK+ueau7OUpiLXkRvr4uBz/IvjoNFhonZU3lWgsLMsxhn
iin6noQ8MKBvyMHyjpN1s2483e5lAZ0+IruRUF50TSkBGuWyhSzwlPUyTu4UGd0wF9CCtElLd3So
7OOCbTDYqFSQqMklxm3su6T176tl+c02u+Liuyb1Y/BD7K9bTn8qjEoYlmvJddyAcCUSi3t8ch0y
gDRC+NEc/rxF/1r90SEEqgnt2zEERAItQggJFV16bvmomudOuaqNbg5cLrk2s/2E7xYGNyhdSVlo
7hXiT8GgIpnGDLCFcUSFxZ4jGKyjQEPCXeTHwFnIuUqQPQ+RBZSwBHNLnnvyNGnNsaYzEE4mnHNh
jJt6qy9Wq4fhzFYQimPJ8Znh2xDMmymwvPwFTY3QM/7EAaWX52dugdKvup6u/FyTlUxB58OEVZWz
yFzXNYZ3Fq6Dj83baJ40jIiLj9H//7qCZPpOU4gD5gdxe28ebea6sduTGCu3UiNdKXLzpKUK26t6
+Ty5+crLyXBSoUXbfNHG+q0oDkS0hN3YNliL0i8J0ymuA8/zacNb/qyquM6Vvno7rEgI1rRx8TME
yWqtzPOyCSxmNo6uZ3jGCJq1F/VZc19EiBR5Iygq4TyzfEDzY1AX9JX6QktjzMUJmnCkgocB8aB5
Cfhci4Ak1iFpUMbnSjnHijG5KI9xL9Xtq9lwPnOtwXrncFW7+NaO/yBexYvaByasmGTxqpMsSsXl
Fb+rD84LpJ0Q1O6xvE+J2g2XPn0P5J1u94Ln9nIQCkPY1zcPhYq3xOamNdKglyCf5/rHYN2F70f6
jLuPzYbGe956XpApH7hLpPFDrid5lGimQCV1icEnUd0uWPER8KTVvQ8bfWv6Fu5hvuDAKMfUgw/+
93xFqiL49aEO6mi2IolqVsbpq2nKLD8+OKxjTRqeWHnmxPuvDrZ1pCiq3iJ3owUD+RUmXI5bxxQm
RT0mCpYpv+cpE3YQSf693pWMGdnQKuWQiN8gck5HSvZn+ubnD4POnt6S929d5gufj945yLYOkhRP
zuQXyrpF1bo/75jYgeLZ7K3VsSx4pWYylBGaMSrLgYktur1mce0uFXuXHBKIR0D9V+JU1yCmdsrL
V1P5hZLK1jjEknkF2xx4V5vT7sMYFsnFOLmZaS3xFQ20GrJw+QtkEPKRS5cBxQ5dwIJHz4LzX/aY
bhFe6n9yHA9jtNlSNFD7PlN2W9fSGCDGlzmmTC37zPq6FYZuz0xrAz9jPBCE0GCmndquQpIAYYCu
rPbsC8chAstQvYU247k0D9jTNDpa7b7if8zcZ+FfTtj05ZZGp9c7ycVeVameiTGQmcyp62iRilXB
G/9Z1EL7bJroqEhwKC0QRT3IzWya+Ts4rOT2p3Hjkd8EOC0yqXVfrhRtFJcAKZkxugzH1Il3ucu/
c2OevU2kxWgbIyWAxXerZHNjISd++SD+WrQuQp6EEJZ4RLLt7/afYLnQzPF5VIJugv9rBq/O8jk3
l8Uo0Q8sHuDKnm1Gbb75pFLWth1Wwc92pBEz1Kb7msGXic42W788xr/T8K8JOTIT8ld+44zXn2lz
4KDj1raPKo8KMghmhZPjcSAthyXXqu9l3YZJo9a7QJVFTEj+Jk8Zt6tWECPj5Qw7vWT4sXHwTpFf
kNfkuDVETu1tovI3XFOvL9E7RujpJfnrVouF80GQNWf6b/W6fEIFTYTBLl6PR/CsczCaXrkiDJsP
0FwZMrSksodyAIqCAcv5xRdiDhht8/mjPZXkWDXXb5xwB5U4os7voqDzH94NYt5FEvygv1j02p5k
e9PSG4uD0Ti2KXqrNKZvpMLeJKeQmxMpKEThaxYQe44RQHSYG+30jkHUG0PZZmjzTIzAAIPq943E
6vKj7qNJk0aryQ5OAjecmHpaIK+5zTAdLmhl2EevG1YOQG7y5Y+Fu/17LeKG1HWAo0yFZIxyw4KA
3ssFQfbbXcwUgISKjGGTym/1Uv1ImuagJJum+BYKr8KM4DQuNGP8ZthujfBJBIi6a0wqNgwUZ4bp
Ft3NxGQdFtYGuR7BF0x5PseX5qN1EziuGaamVsvkkg+CqgelWP4Mdg3VzDRadce4WjATD2TZuuL8
Iwrhf3lXHDvxXsPkMlSWZOMYxn9pt2WxA17w1S/8Oio0jnj5z8Ok/JkBIzO78wnJjn+JjE1H0CD7
T4kGFKxR16GVVKygcXGvUJWr6aNo6A8w3annY1tUsVHvyLmpRg2p1U7goGqOlsj2UyY+qc9OyDc4
Tw2UPKckhKXi/Dy6shJb0TfmWwx3HhcDmwp3vTLoAq09t9/34VF45SHyW+z2tCNo1Xa2ZLE+hPqe
qrK50/+Jd0uI+T88802zdXZWpnTpb9K6fK+RlG7jBP72LRoBboEgvVIFJ2+gxqgtbQ/G7p734wsZ
oZsbwzB4RX8gOyJpv7NrQ/ic480urUhl6FJrwfwGzHdqfRlUVmzD5aHVGmenYZxsxJzxr11eLPJ/
vhTfuGQJ2U5lj8Y4wTIfvfUXABVazWPSYhk2k4gKSSh4HP1HwfWv94xj7hJMDiKvOzmjYZDv4+5p
XrVL8cDEhkULci/vhfeZ4JMjP5XJ+8NjHXT66k28g34Pnj1WTzRZoGE4dw6r9S+kCnsgeOGqCAEU
y4UzTFJYcowLqMMEMLmzeiHeFAnuDyhDyWbNvCFl3JEpGux7hk7P0BdHld0f6teO1x2+f/qGVLzV
i9A46axkIMm4Qi+MMHWbjpM1LzozUmL/D6J/sy692ESJ1wHxUUG5nyZuI1gS5BO/r5LNJXWi50q0
biIRS52aVTFCRYQ9dL/lmv8fvskfk0kdNBfebZ9xUpVZZM0f6QViznX091Q+UCs2QKkv+2GxQBxa
ZBja15UUebBRzQwTK3BihSMXtgKc3bQSZ8PuRGNf2wVbp/Lj23fbsG76ppSsRS7orNODbBFwJgQp
tY5X3O4Fnuhikk/7wELVfWwGGucvq2L1tInoLW7tVXyTx9Zqo6CI2ND3houyaUtBJwintQ0wqUxL
nEJS0fEthRxVXFzC6nN/AJE/KTAqBscU8ImoruFCU9rvJmO6IXbEKRAojQlL7J2CL4Suq21jI3C+
ON7ukjnc+L+GADABchKy94hdIC6wZScRR2tGHC3/13U0VJD/eAnosZW0jPfp6o0nBvyLqDn+iRJP
QJ/Rc5zd9oq2GukCUMw67Vlz7nlfM/yBos+njmS4UgLqzf0LFYIVmaZMkP3wltGd+NS5E8GHoUlp
llaS4WIS3+gT4WM0K0QNmfZhZxhhdrhiIpj2gG3h97Acfav16fYJOHWF8RuFq7KcX9zaOXt/hU9G
9wo6OZrJQlYav7JYIaH8i1QteWYND5kZa4g0UzDJT8mkX2mx/Mf+PC3VawV2aYa6vDkgNuh6nbN6
EPc4vkS3B0yQsSeiRbI+tkFuVYsmQuN4Kaq9nqosOtU1EixCFjrCz0SxI9s4Ri83a918YnXrkxSD
ZeUp2YwaaC01r6U8mV6Qx60Rkqpj/MGQ0m8lSJjPH43WPORAAUf77nCbJHDxzuYilmfQp17FHDUD
woIiXREsZ0WI7vISpJzLef+gpIo/OM7t1w7qBcyL0b8eTSwbVLMt6Nt4yUkAGkrnMldsvTd2O497
FxR0Vo8RlK4IeEJL+s2Ht4eqr7E8ZnddeLGv1j/34lhqSykO8XdNun+v9E7v9eIRR0R60FY4tAMJ
a56/sT/k/r8wHQE1oV2ZplQ5VBiWkabOWwIUcyx7Cl4wg1Hx5popNJKxQ+IMLHLyh4PyK3aVfIpf
jWoIUNsLs7G1ntukLy+kKm8w3Btsf6+zDuXz1XpxRfFSeMiF27MfAuStkWIKm5lcx0SzTCFGtBjg
xrLquHlLkFfhWAYtXaU4CioEOqpnhJsfq3YfbOvjvTBSFiNjX8yVvqJp9IpqxXkxv4iCY5dgTHaH
wgQaGnw7LpsRY8FQQRr/0BuRxI7yoOSEBW1QTBUvT1bno3GToKOUHpCBqzA7QoNq5mXZKzo5Bt4R
Om/w8DNXhlY5LJ4kmOuYmOuKnSJqvDoU53ogZCw86jMQy2+rCD7LHJl2POP3EBE1eY/K++siX+Vb
RbTXmAFPgMcH3caGxFoSINBpyIH/ehcdgTUgDoJAe47sh90NhxtPf1LaMtYolespZd2bR6VcJ0DY
NUSnnQHttrqTfJpS9SsIW1MToS8cIJM/zGZaxfHDpf/j0She22n7WkqfzXHnh6XOh6xnKjEx0nX5
5f8SJ8oS8+pJArXEFB0zAt1YvOYC0uhloNSo+tfqnVt2IhSea9xwqPX14yv5+c6ky8W2kC2rHEmj
CJUHLkqSH6n1HBkZ4aQ4HHSQ6cLpBmlaDYk6qYaGAfpq5WneFC7i5BK8BDVXDAXGNGK2liblVv6Y
kXb4Am/44AXQEwgArbZfMSx2KWiH3YHz9LLSvuUgjtoTP8eu8iyG/lwDBKRtah1z6G3NLA/XJDQz
SiSNKmTfNMHuX7QQONo57j4eXGecjEvZ1Z1XSDL9uChis4A7V3a/B02KYsvEOTZ4UAj7p2qz+W4H
w3ea9OKhcUHRe9XQJZQ10TkulY0ndy5as8HRbh1VCo4WiyZjraycZ1z/RLCQLvQyBOviVFaWGuQJ
sAV9bq6ZEIihGBaSC47mrBER+6VID+K3xLoW5AexLcGDtr3rym/viCp5gZRyRUKRuAD1KAR3+kLu
ZLGHY6XM7qVSySjuBM1qNJfsL46g2qK/8b4RlpIHRh9duZS/ZQTv9RclpfiqVn4/zWzmZz+pGHH8
3CprEe+ySrCZyNbSja01pO5gEAg2xothJCrOq1463uVa9fKZBJnW9ssdZoutNonQckXmqjbu6QwZ
xD63cEWDW2FyAkxRtwiAVi3aDktudSMXdSvTvdS2kwnYxCwuaoZ4BZhwCJCNnnunUPpYXWB/DrSb
6iCflk/qT0M+Q96Gm83lr/+PKjvpslFErAArkNU34tYhlyvum/jnjQsWKSwRhofbZtpnuOEhU6XV
OXwEDr7ZoYhlBU1nbxaTWxZx4jlqOKYqze8Ttsc1SBhHvhkFGQvLfKeFanyQU5PGCIwNmSf/1cPm
an9F/5JauZcZxIyK6aXDnXn4Y9DChFmrSso1oc63uOpyUvsX0v9ImU2mr65PgRTjspy5OKMfV+bi
AaebXD3043yPuMGh2IBMCFhXdy6YF1TDLJ7mMCdgKcYdiWLeU7RsqN8rQp9Mi6JufUZ9wfuLyz8L
gDA0SN31gwPMrvp8QPttI5ay6llp1yUcn/buw3AzO36Ax+36Ww26gjwA9JZokRKoylvVNcNc5Sya
AGW31MSiavMF9DRdTAUWUF3Apfl6NIjpbPO3fkHLr2F+wy1aMFdU7pbGLt2uXkjp/GQPkGzV8+EP
ZeeJ7filFSAra5BkKFUGInsjOlRgwRRcRydwb0kRibFQIKy1nM29whUSFHq4trZUtfzYtHlJkIPA
0E7bPDaJKCiZF6lxr9RAnYjKZNwLSlKJToKfValIXTfnXhh/21GoKs7AtrY26Z0An/PJPfGrm+uL
KxTeSHR1yD4s15tIVhbDsl3BpleuydyTI1zD6+EYIMkzQ+JIbkZqRxKbHzBO3nMw0qc/DxAxTfKC
Oo0w6B7ZpAuCs8UvoMUDqdETsVmAc4o/gXUvx6kR5giilPMwpXikngF2hTAxPxy92WHwk+saIuf1
6bW/3TEv+74YeHIsMsqR5x4o7wXUlj4xsMwuIX5dVWC6ZYDiHi+ALW4eN0jbcWuO131BnTc/GP5u
eIUb0MRuAnF9eoqjC0ZOkH6bHVdieQld6LyEbCIqsKKkiLLP956MASA4A9ud634htB8uHtscP27J
/HYodY4LTU01zQmER5EDsOCGRBOwC/dvh5AzN1KUTnfYEzEXheOdxwlnolGpBFqNfQJWtx7SwmHT
CeqPYhy+kOoAcJz8GLu37KwndjBocVC4Q+4bX2/9wZp0WYJkZqjjhG+HyJKTSBk+sKMsA0wKqXG0
bwxZokHpTpkxA/OJH0RAQTYP4vxiuQIN5V4d08ulHjzir7xySglDrF3q94LSsQSSqZqcNfvuQPaD
WtPFGX24HeUhey+CgihrQJoZykPNCrvcLAgkOwrMaaX+DnfpEivLfRGMfAg/OFSUdp/2kH6y87x3
xq3lahLq6ZOvMYjJ3IsghFVVZ4MmtMcH3gqGqUDckSOGndqH10EavRwILvgM+v41Vqt1Bnlw2zgI
EhzwPRwpQflWMfPavrO7wzv5r7CLGfmmTeeoB6SP3nuBnBsGG+MDIOK55AjFj6bJqPjJ3n0Ju3Od
KteAQLk5fQPAZjMjJiWSRIVE1CTbxoWfMMHhkGK/adm466VpLkVdpmZgju1be3vZ/mA/e9xqwnVM
RwDqHWp8zP7koczSDvDNCekCQRMfftKBXGHCgQEkqTXozgfoAd5bBh6I3dAOxmWxT4QMNrtSMEOV
73O3pRpR62nBiJNBgfbxE9iIQtoczxrk9uVS7dc51swvsQiDEKE/QOUle3jWJDo35Wp6+BM3DB/F
S2SysFZNQVDqK4BFDmzMGt4n6jCKmnIzZihSB2WE2iF4UvZUrjAn5jqiHD48t901zI8m6l68MdAh
9rb23v1Dzp8b0f5UpL6IBG0uDuAdmYXRinYl9/tFuD8KhKLbXlSS5DAf6wiaXbdc1vB1MKgWpnNB
p9cU6sNnDIa6wesGnfYhtZU/h4XW/cGBbc9CGedJI/oADoQPv33lfVniJTYlknDEjQR/t+8nWH/y
v3mXhiBGw/7uI6kTmUhFmJ49UVxv2YzAaPE0KoiObgVxoX6UtmhJ4qfg8sOWhOyQDeYw4cEhjs0K
W9aVDg0PyJNZan7Uf/NXzkV6Fv2gQBZ3Her6ShYGI+o5NPGbvZd6oRCzkkXYyeCuNS0qp6BXCSUu
f8v4nH4ruSDzgV583f7Ly/jMsdlFVHpqbEZXrsw7shLLGgw/2H9h3ACWHZfFQVPGAfWywZmTAgct
W81tMx+UHesqcaM3c1gNJtkA/XUGl+po9muR5bimihRdTcrlKQm0bLjt/b+jPThiT6COlwbGi4IV
tnLJPNhdLKy0A0NqTeQpmnSMmOe42W8SbhdfMnxkGzdFddYJF4PHkL0lc4uH4Vc+7G1Bm+FiaeUz
nhHmJAuDTBO2I48XVec2h4ReYxa1MeSpn9H9HTL88O8T9HB8pgJTrr8cCEvweYGxR3oAU5PrMXjH
7PDCik8Y57Si+CKjp18wkl5994Z6ctIf17W4lKl+PHRCQYG34tulPhnSLzWrO4sHPFkJ+Mvn/Dc9
gkYnwTOn63qoAbi24A3BOH950DlEFAOA6UP61358mp6SYQEh9fJ7M8VSlXsamgRUatwiq+SfOEcx
U4T7v4MttK1xkNTPcssIAJVRfKbuY5Hj+DtkNBCj0tE8qCcozNbZtu5l4Pfy8Wau/4SMak/t43CM
KoA1iV+V19gxWAb0g2/yzviR5fOONNW1K0yx/zNOPymhcNCjQETMVT0IE2oDAznoceYTXvSnQ4UV
6UO+MCVVHh1V+JlG0Xo5XFK/u+jcZKysc3M61Y3h4cKNUGjsuh1iA/R7H0G2B498VSFd0sRONg0C
oAZ0UH7ctWz6Ra1eUb1c+dJGOD8ht4kDcXUWLTm4VpPmqTqGTTU2FLoXzCOlZuWKIiw1JahrQfj/
i7ywi2i7DQ0hoX8x/e8iZT/oVkYkoDdTF6lf0+NmsIUm3CDLu4IY+JF7soEfAmdgO0LtWYwqox3D
xrwlqEECQkkHqNG1jG2K3Y9jFWZJ3B5E6BXbvPc3QM5ow0yv6E74Wzj3b7xtPbre2B7+h3p/CCP9
rw7b26nQx5A8ERKYFyCUyHqrKMCjqPcsFWxQdaDHpnKRTVHNxQpLdrIWSiLmv+KtE5FFperWY9zo
1io/c2kmkU4uer/j3yjVYM6rVA3ffRS1gUOMEI4DUpwQ/m3pwQ1xxxI7HUBFpUzllh9dhMw9dY2q
FJupuMqs2wqVD3nFHgZd9lpaNeRZF+E46EKVZkY2uj+KnvSj77KULxUTHN1O6fq0e+Zh22evLuNx
fpmoGjtiAd55nOFm9iUN6oVS+JfxzN6RRQDtJkItxZrZS3eSuQLMMGl8Wx+i50cBBNuE5nI2jorD
5voVlW0r1S8QLKIsNT0d7pNLaAbveMxLFPOghBC/E642tN7/AbTkNr9v2gLFmv3U+cWabhRrTyea
7E35Ts4qldcKpOLh7IDnBEL6gmjPTGVGSp6xU7HGoYiqvxOb6P4jBvoiVQKmukKlYsHw+6qBTz15
jZXTHww2e6K5rHcsOJZwJK0RlHrBBGs+fksaLXQcyb7uBB1C7g++in7y745u1gsqTRNtq/raeZKb
xqdxkijVKvW3kQjNRRiN75+mXRDzM/g75FMBj4og0EqiIR5jAUyMhEggKblS/Z5+3Hc/BzGBGS64
PD+O9Z9VPFFV/q9/J6xnhPXCU0LLTs9uJzSiBgoPrxAkmaQFnlKU31H/aDSvTza8xAcaP/E73xSX
Ww4rkyt404y77hPYNipAC6TDIHZuvhGTiXMaOL+NDhv52E7v9lBIcRQ2cjDCd7cu3O9K8Xh8bqRN
+G/9E7JzM0D/xG7/CxPMg9G4NVlJEj7v9tdBzkD4jDR8KVb214gwynXgaGUPKaMR58ehNXvdmsUv
8K9iii57gTVKXpgD/6i1G6yZom+VaMGsN108IGzUFmc95+2FpkOtg5DTqWcc1TVRNjSOboaPQY3F
nsWlhorPFpWf9udvQYGoGF7tXPz0OIB4bdHv0vgh8LE0A6pZmlXwl67ihZ+5zG2D8i2pZzIrie1W
ixphTpXbhpx00HcFM0HSQB17ZDjQidVlXt5iGw9bkPEI/ONofIuhM03IoV+Cu0A8+rYCXF0+DCms
yYeaclwzrww2uZ4hrY50eXfMGSg20vwUI4zoG6YUKjHACsdJiD7FhVp5eorP9HbyPfiJqN6DXGoz
siiu/vpHGPj3te3CxLWRjdip+j+Napb7jLt6hvXp8PmgFECD/N+xsy6k3KxbffbGIaN6ZGCdu348
itn14Gu+Z1JWFkLlFqs3sFOW+z6+IgJAAMQY6ajlf4aGgCS4ulPdtkP9utX4IVa4IruoEp2nNnFE
SxX2DZhn08WKjwZHUVqvjkFMXCWIzlrWSsfkA0mOq0ZW2B3w+YEGTbwQrIbVLUCOS7a5dXlGTfGF
rYvufSjfXGAkwwF4Ny0JZrn0C9mhiOEhvlnp2AUTX3ax1Q0plt9ndFzDouqKtsW2OPnUYk1mWg2X
PDXhoS9yvR9jskVL2omQXOfFgtXvVdNvKDC+0bIPnj8O2rxZ0fpT6sjMXg9Ggg3WaEmQlv+C7xSZ
P5cHbjF0unpy1GFea4QWMQblZuvnKBwS21nk4Zj+vTGMU9VrUXDmsPn7QZ3XiecGjNs2f/6iWscW
PtfJWO/kVgO2CtQHEF7ZSWfGMdlIrtLd5zOFo4bpwuRooOm9N5tXPun4qkUagzm7p1liSf81BB7h
aHmeFSLsC766BMQMH8gZVQqKNP5RiL3SFRNwD0RCcm9fjcCHxeU4F+p4aaLJX+IPYLCRDr75Nag+
qOtNBivHzBCyJcwlhYHdfTKCfqT4MMS6SaCXlh9bu6TVCJEg1/nz7hs7wUN7J6rvfTUBaTMWvhTk
Rsq/tWMkgvoP1eUD5g55ZFPikgFcT7L7FW5J7SZzOCNoHr3enj2tzTh8Sooa1yUuLze7kiqCrgLz
W1fjtp5c23lMg3CD3s1WD9RfMeF0hL4ZPp+1b29RVpOe7AN5NZ2H/Q2tbYAAm8fdGoK5TcAyDbyR
oGoubiL70PZYDkHF6XuSQ6vmkTHimqKX8F/QM1/GbTZWuKnD/nSmQdtEWePbFFa0fmtICONrz11u
WLf7s1ghqRqYQY4mv3zHknTvkdEEINdAIM2sP8QtdVTZwPzFSOnADCmb5CWe6D6Q+KMudjI47ngy
VZBeK6jTJI5eZBobER1KHhlimP2DHhvA4v2hSFjaZnS6YJNGEbYnqw3GqkQ+WLChoz8HKCwBRrzq
F21WhKBknfzdpW8vCloXksO9MNu/U7F7w0x+u9t7J9qkOrCD5W8OY7JddoZrD3IDOZvJt2w7iDRw
kWHJEtR3PMpuyexEtir9mdQ/rJXkxsGuvuS9W1yE5ACTiDf3AmWn+WPXV/q+Z0lOuLtqrZMDwJdB
WiQITWMS6aWGv4GTN0LdaOCgSvaTXZZLDkuFFHdI1Go8jnktMPXtphKI6YTYdAEL9wgYjk7V40el
hOavyonxY/j1Cd9JAP90X2ZqCuVIaLzC/tGwJgwRrQCFgAzOC8Clgz00YMoiL+FSgel7nuMFP6p8
Ar5a/PvKjlrsnVSAmRBgn+F2Ma+OqgnO2u4DtN9ss3Y+stJRM+ilNwSClpJf4Yp/HasvqdvBP4pe
z0l2MIMhD3k/Sy8HNR5YoKVjyhZrPUXU7WUDttE1FzYp9cHlCCK8xQwxvslbNp+wdCeTZMs9TH+L
DwnzJzDSKDwhI0NrplO3xgwjARvqWMxrtpU/irUdX/nEpBBtjqpNWBZM2P62hFtFujj13uNwb55I
FOeBsTLgdByUCeJ3kns+cswSiWxCmlbbj/gHPJNErKG43u00YAdXWMAe5CL5UC0xdwD7R7ayhr3D
oGAPYPU4HS1PQOUD+VW/vmvw5VTTVGXGV/eWHRD2zcLu3CpbkkdqHANTosnEqADfCZQVRa0CE9Ix
Q4o2w6hkL1m57dpge/ZD0snqubIAY0J7nPQBWqA10fsDC6PX1XJBGm0cZYenoLNFok2S9OSgnNt1
R3UxQWKls4KR6AOhvN+ofDhyShozrYFTyNUdUu8tXq8RShLb/OnMS2Uvlf0FHFih1M9C45GtZusM
ZD+ltweG7AUhCP854r1Be6yARuBc9+KvaqU1TRiQ/ktHLfu07OydCy11TahzXDyIybIUyiI7GHfm
CWPnWD1SWZ+bK0XwJucZGsXuAwq31Goz52OKpoOeK/fipEYqKPzf2aU0d3MxDzC1JgtMg0mrZnOZ
PwJSQOEdKgRyZTRECnMPM4mYOHrFj/JepC9gUkm8PlABJieiLoBK41O3knJUTMFqnXpvn4Q5V/pN
1PRK045jaj4OXJSAvjk5k6eMZpvoYH+n/GYG3SQZd08KLelvGKlVxo5iDm9NxXFy2BNPt8ob9NAw
g6pp3saMuMC1m3O+PjiCKj3enLGs5qTq51sWb9ZuDsqHjuneJorNKabwAdzDfkLUCuFSstU1EeVW
PZLRjCdIj3La5Mlla8OqHl9KiEa3rBDjRAx5swB6eb8mINuK9rtT/8WVFCxLxK3kD/8GTVTpf8T+
cipTrotxUdngmSfTsNsuSBe+AaC5FALnn3FsINY0RSTkrX0HS2wjg7o02kgqNrEfSZGOTQhr7w2n
NVpoMaiK5iWcSufv5h0SOhksCUWSODYKktMryWX0124x9RI5F7g5iWO0l/xwjCd3Me0RLcB0KvQK
vHbW0T2yv49adtbj0FYerVwdIKgR7fsZZqdlKllDaxnDZzJy1wZUbr6aI5sqINTlAFOdzZSSH+F3
0ex/sDoAJhoESeIknCVWl6YVNaeiZbwHX40K7WRHKXGOlSrnErRYC+vJTaiqbgATLSYz9eR1Tu2V
rl7n77TkqibDvYB9MoMeImo92b10tXUSom4mCdk/mBhvb5AcqmuMaSJAcISRgfdec+Zot4uKA78y
0KNqbNnm3erV+Z29n7vmIYLTvqyihLqw7mn8CRb+Czn1/14CXbvHVLCbj9OMMUWeef3S4NDC7/E7
Krm8Tx/2kdzz8h1xqnq+ce0Em3Y2qeVTrgwnL2VLN+udIWBDzhSMImeXcLFeqKlm7umyyww5Ofwg
aAI66SNT1/InHsZGfoMVCQVp9+kGlaZ5FpaMgM8X7qXSo1tK8LXoQ1IOXm+XYUb0g4QZRmymayWc
uR7JQEPFoWFaZZcTY3K9goP3OShtalULN/ZcZ7U9FKLSLg2WfNNnjv9loP9+1GmtE720gRTWCDPC
f/IPmyUSDt7128Fllrm92JHb84Po5Np8SItzG3pq3fAOV/jRLMnR6wYmdo25Ua5YCaNxGLSBYx0m
A3FLyyZnWvaJOy2PF5AMr1m754dY948fxXSQuetUykNljDaUl/5mb9NvtlyAYZsmn53INzT13roD
8UtVH6mOXxSADWQ/qV3/rlKAEQI6U7LpeihT07XrJu0E8aa0f+lg4es9k89UrF9GqAhCIcWc4dIW
F/dVEWWPaCGzgYZw8K7P4SUDvrq5rcPwMXZaplO8/IrpigildSxVBzq3/IwvUNaWU/UFRb2B832G
2Wb1UFgp6OHYx8N7v7fTLlt/s8ZFYMaDOqtXGpCZk52spS7ZaPFEaEQbSTUJsk+P55E6912lIMQt
OJxU0sl4RHglY27ZySFu+R4F8Fh1/oKu3HnGr3NB3CzB6xUez/9eRWBp0crOLIIQuJyXIlRyye6s
6culVD9L/wfjR/BbCnATqmAyirWdTKWCZk+hjT9Rk/o5UCC0JAPy1mm9a9aveMQdhB0PdWhBihsi
o/vDfbxuu87n71K/0nwj7XezO9y3kp2whBpjesZlcJnsZVkLiJQzIHriBGxMZViRycsDEEZt6anl
cRbVhkbEiQ1LWy0odpX/9ayNEbkoQuC6eZIynyReIp80wRtNK4A6GnRDDZ6U/B+897riOF607Hd2
WOjI+x/lY0VFm+zV7UqdJOLAZvA9NnDJ+ZVJWDfDi6R5xJ4DYSWYn8Bo16QgSLbfmNZOQA6aYrtf
rf4fOU6WXfVn+RyUWXarrhVO5xnRD07CFsx+N4eAEPC+sAqziSRvRIn5Hk1CHFi1PNhdepz8SAL7
X1SpdYdTjVHCklGxNpL+pQh2x8rS/11B4RPWkL/nDCCjKjl9idaZI6pnCaQP/QbcdlLP2XVTLbPR
TtB0gSkOpKP0oclyPM3KE1rL7GcxCd4tKEweyLMQQ2JNZOzKG64fsF1B/SB5YtgAkw/YPZOX+Fio
l0JK7cTqSFgFwIW1JmJIEmOx3aNkI4bguD77Z4jz2ZhZk9jXSViFLMYirX3fMm+Q7whUAEHF4vJh
27W820Xru98bUIOg1l/iOh+iS6KQsOF8hgtDjG+fHovedU/WdZhFZmSDZhvmpGni8O5E/O4Aq/6C
8G+iQD0uCnmjbUZkI9HWQNp3yMLvxKxivY/VccuHgI7fPt1S1pHRpj0Z9kYIjx2JuSrdGHqK7oos
McE04gM79SqjeyF/59ApN/VveyiivnvCdmuxcHoXdBrKGlvrmXOWFt1KgrJnbbt/RDacvx4aCor1
nTz1v0B+1gnbDl5GSRgWL7zNiFpkcg5JUtpaqLPYCMmOugM1iGmooMcwv4nN+2KRZ+BrvsYYeG/r
0ZUCl8wSbqhww9c80Vz83V3k6937+IcmokoL8ny9/LWSNyWCPAwGSPS2IDH64zlV4vq6gQhjL3Uf
7qQ9Iz7xBsI4j2iQqp9f7S8ZQJHR8DSOwWq9QKGLOFCIhbdeQPM0KnX3nsNoKSvOS4kI0rbbgMZz
iBjjvXDeUqCBVyvnN3wgXwpX6unqz5KqKNV/C37Ssj+8MeOuqyOb1CBa3jrZ5s8U4Vuv9rE+bbur
JncmNIFDD4gvA617pMJmJ8pvf8muuGf4Xsc1x/mFDiPpDvasC7V4iO4uh1XFLlnZmMDavv06D8NR
IL9F3020dToqun57vWj7J1ebwtzR3hAu9A6M2NLIIRlvtSpBu272fWYQKX7KmZton5SRSPmnynF7
e6fmmO1nqxqNfIb/5XXzHkU6j3aTsRliOylhLrji9AsfRsA/ZHfYCOd4xo8gW7yIQQATkJj/YUF5
CzQV5WJwSe2NT2z2vJF6MTnTC7RiutYKvTvxnC/NUmUuxPMKlb0zQooM+iGlVb9CvinBvUJPwp0s
T4zRAUxwxyVZefqtq2HcSvrhC/UV+jfj2oSBwwt/4dppSzaJi9S1x3Uhu64zuNRSRN+5AzzzSiX4
C4Vt4jIemejFk8PYV/AyicisGLjTrkS3dVAZB/xM8UCF5lgENTy1pubsH+e+h0o1s4F7U1+r78dn
YoxgiCETUsYx9Xb0uSow26xyj2AwZC+OUgh6v+hDZsi8NPvpsPvicl68JQANHTESNfjFPRTjbJgP
ot/+DU2TnVOl2KngCZ+OY/77QAwR2E4WxcNs5zYik8E/wITQTRjkVNH02o46ZDiGSuu2qoisPn+C
du3l3z+QQvfR9LJ9qqBaw0JIIlTuomG5Fb2xQ1Y91XbgdYu8XQrzhadXM31vAcDxLqc6sK0MRv6i
TPq5g0k3dl+51tkzrWgCuulBRNsUdC7wtY+lohW9soyYNfJYWmGUZ9o7JNu31hkEj5krn7rLgWaE
LbJsVB89EtI/RGdl6Djzlm/GJleAEyZ9Fuvm6CPqkPn6rIzXmDYfoG0Y2FFeU30C6J4MaZXkSbhB
PlcmZljuBgVnB2Rm061cfElNTYKxrjE75U5ye+hBbr/Q7/rLEssgat0zx+SOxgVDykwem65QmrOw
P1/e8QgjE+q1hso4U9hcmQXh4enjDnMfvn8hgltlJwK5n72cWWnUlBcP1anmyRAnSG9byZU+xd0i
RQZPO83oo0C5LJJELi5wqCo+PQLeWj+Ojn0U2vsYl2bJwAz76JXbRVqVI/EivgwKuipHmih+UscT
UUGHVv4gW4uja7Yc2qjj4bF73dBJa/XtBWbQDCQ1zNazFVVkbRuQr4eXNDwrnu2v8NvuDO6AwGqB
xHOf3B9PAhloXuzR3FMV061WFiGM/wqyhAPwTSnxNixKRqQRCg238aE7OozkdPB5ICYac+Am9mLU
v1qt7UFvs6k4XoIJcbqzALPTqYW8UF6J6MtHit1WYhkgKgZ9SjLROPgujqbpVNnjrlU0/s63zWEY
cBQq3Y8UXQ7VRFLH3MKSlAKLIfAAfMaUOR4CmM9p7W/Nh/hM4j4NVpIZP5KN1Ac3ouyPqRrNKi70
prXzekrq7s8Pc1etStUh3geLSguDYF5bbkhZ7PA/HkV7UA2EdIeOyH2iWlqGcoX11O7K4Ci31yNQ
G7jT4zkhh0tvM09YWelkKv7BDyuzPDwurp4+Q/ed7OGHtiHPdJQMlSQN2Ht+Ps5nsDtBTu3YhqZs
BgkCmfX04QWt+JOPgD4dlWC5eHIcGmT+3Qiz+4r+FUVMj1L6qQvUEnJblJzGWLY8FoHNLA47Qjdx
m2YXPQ3mkvy3AZCWzQZtDqWK7vfJMyrC5WrSQkfcN6WbShjl09iCDBvqxszEKeIGG9FtpT3u2zB3
u8FCYU2qlnJwgf20l1rgwjryJXM6h78XPOb/YavXYUCQyeyMwjk98pryBpep0iAx429Xt478AsPJ
9zSTA282cJkIl/h+lcpgWA31j+ENKN3dLMrw9day7UkqLdtKoBDwEhuH9uTI4F7C+N+nS5EB7uuC
iHhitCW5k0Sceg3mLrusLlLSt0XupXpBOM/ssvc3kTnP1Z9Hn5k3c99F6lVjlmCOn286BGHCjiiE
V5WHZT6NeBvCAc05+i9R1cdG5f4R3xYH54av0ZBzjAV+K+WtsoRM6KChVKUx1M4JhLj7WVI76PZA
WhedR0DtcxE8WyWbA93kFuuSMUmA4uEgVbrg3FcwiP1L9VK0TwqTI5RuCTJhfGkV6LyCS4HRsojU
znHnTx+zsN9dbvQSPhf7IGJPhN52JbsXZVT3Xwf+gMwU1b7J9rczWxUNT5tXsRVlZbsnz15tOqMH
rUsMVawtAz2ub+fsS/liy60joBT/AFuNdidMR5LUhfhOlhK7rSTzWzAZuWV6m6GpHLHiUJCoryne
FJS2gxapl1gmcus1PKGGMHmPsCbixknSSATtQGxEe3aeYqh6Vosrn0fhfBTHipcfSjOPy1XTZf9f
P6mmaWcvK33IiK/0ZvXoDfPN+mbSU2OB6lVAyVISEhQ0f3BvEU0+ZYoeZo7q5mBj85vq5XdO5LMj
lkp7SJ2+VZh35y7iFg53wT2Gix7vabd1BEvj8B9aNqwAsYB+8/gmDvGbywJf+TlD1euUFIvbKX7J
dx/R6nM5+uhC50BC4lcQgzSDyFzHAocwjR8KRKV1EQ+tkrlTo3kLrPX7FsMb1X7ktFTm7dPLx47h
quWNLz9Mx2caJUieo1EuRYl2JkqoZwTIWRCc2QrV1P4KCWzLQaR7ssMMAt/muTFrpOlMBBxiptBj
pfb3yx/jS1H7FlF3ayEBFqnS142UOBQgFcuNBDzys+v+eKkT638PT4oAfw+Cb9nQ0vzQUmWKfPTB
ltf8XIy5QRcaGYLH5fXE33wPsSMkpMdWPgMYjJ1nNoQdyvWc7SIVRKnTNJJcM3CJuOMXBkQFlz3I
9Ob8RunTHfawe/q+AsThujgyWWqG7CbQ0G4VRuzdRGpImxTmRwz2oPzxxpR1FOzegNQ3IBu0Yc6F
3jXFrgEB98L2Lze8wI7Sj8WLtMyc/4Z1ovNB2qWUSssA6o2eRG63LepLOs1qJjJgXxKxnTitofXU
Ko/DvYy9PIogyFpX7BBpgIyZdBqrnB1yNdCkMcS6mdOlMu1+Cr65dtLQaZPhZqBHb+BcVRtZnNxj
MzNKNoWXEDB5bCzUpbvDmuI88HrfaMcID+nCCCa9w12mHovnv6c0V5YDwlcCiuKejhD4b7h4ofpc
ICP6GBg6dNtEAmKbm4apJF3O7cvLPm8IfCSsamCD/AvoAug1o+akDh16+LBRuJTSPGk7N9ZrX6Sz
vGiYeLA2w60tjqrpFfH/n/eqwuXy1EF07LpHbycexGM7iwqeAYKNczZSDS6c3Sk9A+FJPAzLAfqF
SFIvkfNYca4QIdSX1EPR1/p6U+e+//E54kMYZabDGY/VvvTynNgH3CDqnCGF9tnrD2oU1Imdgc3D
/CaCw7rNVbMekgW17mv31WY06mmAwzUaQU6QPn9MsxWC2YW6sDuHAwDzaD/hGgo2D2vNKLBqBawF
DOKb3dUGKniEiWVIzpF5NAINiKqguWJ8+yRBPj4s4ezXlYJ1Newg6/TcUgro0fMtSathcxn9w/gy
VyWcsNci7/e+G18mN9oU3bKFCVj95unSdPUepDmcXJQIW72NeaD8HMQSkqZpOeNvnm8QJ9D2urgZ
JZxeh8qQ8PbfqtM9YwCA+n3vmRucAXXEJfc9le83ow03atFJeErjeVyLe2mM37khNUwPjMfbjnSu
1jctZPnKM6HZQYkKpdHlfVm96mHTdtHUB59yULrPM8eyiYAr9KTLKsKOt99/lYpIUMvw3/8IqUvM
vEHs01pRk3vmul2A/voYlBFKsQmFPK+81f91or9ZxBMava5C+G6UScusNB3QSEC0/V8qfH4bE8um
KAIlEi4EA4pwy8mm0Z/0E2mJ6qaJ3wXva/fQSKvGFO/GKkB8EuQr9AVagAU0Kly4WEkA+ZzVtpwp
qTdi2btmbwhggNu/rEFxcxoh07r2dASKYHdTbIoAGWdy7rthLC8ndVb8Fn3iBxamASw2ok8aCWkk
Vzi7TzO2SZlcB/p/60jmquJgPtYZ4r5TR2Vj/z8a7eCxqhOWZfzWC0tL0MDiGfV/c+SodTfDMh0J
fLITYR+c3lBRe65HPGjEQ5g9UH/1qbLpEOdk9FTlhDcUjgZOPg2vPjZhx021OEemiSEJjIqUj0Sw
qViRMOUTwEcGPHVKxt84L2WxRVr62K62H9WeKYyT8erCd1qmzIrmrADyPRh8//MtoeCYwOKXhWXQ
jZ1hfhlxbBucwnrgP9pQ+xUzRMC/W1gOFRfYHE6B33uSJEeFJlSUb4U/48WwgErnOwDEjD06Tk+n
qP/6VjZOQscbXbP+NZM3/1dgNphcXIHWSxuvqEY35ZJaRgP/Q1wN6ae9w15nhIHnKIhqrEH0jgQl
//Rc2vEp+jvNn9WQnS0kQDI73LzReev4HltPuJ76iva+01QINLNfuzTCFni9AfAAPOqqPlmtzG7v
Oach4Jd5+I7EA+abKLzhtdAqMMKtWvktgyOyR1G3SYxitMc2PT4bCyvWd3fhLVW2LuTayrrJiTlO
LrOM+l3yRa5RxBE9E0zDcx4YIhNtA8flP2ougBdGuzzB37pHIiTsPhWQ+ozIpQ6OdzdWRQmy+9UB
UnPpRVtHRewiObIrjllmD4fmr8cacHZDM4ofS8h8qtjf6dE72WS8VmzHKxBzZET2BmqaRjUTKmsQ
0omwJPQKpEgFmd1v+/SnSwlV6Og2a0H3it9+vUbm8NMCA3pHT0rg/XyKbjMLQ89LzhpGcizh7r+S
mbCY/wvCevfVcscdGP+i4LEPpd+I1FeSXP43Mg9bBjUULL3DZD+V8xkup+LlIsJ2MEuDVjQxHQv3
VJcyWyY+cfpzzgdWNCDAVThqf8DpWCbePaB+SpHBhOpC/u97CKMibeoLXEo9zGZO+BkWOh2kFVGP
TCZRXtfVMKnfNfz1pxZmR4hGnVowq1+USD7SmFAjYURqBW4OqwSnevR4DV4pwjLGCYLeyS8w1tOD
qtyyo14OkOiuJ/4qREYvAUFHEnRMy0uGYVOnt6az/eQhztpoIlUa5CdlnvroOCHC2mCbmSaHpYaU
t0CTQDWmrorQBlK6ONwvxKw7QUtsfrTR+4i4t5mnHDsp4NIiRbgf4UkeiQs/bDEbZLXkXdee3qvg
0YZEAIral3fNzrLi1hRbHFiYLssfWf6phJgOkUJ4ZkyCXv9uYArQuPRubwe9amfyN/HzCfqlxdB9
dXQv8V0kdACeDltn4Vki4U4vRDyb3gYAG6wpSBVv+rB4fqUWdaTE7cMCjwTncX3PwtJrUIUJl6K8
v8uSEVRzuHeCNosrrfkj6fBjFwSbZTTTxZIfStemF5xPfRm5hkeDFNLVUAwd/+/L3GsM+d8AV5iM
/lbN2zPO+r2uMzq+vUU60jcz63s8rmKDQPfJlAL2/6dahE/zfjPz9jFK0egDwaKsvTKfdAqXIvgX
Yxo9Zsf13gg3zfuQCpCqmCPdQuKy1ZMzF0SLRZTNJ20xrWxaRtRZWrx6Mjkt86Yhq4djMmOl5owv
jeOKNjxS07pa1I+groeahVetOobnt1k+M30gjjWAdUkd4MDyqU8mc7TBUQx13h95JOi2O389r4Fk
IgCLIHvDg3njQSultckWLSk7Kf6687dRu1PF5+UFCLhDnZnVFiONW2wcIOlPqlrULZO4RhhHPZOK
nBSEhAL5fta5Qs7G2Wp9lp9nTjWyukvMY0rWvXp3M+KmhyP3IQ7lAA2ADCdsapNeVOGNUaXlcI2t
XL47K0/LFH42hUaubimpmNNQUie0rdrRysgaFTG1U8hl1R41fSaIhBFzVC4yKgwcZwNfecFFLfYR
A95jWvnPG8QWm4UPym7/cr6CdoaxGLyuzuEw7oGyip1LPBiaZSr18bFV9XuEWXNK89c+cc0poDd4
6vwEqW9nx82gQJWe0yfLFe1PeUAcj3Gv+HcPwfYrZcJ9l0PewYqEVfiwBqYVIyPlIaa95B5441yr
ZNvaW7Km4gj2Qura5gmK8zd4lnNWGGZW8YQEJBgrE/RI1MowO5OOxJXV9Jue6EgPnrofUZ1ZalPh
S/QhwdEYRggUSbWrmpBgEAlW/Av+bYPuCIlDxp9W8UHkw6URo6KHKr9bgFf56KQQITHwGAlwrdjz
qJCJ5VK2Zj+NbJw0VLGd4BwrqQ73ysqSqJhS6VfP6JFT+qRIFb0WgMM5cTJ06DtAbPuijd3zXS39
q0QsY9QX4SzjXrVuocb8okZEAlJwOxvemPJbJ2maIPgi1T0OhFR2Uhed5CJejyWVAfKTb7gndkb2
NJ+iUKpfvoZacWwIoPUC34PY4VeW6Dbl7/uIv70ZYaSFAldYy2lYrdWYwSuFOz31CnJoyQCtClsd
AYThUO8dnlfJ6iP1gOXLIBPQDhIld4I7liBlXVMAeKAe8ehk6jowdfrHReGZXAcmqNdm+578PTXb
IxItsaIVVsGuKnea4poSt2Grkpzb30gk/INgmkgst5sZhq15wqBk5Yfjxw0mWhzYFuObixM57PbE
NG4sYxdc+TeortKTD6dpAR9DQsvL7BFq80TBwCEkdRpkay4qvh4TuQixleRR+NVBfcHdby7PkAT3
VGvWYtUx0TJj+6fgkSHsqacY7vNCMnYTHiP9z8D2N/H487MV5M4E+15VZXIcIwuKsztOonH2qprQ
0qK1lX/0Hn8LWBCf4jcBZGmwnx6ygQ7zZ9WaCbyDFe6YdliJXzXJ/nFpAD+TGhRWeJmjTI5RB+6X
w0i3QryJy3h5GCshNrq65g0XYIZXA4GBjpj9XwcbwwAJeULVueS/702D5295g1h9D4vsTlH5pEOe
2oSI+b9GZ7EQB30xMWI6/bO7fcBiTtrgbisezdI9Z+ZbCHiU2KtYA0SPtrv8afJanwxsAhpk9x1T
t/GARRDdFQAy0aj/7opjg1kn6ghtMkh5Neml8hMU3Jt1+uqWMa+jCY+YRUF+h5WJ0pL4qm70lmCD
iFtwuh5qgfw20L3HY9ccviOgT2oZWp9llJni2TcyhCu0hz4N+tCczugizZrV93Z3AgoheWcFYyfz
TpGLWSrn3UVGP+lJRcMVW8fgehcqHX+XzhsMHeYqQ04Nbyev8foMlsHN3HBuAqpwL6lNXybBSg5/
yL2AlAgNiSZHIPJ38wDhSlNFZPsbVIQAbaUnd2i9xb8XUCFrh2DSxB30iKAj3bHPZK9bSn4OHLcN
5fpMQXp2QDHnnb+bGR5PzBMngc7PimmfvZtVwGd7OXl3lhXIDTtVhq+UXFugfWH12jee2aTIX1Md
45ZdTBEi8HiV4ZRxH922WubApbRjwsZCbpDpaBbfcOibJUWe19BQMaZbySS10XYhfvHxzOOKmhol
bfuAHlB00V/cV7Svz2vwqqwdNin/d2xm2fsVwKdkPbpH8BO07K8nuHYEiXC3vglMmSBF7254Kcmu
dRu63neKtXAT+Sq8YsBQPro2aWy5BZ6sMGfNJrfZlTJF1nsLTD8XGh5lj3qcxRDWw1m+u4j/waFz
7Mmvq6yo1ERrR5zOYDtXgOCvBAxqK+eULbCwm38Y2n7XJwQn0X80U4QhdS5eF9ot5GTNUjtxasTx
k/UqVlvYrJJ/peqDMOg/BztL2Tekwq+gBktLLMNSBXgaQcYjxSot7IwmTRaf1BlWlrvanBWKtlkr
A3YnSWBXMMj1oBdQyucSPTZFFalm+Y+b05GNEx3pa72hxuuAeSNU0LM6oMx9H8pCRRX0XrlLh+Da
UX7x+7R15ACZuOv//YIw5C2rsgORqeaDr85EGjseDat/IR1Munta6Z2moVo+LNMxrsK95/ZmUaBd
E9EkukE1zXGVcChf7aS6haCUu1g/NmX6mbHaWtvgQcHHt6eSy2XTlBvyen12TVoxqIDvm47Suq5e
WOPiP1X7hI17/qAjHy68T9UZpHTi+IvG7Pfb6RgG3ZlITKn4NQ78DB4TBKHsGM6zGdI7RyhyOaE2
ltjZDS08VHAUiU7Flzb0QX4yJ0VJ432DdnQ8A6DisHorrDtTuvLEHitkOwS/FAu1EWTxk5iJzjnM
fX+iUBdebBPGHYFoW7/8aGFhM7FIqBFFxRng5Dm+TqHJo9ovVN2VkgbqC4EG1Zlk/ypy0w4f2qvK
MkV+ZWd6fuZQS/vkhdNVWEiaHCtaDLq9QZinJNo/iwgEy09H6ZGWwCXyFY0L4nNOYyu6s6MZbtBU
ke+HBVL35E1BpsIvF6B3WXMnidelexJ1ye5bYoh+kdxTYbY61nhq6U8ypFCObM5DRspDoG/oSQyr
gOoRbk7mNZHiYrM81VVOdOQo5yT4ZxrIcEVW3+terAP2JX1XeyzyKBep5QaKBN2UiT6xyG4SoO5R
XErZG7DnUphZBn7JbHDXtj5IOl3I5QrdXFyi8EuGhMxWkUXE87v5e7NTarNeG9QSAu2uESiy7KF2
cli7cIP66O8llXbMJTydIj1d1ymMJIXPKByQ+cQciYvk62QqI8jp6bdbxhzNLoycwzROgcu6sESA
0qcaVKpyE7x2Z8Tp4dVL9F4bvMUOy6l7ade4jqld2mbt52QBxj2IBIOYa5ScezI6An2McyhINoZ9
GJMfCZPC0rQ3AbyhXLrsD4cN/IbBD2yetQd2oQFp4cI7scoWFfzV+EmtqrXC4CVtOGaI/aSLx4Ub
Zg3o9BUyNR+br/0fx+eU0ntljp3Uy29haIgk+ikP/e2uaB7GlIReZ2fWZ4N1PDIHbjQheJr3OFH6
8PwFo0ySzWqYMTU0CE30WirXkKmQomXpmH4msuwU1eF7Svt3MkbG6GOap/j7hdPWGGVeoQedUP62
mZLGwCCZ6VkQyTdGhcASUqcgELAX/L9LTOpU9rjzAsabvHujnc3MJ0SHht/XlDPOGmDCe47xRi+x
jSu4zjRCABADQJlqawXIiG9P6LBt7kF8WwXUvTokCU+VJWzxNWMd/wTw4JRI1Syvvq4imyIAISgE
B46njKQwqs+Fj4jE0QwqJqTrItkPYk8c/fJEc58ZwvkswhemmzCDcp44zkelqIUgDfIITAOX+jMJ
EfRc1BJn8cZqW45p8O0Y5NVWOBQlXKb/pq4xMBudRHfNYXIQNyCdR+Tkwf3fDHv60B/cxeoxLXM7
WUeTY7s7zOC2nqZJIBqGnzA4MXCzmKTDh9Yzmu7i+Mgk6x+iWLqoRKztC5eM+9joNrwZT6cjmg0s
upSdWkVZyIz1l9Xy49yDXYPDjj23ou8vDV1MbgCpIH3AA4DwdEIw4xWMLhsNeFhgLu8nO8JYM0Hp
bNi0hKyI5wJJTUkLbVCmceneHlbkEzKGH2cqA/yeLpVz13+zWBsA6/IVmia5a629RYYRLJSvRqE5
aw2qUt66+U2rbk/IbeYkXPtFm3+Yc5LYOxv3pqMOJfIv91NEnZU4fH9nG4WjNecqY4L8FVzLQ6wP
cmG5asSVSEtlbaeGFowxJQaBEIMFz9k5wagpuUmNutH+P2ntNxSkotrqtFlFqSBuuRyo0Tz+V/mo
r2PLOfsWybIMIKNhKdcjSRIkTrjLpiWhhrAxl2oqix7p1KVndr75wynqiGL3wVloECOjLKmYFX94
Gm5TrC7m2wDV7W+sXQ+jWXbX2Cj1ZeGs8hYi1hnrDG5QXuj59GunJH3FD/9p0gN+6haXkpCIasmk
P0hxlSRmLx6qk+U70aBPhfSd82OT+BKz6PKsY4xgsKiU8sTPKGmJ+GHnKcV7+DtvwwfcaWTpwR0J
wapMkfHUVp/rnVKEna+5S/QqXqOfqou7374BmDeD/RWCg9oGNLFF/LyVXL/7KigWT5nrDWu/FcP1
0ZkFgDQUROnwIbtImB0ptkWbHDmNpgJhSG8IHOLRW0y90kTKO7fEX6qc8zuRnoCqQrRXca7VF8Sk
2+kNvFQTeSyDs3BoeL/mvw8Q9C8BC48Z6SWbGpNnATwwKuuEnoB5q8UjEtoxCxYFvh4O+niOnSpf
Q7zhMWONKdkvY7m6QpXRrmoPCa+FaIxJabwBIQ8TFG5bZC2NTftS+LAQIP3khxfR+VWYUYO8rZqQ
DCuL03qY1sE4D5P1tdjqsXVVtTRbe+ID8JlMSv/1fUXqdkOkAettQwe0ogBQlSQmzlVXLhMH2Zju
WDkcYFU+y+mVvpylOMraF0oHTAFa3tqh/hLzfeijmJHW1blWa+K9VBXTUU50CK8lP5cdFuuCn930
NtjDUiK2JQsnx1KI2KqFadoMUMz6305G6rdDzu7x3qY722kCFAiDudf+bC2fpE5iT+Xsg0xgnHWg
6RsH9sgkr6fiVQGwAsqTzeDoQWKpXLU/wbP/Ynp9U6d8s5ZL25XY5nQKK0nSt6XtTaBmZdRKyJVM
xuSnP5yP7X0WYiY7x8iXhvEKkKfRr8pYvy8V4hE2Tgha2AS4v14CkrJ1Rs+l1XTQf34e0kQgjVeI
972pQu3H5X1NKtD84NkBx1XQWFDhfVC6/zRmR2G980oBfq1i+Mu5CySLevOwsJ+43ir08L5dobQz
GS6UfScXTDFYlma3BX+ZA6vHKVHi9qbk1ApR5iFVOxKesH2qax6obDHq7RgcZ6ANOkm/RtigitVQ
5FsyvO6KoxB5pLWiXlaV8s0ucJE/Vu1SM4T6W6wg3YNG9k4cjduAgn64Z+5F3KuOZYP5QRhP4T4i
455/qQDOwihVOjrqhGsJW2gIK4gleWEOxzsNhZP4QzIhW3M9DYuAP0ANgDqBSJQQb63V68Azp2B7
PT0aV2NqKGOt5WAvoE8y3tcY4DnAEHLAXjYsHT4xR4Z4GlHfMNQwSmHD7RkaBTNzkLZiTJC23MGv
CURayESScgMb23w+esJYBHEBl3u5f28B68B6XZ0Ax5QefqqVo3mOLy+OtfSbdBC3/PIMKrIDZNYM
ZB3eFWu47zCqAVEiupxMHoohf+qJb0wPke4xB6ISNLC4T6o0hHvVPCe2JuaAv0nMEB8aMT5e2XvS
hZ1lYe5Y8yfCILWm1GfAIpqydUTgB45jA5MPWBRPkALacHG2e1AirXUvVOysmq3CfDMjG0/dfg1u
tlivZPL//egkch+UuN804ZfQjneYIYQoF/aGi3PyrTLmzW/enkAoytrD2h84D9O3rUNKH75fSu1P
33NZhVfR9oXAUgA1twUD5ooU8VpI7jbd6q6wS6gOakxHj+P6zQEdveiCqeHxK7QI5+XMl+bnXw/y
6pk5dJW4GghrytQRU7A6GLR3QRFVKs3SGEpewSk/KCxeSptPmjlkxfzD7wWOGjblQYy7dt2vkGLn
wlP1lkDc4eahplo4CMYX1mWLaFn+pbiw4Ubsz7FQ0eQ5lcM1Od8eqtQVgj7Gb4d2rjaDDXFprZn7
mXhLaGlrVJ1tkdrBRtbwXeXX8J6nmftXDeqC4HzvJaiafqnB9jCA2KTKeISyPlBS0iNGfInELPYx
PBZDML6r1FcU8pbQfnNBAh3TsPZrFBSlbMcSnXXK+Fmh9iANouhNArKRud25+hYxxbB3jgVJ5thd
xGW6gIx+YqyMRt8imqrXj/2meaDZh0imPHcCTraXun4rwrR0VSmI1UWY6a+rStUhD8wxRHDN1sus
n5DcyHdUTOCbZfJDFjIfE3CpNI0o+0/lxaNNzQPPPwJN0QJPatvkDQksVHjQdW25y5KwOvEGDlHm
UflxMHQAMF3akMmiwX1Dr8z6nzq5noztS+rVFJenz4lv5C7BZTqr2jLxgI5v1p7FVsffqqVMmySR
24qDvh846ymB5XlQqByFEiAk2tbmcDtqivOciSe5Ct7WR6HTxKuAxtww+YoCkggXsnQbZSlhArvC
1RZtUs6XdERaKpJ+4PSvY99NIhqsADhwHkwRtEzIWXkNup9kzb4ZXhgOJo2C12OY0p90UrRmqMzZ
r1DnZllrGCBjfjLon1V9lrZ/ydX5H1+N+XDOipFb2BR6EIc/p3+jnMbFHNuMx6yjxCwM69tourbE
IVrsIxyScd73lCXNdcYBNZFdu6603SRFyRUDXBCOjw4X8tG6bJ6LFfOdVxdYjX8v8LNSszOd2/dM
sNRRjk+QWM/GXUn8YuFVqdmQJn5pNcdkWz6EZ5b1yDIis0p+LYLqmM+T783xwX6wtTYnpBnDeEoW
7mEM+IBI1t6zpZ2pCRxod4omGkWPSUjxiTaWDftzGhwUjAqRc2OpEqVDTT/fWFav/ugV475Y2ZmL
uDMdEgGsHVWosLWi7h4GPIpSoYd5DHq3/zVeT1pREgsrDV6jsouIKW66Go0TAh3F7WQCIFCJvkXo
5z/6sSiJLqlxoDi4VsMPxeSEItArqWkGZCxkWiUyS9wyLmacT05FJnWkr0BNBFoPjkTQDH7G3A0f
ZfUkiQIWjla8xew/09kXIi/tnw3j1liwDH9Vam3dkTgJRo2IgAGYlfRq9m49/iugxjiVMvug5wgi
GY83VMjF3i63LMJnbDNsHLkQwTVJ3YOEDhNaTvf5oFOxDtGnJ235Wyzga3jku9e9OYLpYaKl2cTr
/m5mxgHgF3NLYjxA7QVVo2cyjHSMogmkdUACXEzH/0kp4DFFAKZbTcfxqSeG+0mg4h0Zk0kJOfPO
WyjyJCIg/nc/eutaZjU8Z9z6hVjZ1p5ANer1jKRsM1di110g8gWC19rJxtbVijrzT5hCj5B1aGlc
aW26AR3z7e7LGxusZ3Xm6wkmetHKQ4BjJa1VLMf7YdIkQph+bjPVgFhN74BAl6i7n6ru0yAgbfLP
LvM8wZctpWIRmnX8dv7shkWLQuIYwL09XA/4g5T5RQfSjs9sTJ/tyOXAEYtlV3mvr7LOqSyaMpao
UEBdnRyTAFJJNVC3sIW5IWQq3sNNasDko6EG9xW9QooWH6eojSth5f0z7oSSp/ZIAtYkWSUqjKwF
5lppNlUg/PJhxw1JeqJxTA0urGwQl3a+7z2ty6qSiX75ZaZIfcv0mvvd2FXccpFi3p03/umOEUOf
c9syAEIJPOLt4xEmYq5pt+3z0WX0MsHKusPTq7IvP02Nnkf716AHYKnkSEtvIWc4euCbcG4NJpzk
pw//8YDYx1G7Dnf/xBlpeXJeEaxU26elV2t2Hs/Gak5e2sObTnoY9gUa5RVPNwUjyqhha3x/kTXS
3fWnpKySpm5htevbXNI4a4BsdowoU1PHE/4/b2gmaWN8rAlX0eAvpd+fqtSkIyLvySSgZwjLHW9a
s0ChQi1dkrb9/dtRBkykALWKmrFaKy7EVAuROf2bqh+py4X38swS1Xbl7OaKLtIWSuU9ErirStKn
GfXuHTKm6MCfv4Lg627r49Eybo4mzD1awO7kX+0aPQukWI8EVPUjVWgDLmdEpbyF1SOLjEWJqKY6
KhKjrtbw5ovX/WsiE1f5lXO3KVJGolKq71G0scpmdfNA2eVZ0+LbT4dJO8bf8VKUua9EPcGURVNA
+qwX1WCDP8hSdYs7AHtpgYPSk7CEk0Vwv/OK9Wt94gNZKK8bK1Mgzx4i55XNlpVgPsM7WSHKWRe/
c4645r78ekUW4Q6/D1WdOHBrKzmq6boX8P3W1D86GlrFx8KaDzTVwTVxhXj290Rk+5LB0fID3a8m
JBQqzjbpgsoCzInMijuxnLXueQO6MQMwKfqyrqpVzutavTziglswVo+InKHfgOHrwxeoiWLOAdwb
8Z1hIeNnBsyngPHO85ArizHJJMxM9gPUigDoEasFeqde3AmYCeFikb2c245zUkUY4Q7oWSS+mSwb
ToMADuJLx3kOqtFE880r7oF6jl9Mj1nukr+1fq5T3+Ad2T/tpOz+7ZqHkFwnPAvdDe7avWebeNGE
rLTln9VrYCtq2X8VAUyOcPWfeVrTA8hkByz0/ZKHQF19sXQSzOiW+hj+5WMDpEKcWujvX7ytYgGI
DnPm4Iyhs6V/VhuCqj4PyOBHXq94EuEk25zR37q8UDM2sU4h/uKEox1FVWIq8yrJeXAFkIWzDmhh
yip2uUa6IlqzFlEjfshMrd40mclybrgqGzMTtNunvewUdivbEQS7VdcPOAAytDx7DRRTFEs0MzyN
dUDdD8Lga7xqWp7Pxj97eZMtFQ73F84Xk9f84I4K18hO+4KzrGtY25yG3ROhhhbvEOL5empcoVI9
X+HsS2cKMaO118r/HQjW5nBv1d1RPHTrHTmHaWcDW+Kzsgc9m/7mGS/SYB3MCOFNOAX8QSrk3eCY
OmTzXtAuuriR2rNaTFTEAXGW8o9ABKFcxsp5QxuuVJeap25YhCw25bxRGrI5NHAGVZWMoUIVHwzk
Xq9lEz7ifKXuvka/b5PwyrJ5MLT670RwcEeaRfQxTnkmEXeycht7QGRFHlXEegGFpQCCLcIv5KpR
HrYoE5HmhpTL3EgLwJ1deGx9ydW3YrK/5jj3MjmknqhV6WybBwhMWDUNzftlMWsXjzLHwaMggNZP
0vtHnYqMaDx7nGjlUQDJNs7XNzkJuEetPZsHQLVYt0ZJ7S3e0YB4tUMXHmcTQT8rIdpuVuXCOlhc
BG66VRmOXtNEmXWxvPKrzS/RiTI+pNxN4yJkIUsmO4CZiMZpFLDgJ5DbhYqBJaO8S/vQY8bc60xX
STOjtin6beHCCVkHSqMRjFWhGQFP4vMz5NF1SWKzLfY+Awc8fompfejBdr3nARsWQCfeg/8xs71z
KJiWzMQaaYQ9b13BuonP2b0GSjUErQ4v1hNj1JydeoIl98kctVXmhY7if9YcxwUfDqmXGX43sOi7
vrVaNhtAXaEfbF1EQwGkNGb/5TFuauJPGVL7IdLPHjXyJKmwvp0fd3z8BlW5O/LaER9bF+FKKJic
ycZtPFut9ME/XevbdfrcTDuv7G5yibFRpdIh4O2YaWSaI6saPGSVl8tSBi0fonjT8TSqPufBP9/i
kzcUSA3j7Q9mevpu5bJrGAYMd5/g8eu+tbFVA7LbectqncyUyb2heMIjtXyR4zP3PRH++McRXZ/g
NZb0Opb6z1E6MV7OTPiBt8RSqeeTks4y2fOMuFjVYnWR6yFdMAbrc/f8Of0RayYo22d4JSEQ5MBT
ZYAc+SieUKKLVfLq6B7MAhmObFHDaUAc4mWy9asDaF+TmPRdR5revv9nfil56qDFlzxardEDjohO
tjS1os3jfGZGLOnX/xBJyQg7O4mW17GJJqdSUzEvrdUB6Duj7fu/KJus+jq5iHg6MpSVHk2t70U0
Wf8l1OGb6TMzbxlAvoAlEtvpCzJ/EawdEtpj7vSHaDyu/cYPb27wGgnfpPvuS35k5x6idCpIXkre
uq8f2SmZUUSE3DmJqs4rBgHbR3PmIzVQDhsiW0mcRQbUMlfsiV53S8xVj/kRNL+4VHVnD8n/Nr/X
BNGqijjo3pwqki/6f20AObyjtmTu9mEkO+xFdMDTmRoSVrSdquJqWtzuA1JXaOoviRifI4SZvqEZ
7Q5Sa1Oyy9nbIXbkihU3g8K7CHb6AcUmQ6hjI/WqQY/m/76omNC3CEN1DYoC+5FnHGgMMwIxzu7p
dqlhq5xfZQ6lvleorHge2V6CXLfDZr0ouUVe/IRLBsrtW5FrAxQygkJavBrQh1sxw1KIDagc3Bt9
2MtA3rZL72hcWlRuYGaLB1ZP2xtX7v2WlFl/TaGzWANn8y7jjZb52zCea5shByAXs2jv91sfogvL
Ag6WYEBaVPa1lBzz7Fpp5rrnijVG9lm0NNiawEsfri828l2O8+QyNvq3f8YHXKhovrs6WrrFoGdQ
ypubIsAg52sOGgO7+0PIuV56Nxvr8Bpbsdbv7tak3lJWOwR7Nbb+oONBT2nWpCaIo6lETM3brnOz
WY85Bid0NqWbrVC8EQjO8/BWv0dIKjxqtIegQDMuFxdftwAVz/PXrPZdyNyUwpP8wKmnALoZG8G1
73FRKhCI/7YWnW2SwhEqcm4uEKU4q7QXJWmMbq6WLzYsESek7egRj9QTnXONz/EE8rRpsEW7fxJi
wSAEq0kYpEvszgQQcrk88TYxCy9JQZYWeM4FL5NMQb05qr6c4qaAfWihi2Xi2ufNnBoJ8BXwbmUL
pG3/B6A86qe8HPdPzgnqGQmjXGfvt44WSuBDH9w7Kfc4MQbW7bmpENCFxueyMfFjXocbDUjkU16t
0LatGQ6+6Q7kpQbymiUGcC42Oneslhqw782qLDN2A+30jvzRie762SFJtzqHStnIKbGKnM1/0YtG
zLORCbs5B2uzHATCTX/BVpcfVZdIJuLPaCan2D4TVB6Po4a2+hNRKVRGH0qfawcgDqevXVtIkd3H
hAVt4M5p5BCO7PcltXBwhuzDicTMYS0NIfUtUwi6c8ardeDHRArCU2nfoS4k0LsBW+rziqadT6KJ
kVC74OEg8MT/sqUXyEm6WhaQM8JHbvhbH0zx824L9NM1yvAlBZMrvSRrJLbAaroiO5uEUL3fYgbv
2o5k2S3DTkt8b5w2AIwID9T7LjXRAtDfrhKYWxxGYy3IYaansU0NFcWMtgEuoWxm4M/DPc2yVOqO
qtSfv0h8FubH1RD02lY2BoWpqBReGPScpkwgK/D6wlDi2yV+xJ0yiaMqvNGWDbSQSOByogAJ3lH1
WhttX1Q/Fd1CxPexoH6O8QyojFd2F5GDgl9Dgzgq2xDR5XRPa4pl/FnBN7uNPHWGjS6Bm2FAWH11
fyjPjnJyJA9cXMEqIAEdXVbUwy3W/U+OiHoDaa9KcwGZD5/ek09fzbOJjFM7hvzTJ9rl3zdLfCPs
mFl/xv7vT+bXrXSdsxGBSh42nhFo9f11Wx2WHy4otxkbNocoJN6hzjK2QzT9DxaKTcFPxp0yOh0u
SSbi+it9t46QtWECfMu1IqkUN6D4F91RjL+zfRuGfdmt34x1seWcId8hErVH6M6csdJivFw1fr5w
ldXvxY4BSPf9mC+OtTyOYvAhcz7fyaUxB8/tivfwj/ODa12yEMpNFjcpC+B+vAGk2FVV1SQMYSAO
OtogMIrIN2qPngalMXF7KXu7DC3zRLTSRPY7YPs9MgJO+wkaSJZLm9xMUB5pnDw8qSjBTufAhkON
aHprOu0vb2GhdCHMlaTnHmBcQh280nQDv9S9cDVhwfUWRE6XawLMAi4ZF43zmelm0vKrQ6YBqniZ
c/uMygRcZqY36NK6K7p8qnKmbepK0ly/N64wptCtHXGmgDaCnJb+bY2fKB/PLztgXpY60YtFITye
4kajG6b8PGGeLfzhof61bGcPfXQVDnkO95eSB9agPgHkPrQD7EQ58VU9bbZ1VpRGTU0y7TaYtqyD
WpP1jkkegfbYfZIOq/QfXFZ8AcvciR3NAX5FEUaQJUtaV9w2N1GpJyG25oL27SnIq3XtjWES1YiH
l2FGmy72JAeV7owBwVDuWJT6VadHL+9+rhECpsW810KmhbWPELW4NQzxvzbLTT77dpGAf735tGzD
IV0Xi5fGZtKONxX+GzoV+misHShR8m6MlHMKueY62FS+XWEBie1AZXI1CMStuU2fVqOow7UgBIZi
mtZuIdHl2SQxSV6v411k1UV9TCbHvnLZSjSZQyPnKahLFW80ZAmnGo+msZvbtbfHYfvq8vxn1vuh
BDrjFnsgbfcmxZ6l33BWoVfiByZLDRXzyyxyK+F4vsGE84up9D2y0byJugZzApVNgo3mnaGxuwZg
7wziZeFv4rlm3axwr8MKYSE9mz73KakN/9A3CQdbtWaoJAmNCLaOIkoH/IWki4ybjMRR9Gg4nqT9
swaosoHDXyVu1SsQt+lyrbHsnzqT93O3ZJuspzujPNEpki3ddJZJ7WZfNvuNIILdEMNhvTTWzjip
pmu4Mq/Pq97Q/O3pSaT65HsnKCS8qdDGSOhlaXCWFYYPvQwY/44J6r/XZW5qqYepucNQbgjWKyiT
RbzEpmrAAxnPjeMvXDj4OPJ+Mx/cd3C/KN06Eqk+a9i3a42axtFcAjrIr+uhKEQuMglHJg9T7jhe
UC6LqlEBQfVavR0PNyZSciFnkKfJ7kpsajZNKZrvCBr3W5RP12k8bnS3Oise/A32bUxecPzYsFfo
0IIPVd7PSkLJpEuWq87Vf5YQpBW2XQVrrq1bzyJOTCNI1lzfXWBbln+V2H9SHDmOSjhjFtqOJdJB
EgKsrujCr6uhpTqdMuD4RAn8ZpAwZvRP7gfoX8iZflf7d+SXaa5PzCSLeUcVHmSBT6J0PunjQcXq
72tjgVEV0OnfrRQLiPbL73Koc9yPXlWPmFx91Khdk6Td+GOBc9umU7fULH9fh0Cw/j3kFOG2kU0E
ukqDcSAghbQp0cp6ISzZnvWq9D8pyr8vodMuHCfjeKR1e4EwQNf3JJBSu5S+pFOOxxNNAl6zIraO
5R7RiS9E+2pnn1I6znnNME23WIPdKV2lwVbp5CYw3P3BUupCg87b5ccrGyDK7A0WVaIcLB7Jw4rm
irsJUjrZQSwVJxq4ZwrySyWfWwwB5UxthxFhUc9MnA3DN9q6k05vxqO92LdCL5W9P5VlBZ/FCpo/
f2yIkHvHLFF2ooOD8TArp4GQJWY79+P7+RGFXznXdIaLI1t6Crq83Cx7xHIdGjbac4RIVZsk00RS
6sCL0vDMFysF++KUEDoTg96XoY1NuHh0NDeU1DdBrSA4lOv3B9PKeLk16GJM0zG+1Nv4l5JQpzoK
o9huJewyxR5PUQeixKFPMKkdB/PMcr+Zqq2v3yyHjzlMd89qWvyoq2rN+2cUyOgXHOy791YNFILy
4qEolWVuojXAJRvxQT0hdDnQlW1LBtNHzPXeL5sev7Tff+xCpFVv81PHcojM0wq/DB3B3GocaPs8
tvzAVFqzYFrWum53DA+8ZGNY5JJutrEGDxGfJXQlDfSEL2hqqTxhBdVfQZi5+OHvpa0uV6uyS+x8
Bw7TIhXS2zY5ShjzHHIZxscdqby+tO6/JQWxzjlwLS+bT3CiCOs66l3KxGVdiwU9LAD0YhhMEHnU
psettNhgQPp4dLKZANjW13PQhrKcw299iasugPuBlPqC8adyWHQKTWSZs98WmlkO/xpYxCxe6INF
/qEr8B0KFuy2ZtY+TlT0cHFeI6ZGZQsYrkosoas+AJpjavdTVYW+WGikwrbjL8GRxPINSmr2ISKh
j1kC0NHER7rNHyFWYZxli/D+FPeYNaOFT+/af1ym3GqbjoHZ01sRDaU7uBni67dkUo7IBCXJ7f1U
dVnx065pM0dm/EYCca8Sw8DDemDQpzzMysoBZdGiMQ+qSyXjamx5RikIyGpDNSDE9M1ljvXm1r9s
x3PUfJsEo5hxAZ7nJ3nICOYzYhWMm5KqHgtxZbHp0UhhT8ykOLt0KPlxh5+gLQugCAPxCz0fyy3S
+sEBL6KaznJPXNnYjD+pLD7oNDcNNsdio7aan/McZw6DKrXatMsXPrPANoFSkpxomyijAt2PinO0
C4ZWtQ2P2ogxJKRwJ0anoroTu9iqSXkuiN5p1ywnYK+80z9eJI9XfqdBoYJEcvp659S8zrP95jIP
4wbJliMPEbfJjukZAfnAPFCVz2hWNfc/TRL1MvvzEF5rLDrlFWPaoYXx6GZtwO51HHEUs3pRSlGE
uV9NGYceCtBajcFR6srkPHCfDrPYFNzZvakS0LydwxqayrrqZ0PGgZKPctg+oebLH5VwW7FZ6wH8
eOT8TSUfahbODDbZhQ6VidikK8EvdSPnpB1htgDPgMJRfP3RDLc63+WUuBWNa/C6oTZaWIG2JBf1
xTycqKTPCfN7VNWJhnk1R/ESV3pbb64F8O0J3fTSBe29nPbwduoG7pSCKOgESZn/d/dhv/0pi8Lf
NOOTwSMj7S/ep7qA+KqudtGq+/OQDcawGoa2nYMk+XNSeDWEZaoQ1PRSxD1qHY3OBjq+lq93cBXw
I8UdX2NWVYC8sA9twfKfIOunQm6j7NwySoKCdwUCH8zOnhCBJOH0y4huF4FLbLnjv60n3tUnXOlJ
UdNOP1pwkyAzCyNHUe/0ZuP1x4vQtjP6zxOI906AaYC+hP8lB7nADF4NQSj02TJ9e30BDhS0pLSW
dpr9cdbZIF+7zO9QXgW9n3xlqlw3sq0dQZxZG9aMffI9HYUQdo5kOzVtu3zAFV9qV5nTcTf4z31d
nUfa2L3e2xqlYdLOjEucF9VCHzR8YsHoF3+n2UqKGj4lN3pbAcELuQ61Qo+EgnKnzRwwgAajqaFy
zaMyWU83C7mZIVkcNzXvIwbbk67opUC3xIMpG5qLxLC4aq38Xg4WTR99ZtoCz/6ETZC1FoMJGlY5
/pIeC07CWBkxTN3k9MOvWTr/aQU08wX7CetzKiEDzcAMuwqe5U7tBQa4VOqwHlNCuhqp/CN8sR+L
jtLnHUKAm4EUzt6e/zG5E/WalhLJbNgunUCdnyWXU41WVlJHurIoldIv/xHjHsEFY96JEnU7Lfo3
zBRUv1worBxO6CNMxua46EDD2eHJhW3Ces5OATZ/t5QMGLCTI+4B5kFVWY/5QGpQ8flMHwQB+jBL
K5WpDmOpm0g3xgORGKKnjEhwwGcoibyk5vHsvIHV77W5yG2IUmdqQ50BGZBA/YKhr1Y+S6MTUodV
IxELK9Ms8e7KG5ig9UJ+z+RgdK7G7aTLK25gJHb0JlNQF5Yrl2+7/N569BU9l9k5+eKTeXxgCVse
++Y3+YTm3/e9ZHIRgh4dpEtaRYAXUQ+pwO/QGLJsrq53r/hDZq++5lF4xKbRNjqSLxKkxVw/Vhkj
78Yw4lROGoG+GQpOzRRusmpC5QV8Yw7fVU7bBxTwGUo539Z3FIvB3AS33O7kBP7o5THHuR0+XlLG
3ZGgAPl8kI0RXCefHWbEq1VVr0lm/BgfdHZyVb7qINqLxjl1LegDwD3YSfJUgIe3f95mG9XpzVjj
u3vvsUBI22M2Yvn257UzBwi38cqecXZPrRm/1yUNjV3IoLyIsv/vNEZToJKvnjxSuYsL65m1Wyzc
VRbeDaqyAuMliykbbPOTsj5TGjkODYEelaf7lHK8o9Izx4RuTSmG89+bv1Z/D4ZgmKPMADaJhpRE
G5Dee2+dea++6tbyaGdM+rfx15iitrXVQvGRtYyoSQNA4G+Qyf88MsBYYO1rBGRWfQTDfl2KhFuE
3LH7d6KlwTQGhuDSMAHpHwtwY8utK4KbJ799ruCXfpnL0PCt7yO2NurjfcfZRQmV9Jh9vKwDY+78
yo0bImr/49etxGLz1vg8j3buOZJawZ7hGC0aydqTm6D77lbquoYTBq0HKGTkVDqGhczQUYq75U7X
pux5VY661vXEJuD0M57Z3HnD7xyamh2Srfla6Rj1fV/bsqvIx+jckB8d9WC2WCYHLyluv4d43s8M
+OIOWFzbOYH//NyMPpn7Y34jTdkuKPp91wlZD+d6AKcGNHlAVoFyl9f9rVgHUkbbsoXRVx0rbD3p
Q/ozCqGJaCKLsIDtgTpvLCqopg1z7UtsF3M88itiwtob6WKgpUXZGFZzn2MyAvcp4mPnkNTGdjC+
cGU12ip0H3gRO9bigOikAfdtbmqrhW9xKbGDjyGQ14i00UGG4rMgPzT7g4qtgEImrQ7M6EMgMIa2
xxGH6xNWgf+vhdw+uGylULwEdn+I+IQhjODVzbQIaGo6JuQuIGi8qjNg1mMQY+CgSap7mQSWunOv
lU2wkTxYE109awHSESaiQZQf8S7waJFsl6uCLP24CVxB0ZIWlt9Y8xpL+RsXAYNtroFO0GqRp/5o
3p3iVpkNMVL1QD3Rc1lVG4iOhbkoCajjXirIE9yfsYyuAX7LGB2L+1XjIKvIFLDsdFAkj5Hnu5AT
NmzCiKdG1Mmudi6K/8DYrOA664NkFhppWByRAYIpgFZYmbXVpzwCr6ssBBMIsseVRY/C15boNi9f
jQqD8bRDNcKrart46rclDS2TLnKFevFiDj7JzjhGtgk8usAFiHRQLJPDGhkj0g+UePRBL9CR2eA7
cie1EWPY3G3jNb/0T1gfP5rzDxq2QzuuDBmUt6WmgwgP1e3YZ2ubDaNcjO4F/aB9kMvOYD5MB7lc
NProzocAmGwjxabzUSAgJ/MvUH3AU889ZPtsgCBZ34BGkempdAZZQp7DiKzrz478RvgRvCoHctwE
bYYpe4KSXtrmqH54taI7aDAwW7anXkQW9mfFF8fgNKsWmC/fWZiva+UhfS1yCrKptEF0qhOScvsA
IrGoiFTkMqEoKOEJFAv4Fir3M2JOqRwqY14EoeHbRmQsUXvvgGUi1YEQ6OdlLZ3O+pKV/EXOzaIZ
efX2E6mNDZfPSPKTqbr9ih7OTKF4FgONlmkpqJDBfIN+m2rMobQWhJp/1J/gNSVEIRhQRu5PcNWh
pOhqAUmM8anexnw3MJImlRAHSLStyJ56mtu67El5a6GnUCAlrMvfzF24ctyfznIB4ZueOnSplKqg
143VySBhRBXXtjCtGnDk2DNJJH8Pj1IfToWbjgMxptMGeOarCBUT/o20xE56nmjnwALluXBCSqS7
ldWJuxtFs4oe/bZXlEO8WOi541FNLhUJ+3rYW1jgwGWm/xVHZQsagbYs+8GEiGkSimvi71toOCs/
M8/9SeGiiXaw/VZ8DlyW5GzbWyf9/JIE8fj6w5EA8skK4wwafx66UGU1jZxW6EaWa1+F1P05TVPy
O9ZhTRnUoiFsFTQhDkcYqt6xr+kE+m0Qej0j0VkJvctxLGGsT+uUsHxlQmHHhbOJiU/DfPo1Py/8
Z1p04BhLLpXWN/qOmkAWKI09xRDReVHqON8vEuE3SvGBdioINWmCaq4s0Dnarz4VKNNsCh7XTc4g
bqV+qVoqzviHt9IgdTLZs04qZEN41rjpM3BmvZRvmoTWtAJl8Hw8vZc3r5V7okmq1H6jzVUlSsVm
r1Vjs0VZJvzakVVAFwWwKfiIcv82pcnWjzOF31qln+PzUb7E6TBBIcRhLGr0PCpuO8drktNIYFid
vEKKdPt5XahPG1/RWfxe4i32jRuT+C2ZFXsRn8dyX4rPRJ5g5PlAgAqi0ijCGfrkwLd5p2q7pexn
P2ge3RdbptN8mGdjQTKKEAMFyuEs+wkWzxHyaX/TFQGdSkgzShqPlLxNULR7e1ePGf5M8dHfBa1n
Z5yI/mFPWF5H2OtifqoNDU1D9aXoz1rneEhH/9bJFeOEPGh3AubWDvrOS0lzNh1HOiSHFNPz3Loa
c4KM5qvwy8ZyR/G/p9wySR1tVIYbTZxc5eCF36hjHEJKCftvzBsqSiSJ15niWAJH5b7v5W7cEcIK
kaVFh85TA8xtt6HEZC+NW/+Opa4Xvf6jwKZf+1zkp/unfpCiEWCGVCF4s29c8ZckW6OlS3POknBx
oR6t6+cDK8ezBtq+gMydlJLFzkcApvD0rLypf/ZSkTn+Rkd0RpH0JVCZK3qQQCfXg8Nnc4XeoOgu
sNbmT9mhRiaQYg8Xw+wjEKSNcR6bAqVykPuzNg6thGgcCsiNiCeVfY/SAHxZtQ9hW4gttZFNel0k
051+7Yf7XiTxegGM2ub0mySqFFNGqQDw+KaMLG8J3VkPdTa29pqg2SuhLEnQcSXmBB7tWxZsIZUt
W6m+C7QdNe27oOVgUSNpbXK2c046eIpnoRiDPsy+jUeYq0k9yp47sEM0lTC257TGOv35EtSbkUZi
xGPjutNrO/zu7FWqnBe749qxYfdnAaftXIN7B2mK5IvvlQsn93cGEQMzMPdg5mob+WcbPDZGwTa0
2yT4y6BKGK0iP/LsLPh1+BDg/GwowbLFvQRYXnS2TlGtzyPqD1vthOXcPQ5WFjVB5/35hOlBxelt
pG3BzUElEZkdWU9GkeXg34BH0Bu7hu2ElS2WzQKT6I+utkcJN9RzbRkZ9E3FT7nVOSy1lAgfmBFE
aW4+a8GS7eUD48x5tABiCj1juEsFFc9f6lT5hep/flXuh2zPhZlRN2HDcAqtxXSbZlTSlDvc3nHL
rm30syGnJqLGZ0SugheJJen7P5y/wOUxSWtOyk8TCOm7NWvkZ01hmRpDv2rszZgVjP49M6z8kZl4
2lnUnvGjPucL0aPrEww0NUZwt0jg/NJKEQZAuVvDaVp8kzmmF0cIr+glIAM6XKkckJegvnNru0zC
ezoY4aGkAvihNZ8jXzvv5fW6INH1FRYHP54LmfK8R90/PPUFsf1JsOlwymtMvhTP6p3Xuxp0/6mk
tROUk+W8nRWHoaa4duffmY9LLRo6L7LG8ubHf9TCZ2FVf02hgDGXBWkM5XKXIUEGA2x3Poemi1YU
JTnY7BjaheWNTJWi7j+8ZO1OSo+lsf05QOVocrVOskgt67wcRyW7xLXu3sP334YWj3xdMicnDFz5
k2tGZ3gZRDCCZl2PoZ4WRD4po1yeRPihElOcBvYILGfL3qu8WEaNmBbnvoSzMY5jUM6qHqYwh2XE
Gsc8w0LkrXSAxoK9KNuS6jMLSrr6UmVNIS+j4yCiXq8cXQTMmvL0elIHjqP/GBfozhdTUXbt0XZs
aN6uyZXLpjFdKHiJxZHM5+L7U1ejUx7uO1bs1LWehZbLoaMIMAd2JgCOiJlsYXCSIsuLR6iAXcxM
YI9bfKc02JS9MTgY/jyNzduqkVRFnud7Mu9feHgzOgSb6kI1IudZwdhRlW2ujt+zlTnoalIYVfgf
b9FbofDRAb+DZCR7hPSXSnDKmTfUxewXBQNKxp9QoR8Dd8wgewr5//FDxzMGFCpNevShE7dz1Ihn
GoqfLJsC3quOoot+Hq595xs9BRCHsbbgc1NwgjiQGFvZRV8D0ruV7dKUdGnIeT5cKw0fwpVAd4m9
vMfSJr1tKcpEEDw1JGS/ar+OHHNco7nDwtOUa2PhkrFAboO82m0t5ztgBCRde/kIloFrMbOkF9KR
d1IlR/5h+Allppbl08pY9JpNd96+xq0XA3kMSba2+Sy6VoGzp6lZn9gcNIB3XQ4+ykw3h3g8O7lC
5KLPxJ/3OgAfsMd9pW7Y7mkBEu0nhmnxHBYYCnFWv0CLGPFvLm161Od1mR3DN9NmKuZ28zR/fJga
D3kn2s2lwqz2iP9lCOZKSfnAGo8lQCwUlRqwpHe0OY+fQ3dJSiFwQf5NPwXlhyj4xJZ33Tr+MawX
8KgeeJe6MMZSetgBsAIpVZxmHSfssVYtBN7swZ95wX4N5zHCHHKfZcgGv0CsOzH6hBD2dWviYPQy
E+BV8Syuiha34bKZXm0dt4yE2R53DY87rPfDJeGap/DA21Qjt8IwviyZerIZTteKbMQpEybQvC4B
43iSI28WGpCmJvjVFcdtIvYCKcAoytQrCAMoEO8wXhTgNUBtzW6C3qQZuTCf7VahhRmVgA2f5RXt
gPwXS9lQASZQPxs8VGUkzuFkUbuXwvaJC7byq7DBNQ0Z4aQVtIWnXZMYg7sCZDXB+1byrdTb/wsv
hg1Blr5Ow/pYbY+Qut1CKuODoWOo63Km6T+w8cwE+bO6Dr/AbERK8NWkwEvU/A9IzSZR0sx+OAqo
C5x/YN1QD8p2Xiq5S5XjKHNJ/iiIhdMO4UuGKxXP+n3iU4Tqcnaiw8aiE61lWoKGxSbBK2CHkJWq
S0mOGc2MlFdW7mvYoHghPrt8TGPrjjTixB4LdGVdt8oECvTZnCIto+EAG0xRSZAiyIm51YNQ1P+z
KNnMoLmR8ScL5ba3gAsbVwPd0bJfnWul8hDOCyXBEY6/4T98kbhDvQirxI4kE7hEwWLFjYqt/wTQ
WB/pc2Ri0NY0MNRF6p5ocJNNV3ZoEHoZE5XshS6Z9CWNg7MnN951IJF81iVKcsl3C0g7+5vhf2vp
D+3dMaNCgd0FL/PxMQh6SR43rLknUdw4a/3bfBrzq4gjgHHpiY1o0k+5iYvZaJE3WP8Myx03yxL0
HitMUV/7A4N2o6MHifyEApg5ArgCTKC4pAY2c/+msweHqJKwJmiBcsYfFHJHBxP50ZlasKCkp5Da
RWp9pmBWrbD8Fpbw4nDW6GVVKxLtPNNorYJQZHZ13KwCfHRl9PYd2fjODSLQsFik7eoR8D8R+6Zi
LVeuJ52/mxdM7quoanyfBObbPsThIMcC/qdnr1aq9mHBvHokGvEF2BszTqcJHMaXE+TQjk1CVvqg
6cmXs430RCsfQjnCSRKrnHFbqHl+0n0JJlCozP9oj/ddHguEeRKtDyAkT1OZP/H2Rg2rxjP1aVye
OeY89IoOiGgA33LvhR/PvQjNdL/TgH7ISi3E9LgaQ6WtOLhWsx0xKLt1h/7i4YxLiUezrW/wbrTq
WZeqD8L+9edARHuDacxc+dLxgQABELpfHC5Tu97bIoSOinC7NipkJIrTgvVSLfAp8d9LCZZyHmDg
F4YXSuAXZ9OEuevd3HGWrRYr0cD2agnPwzVF5cr3kvrfAhH8YPIrASlFabew9q2cIr6ZleRyhU+Q
04/dooe4vCo+ND7wYNiIs7DiF2vhu1TLYHJ1ii3eFxeC7rPzM/Brz85LSSQSPK16bUHCCnGFdHrB
ZqLwchXJ92A2nYdk1e4t51V7IzOrW4RaTw6B8hyKmEZ7tW2S7bZN1NeYDFK55pbiX6h28LLr1Nzk
RiEfRJsGVuSETD+PDaOcacOlf3gE/asxUIKVx9iXGcmppUFsCSSl7A2JoW9a2mUsZ4EZSma5UhKG
STYh66Rea0dAxybobMISNqE/avxoVL4zfElmkqqMk28VNcbt3LT0HADQRLyldzJKlzTe0qKZVqxq
np5yfFBiBvUalCcfBIkNWQSuIE1Hw4d7nTXwnQhlPvUdb3i66JFJCSUc4gCmmy0LDTNwTLwtlUUz
DYdaUwEQopnaSRgUmQ/+eE9wfs8JEnuq93hGF61laEhOYTFw0/qSNa3X1NV3rjiTeeNaoOCBzyd2
pF/DK31FvcPwQV8jVDL0QqBN18zmlgb9fcoGYWKSdCDDEHgKl4XAK7mKFKjnI6rJsBCFXoGfPNqy
5Hy3YHHC20elM6peIswXydijKtWpKBjzXIguINFhX6dmNCulPgMeKEg7djwotqsyBZ/GvFJ87ejX
2lXGPWlCKd1fafeDSW1dlo4CK0GPDnrPMCB6Ll03AMa9AbYpneiRKXdultyJ2MJ4FGpl5Xz9YMvD
gVpNQE9QmDyfCS0+uPPidZ7z5p2hS52d/KSWCS0xlyTn+O5wzmdc7kgaMdFUeHuDgsQLI0S1dO8o
CAKf3O3bK7VoK+IMG+ZFan4Ai8/SW90ZiMzK/Rz0omEgZA2qEvD6J18gg/CDCVr8KsiyGRuMpL4G
lOqQOQG2vUnPD12Oj7pxhC25z2xyo7BfYlSIqW2mdFV40jAuTMBUzQtMOh/H9XJYo8Ps3sTZLTan
DMyUYJ1B5RZB5Xz2xJQnJmyZIKRdNcPBxi8aCWAyqSGKhWVYnyXwp9A9e9aZBM/SRZcRce41vMtI
dC2L0Mnh0ZJQeZbzKdIL5BenbRHTAEzs4te1pFx9apxP4HEoApMjeCtSkaD2bOmN5O+zXEh3LiEi
CPesu9oxde+6IHPeuOUysbKYfIHLdwXtvytm7mX6iN86rZka4JbLgj1YXwBT0jMM0WqMppAQ0VWi
tCskM0Gu2meJLANec0nsL7USkAWZSkusQa/3w3MXp0Rp7/GeICg63UDeQbGq2gHoI2X1Fl068MBL
EAT23D9W8rysTp9I4SrJrptPIOEF4iU1Gskanh4hE4fc9teQlkjzRXVoPboniOmTk6uUeOtrPzZ4
DuwBn9Gu5e6kl50n9yiS/K6Qy8tzqDczcEmP4karsK50QMEo5oq81xFbEhzHI5SmAhOOdSkpg72J
rzj7egS+3t6SFrWApEgN7HwZ7a1xmdY+WObn1TP638BBf6MPnMFVhTk9LOZAxvXcTreq/n44YX0I
TvRMOKCbgHBbyWuplrdk//LCsy3wPIlFgT1yn2qxS71Z5QrYdUgo3GMVJdTfGumfVQly+epFi4Dl
z0Hbwlt8+zpAsmzoYGa5lFYoKGguI+pIlEKO9jPzYceKGYMviXuV1nKjS5iLifCWR7Qmtw8KF515
6SM7Ovi4rN3rrDBDk76mj++Y2pNHfdgkDoCJLYXRisY33PUBxQbFu02tW304cVBlbmjz3XAO8MLD
veAugbeS3K9zopebtDOy+thsCe1IFyOhdARyqk0PAFZX568pk4QYRoQiL0uixK8S4mHVT44Kte15
0tSCmCZqQ41R/BEZfBDIkyZfStzpLi5QU1bS0D3K//uFFNUF7arXsuYKKkqpzXWkz4ljtk+6fu8p
NhhFTO7RitswLAvv1QmtO1ktKGpd8+m8u39Ao9Ke5I/m8pIUUQ6B6YjoTgSnGlMKScmA/bMolCIv
ObYdZ2Aulg6lHJz3Ggez7HgSM2EdPBfN5ahC1oFNHql1sci9sRfhOncqLOTKvr2K3l7akb0gIkLD
hFDsX1CELesjAOaJ6UDyMtyIEkg7zJWOpPO4rgcHrBNe9akBNVIfILVvp1M/7vTkYecPiQcqc4hI
P1SqumgHO+GBbMnMZDvsjnLUsHRPIwYBAaZq3MfsR0Lbl2n+cZjCCadeuCl42U1P/oy9OmHrJF1F
k/L3AMAO8qZfgrRWsfGSJRNTpu1oCZqq0HoARew5C/3VF9yDU+1Lqq9Jbhpbul6BgjoRYXsSAUEZ
a+sxyqpEsIUokf9p0gKyz1FPiNrvu7qIYk8hsgeW6JV0Vpno3uS/rGZr8F9Yi7LPnmSrTl1olHnS
4NGia51Wa/mwvEeN/uU0pb6UdM1ZvRrrbuHTaQMXO4DlfKVW/q0rGuJ4H6PM/BSp5QRQckc/vCG9
mP0GJYXajUrm9q+lvVKh6tAhUC7gM3O5FW/Uly2DlcXAk5TExka/3pKl7nIocoiJk0vlfgQxcplu
WnEmR4t6krvx2rzWOBxG6G1tZomYkqRJUvbvdG9/7o/S1BsNEh82WU/jW4tVz02TLh4KoLwzGRkg
UQhsD1lg0XIqZKo6xHhGE/fYq6kNILZQie76RwscSMFmLnb0wN4rJP/gSr5DPSChsnS72vvRaG73
3w6z35NhTnj1uUPUuuHHXbB0lgsr/ojfTm/Sn3E0zGGOFnkW31b2R80DOX6K0HtR2gCbaYCpwNDX
Ctf3s1uiD9/MtihtCwRY5iHZ8aMN4tutC+tNEf4Qfw9p4IFgHGluJrdhT5dvCary09EnQWV8FO9f
UiqfJ6O1OxGbJ/7WOiZDn1I6DATmCu7k3X292YuTozcxIKJH0W9N4He1mQrHrye74md/XZBMh41G
V1dMD4s2a4vHV7mz1Qy7sguH9PBSrmpBH99FR1pUAsvFN42raZdbi/z20gjIXPTGjhq6tyHArDw4
Qz2fCFsZjFSex+5VC8OYMgdVsTYNiYRb5m/bFZKElserRo5uDoyDr0+nHr49LkCAbZJoYsynp/jO
Y+b3lU2I/VR0NI3cx2danpeuz9DDF8k1TF2w1/pBU2Ir9GyNrCPlBKQ1IDqgjrphK2rbycf/z8Qo
XRhGEBdZJWUgCKjbo3mlxveUTbx7E7ECu2Xu1DWDo2FOd/BrNVoMVyheOVokDt7LEn/GlsyIJPLk
R3HNwyL3g3ckxlKcSmTBpzzR1oRSQE4hfCeHJ2IC34ssSm0DBh+gm9BcbTfvpyPsfiCGDC0IfNHR
H7rWuUeNkHEQv9leKXMvY94C8k0mCGElIFoUJqamgKTvnioC7M+w5tUHBPfZnV3EEFH/skJcA1uJ
Jg/eRaFnrVUbJWmy2IahD8PPN6LMOYH+3qe9mTen9n4cUuXPLb20QTSv5pbOeG6gQw3NNlov+LCN
L5k6yvkhNQT1lR8MFczUufYJ8kdsXEAHzgPJo4cJPkYZXQIsrpZdBm9dzr7tPR/hDjJ+BehgLE5N
9CUXTajKV/C46h2tZWnlT98oaK6IIgrtczChcGVnwb+DifFOBX0fF6A8aP0iPT5IrMMYKf4j72UO
K9EeQJzNao/bUxGNT5miMTk2pmdhTxLzq2EG4ZuCmSKiFbNLX8/q1AsHU2azHBIM20NWdWdHBz3t
u1xtr+eiYRNIxWAUBUM+cJyDZ1SFVxS2RYr2RYdCvbfHhfrw17lpxB+QaGn0SsQ7hovhBbYmyK0w
mkQ91GrQN956crf7FIczPDClV36f4wwhAjcVdhsHuIN35P1hHZ+/DNzf6zzgiJwwDt8RoCiQHXMk
WNRCdxfnBSLJuJdTC593WQRcUaVzzVN25iADxd4wELAliTtmZ/bFWEnN1l2QifAaGXHxd1NOcFaS
R7SkXnOXOwP/L/BCVLb6/CVN2C455znu4pE57/oiHvB5dUlTgripYgsbAzcj2NvyI1wIA3LFXRzT
NzuXWkOm1FBSwOTPp1U8o/3XK69NfQrKc+maumb4/8wUNbijfFm9b7BrUCNjXbsYy2kHFVluYW49
4m8LLM56d1vKkG5Ay7C0VRmxceXskz7zBJR0G4dveMO+vrP3hDJ/j3WHi7QA3mW9+5ALPuhkGUW+
PA49YFe6S0AcLXUXhBjFq1fx/yATWsEuf91ldGXGxV7v0YlaJ7m/cWO5cyyu0GotrVJTIjjgVKNl
fP1g4NbzYyqwhUDNBhKuBVM5kWgHcrTv2+B7a04mIogzQBaFDYE08QITtEdQ9PVGtL+zOAspL5DX
LjWpyPJrJojc2JT2vsk+C3+yorMyeIFXk2kBEctSZJJHkzLro8CpNLqsG+qU7I7RCAos44Y/QnUV
WREwi/CoDp4ODGOe4oawXSweyWrDS19XJC3iahjQXVYFbtqp97WQK1G7qthphx0MgphWLTtC+YNp
mPdzllKcaqi05cVO0YfdjRviRvHYMxDdpUkbaf8Y2u6YqJq0v7zFB/uR7fRiiBjKPwj6YMf4XzsN
ZGEVrmt6tdHSvt98Q/9iaZVYnyodpw0wKeUduNw3JZYVrtshFBXYlUvtZ/52/CSrIIn9Hk6+h0bI
yAER4gp5p9bZUjQrE/fqm9rfC6ZI61qdfPnDZ+Hiumjf25adLAm9RSUVCrNHBU681zwX0gR9LKcj
hIN6iOsxOefaAbYiP+XkLZvCaLyMCE303ihcw6QjyWMc7yfY+CAmQrWv5dilXQ+xEZ/xRyIuHf52
lutU8/j+Ax3LllTNflhl+/ZjE7sxZenzB56aNNtGq87O1SkAdlQk1NeYXiVSK78UA6tNOcr4KXs1
Qo5EsjQkHPdH2SHPdQRX35qhWKtgXKmq96+OR++vJCQ/VxPiMlbXMsP4vK2XZom5XscvXp5TZBKh
xEqAbBMfGFh+WF+rVwmhOAs5v/5ElsImcn6K/RfvvWOYSM7l9bUrvcU9INyHajPro4RWey1vuPcO
859lpcZHj9L0p4V6Yhfozp00YugPqrZKopTduAF4KfeoGPHUP5DorFx+/gNkJwq0yd9tJ9GZNiFD
DiAjeyJ41gHQXEuSyf6VPPdEOLTd+higntMlHSnqKvw0xzLlklrvRxylbqSeFLL6xo7xciKvkaEE
mzGtpNnkCeBu5ydQib6LpAP03M4hELAg6lbB4LheIGzOOXHjpvb6DQFv6IL1sehV8mCqHRZqfix5
5q7TALX8wFB96bJVikSwhB2T9ayY5wIi1cCwNhP3tZW+A7Udr/4r+ozTs739uCpm1IYaxydCfvw1
LStgn5su62qFqvXTcrXcS9XfswJjmrbRmaHkf0RcmVnzpKEDJGU8hZoAyNSxKBqXvSZXa/9zLpFI
4mLDQKHMyfmslvuwsmoMvTBc936tVSh+PDSPjrqvWXM6JOLfLTYrqVabodwoocKGKUFiIpWSOzW0
qa55wCcj4yGVzh9IkDa++iCyxXWS61e3yyLf7EbfRWKJfUBT8m9MjQ1NWOvXu29d4dg4huySx5js
GWvyZr2nLSuT/o5z85dOszIosJEd/hpNFdaZu7W1g7uBJ7AsSrcu/WkMHWqVqdUnV9KvmkO4hpCe
swnPDjmLauYbnDAPQMR9Fb4JAZg+PWBFCtP7J4yy0cn1Kr7Ux6CYTBh4lzGquq6aFVtu25fXCuqr
HmB8cNgKec42XIvQAHb9lyNhiZRpwdtyCn4CsVfJ3LBp9rpLKvuuoe98cL5TWfcvqmKgDmFyaAxp
86ifWUPCqjZBZd90yHBCswz1+V1lIWbP65NZfqKXreLezVur2/YBvft99mQWA5e4lwxPi7MOR5Sr
wyEfMhyJVPuIi2DVLsjQJdGJWwc+S1mgksWKRVASUZWJP19tsze2L8YdXAoUd3MhTksdD4zU3l72
WK8VmMvKiilp/Bo3T72ntEipmHyVgax8opYEnuje9xVQj2A+dGFWGVn2T5eR3SwfxBp2TkRGRbkS
hVSa+TNeOSF162hlCM6YQ22NQ8FRJdjx8xybPVV7GhC+uHSoW1HMYtkWX8xRvWJHl8WLCP73YSFQ
FVC5tOdZ4Jb5bsq8p4nHlyl9Znb7SShdZ5HhDQxpooXM3cPpIv82fZ/x/MpJ/nhEzXs1SWyneVPv
IocRIA7+CuficI1Ut//ReShJQ2CTPWyk2RJkNKXeBl8eRHIYZAdlBZ2PmqFV8pe3JWwM8IajG84V
blIQ8TX9QusI3RkQ1E6GRD/q/ihkgIcqiE8+lmeqnD20Qft0CFGNdwVRQK3Wh5jQG/M0rsVcPGVh
GDZv8hsgdW7c9dWW+AtbbCm6v0rBU+TB170NUh7dw5OCOTiMzcJCEpJInQWg855I1m1xDXWWVobx
JAY5NrW+Sn/k7WBbUvDQiBRb58T7HBVUKTxrOss4vpkYYftoN3BAErz8Q4siwHyAwZ5mEYj6dQ6N
fOMhgbZUESJxJr9/wTWuCVAFpu5MwOiJx0SvpIan0dumZ1CjiIydoKWAcUTf3yX8ynUdi1wL0Y5V
o+wb8TdiTXdq6qk0MVU1yZ+awbpi9AJBE08tXYBazZBZQklrQ4LIpL/Fn/oMQZlUh+hyaebgrGii
QMDC3/av9IzBYXV63eg7hQpVCRU3tvPrOaWCOJ8ZUMA+tqqC9YV8inRVxyFYfNyslw2umxWmEGdf
ke0JJh2W6dQfeSDQejECof9eHhudOHZLSeasaLl4CIfapuICJwDQ5Xyzqm3lwMoLCbUhPUK0uva5
d+Rl2xEMz9bxqRwlTZwd1zwqBGpjuwvZvY9DQCdTcz2ka9+pbouiZT9dOcXJdKRPp2FcH8tXrVeG
2bdT+0NhsgiQuPau182hFgp2kk8GIogOEiEVtuWLyDfxQDKVDwpRshFBiRv+j7sJBCvGE/KohAE/
AGePpq6SPqBC/1SJ113EirWitTcQfs/oKtbAtZGWamIHDajbibddS+rcllfnib3wGcvktGnfag1Y
eNkxvB7CicmJNXgd7zAj6XxsLKYAXTIHtbspwVDS995JCf+702YGYtXcfMjskNS69j0sLoa1v0n5
L53l2zRLqdzwfylshyeYU4a19eDNnafynGrlwgaywIK4ydMz9r529A0IwBfSRXnqzs41uSwuS1PL
035eXP+ty/C9FlTJCBap1jfjJmBGWcMIZC6N79bPYoNjmR2eNeg2L6Odm1g8m4NEoZ9gnml3GMUK
2CXOkV5chkRMx+jzphqsD4XK8jcVOu2PhV7IKAILt+c/Y7zU/gLAEPAakVrMvevQD7Oa2yNISMQy
nCbESWxREQUF2shQlbexLB//LG4qy10hwE990i1N9Yz6N4bSCuhxOW4wYflze56qiLMy0KSry6dd
94r3SCx+Q2kUgJO4cWgS9JkwB8U7qLPgCR9tn8YdBhUSQvWa59e6hcYfqUbHp7aBjhnI4y8zBaPT
asOjKbT6vIPS5IKif+ddLzTEO6uyX3ASQ6VqzQoSBnpWXQdTXAayMq2C7s3depDQDPUL+JDL+iDN
5LXz+gnemSEY1iCIFlqIuxnZvXnyuQ3V1PmYHBfOMc+Cna6vBy1DEi/2sZ2vsoRoZGrh2nhPdJcU
+GU0Du1ByjKxQ8jiIMBk8KIiDA8xOtpk3S9LUib1QvexreIcagCGY7eI5w/2TxWG4SodqMNkUAeA
O2gJ+EoYcu1oENrFnAVJ/cJrdhOwYQQ9oZ4THtSmhAlhO38SD2agrvGfmguYSI/Y53yAnfsx6EPe
2S4hMDfPblA5DnwwDEBikuz+n/gUweELJcNAkifMM0AIa3V8aeOfYMOQOewIY6FXcVoWS1SKPLGo
7V1dnwhLuLZS8AH21hCuYgAlhydyokYJlB5glyapZj9vIUjjoGSIfIml1u4BfqwtbDavER+23WgF
CzhQV3hW2Gk+i5JR18OSagWSRLDESbLHC4F1dmRybXSZm0sbr6xxg8wT+DkL6F2ivQ6PpFT5duSR
HMYvVgr8RrGNqIisn2S6qPQ4Fcmns5PgCrS9pxOoPZPj5X/ezTvY0DR/uCylN56IomtRHDmwLF7L
RPXS72fFgzYytytaaVVH167CuUgWYK7FjSsr0rgqUY3qBV4HWjNfDYdvt3IbhYzta0Hf5IfyUHqu
6YOUQ/lUeYm/QkhplzUYsHBTcur14nUs1XAxWyJyuPks63IEtyJrICRJBMrzIJWu62Aa72iIvl6+
wKI0iXrCK/ubW4okZjfqLMXCSopn0Qqpk5+IETux192VcpkMFBAMQiJzmsdrQf+rSrei+LmoZEV1
aDPyO0QSepjzh8kIp7HFDl1WSm3nF78YKHZFcaF5rDDw4QC5EKtRdbBL4LwxFrv1vUDMZlD9KRrF
uAh5Y3DAwWz+IUHvOppeuaK7Ww+cVPwPgCX6sfFIV2PexYS2z3gPuXmQKTmE5Nm/zrxh6kgY8uBr
PbUqnrJepu6NXM68qj30QpT20mHc4dqPenpZ2KNR/zDvXVmMU6NMhC8SY8SO7n3/UpTy3jTlbm6s
bV2f21gwKi9SsfUoIUNRPkEnQs1qS60LJykvhyDwmlGApmG5/YdyUToJ6jEfXJQvYmkac9JbiCyT
+ziNVD5sPnl4377YuYdSbNIt0OMRGoOySXuvxx+/JUtB6OTzcdP7vg99xCd2rgUlJg8UjwSMHNe2
+WWHKOhUVd11HL/jFiOeLcvsy94WK62mNuB7c33rVMrqPa7weEfzCp/KinwCV/jlsvci26ZSW1Y7
OAXUxtETbI7m+JMwTGfuSZGsylhAHXJZ/AxBv4LQ6HpIDsyZfIIQwXSqPx6PbmMLZdwJli74ztoV
Pk3e1+OY4JQ/dy3igSYMBtGNyg9yNJl2Ll9qWVrK/PXE7g3bPI4jKtY+YVN9YBk5S8bWEvEcp5c0
9pwe3ZoSfLoZzZbTJqt471DB3iN5zz6S1GuLsktJfkHe6WOQg/zDTKDcIcLSTEzzhOJPjSVEACBS
rWuHhcW5pdF1aXVqRiL3S1vTsXjxDs29cUIREP9T2flAkHe8QvzH983khPROIgiehxd6eyf9pCFW
X1VAV8GdM8Qdfd8U+CS3pmKnwfBZFwY9/2gmvgiuI+vntFW7TkwUHxs9L3jH1aNMKWsFCxr6h8sd
HgqZFix2DVvqQ7AbJ3laCTTumqoGR76va+dqHIJNZ86z7GwyT0Rw1dVOaUMpscuD4nGG0hTQFCo2
Y5RDSPEksE70wePnQkUutg1KVDGuRprgcBzCSASM7MFY9x5PRP02J+wHh+JRfKRBuqd+lE/ThdLJ
aDiys0bi8skzRMO1oAYuN0+DjgVimZjqQByFi8XzJnPFlu10nJMo666V77Zud8mrUr1aQ8XQ/cwD
msi5wRV6l/poUONCCE5zgVCS7E2QuWfm/QD7xX5ihVezJKf4ux9vw2RhtENsOoPGktjrrsmSXN4e
3DQi1CJtKsxDdXmpZ7LzSuVdw43nna6CVTCOUJZFh1aYs2U8mA9iDlu1duQFNpa3jvIWpnib0YtM
hDd4VGKgCAYOgBCkw9xME9cg8PHphZSwlUlnOA4qnkhGaYDARQoyUyDqe6wduAzHE0u7J1oDvFrK
w85ePFv17biyJM25TI1t85uVXVoSAqfewb7bs0M8e/f7/2TM4TeVjiF1IeCjO+WIwA1mEpPoODuH
8VWxXHOblvNvevT3ktZ1ARNG9Z1IRXD0VdYCmhjwbM5w+7yI4lM52x8Evit7Z3favKbfUeLwT06w
CyzpfLbSqpaAJ/OhJEdMoTynTyxwPT1WUWk1WwqoXg3rSeBDtWWhsacqjzxcs70AsLw2/gbBvetz
tRnE7O2Spyhneiw3gtqmH5+Rq4QvRKfIJ7YmtIpgwsnw6YXC1DkcadoQKAlOnmtPgb9oRBSBJWGg
qKRFE3o1x6EqOVVQfSrrxBSOk4O/2oqqQs6aBu5eTIMVEbTGXBgzww/ZFquEoxm1zV6+ZBEUUU2W
1jXB4jAX2QyRSFGE/D26xh+nJX19xj58H5Ap6q4ASOXwq/lMpb7nZHrPgq0Jf+Fpwhk6y4ee1y7Q
bA0OQLfE2NT45LDH9EkvPfOx0ReK53SZI8cz0A7fDuYpTsStOsO5QP6hzfN/N/a0G/w/WkSw8TZ8
DA2NuCHjlEe843U2G96dDpYG/yDsjd9hThnQ+wV80JaVhIy7a/U2XgwOXkPjLaRBq+CV7DGwIddX
gbdnlNSu0LcqV983KeYTkBN5pSOBotlZLGa1OuSZvMM48Ndg+1+uMpf3yR8el4Ig9LohHVw8oWUg
3ZLANOrYRRf+981cuN39DvlnuJHN8dMxLDjmV6of3+VWtpk1u/McbLpzhyaz8wimVkwhsE+0yARY
jdfVZFHGflXyBiUPD6QLyAAkBhyECWM0Rw0XfCbv7zgtlxgTEtzIPkbuHEAbY08PVFce9990xEEi
/KgtHRluiRnCVaDZNpFlG33V/YnbEBjH6RKUbl4Wk/IRT5o1/v6zFRL1tbxQVuCSaEs8RQGPULzn
4fgV3dBcM7uV5n+sjFnHoW5+mbse+QjK5+irWVwqZmyAeNIIUBZGyLrdI0P+w0QnFTyEgGyGxoCV
Gsdmei9Ze7prcjWYeCBbDuhCzSKye9ZO3NvO66JnXUTOGBRDGAeVYTwlf8wEHrTr6J+foe24m/DH
yhUmot5P6odZMkRYfXWUgKfSDn7bHmA8zbsXoIBgk141d7tLHOkxIOsnuNshz3jgrp+ZK19O7/8+
h3MnMtmDl8rGTDg/dugx6Ij9ZrDpWcVZEKOFnY5JCCbGRgf4IoKmI9/iFUgQLx8Q8F2em86jXTux
zgiqRZNObEHKWDnT7Q3RPXH3w8v8B8ab544rHB4TE+vc2XQAdY+OwytDaJYUm3WGskVKwcTONU0A
wj1tdprqNTMeCgbgiqSOz8h3XurZCHRx8MihkQTMucvqS3Fiv7m8WGvj3esjlhYoJgzXDxrTdadQ
f9hhffCrYI1giyMmvbDJz+rOa6de5OwDxLZyCKRh5hC6O9HbR0XmwmeSVmN1Ta9dV7bkQDsVhglt
Ib5PfTHwhz5Jv63H+g8cejofkbx0faAtOoREFQuDOhT99a3x9VZy+4z1TI30b6cmsYx/hUFW/PDh
HMneHt1OrN5o6+l5RII9xeVo++twVLKnSXUzU0o0XZJtWHgPAB8Fmuf7V1UvPAZFO/nVDfcQxs0S
rZ7/KJEcbfTy4v1PDD+ZVBKh02ctbKEgHROB0vpgMGjfv2C+//OiaPokwEicbC9zLihtMg+kJBys
HLet8XiBmCvbxBBV9xcbOgDjJIwmdplGveuz38u4nxtP3foZAhMiXZzXuP2/hsVPPCHYZ+bWsEwp
rv29BHgKNAnrxImKmq2mM5GUKOOkIfwa/qnIJ50EPOyK067pe++3rSEtW4lDg7sKkF0bRgO9ToVZ
/DemV/FrCxI/ZS8MDDjJ0ginui6j0QBzdw12AicbXEfAD7sS6TsTyOOKux2e3LwN3hgIcBmo6hAU
T2Km+xqAHT2q1KNGz4QiUlhWWBiTZfDKuMMufQZ0wBFBSzTXpLFiipYDnQYE89UCgQaUGNqIdI3l
1CJpw/EFZQX9cRQC+AO3qV21PbtV5qduV1yYWDOZuSse8BSus+LAzA0wf2HxaUIht7BSSqSjeZzb
QFRcUk8I5XK+A5mugXxB931o7lJoyDNsmjU9ObGruqH5YqPZGAH6j8NVdcd3yuNtLU5xrdcVAP2K
HNAteWBYoO/m2igr61DIkxls6ZGVv234GssUs8a7RRxw8NaULhY3pCXp52Poah2v7xTf3bhwqJrJ
LgItU4xUozRYUrCC3SG/XJMq1p31y1rFxItJBGnnk2OuqSZrbDnHXOaRdBIHcR/qYJHlLiG3ooaD
zMlOMF89L8IlA7Nk3DVDsTIHTObSNYYcK41m8gOX3wErap5+6KOEv2JEeioUYzd+wMY+8zZFOUdb
4EqK5163WugI0auR0LgvJars2IOyZfx8l3qE4tdJPxx4Hqpl189rZ4Ccyh1Z5UlMMJDOUe/MHyja
IWt7VVEntSneqhSd/z30FLcn6zrdUq5VE9t0qgF9uX2ZcfR5QofBSCX+VLuuJQDg5MaxVKcfukRo
36mYAMtUWM3yvNoUt5KG/X85pAzQMWQhsapQaaWwCPwc+OQsJ0arSzW6/OnsIGw/6RGQDfIBs3m8
J5grHIfNwpO1Br3tiQL3x4Rf6svpEGIuO7q/rFSOAchrL31Lns9aSBMBIMI4cd46DC7Dui0tcthZ
uN2CdP4mkg6ccFo206bYQZiuMu8ka0DIa1grqZgUJXWrpNnskEvAPXp1wwUBRdOEFnw0yJRepYnK
7IugSfTS8bHte0VJZ5ReSbyK3gWoRP7WeA3UlpTHH42w0dsqjI3brL1pP7GbKC8Xk3lEEDeA5byN
2dgn/TjjC9xlQi6b350+ErUxNRx70RWE0FruUgAhY7dW8vXT9YiHmQUzyB482nq/eN/s1+rphoUw
3FD7xmt2RxoOHz7xDjKQI0EBd4rMquevkU9ZHAoiA/W9D3X30e1UzOIyyMxRylL52GjyZomVqim9
JHfc21DjxWpAZ+3sgCvfZszOFKdZZ2lVSoSOogUyCOmI2ZLSPl73YJMLBYgqcGnpUI79TDuXETGe
u3/loZ/HIb+v6pdFmBTmWTYuqUcUGxM/Z07NPIfCVUVO+jIJpwzGDA4mJYq9aVTs3p9dRttSKMQG
IfDFe0gTLyOgWAfS/hQNvfu87aLzMBaamcvEFUEP4xs1itbFCbUY2Xr7tKg+coAQ0hXeWy71Bj6i
T9OsKeDUsLJQqN9Od9y9zcCp/XJ5uza69p6IeNLYo3DNGjxNLDmvjzRS1eZUnkpyVtxemWDarwAH
vXb7r7U23XKlNokQHIqufEDS93xkfbC8cQs9sivk4emaZI3EYNAtd1T/qbmaqSxKmdmHQkhxkC61
dYxsRKvkHoyJwRBbsrcs19xtbU9M21lhfXMt4t1cOZY62KcihLMYxzDzNkW7OncLFQirQg4h3H+b
kx7BSImOQ5izaYBKZjnMSJ/1HYyZVxXAPaUmjF/d7vxgIw+RUs163x5HBccucttSonWd0f/iBuN+
W3nbKNefGXTkemOcQVEem+o/FrhtMQhSFmeGXVW9vskdA70p9NjUJdLtsrMM4/MqDHB2vnk4mtJM
x6e5lMSl6Y82E4Ani3vbaV64epahiFiMEHxjXgmJTu8IZ7JYHYvNSR4sq4X7gE18a5kAYkb5I7ZW
wb178GYe+Jq+n7ntNaI1LwrmLchnA3KMsff0S4ouc34/zAvRGNCmsohRCsz5DbUxB5zmQWAOYVZ4
MPMIVrE5BJJfTB5pL1CVKQ3Mt9nFX8RwC6+Z8WJGf6xEb3eL6Tyz6Iepqod91M4RB7wo9FWBtQIM
BVRtVzobYxILpZ58kR8oULwT9/YQklIdJF6NPiW5TezA0/4ntmg6njZe5+n+DNLkMhi5zkm0ONeQ
bxu+Z1wfCjDxCuWHmGz++85fzPyzr+0JzkpYoNwHzoGFuB0AHOOrq1YDHAzXxDoYAwp/Pg0LkG/e
eDEdRNsQv7efjlL1g4O8xTRC58MQcFOst9O/qcupa2dv0QfLmu0VCV2oPd9wG8xgcx9Kp+LoSH5v
6ctc1yETGFz2OQnF8Q40R63FzYuV+WUc+0I0CPCRE2VsBaOqGp0EZuPnjTEIjTP6k3Sga3+oCPHj
dcBTwAts1dHjkRn3mShruZZDsBECw0CBkcW8kiXEowEbgkV7JmzzycAFwepz8/NnYSCr5fHJEX8y
Zf3wvoEJjLvsVk7dz/viv/JcoE2OVr5lPTuti1IhFUx0kPpGwpC7ydMrhGY2g8zqsg7EDU9VIf+4
RCx7DCT29MNKsfHNN2IRWxGZwG0Q9ro/+xbQbXx8Rm1CFGi5yBBOMwWxAbjYfG58C/10UuVdusfM
yIl9QrX6yNsa0eEZe/OpNn54aXpXDY/BQJFcWEfk8rU8TleaeAyWXwS7HTxVv7sKDpV8w2RlvS/D
He7eiVTjRTAat901JJejtgkFoA7XvG9yw1UTNfCGecXGTXoTF2au8aComrcrZa33OriNAnrxZbRa
9Z9IQ0Qi0jd9wxoyHHPNIF6dWxYe4aGqQOZefdOgkIOBoGCLg6SjMOfc/ZcQa4iFxQ67jXIa38jq
xnXtYzBtj1wjYRYLEHt7eaKcjb15FwdTYk0Ro32yzk2vPK6L2vV8RnjxRUgj5+4j2F1/oHUn/i4g
19F4PpyMzoJEFjr+bGTdcKn8F27IHLL647IbFn6SIhYD3Wwi6La8uPRXpf8HLLJzt6HOeKGmD+8E
y7qsObetoH/yiShz5QmonwoYFIEW5hqnhJN0C3ZWupjp9PL3/YUUwOHQpcvNmDQIXAinUtLHdEzh
fuAq8BSn3g1OXJfR3utmFO3FRn/G+njU933rlB4scC5IN7mP99AvGDDMDcsuoliGPrZGBDOhJ2Mb
HT+rCKWzYnxBLpvu+wq8RUP7Fn64p/dLt7VgXWoK9iOCyVobuQH45+m2Cr02+EiZIYmb3OsLpaKI
gWPbYM+JwTWL50wu1337jLTrpJ1OOwwl7p1AWCw1qV6K/Q0VubO1xxkYXEfd6zBl5LPZGMcHVJjN
I+pYkecovc/HsLk2+VbvtojHQO3uvBb+IkrTMqp46+B75Ev/EipWTEZoXPv77fsPpDFXdI2yvu2d
mHtZuJaWj1Ik79XxIlp9U/atY4IF85JnyN4WbgPFhpMrTk5bIk9jd/mNvvM0dQmFseDn0nr5HiRX
Pg0EXOgFWn4q+eVUFIYN0lG7RSuV3Wm3FFyLddG2eKiyeXm14LmLCGgc4auzhua0SYXRi8FF8v4Q
qmwcoqSrvOVuA9n5m2X4Zw2iClmcRP499lP9Y/BU4EgCMZ8Y3nHMqk792clZ5W4uqfVFbZqTnPND
PaChr8A1ZMwrEJ0mTJTqwpayTzUk0EaKVO3bSn+qhwkstHZZQ7NhNwcM2VYNRnXSU5FDodskOtK3
ek01N0uez8XoBrBi9tNStN2KKjjiDcgCOdVrJdZvxKNCs+x6Z9pfFjMH2b27EyJOs247tGOCS3c5
mI9pO+inGYtBZ7ogQDQClaETxV4W2vEROZNDvpCwMVFXXL6OUFab19h5NTjPR1iRPaXpJ49gBAzU
Sln3KpOR2mK/qShEpQhpVL7oMSgycFqOBaDMZkXs9vy79ppdP4qECxJC8L7r4tnWEfYvs+1adwYl
Smuqit8gFRQsjcjmC4EAaGap22RzVbhxuhEQfJ1nW66a5bDZC5vQ1iHc5Whx4rhnp7JUPLRtd8uT
ph4fzg1EbFo0qPJgQOp3/ZKDMA0oaNem7QaBh6ZZ2TJMpzlCszO3Ka+FyyUz0uHxOvBN4RWqtmfQ
mtJ5mPwCwi5PT9B61ERoSvl/FeH2URwZXrF9kvOTUBbg74Qq4iumg7ace1dnEyveIGK+D7wp3cdW
b6C05gZqDuaHI33WUaNixLaVCut8dsv9EymL4roMGH0ukZdKxB515xANykBKiyhNXOmk7V5LKvl+
HH5t1YCsgm3bLNyWEyhsnRTgZTGqPg8zFbqrXLnCDoV6fSurlWk3XbMorzHzLbSon4ILmx2HykOd
1wEdU1SV3StzrkIjkKk91Pzto2B8tLCKxRUCOyseZQnzEDnnw6mjXEJpN4yzEsy5P8IZCP8hAmER
dBdxhQ1Z2ywoFUt5PkfLkhJvanqV2O1EUmZSDu5RHd3j44NbiLzyp8gYUEyScbpk2yv7I6x3xybg
ecypsNOjiHoJ9/O5crv3Fk4B9Ij/xDVccB5pMeLYbWo9eX/1tsLfHv+7vWJIVUettQzPjpHI796j
c+zMCsHNfUyp5TL3eSNjawdvBGBqMjlCetcGtq5fcY1ylnB5mXUVj0enftXeRyIpV6CAbzDt25fQ
zeTJeGA+kKgcVLxXsPJWIQE1Wgte3jqSa8Z7bk8XjEKPihMeb+aMWGcB1CfSSPqhJ4SO8P1Ft9fR
sfwtijoS/jvOdjSXW7eKKUH4PcdEPArtyjv99mTgUFd++97GrKotNyy0enwll/49HszpEHwSZ5ch
MNL+HXA+vscvSyDPfEipR22wq/W5P4N8A/6SWAQJXbTJCnN1OCeCjUU/r873f6tvNIfQh4pVq9AH
5t2JKznB1eF6tma4vGp+ikQwvn6kuV1v7mH+9k7rRP+eleu+iLRiKSqIp8nxIKkFJauxx9xLn2en
0+e5/pmp6Q99XWaJ8oNZwh8rlzS5MRuc+5SRTWNkmr7rdy4CL9p5DN3P0ur+VZVRanfRordBu6hV
Z9LASNiOPp+7mmIXhlDILHvTEP617fBuyXX+ww6IBd4d0PWLcSnmI548a+ixendC30lzmLnF+j52
gEEWnIobtSqJKBu2kCWmwmeoj951u5S0GzqRVWpva1mQMEDN2Xvqg0uqSoEgaeeKAYbT1XrB6yKi
MJpb6SIt/RcOTL7/3YhT1ykQXr/iilr12LwLl7vd6RRMY/Px1wNaQ4FYXdHObuvjTidgS8ayvM3W
krswACEFA8dlHnU3e65NK8ENr/+5Q7FG24pRKbcfrq2Eu7PUaUW39Bs4wqMlKgiRJQPGNvCT4isT
HH6mCCXXRej95hfQXLMWbvLp6+iwXqhdqZwJYkImlmR0PT9PPkfpKgVu+0JhXRySxoIaC2+zXoY1
YiD2U5QOdiZXAUHJHD5yGnLRIBopdSxnEMPm5tc0B3swoC7bgNFY+AB7eKD9yAV/eUFJjFMIyUhN
Rm4PGVcg7aSpLUK8paxyKsMsSFdTtG3jvnx2oiQH9pzz1W8hX6VrrYi6F1O6kUJQacD07UIRhclU
E2Tkg7LFpMYqIwNOA7Fci7Ivwl3QzzRbhXGi+l8cX6XT/OKnBztFHmYjXNauZgLRygcIwE6pJCh9
7abwOEdu+o0l4mM7JrJNT2MBb+Lu4/9pnn/pWR9afDE2+aIpbF6kvCzWKA9IXQ++qO/zyAUmlAr2
vdaQs2MMRUleALDpnz+j1UVjCikoQpOvYwMPMbpL2hnMFPsjegGYteS/DyhjIjI0iYAAyqBjxXop
VXbTRHEMHSWmZM+GcLdGZCditUH/tlFydMSv+d2Mx/QQ4K5UcXcRsLWkaxRu695tcLZa5IfH52B9
s6QApiIhHkEAq+Jnhk97JDnEdjGa0EjOQVAylejvp0FLJCjTcs1I/sCvDzq46eiHDRllseGSA0GO
iRzQQD/8V6ddVl1jiFWCvcUdRvKWT7kPtbLw9/rziPht1tMFInvODHQQba2SGb7OZ4yHe6mgTMWd
Hd5OnHjjr6saMwmpyFlP+RD0MvprFPvH+mtu8qUJk/VTqmRlKpUub8zaHIOg+meszr4ASvZ79xmv
nkb0uHL4uCYvh2FAhWOJI6Sxo8BY4D/RQkCmLixyGFztXOsLGpG90Pzol+z+cpEbwEtXjwC3Agfy
ekpb8qCohsYxKbskiF9pkyD7VPUGwW+Q5WeZGQq04NTIu5371qi03PcIqmQbEC1vOtQHkCyln3p/
RX4esQZq1G3pzt6GCr/gwlJeuM8jBIoO0/SkLOudqGBKEFarZGRvvTIIDC+ZRVz4kc1iC5wKj3X7
46YtGuOfzqON4LXP+/BkuFqzLBZPJMFv+BqeDT2j2R1F+Wb46RTtl+B2XVDSx+zOWyMJ+THYnJgS
Haz8hUnJyYzlxsv1JeHhK2njMqa7b+Ti4gDTYxqz34roE8af6oIGWqGKwkAs5eKzYI9YfJTRu893
38zBbLm9qJ1pvXhpfhjW4kOnOUggW1mewQs33/k7c909reQAVun5H3kLka8nRIA0PK0NcFz1YqCc
n5IEv3ynsbDu00An7kBeFAhfHoDKtLkQaBeHgMAaZ+o88TKkS44KAih6Ckm0jKZ7j+NrMpWyeUjV
hY4J9XIAmWpPvEPucOBr4RCGCkiBBYfoZr8bEGBwdxjYZMCietTu5aT9q81ZvMj5rXo+iEOTIccV
GePtAq5UnWvGLVAHtJc7nlQorH80KJfe+/7Gdw3IpOyBSn5ZcGJXgepqT2YCP2pHHm+0u8Hd01s7
02f3VhOSbS36TLU3mvje1tMGEV1qCkNvhMKuf2fYT1zTMSRgX5sEbLpwm+/W1WEsLZP9sZx5yZbA
i+q2AXLJsHE3SIW601n2V+PjyYGoBK6FXCzEFobnN9ivPOoCxxJdw3J88eEC1Fv7mnVtuOHoAzWG
o3x4fEfk0klQByYwRb0LUOmG+vTjsaHwq+fvQYNOPYip4CscI4ugIMdZVl+sYEX38MF/AV7RYYoC
c1VxcS0ePcqmVB3e/5npmBu/nK6UieE5hlohH7xigZOuqRcwrAnaZTzH6ZaAPqcEQ1V6kx5CqkSh
nEbtPyZ7dgVxOQqP3qmmA3J846VC7ibsU0D7ecY+LpJSqzJ7Omd/VQk7Jq5ka6MsgsXEflCJ4Xu3
ywpppJDy4SoEjuNB4Vy22dCr1W5ebs520XO//IdjCCtw8lXvOTEzoE1mzwp0evz6icIK/sIFM3+K
ZjE+NpcudpwdPO05hPsS8CIy8ooaaR5zztTdXQeHVopHIrY+S9a3lG1vrL3LpoOwlyL40wRvJMEL
iT9Tzf4UbO+zbHPQnjLRyDWcjt4XsKVqJ7bKDapuyS83K9PnlooZ47El8wn7NUt5kpdA8MrQrk7Q
VPPn8IApMUKo5YMU+yDFtbY5eQruA7xjG9js8+95y+EErfiIV52WQzBd6ApZtgMcTMqKKkCCUV4t
dIW/NN5RKusGG8m6vbmvVD8N7t5K3gqcY1sDqOkLK3UbBIQFKE45Yh5S639teEAtRwxr1JivnbVN
xBMpZAc6oCBlAe/bAEaFjg7M6d9YhBmz84nqvkAdh6Pt0HLVI6v4oWvFtnL6OIKZLxkbTGJmnrZh
2t/3eGMK4jRQsg/4igBoXK8oQzLWXIaI9zXCsRLi1Rog91dnN33SEqmiJP3EsDqI8EQ4pYmQl8Q0
NAKut06lV3jfM5lMgnhgCTGSq4X3KQPG5W2q0GHohv53OV0koEm0hE6SdypVE0DtB/c/fzEeRFuz
sbtw6iUmU9Cv6DGnxOro7vMcGTyFd0SSKOaVS9F11LHnD+PAixYXxzVvRSDvsyVil5wt375Nb/0L
qrzCyAxX8MeXzveRlOl5FsBKeAhF9JpgbKfDpaZK7hg8O+PhNLuVGWEPdrytqG4297g5B894cC/w
C0yhPR4Q8w9Sbr1XFy+SsNoieSFiK2bEwFYdDwUxxgAQBvTjBjw60XRLlSlZtWHwjZ3OWNQXh+8q
CiX2KdTeZGGLlJNxHXVQp3Rwnzmpoa5emy1jC6QJ9zoy4CwzZADdhQFXAbm3tKhmhWukXQInilsD
rg6i5khvGgMVrvhLMw1Fp2csZxWsp2oMzYjp/0dadvU40MNf7ApJEGzrTLTi+3chHu4sMJ/LSJsZ
83yKotWvqLKd8NJT1+2fGZm6zPrd68ZkdTPbk787KLJnilTS8Egnaf7rkJeoQapoyIUr5+nn1Zsq
lzAJOXeJfhXKN+PeB5JHcxt8H1n0DrPiEg/FvCXkKQToEkvO8UTaatEZfs1t/nSzfKOl3cm7tAE3
AHhoO+7Ssaw8pcaJTGW8vFnJhZOaGdgX4YBE00VLWU+zJMsCTQrivF+0z2hnF8UerQhAm7JdeVJ3
QEOoadNO56L0ZUDkjco2tirUyUWSmiqfu9dc2jE4f5PwSH+I8AsrH9ATNfsI6ckau/UWmyTh3Aan
MmeKAWkSQw0Y9ouE90j4vwFnBkljrYEG12gW5vdcYKuEUExLYK7bDXcyxgRVt9F6dT5RrDes73dC
5Xqm/is7msyoyMdenzzMCGQgZbFHO9TfbwkXaWz0267Dtj7uluS56aX/uJMzmMMKcyK8LpTkGxGm
Wg6zsekYlf5o5f8jbXhiCB8peRkgHVdzmNSscoSLvsZN0gB67zeBn7LNz1jv3kenei1RWRMOYCA8
jbsXF5F4UH+rPx2W7tl7stmChq0u9IOxxZobe7K1KLkyl+vWklVk3GnYjOVYI8SvIMnATJNx4ly9
oP3J+TsL8X42fDDrfPWb+8dINQrqvunnSQASMkh02eVjB3Qrp3gGh5ZqdlYNEFIo7/kRZXp4379q
cITYAuZXtCmVhUCCYPIYnYPuxk3S8Vj1IrefMKJfWlZQ84MRGRGI1OhPhI0hlXw8QjMe6wgKuyET
UnF/fuppkvYJftYDbIpWe8A2WJJGDhLaYc6+oUNWO+uZMlwLWuyzh4whzw4HpNmNmZZBQeHBdf5P
Xxf87q77GKazXH92d2BE0yv3bJsSU2N8QU2NRon3VDxhaRTk8Lsbe3aJUK5FEnvtNyFJ3raObGWU
lg93GbpTZ27yNLt5NewakTPDVdcVMZM8wtvQAJo5JevoIQ68r5wHiIb6QnmhHq4g4wRmVBpnzssF
WUPJMm48to3FVAGB5M8peMl9Q/RZ2YRKMrUPoNeUApUMsn5WMCE7548NfKgPAmDP2cU0EYN2zICg
U0dYuPC5wsXglPacVT/toL97bwjHn4yghZ/iJ0p2ajZT9i8IIknYonpdf7jUO4KF/LKv+ih7K3Jd
kP+Nh7m95RLC6p+0Ow/xsW0h/Y7m6YJUveBnymmyAQRSjx3MJtMWKWcPmXpfIYObAXw8e6FrMa7j
DNUC/o3hvg02KZRwW0pdkdhjgPiZ4HYV5bVICsAuaun4feklADPi5qs0Cdt3
`protect end_protected
