`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73904)
`protect data_block
nvtpb80h2zEjySd0ZXxV+xKxp2Wi43NKCupDeRYb9uyxQD8bifoBH5MhCGnCzN+NIqXa0vDCfIXt
zIxFTUQnrzoBmc7tHTCEOsaCG1cEg3cLbk2tDp1la0FaS2D+19BXg+LLhKluFp54ewzlSu2CCEa1
9F1CNwUpxlPYYiBJxcxfIrhY0Sqd2THT/OkoPmgFKQjYYYO4Tv/oTZVVqphEmb3ptByJWU90e8WB
Fc3vkY0MK3y0a8fl0uCYXetE2fWOnpenmDmGNxJFK2b93kDe3qcEWmptfaoWr7RTnhmIivX0a64x
Rey47N63uxb9ts9p0PUV0+t79aIOU9B9fRJgD3VubX9P8+eHhEFaO3CnaXElqbjIyypNCmH+lDhg
uq6gYJRqsfQQKJhd3Qi2yxtRsvPYcRXRz54O7+HI3QLPKLWNmHqr4QYtyTQ67eKNcmOIIHB3phQh
rCKyYPyo8f5A3rr3g5fmm76ZquJyDPMGKS6cuVYxXkV6tI6BOVcAEM2r2wS1zzGWnHIykHA5o533
gOP6JoVXHKNL2DTMisKgTjttyd9Pc1oOoA4naxacZ+8Yv77rAnbDC8SQjJg6OyWuQfg3j35nAAI5
kQqiWJFRprYxKVCoWrHrYHNXtjMjTTwir8yt/ZFkdByONmB3VZ0/hO0qjpBN1BhBjq6cZzkVEqta
P9yPnXl/bBfbsVB4GqjbezTGGqwpo+cWL7BhaK3aCnvrJfBh6cNkdU37wO9q3jKMBRmXXJwPAnrA
NdfVF8ATEwZNuBwZWBGWXeCiYbOIvLifJe2qSU7fj7PJqhiod00TPTpcbGtVHZO8UCfCv7dTUZ4w
qAmwLqg+B0+MhIxVIHWlYOoV69DPmAUb0M4Em1wMTZ37zRH+B59j8Zg12vnS3iBP6OiIs6+e0A73
XezB+3rsQBhAWc+jSJo3zdOLEhWnN/wJzHmw+DAqjepROilgBnzvaUY1AakBWTwTB2yzovTlVefl
tS3FM+61roPDN0rc5vK8LVCBd7QiMbrahW7VUx4BqXpNfpozdfAzc7jmvx5LzyzpNNa8iY2XTlb5
rwgJCUfkQOETCXAl3m8PVN1WkuRAwIjtugKusrP2JS3NP9sywgAxYSy3EMeXU40Y6ficEEgqc9YO
tflw6/p1Ww7CTyf5wSRaxQXIqrxewqyXP7NIUUJVslOWD+s5z1C651qPzzJ6hpoEBEUAfMlfmKE6
iudoZQFG4iOLmE1TzMDknwS2x8moDU48Pn2J4h2yDRaE9U49oFbmztdjqCWIIbaouBCits/4ZhkL
UeA5WlbH8Ud4bXGfgp2XH0TLTmU0ZDxL/W6FBQm4l9m7COrTNxg0fwz1hliXzS2KgptNPJhHnKC7
2ZCrWRsEfb3rOBCm34UNTwLKsck0QJB82fZ0vQDdHWYthpQ9ReXubhPfIdyKAHvCCFcvSGpPStCI
XpvYWDV9LfggpPavZA9aZW0ENSvgiuZauaKpkoue4mjwg5/HrlhiexcAmMyGAd8KsA9B//pkRc1e
0GPbsBPaTkcygEVotE1Snj2zAJWDnQLElwMEzsPfqukJchVcnU4fp5C0q6X3YWV/MLz7xbKG7HsG
8PpBh7cU6OutslPQUBgZdg0VGeqPz8OiEvOheKdBP1qIjoQ3Eo4H9dmMy50Ltgr43ohO5faUiZwQ
zBjSH4TuMgOCdwGUQEVoRSUhuLRKBtY42jK6kbV6s2U2K0hHYty6kq50EdGTC7g/NiaieZa8szKG
PaUNmAEd2Jo0dEchzqJDjzF6lEzA9BMRlnRPr/OJ/gsnzFC0bnzlPtXBM1QxBlEKNaJB2VdM5MSO
Kba2/xcwb4aqHzvBRVhSe/k7KkRq1q58H17oi92z+ayl6GJgdjFiiKIQF6wdAwwxSJRnAYmbO/04
St1DbPkWY/yEpUhTGAqmiDVl9pdaKlfR/SSoAD+PA6f87JYJj+q3G09cyrAZaK4ovDS/yw1T3lG4
LZUWOwOqjH8wP+rXs38tmRiqzqa1LmnebDrfdoRs8OL8ZEsY5EP28ZB+3mCuy0IwkNNqTcWp3Z9Z
l6arl2SB2mb1HZx7kVDHwkF+qOus586PabVzeLhlu+OxdagX2DOCyc1biyd6arSRBf6hy9piIv0m
G7jkpM3k9T91uWDgK5NHfDaESoRPuRAWNReCrxo10R0GZpeh6aWCmpXESrr+g/1S+YSI0Xv693K+
pJiZ4Fo0xObPFxcVwz4dAfY5c+ITfUFeVwUBM4CWiKIQ2cQC1FB03y2nkVotojYGJQcY7SRLL29H
cfuRO90solsZK2kOzbDUnzwpT13Uui7q1GvQEqg2yQAiExbNbQ9EzZAwEMeikomRyxm3ZUu11J3Y
y+MmnijUE9Q7y/OhKp36WvCpD0wzHLrKICnJg0jo5DhBd0llpFezJWzq6epHM6vTrWOHXuXnlZFv
2E6i2q4UiBMdfPKaShntJO6s94q0IjZ2kTqUzOP7UdpF4XOYnmUd5GUXS7zoAzJ8GmlE+HdvpntP
eRGVDcJMfu1n1vL/lpf93gxPGPcuMwTQ1qxD5NThaQzzcbioUnWG78RcfSkiHQzDWxW25z2WZ6pb
4z1praZ9MGX5WLaGSZz9EoWJ3AlUrz7NAIfwrMTTpXZSMAc3n33c/JgK+8hThccrYJvprnZcu5go
NcMX/vatpg9g2OaBvFdXRGCAWWQpuv+mlUrejPre3Og1c04/cxJROq0cEONhsUr+OuTlTh3+pKay
pJxFNEZTH9dKzAl2a+drCKd+8+MOide7s3kxlGBEZAlP6Md4nkjL1gOfr0Z8uf0qhhyEnIYoyFfi
1z0r4YT3IIcDGhdsGqtgcE5n4gIQ/IGF7Ft75/gkBzu4InXtmzi+asPX+beI1Dq22gtjsaPeV4SX
OnvsvHO2JgOzeSOQJryzRfn68ENUohdUBUb2Ym00VSQrdc8E6y1Up1jkakMjv+vhrKqHeEQ8WEHe
D/9wXz1NxwgnSZvu/l50i6Zh1PsM9pM62su8CbtVHnfdR5LZ3pD/N1blTf/QOMwIpB/bTCmd0Aaj
6Xc0v4U1bveyqqWOiozMu59gcdcodxXPQzqtuEPBRgXIJGGpfp7LJoRxz1/h3Osfu3+B24yOOk5F
UOTEHMxhpb1PBLcwaodVWwCSijOVywp1LivL7CQndMP0EgU8FnvblBlrEsDsI5iMVeROcD/VVo89
xg4iYYylz6f1JwO764r1H0CdildniuquL7KoQTQLRaS0i4Ndzy1wOIN4Z/MjqYCKlnuPU9rRzOfg
Gg5vl4mnhoJgRcEf5+u+TNkjiqMIOv7LZ21YpqCaGsP+M045vpG/YNrzwjjaUnxoySXr6xHTVh5M
KkLQFQRy8mFiCeenBUUyu3YmrUhsl/ZJOQdfK0osTHOIdazWzDv2+reAttIBxTkc3zsrhUueOv/x
XaVtWmAAKATxBqPioYx8PB95y7QP6h7OBKelQgSwqWNqtkml0nbKYPKu4e1vT0gcT0Rsj6FU1ihd
V7cNm4/b026l1adQSQmFbOYzmLQXbZ9Q2xwefuLMwyKYxjtDS72ghv2qFa8HJcJElwwbwu4W7jOl
sDH4LAByVRjoZy9d+GEnYCZPcOwWQsHm1M5GLsrAuwpqi6QWmv87umE0QCPR3Pt9J6zHBbPopMYI
ILnE/A5mUjpzc/wD7o7SsYTmyGL57X8sLGSNNWFC8VuEFyuaCSsrOnWEbVWV7vbNw+dxgy5XGkUf
3yEoZvyQGhPmjQBe65U6BrXN/5lFM2hns+sCPawnBlW06okHDp9DjRPw7vUr2Ncf5vwD0o2gmIW1
ytz4OFWEkBA8KZC8THel04H4kwjKN4pl/NhYBUuVr0t+0pJOoNYlgQsMpWcpMdbB4QtJ2K99kxIh
eRe40+56jNnN5JQ9c2wDmIak80Hq9n6NkjBo56ymKd14uLtQ5Meg6s5RKkG1NP9e3BIv4CNPq0ed
BgQrdODfj0o/fIrxq8sJmKNNtwM83adHUubm6NK3S1BW0Wuutg1uLqvyHwn3wUtxgVYm2CCGQp2J
2/v+9sTSwTgemWu9n0/3sIJVgDSC/txrEpqCrYzJ/Hbp+wh5SmcROikSKpQsB+y2rf0mJP73MZjv
q6u38UR8cffsCAZVM26Lhg9pCK2GZWt7LgkJ22rmmdxkKmTUMy8yjcw5kb22pTWULWVyl8lf2fcq
viU4vMOhkEOe5/b9noHlZ45rU73shCn8dLVPTunKeWauFB1d1EpFbEpaJ0cQsPtm1b4a0PqESRQV
qlVn8MMVD/XUa5fQLYj3wm+jODO8n1a5aMhH/OxD6X4YfLFcIHscBm73RNDnP4ui6oHmoom5ssFd
36ytsJeNRlndOlNQi8H6huJ6FsiPxtsdwnJ5mO2/0X6OMkvyOWRljjJN9HEiD/XopWAXCFKa2lFb
NJY8p5ElkaOTYC0q3vC2+21v1dYJEcrt8J9iQuX7pwsp3JjEmpNOT38NEOvfjfwHE4/gqEPc0e+K
YWWDvUzyvFoSkiMUijlU2OV9utmZWhaS6wL761H+10WbUegyBnvAcxYiAgg6HEzonspiFBs0CEfc
TNqGuFfJMuumGIXsQo5zqWYzP9XOFZe2UkiVWwQ+4ti8KhAd8ZhnZkBmMu4CZfZ+sEvcRjs+EPrz
ZXI5dgOkibQCjNsCqqUGK9hrbXvCMHUhKoTOY4F9VEKCzBNrHMGI0Zppb5DkteM0sdlWMt1Ze+S5
f1ZruIFtBNAXhH+eWKzice8wxAWLnzM1FcGT9fLDBLnNFeUVrvg7Khzz2JZQ2H2zsWUOyzOsp54F
/OsCYXPgnCmU38EidOlqIffoXe/Ftip6LUN1cwR2lECRlfIXiFtIuFqg59xlHpcSPVJtWsIa2wUf
8D5KruF2ybgd2BmGYuD3wi9wOrB7Zlq6Cph3dW0nP2ojaQreHNqs9aV2ijufhNPapUcXrIFZc6o2
xvzC9OPDodkbMZ4tij/i1lWq6yxFVuDHcWNHw8WgqwSM+eLxTIXKHZds9ddYL01rJhepnOKFJTfP
RQXt8mstlLEnN5TqByYn3Hr1poClrwJ9WTci++b+kifCthaW5YAxTvWHSdwJFNrS4sniqo8JCcpo
MZ0t7ywBlTxto5zllbeVPwNPcwDdSBwxn+CFUJZrO4v7/3V9agsS40NrRyAZ//7vHYHzxFsKX0kI
Ytic9DZaU/wz8cktsHtSTVNCgwgTrNo6MjvBj7rmFuh9rvCBWJM9n15qPQHEiG1uvMq6tyw/f0NW
esmNnbVMB2ebxpOjcf+A3eni89qJgbJu5SOAMs0sGFILkBVN8f53QpzTvdV5Xy6R6ANN1gqIdRD/
uNb76Rtc3O6wIlNuG7LFC9px8xfpCGmRiBxOoVPfSwmiNbhT0rRS5pExsmyVOT7nm4nUSG/nsefW
4q9oPQlrJeEzp27pmFKtDkUikJnNlZ1rmn8oT+OLsb7ni0LhycZpBVakrIR7/YvWjL0AxetVf3Ed
Aj6gDkxvBDKacRyWcwRIbj8+YxHNUcJEUEQo8ADqOMp8z3zrGGoHEYxQkQd05QR1W+6RPjKtIKY9
SPHPDtu44cfr/1nE6ZuEDUFzy3CFl/Z767MK5xnEd63whWuIE/nspKuIzLPvJpf5/HH6j+jtAdpj
jYH6oFtvSocIy8kqmIKSGtB6kVV1isV78nU2GAmiCzOfhj2sGoa4eaAGC7ssCQmDp8aAegRqbRA3
Hc360xCm4t+SKAG1YfXNVSESeYW7yuyDghUInKoh3if+KRYIBZd3hwjRNngPaj0WSjEwCxwWN8A7
5zJJptEs7VXosFfZ6decpRUBCGk7ptj2lVqMZdGrVdcYeMccfETpYQtjxiGIYjfjkKNKu5C7nRZc
jAFMVpDdYmcRhztEic9xaDhg2pihS5GZDyxxTei/OmrXrMwbREB+GmLtU/jw4/BI1kfurk2mgXEa
bQqMTZnOTWlhffBu9v8fDKxMygBgXhg7CKEpCiv8SnNZb2Us/jlbrC2InFbq8XfGM001PpKAeSA3
Xa+3ZwQ7wTxUv9R+r/x2dTWRZqNcDVtda01PxYoYJDwMCeqIRVgCmrE1EF6+QV3XCxjALtWXFq/3
YE+iaixl+NgL081YrkEkOE/0n31LH73jalJwAJHPf1OuYAyR2rW/j8yjpv+w5Ru3fSYzhgUgWhZR
ipFJ8LMp4jrWTl6aJ2yuTRVxAxOTHyoa9gHfTVmKitLrKHbcS9MQM5efWDPjqN32ZFjc8GVi58Mb
EvjSvXSkcIFihsA/PMHDZis8zFdQTSggR9wSAIT3Im9hXh7Lt8T8rU/foA0gU3Ezg6MbiCbPSPDA
xz3iYcj8+kuXOoJg48Mu5NtMfKwzAo6jEDLNeke/MmrYZgVglkshP7/JSqA1U31tk76p55JIFV9J
iedl5bltpTWRfJjXtXdJg1kJgG4HKm7LYhbzD5+M5sl48nAqa4scJ0RG/cVdnz0QB6vx6jmUjV02
SKVZz06dgK9cwUSRyMIUvpQvEv/xARTCv7xTI0Jyw+mERCtb5C5OiFxu4XFwaske89yaOWgNs7WS
aoEsoBXzu4skuFyrHO2gzTekCiuNy3hoZWN5hLXfrp8c21a7ZOFA+pcqRiTV1o5XXCpwQjRmAF81
CcH6WPp7bPJQMpfYHC4OT70/DMrroFNT2VmrqdqMUOoOCpV+zWynfkROwo8h6eghRyTvERc6S14g
xwCuehsfL8wgVre1e7CR/zUx7xdoLsOOm9PS2SC3eSzpst6P4oviXZc8wS9kLzOt4rUIbOetEL4T
qY7p7ER6Q7wD9/x2/ldIS61nE6vhcZBht1QK4KAivEh4Zu/U5+JrF34Ljx1CQNJ1eif5TVpS9kiR
oaOzdu4eATKqL+u4dznrMIvvHzC6PqeCNL+FKJ0gIvZhRu8MPiPhfiLlTUbK9AN1eLFRNzF9S661
Ps3zj1b0h8/hfBwo6PKQ3Lq17sJivSD4LoJ3iN9/Qt+xtiF0nkSPk+Sfi6/MUPshXMzvPoG89wDi
zwE2fBtuy/UVnL48fvyAMZacPxMv7yg/0l8p7x2jdGMUn4OkajLtkmfC1Wqa04EVZObDuFU9dBsi
L/97THtqCYu9tYkZylm+JoMwJ8Q43eMK0yKRjWFVoFGW1uxczrsf7ig3fxnGsgcaogKWXiy4leqd
NjjSwxxVX6ED8qPkXQV1+oPNXtMW7fdhppeVEIbOXGlGGAETr9O8ubjGJIIiFZpq+LgJLftYyJ/a
rJr6P8pg+m2CP9SXLzwaLKXFIB9toQyMVTyajysMkhy8p34JrXF/DU7pKLNMhA5h5Q/loOpy8BwU
bFIsFRsgEYAZM//hBTzHi/EI8LBqlHC+PLuV60CbMio75wtQ9cVG+GVudV5RS2STxTqqk6c9ahls
dmf2MWHB5JZ1eP2KrjD0uj84nQZqUIoZIpVojjWFAGe33IJSm06Og8ul57KQtrRoHZ55DBmbWoo3
wPu55eVLu7tNL4W96crkGF963ESoVZSpFb/AeS1T8BPL4MPlWSYwSTMn+XrrWXRAe5N7d7VZSluF
hR18rrhAjyCAjmYfVx58txkCZ1Il4UWyY8rCRwFYfqm7mNyp/TFjNnzHmeT7+Fp7opgsi4+pvQha
Jsv9Uv/Ajps8WFPFoWGdRl4v7JtSnRiMDqtC0bssIetwR86uCiBvu4ndIhWUGUNUnS81gcRd1dYH
VTTXD471dgPRpdfnsPLT1ccsNqne4hkTQOuZwPumrPk3ZmSxYCjVGTJBSqCkCWcdGbr2/bMz2ZSe
Pc6QdxjC5RZOuyygrF1G2H9Szukc7QcmMkvkc3zSsbVD0Xw9073j1Vay4Bz1DuC91nx3GtPAqbva
mIXtXayi1n6hKa9c/rQAqhhbE/XzqHShLi9Bx9rummoIPeU9GTUqJbfD43BhT8nr+WPI03Zm7OWE
WbcEsUNbCOMuVWHQDSqhWcggZNeZstJSNeNWpMEfwhTrc88etKMs7svE12Z87JkwldXVIk/PDyLR
xfaggkn81aI2CqgJobqDDcwibG6x+EM4Faq73gNt/GrPd64/tr0wpRNu+DJjoj/NMHjXPHC3y93S
AtMLWc3sb48WD2EKdJgx0jl9RujqDDltua2jkPUiVvcnHbREYzoFu9E3w2jRzieNBozsE6kM1hL1
YKU6Zs3Ji9K6C5Ea5HjSU5YasSJhldOihN1hAGtLb0aUU71/qDg9TFGTgxZWOGqdUd/LmVOdulj0
omoBiXmixacKkqxPxYtE/lNKJhCTz0mCwbm1VWm7uklUQeDr+emb45hoMkWQw22ZA95Z8btCl7f8
yB6f5W6q4TSG0lR9gV/xAJZHvPWN+CJHbzAmx9tFLSJ4BKTS8u1YTWaPxZ+Lsr+dy4n0VjRv8yIS
D7gLXo5eGxDQvBlkFS78d5IqiaDh1LzMI+KOhMIVKZOggkDPzPUwtm0L+Kv3v+xtHx6sT/7HAS7U
87GZLHIAPpgnE9FkQZeEQFb+wSiLHcvjWTIFy655r40EMagZ5B3bKETFvhDKO081VWhpvO+bx61i
fxVqGVBr9n2jCy2XHmZiw/G0zFetYYObRYAEQwmYLJXkwe+KhEBgWhA4K7/RDfCIhXAMHRDrtuyj
o5WtoqPkIFHH4FUSU6xRBy7r+dJqC0psIP/nmnBhzdOyS6wDL+T3wlKQmS/BsgGhveiB/dkIOLv0
giZWZBwdPCAfi2UIsYMOg6kY2Q+rJ4vVIwzCAuqd6R64oRPh21oMrAFHGn9BORMDRuY1gjINow9p
2cq4j9Miqz6q1jKcxXnsfa0puQErIYiRKyfaVCAjVm6/MttiSiIjzHKnirguKfq4d7tENHUQx7T9
REnMDxYcam5TzZFK1/qy3K5OdH1kpkeNBCBtdFU6mF1qDVMjazLNl+s61MMxqzKq98eoRewlfW9s
ZJaK8y+PJn3duGD5MdSopmnhN9ng6DgHn4IsymYVic32mktSmF5FZfYdNjdSVJbybFmJqP7BV/5J
ygD7RrzhfwSwkBgnNMFxKfFtRRZU9HITQY3KF/boSZ/XC/cArTLQkt70QwOprkooXgW0wbLT8uVZ
z7s5dvumrnSH8BTbg1Kn+E5Jn2sSvL+XsehGug2RuurjsWPV6BeamkGcuJFKoQsOgoFdK+Bx67vm
hiJXcSkxONWftlyIP0mRBOhg5f00LoUf7tGajvQSXr8BNX2b/3hSWPLJewoqBlZcslk/Gf6P6Xqz
3AebNfU1UP92ckSCLR1iIXUER/dcmlKC5GYkLgEI2cJjAXeuo/AaDfyYJxIm/KyYp80ERGuF/2+H
4mCjZWwdanIYyMKJp3KiTtiij1lLb4mNjnWWzrx1ONnLUB9lFft/IscTqnNItrzOR8SQfDWyn50Q
vRs11s0UE3FhqWFwPjTWuW/vlLbcv6Ig+HF0duSUrQaxmVKQ9S7nrneUgtdKzfm/4rac5WKFkudw
+ddKijn5LoYBkk7vqy5Sbj9rsuhFhuGThT5k95x5pm0iYPFvMvD4o5jLinErMz3lpYNGr3OhKOFL
C089G/CLBN5+Fs0kYAbKmZ08IiqKkL6twdZrZLkgpmh5IAHJZ7DMh7w7YyeMP0K/71DOgIkSCLOM
VXihhDmtQPpD61T6w6X6ewk3m3ysOzf9IiXglSNTkZaNHulo+PRorHE9EgburD82fVbyASORsOHN
EtXlPCzAgdDeQXYZ7L5VEcloeyq3zllKRFtIea1CMyVOnne/d2f0TVXAvrPb6VZH/OqvL8ZNAJOJ
QdKiOmL//dV8dv0sCuAnCbCc24+SMJJUF0UhUx/o+sFv/zz6LmfZgc8+o+hOBKZRxD/uDaDlimp4
h7XAAkAhZRkf4odNcqm4AXPQa4SnnwxDq5kSa+E5JdGF1dNkH5c+fXtpQv0QgI4JvQ1k0F/bFD1t
92DVh0wIFqgZ9o+1F/H7ajwxsdfoeYQp2KSLvG+50OCzi8Enw2ghkbjD5tG+SFOO880ynqxR8O3i
pq1l2BRYkM4XQG6pGS8deoKLNjgdtQqWAQu7PY61oNet4ggxJGh0SZIVStqPRVNCNM/VTcWSbEgW
L7twuCGges8jXZTZhDqLrJoE0zErT+PtZGaCpEPAyrmgvhL3gCebV3SHTBLUhUR351OjEEx7s+Kx
wIvmvQvWbzEKdQLNWaxzJGgMGL4oVVQTxtpqDcAflt7986cKWrog2BqQOm8KSMlz6975mtUGWJ3A
M7Cj7SvYhxcng19yytxlkf/Y2Meen0zEV952SFrZx4UA0TRTgKs9pgDITguuS5QsizzRLPgG+N5l
6/B4eqaCmjqiug01p1mY9hp2kNIYWKuIAVe56fQyYjy9gWzEofoGIFDupQfTkxJdDr9HpSIRDFK/
5qKnfMFxfb38zyVvVrmKafckNuNkbf444gysVgIJwhId43KtMyuAvInli+RfB9nP/grByz5/ZZQy
SrRMyZwpXUoFmwpJHO8lwkyGmk/JNk+tU3rd2askorSHZLKCUymaduHQya9bPDBmsgNY6q5NsMub
AGUoIMIZfoeMZZsLUrTQjXxA8CwueDmALKjf8ggPvcYuIk+woEXlihRv06TivktEPdwfcFLXJ/zT
9GD9Tu2pein/v0CaaaCgfA5HjGzmld02ffND21+ZCXHKVFqEbcUqxLVJ8wfMfalxVZXJvGFKgvS0
mK6BMdmwzBwWwtguv3kDkaWt3YypEnFbh+KtNo1f3eQ5gSyFyfO/3xYLRufZSm3loKfFvf8okgAi
giS8/uA7GxK88tT5xA/EuVj1wa+ny3nyuzxZDiIlEOWn0OTI9zNurybj2WzNx3AOqrSa26F8yF0W
rGHmFODR8DHcJGJD62KCYXOnOa5i46thqDrZpF+q6CjuZQCNifXwtDt7sUhSy1YTVfhq1QqBy/QH
RYpISB3W33Jstovxk/s0dz1FUwuksZH6ZgMvImdubNpjXol27Sb4233IcFvcGiDUwGLzA64rCla+
m1uxgfxMAeHsLIIQ9pmnsXAJ35K9qpDq+IflaFx3fjQU6SF8VuJQ69lAw6S7P955KF9W0keygyN+
SOBRfM7sq7EwmCfP4WNKqFVVUV5kB5/bIOEWc2+8Q4/FUO5Np8vbFvyhkWZ2cvyjdAZq8+iog5U9
Vup1thmU2m/AKNjzzgps/w+mfWQrEJZwBo7XxqAM60AjVgeY5gJm1My0+NxBqkSZRR4D+o8ZFbwf
iCuKnbGky1HM3BtpbZ9y6WJIRoYEMw8Wr1fjoP7p6WbSl+Hdkc5s5GI6aEzZgceYtYBYg7oZ0GwX
z3vKXX/1t+VSqOahpOsAYB7AI2PBWX9UmxhqQt94S7DchLIaVdYtGsFGZfI8Nd/J8qXaPDeN+QXy
d+CWxFk6gUYEwez0EGfVOWBLSbR2nf5SAClPOXvInXAXfzm7ymiqvEtVniH0hwNXR+6MI4P4yJZQ
0IkJOJlIvNVcERU7fto/odMgufjx7vx/UOopswBFvehJ9sNoaBAJXrt08Yhdtu2iSwHUyocbk4M6
5ED0KeeEW39sbWcX2mU65pj/KW8rBMk5gb2E3pqdoBZ5AzDn3ZV6k6jJiBlnaa3MiQheyFPwU9yE
s23Q6+9E2UWziHf49HqY+trYqIOeHC2ucZB5K4MKmxM4+56FACxIighAknzGQ6ZKD7AQzT08kiQf
XE+wLF86xV7OYUknNB+KmCCZbMFSUpYc7yjn7J1DlwymNoA4f34d22gQzwbbckuKkXh3X9EcMRT8
SiFbIX+2DMiglcO7OtGTo+kbydJ9KhQmNw5HFUno3W7YdNEDTLKbpb1OMibOlbNXECoZQGnwujSt
VLbpkwRHUDT6Yom5CiCJMv5HvLdXHuraEEWKw/tpPGagsKqAO2uYmQFP+uq8p5xeAq6QhRT/QyDu
rhs9Wo59bD4t3glISyW8punQdx+GYKKrgoIba2hzrj2PMvTC7RF3r1t6YuEMxNWUL64CaFpxfQw9
tAYNa/frfUswQ7zcF6rCFEHEaxIdhEoS6jGpYp6dfww3r079k4q4KDpIxOB2qgnJxlSUwpAjDsLS
AgvB9XrGazHOM031UV6ABRPz7ibau4JLZ/LkMxSzTnuZH2eiEkmyU07ncn1zJSTgovDNlEYEvR9i
bi6edwfYKQoAO4plvlKTTaKo5dHTJs0BhWZIHqvIPh456mEM+evCOkqaz2O4Ay5St1zLa0ta26wa
HrWpiypsr317Y+KaV/Sp6Rd2Jjix2mn3RQA5y8/4tdI1gTTDfdxnGodbQE+W84T3XjWzZxInYIOD
wnWeAvb8EM7y6iFf7x2iOreA9I/ImhLoLsatRn1XwIZpIjzbB0tkzt30xUpvVWRi5O9g+Gb0JSDi
+EJJ89DeZsUjSh4FyvCI9VF2iLVqkqzhMsMcHfk1yKNlkaa+728YvW/L+F/2ILAq2HMmLCS2NP6/
TBTAT7/o3ZgmTdJ+DpeqCRJyh1OYffA/DdinOPT4/jyvmyVTWfMfn98JfyBTKJRBmaybM/in2rtF
3spC2Nqu7KFDhnagjcP77g3t+A8AVB6d//Kfgz8oFc+9hgt5DTXw7nuLYvRYvrLCEy644c16isYQ
OPbzOGzeVjGzGukDas9npraHh0DVGIQ5lxRLEXoYRGSWsCvCsWaITjx3PGtwBCLRc4/hgnA3iCun
wYy1GYROf0rkTN6O5Qhb0tQX6vpxI0gFQMs341/pjnLKAE8Na/ZaQWNQ/T3zLww6jbFfE7doEKmH
uTjOa+7Dsf0bKcj97B8AGL0QbqX/Ak3NGQTloITbSa6TBFQOLRJpvbgI8pX+OUhTALGASwiysuQH
r87S2VMl1Kl9xLegA317bcPpv5NuSUakVUrpDIPiFlr/Ie6WLvxRKK8Ycot7qxIHN8kNTdJ4Whtk
tXwne/gzH9n6UVoZtUW2lx3zmgqaNI4TrXf+RMksJpf9TbuG+6E0YVoyMBim/SRuLqsU3VmoUQhS
lSKOoZXB+FckeFbYlPCd7AaJusJVyt6q0bDa8gHNjRfJJ0R7LEPnSNX5KKAsZX251u60VWXZMLMS
c+7S9blbFbwMLMNdv+VSAPfXoliSpSbElsBrVWG8nN+Qpgn+FOdZgf/LvyC+zLT09T2g2C4pKHyb
QXPQM5DLWonXyb05wLsPgY3vHF0t+oT6Q7XaFMLXe/6vFg1vpW9BubYFsaZbhsp3yt09JKeTHMAk
fn5XrxJ0MhvbJrdJv553umdIWkjjgVBFzsVxjLUChT7DB3/bjoSsg8VtoRpUcH90qMvui3LWG60N
6cnruEYuIqqiStZNxQcXxLzlKLNPurEO3Xu8guP7NHTMtJOMhHiJZZ9lMA+9oJU40yY2jqJZjuqA
vwavIHFHxZgZbLjYbYMotauUHahhclwx8fGKRKDPgxSpiRNGkSilN5l/xKZrO4Wy9hUMb+201z0E
IneF8vdWa/ZAAv6xd1VqUJdpTY5JVMIFpuoDmi2AP5NDjtuMXSoT9RLDRnnhlI3OmNSiSl+RzIiD
E7xsaRAR05fFQNiul3lpm1edM51vC9/f9djdz7nyQ0ER1GVRf93zp9d9gVPcfw3Lv69h86Bafpo3
y/e/mqZQBJrV7s9Pn+o2Zi9+NEt/4tDYrxjEn8Myx6UefHrR/WfpovCMVWnxFhE7dT2EVshvQN3i
6oBHr8bJA1O1EJLY+80lQ8u0BAEPM/Ybj4f0rKoCR/DgnXVCsYjAcElk/W0y2FTlnS9VfwBjCyYD
G0aXtMpf28lEWDXHwyK6m+iNv0cJu+H3X6SZOzGCZL5+FMv6Kb03fyL1F1Cxr1pdLyY1ifQY/Rxd
PqmVbEgrC5FJ8esLAdOC9bgOHZOWFfJtHsesLp3I8Qg7CLiqDYzlYmZNX8zkPxHmpjTsuwUlnPyq
W8we4zUZf8galc8BD4TfmWHFJmBmStITZ3q7B8AVpYwPFpcNge4T7NvidsVhmCRHgtkqZm25sJOD
uMzcmPc6DcKtmBj/ub4L/i+o1uGLaAMmttrzElJBwyHNf9wA5lICVVo2UiCqyK+oC1ajiLEzJ6kd
ehZ6VbRY1b4teGfHAKtH+N6Nd+Br3y0d6OgmyfoH4keyFn4hVR/CDWwyxFaj/1h7n5gKTRZhj+9J
Mt87d4a5cajb0JifG6ypcc0iFQJL+zCPB5L/zSdb1oOX8qdsxq8WwaeSLggY08uQj1mVTc15nufe
UGrWcSXxP5avoRf4vk9qDh5cDnVXb2hazIqfPPSJc+18wCi+hjsBAI3GJFRYVPC7PH7Ajp6P+fpJ
YduELPaME3jKjtlGzPJTXLcf8AyUxROSXIugEOjZiJoA5SvsoqGwDSialhYxMyJvgKBJrOBX4AW5
KhSEc7uhx94w7JJz3H5TkrsU8CIxGs86qY5h1COy/+v96nGrb7P6ge+t5XqVmOUWGEwUKYdSxMuD
j7kI6lK45I0gXYiRyI+skz41bFuf0tWjQ10ybxOTOb7JXswI6nn2py35HnlvXUVRFP8EerHRTe9E
Xvr6Uvjq1jlDypxahq1A1T1pv4ai2wXH6NIZINSdjRnKRbXY1ej8VmcE2uz/zac8iHU3Rs3Wl/zF
SMLy2vf/7wqQJSZfN01Kds8JjmHcmqsnqMtTxzENba4GiUK4W54DN/i9T4+KU4BBo/pt8IOq4CS2
huEfQBTsIsYUUYuzN5WPKI/y9nU4whWGGLJbHr6YsXIyy6dEtawN13/0/WiCYsLYsKZbTR6Cyzcs
nXrXUhwLl8VzKmYmHdOrGqhGM0hAopE7t7afgKnJeGHF8yfxXpfn1ql9p0vbhSuPitETqsUycsxx
uQjrplDsEHrj8mlDDZ6yB/kvZ/qF37vAxIbcaTuw/Nj2iNLaV34IoA6TlTGz9aQlFIxKgTt7HGxq
efPX50tW/fsFu5i8cx6Nep3M6IJss4egciBTpOAfskSkqBhBIfO987eHeoDm8dz8m5G/vRLMX/V3
JEl0xfsZJAISNWGxV5gMz67YUPc1RXFgfUey9yfTyGvBG6zW8DQOx2P6y2hhpJtYh36pXpFEsIu7
riewG7CTrPnAqQwuMhu1mhcPupu/DyaKRb36ZA3wh18auAf6kfNCrSwbz/0M3OanwN+l5GccsD9O
SFBvd/xEWV2NF5gzxso+Bh1/DL2VzGgzh5pbgFA+pM8uRF6OtsJoZkWSlPY8HW2GCnnwhkrfCHZG
irhWN0s92O7i/blo3bxGKZp/LAhjTK6x+R9mNB0b+CwUMJtEK2MeQBKmnylvcKV8WkUxJb8V41Ej
72tBsMnNmEJ3V31GMBC/vwtj0sZBI2igoLSVE8ZOH2FJRMOcRJHF4CoipWjgBwh8Sg3hlzw60KAg
nH5GdEcaUB+MrAdq8p5OEig6swIY2PxLl6wMLe6g4GyWw/4EedTN4tZRpJIS0+Jus55gGcC4fue9
QwUP43ValQ/KtsXxJCxKAAi+UY19a1XCAOJa1cmA+7klxFBXumzbtzvhxkiAgN3eo41qV5Qk/lBo
wx0ZrOJxbc+SEBW7KBKse01gM4TfWYcduTkP1V9LbeBsukmKF7Extlh+7VYk7r8P2KQfiLcypBUI
bQQIwczGjrp9YiXlsiHVbwNf+T1DjFw1V4ZRsnjFK/MF4hEGe71hOw0BiOopK3AJjlQOJJCc3PmI
c2ntPb+JXLF+XjP3dXmh9OS+wwlCb05GDagYWwIN/HESlPxsCUtwjjYZ5b61cOL23MtnoaRSXQNr
CzxGct7hjQZuWFq4rIzYZ7lzZAGpeOw944kCphzb7W+lvJ+vTxnfbl0USjJDAm6IdqE0V90BDeat
XXQI3UGhMpeTGh/BXrwG/BoJ9K6xC6xEtm1L/tvfzNe3f5CrZ8Ivn/6N3hbAJPZbns5PHV5I2zCX
9LCIulmpEn476RrZgILIizkIechcTp1vSliLRowfxXa4awz1WffSwcpIuQZnvF3e/LIeNwyin5CY
cNGJ281F4fPRtpBy5gqo/hYGLv5BWO3D7LeZvO6cWEhqC71jrPWYp8Ru1Ps52qbrQuIvjdCsQLyZ
B4+PKu6ylSSV5b09WARibLQPTeWvBtLRubFOMnQ+NDhL2WtzSDul68AeXLe5EvG9CqqIS5/dEQCf
FwFVgaZdJpCH1g7tRHd8GksWQqs0mtnXuM1RZki0OH71UAb33uGnb8eEdKCblSqEWlkgzdlIQB+K
6tvjBER7lT0m7XCff9qbs68m9mcqxKv6LtkZVmpkNqzActgWo1IoFrgLLkYe0mNFsdvrJ6SISUcH
9m3RQ5hgYNfKy18xLx5lthulNihP2rxI8NCnx/2J4YubbaZQNhve6ENezSUuqvR79UyrHIWVG/ms
kl5jMa03y98e+YRAiyVwzC0mWtNuHR9tX3t09si7zszwr4vu5Wiv1XUhBgqL5Fsek2RHUrnZvPUF
NEaYXx7ty3BMQrlS8HMGQTkC78v7JpQKJJ0gjHdHRI7t4MXSYUxloYFAtQ0zLrYFgPJALwijMSkI
BcBWs7wSRySnKPE1F0m9lXblf1tiAV6O4I4IbSHfUtAWK/CWagUDA3iF92f4+W7zO6egJoz8TkLH
lyQA8N+67d+yp+nQ9q9V+IOSVT4AIWEURcz5PHCzc7uofJwizaE5jt2rVeKyPR33WFFSe4M3z+en
F4zaUZt/Go/kOsv5DzeVgyD4SVpZRwOLuSJ1B89ehq8+vNjBvujfVr3u7/WsEdpZbNrVyqr/Fg//
Yy8WKDnuHCdJSVYm9csixn80m9ay4ae5G7Qc2mD9C/Xd171Ev6EPF1nci/LiUI+QWrIm9i112uOl
Qosr+PnWIUd5ZlNmnIi3zfRAxaqUMr1SFyF+wTAcfBp/jy/jIInULNFBLjHCj6hrCzSz/+miLX7r
2tZCvvFmrZAdk+POzXQDjoXWX+Xx4Ptxr+R5Txs4zJXpNtHKmTwoe5SGIrXuj1dntOVjo1+DldVH
wLBnQOa+mZPoT2I2Q1La5ISJqGlwXPrYZjPReI+aQMVCCsOkRhGHXcpL8aqen1UBqAiiHIhG2i6U
2j6PRfs49g8/mnUeFkyBdwyMQ1jLAGhDhGJy9oi5yuNi9MGdlfHABkGwIK+uWBh4qqKioBtdkPrK
ArcZxinR3kA2B5SD5AhOtZ9E98PQpEElMJARsNb9NLlrLYu9oqp60HO2cqIFfMchrckcmM8vNf3f
eG3EVj0MpAc7dn4FqtsVWO0YtU6bunAYfAhrqqBwwXp3bLqoRgB6QlImvgusFVnzd9fSRthzvTbs
uh0QaIi2IuJXdDDGDxS4rul0Y5JIomrJDBZpXQsnuOZ7zGwI3V0VaEp2z2HVpuh1cCzH52NjTgDF
qF2yAZoXTilHA4g1KubR2s0JAJyT8L8zmAgiweOb2LYHa2WyTK1VpW6MqdLbInM0Uo/IAc+hpZ7h
s3IFx4w0Ylc/nRHALXJ5tgqiWfCq8lBYNsIgfeC9DN4ltuz1wKPuiw19kL/yCtqUewyJlYyQkQnX
SKvn3Y0U4wHS+OrAWsd3RRdv3S7mvl2+W8BujyCOsraYgpwU+JIml8rtHU1yJyPU66AJwCm/vTV5
jnpnEDWlOPAa2bo1x485PxYfloV6UrMrcCQOvyNtPups16FNTP2ClQHrnvE5ZXhKqhCjq2nOryRM
s4HAQlwP3xoLMND/tHYyPaNgUH327ljCabTiZ9c5aboWIuPGqMZ2+QpSCLubiuz1lUQYvpY7uTJ2
hnPva4lY8/v/q6em6Yn6ORPwaUkPs6Xto60aLI5mzHkMEISPjb5qbF+qcPZs6E7WLP8lw4/p8If+
78ZvfVbAwjDqUcb6X+4zm7lNEWbfbJPnQDDhno5NKL/XkkLBsyNpJuFE0gBohz29YJB5yhvSvD7t
Y90PtD73qUBqiPlqCQ88p6yEU+8/owEl6HHvSW6GxYh1kYXigNycIDYnYYxNVwLv/97UUbj43vkg
E6ctShcE4MUyWqF1DC/T3kubdEh9ToKfxcaFzQ17NlWkRINE2FgVeGDT7xDs5TiDULCMyBO0ApO8
hFN6aZd9+yl5lJaleGVrwzRPhNOFpPbXz209rxtx/S/sjgc0IABZOTFPUjEE0UYV6R9LKx7pLdGD
hfc8Rnb7msT6YkWJCRNmbk/1yvMsHWf7t+/yhfvHqVRFvTWZ+2lns3qVjKX27390dyhLXw31S+bz
LmDUxaYNIwcTZTB5YmRoxVqF4n5fRsMDOHArpHZ2z7bNUvYP1eFIXIXY6otQNPHXa3xEmFrLHQ6V
SD3E+f8ot5VgKesNzYFXwRxk8v2/3gfLmjhXPsQv3B5VmPMEvw2p0jobvxwJrh7JBSLk1cjhyZ7W
+ShLHs8OSk0KL7u4r2tU5w4nwXhW+vYuxTjN5IOdC7yRTXL1XH1a/pw1AZE8+pCrxpK6Y9w/poRR
HWcwj98aArDodDNx0ZIZWLJkPIwdjIMNP+Afmunhy19BBfT4jyzG+4YzimQR31z0IigT+i9O8uDs
CndESWVq0Ondvu9ZZHREEOXTdO+tevI3bODyn7VfViV0LjPqFtnc6t6aESZDtRCANxvqb48LS23b
vt5BsH8Bnkr5C1wJl5oH7hyrhvWbEMM5AsIlqgVpKvi6CpD7TF3wT963FdywfhhIfYfEuruEGW42
BDlLxPHs7fo0R2uAbg1vfA9iRQp62UWXykBAiwoviR9lKY/xwo/MJINbc3WjClg7PTeje9ISBwlv
Q8SxUp+Fyehm1yq/Wjdo4TcgcR8yP4IrS8eTDUOy+NWea1cBOAA7XfBcAvhiwyY7lyGXoJGYZ/FT
Gy473l00DoE6y/HXm5B20Y+M7aG6D4/62VZUT6qeMYBJ3AOXcLqoYIJeYn1k1Ek9TfGBW79w1Duk
CBEvUTL1BtcO88zyx9MlIOxNU3jac0vpjN7lRYLuxKT65cZTyZhAJpwlari3/PkyJ8BBs/W2tFzg
J+/njsfe8CB1VmDzV1f88RhatS/wa+W11Xf8oap2c5bJGGuHgoQK7+FeNOukXPiKYwQ16wzWHbyj
QiNmus2khup8+HWVPhks8i6rGq837On5nkCQADNKE6hUTAzXhGMkcDoQqRG8Y508A/SMQuF4++aD
GNdDI6/pi4MpR74gHz3vY9ZP7kIuZMMbNsDgXOqxN995jonhGMTDIOE/yy41IK7yY+F89V/m6GmI
tCbPNiGe50BBeG7zK1m9wHKyPnsu63DPKYCyxmceaY217qJCCliUbD2JlcgJ0ZrlbeyWZEIm0j/F
4IqPemJF8Hp9/Cik36ZYiwVMBOX6bfilLKqe6k70ZImRtw38WzIE8YCMUX/terxZqfO7wstI7Bwc
FN3u63C02Z9PnxfPfY6GXOknPnfLxrh769R8xYEYLOkfMxAwZgYtT6z5PBCJu9J4JBBQXakw09q8
wmNV8lIgKrPEun9XnN7zRAmWyTQt9t1Lny1oa6BFgs3/y7RieS8UtAvsNo+NNbUejJNXy1wkUSFj
0qTsyiZxYgKXyaxXMtztrQFb41lcm68vD0Q9KGj0Ic/uIF+r3IW43GO9j3XOW8pJQxPWgmCXhdWS
HImuLKxntflM0FEiN2V2mnivTXH1FASBONtWx8oQAY0YQL+k2QFseLuBO04t4mW0CLp974pMb675
HfwgN7RnmshIj6JX71lFKn9QQX1D3hcQJerQ1FgJ6Vq5hKxD3cYdCSVUU9r2zdIyNYnE7Ja9jAO2
KlHVAjGbzWMNQ8IMLs2mXo9fuMUB4L8LyrE57dWpmLfNqemgC6PBk4TYiTXP9VZuKq+UL1laPVOd
STewB6e4xVAc6DHp0UUiFzDE/77/jb4zCyGeNJw7ZF38l/7rv7Qa1Fci4RU796GPrJ91zlseTvEf
y9Us0qEZWaUfjOQE9PMyQGRs8hARVk42JBgvqhqOvTTR+vucUAzpvg60sLdd+2X2+ikcKQCVj217
nCSbrcw/YJ9Yc5NeKu7zHqYdVfUbWyTkFItUeKQ5YFUYKM1RNQydYRLgWBsHF0v44m8UMkNn6oQD
tSuQE6pAtC2T5/PQTmx7A++vJgFXX/+vBA686K3FnurSKeAqX/U0epxuwBPiQPnDkRxQ6r2T6tjD
JFoy6q4PrW7H1sBoFEEM2hI87vvQz51+ULdAaadMejgy+1ivr49tajrqhPt5ocWSnY3NfYX9phjG
K7HbNtYEGPyjkmvXYHoCnZaX/EXkrsFpZoG04HFd3v3DReScxmzDQv2vsGvBeY331N6mZTcdrydK
MivykUWKYoovL6cz+OcdIfgorJiOqRK/0TJzGgvqgIjznyVdgxDCgkKnVAH60JMq6S0dGQRH7Tia
phNcoTfYkqTGvdrZhMvNybnqaBW2QyLu2j67HEga4gj2UkKC2M5kJ1330LM/1DkRJnammhA/+jfx
/Ozc3wbMKQolC7lnZPp/aU6yIIOY/qMb89ac+p3VZQYGxwi9M3vnU4ZUzSl2OC5zrZGWMUfztGat
jceihFPYBI5694NgR1iSOy9XN5AnuCfoqhlfE05xA8B0mq1vgHQ7EM9/32dVyacWdG6vAkY+eNJU
wOG50D8y2quBgYhL801SIRVktEjmWjyyrL4Rb3oHHvRxDnLPC690ObsdirCuZekRxXAphi3HFDF2
Wr9fSyIn4BUbgi6pQERjGjRzluuwSBxbFPuXfRUvTCCpMw8Rr4wFH8SkyRK5MlSdwmDEeqRYyoL3
iy8BJQZucuGaNbbZM7/dUMbib+xiBg0vzKFP2Hzl9o6oqGjbwIhsX5dwhhjer7c7V3t22IK4sY7J
bMw+MiUjcPiEFmuMjrOqND7vPkrS6xMrjg6XWSp5lzsFPT85KDiYSUGftX4ZooRRliT0iahYnG7t
pCqJG+1bdDV5YCcQfu3sz0Kt28kx/Vw87uEM0C3HoXNbqphzNdRW+kKaAjhfVCIYsLtlXhVlOwGz
Z4D/fdxr+AzwBdXqaCJXAXfYP0chQjkKvIMMV2p3zTam2liSmBxF6mtPlk0gXuDUpwQliZerViLK
GHTtkAojPh6vRsBJF5lE72LQFTM9+SCFFKU3TVeOLHeCT+4eexAYeoXIHaJpouU6HfyaZbRjcVZd
j2evzWq/1n4OvCoVA6qF9Xrd7yNTbNorgWpgDC+rZRxbthncGDYSUGWLyhCZ5lAHDozKmwu9oQyP
i+ZZcwnAxYNmoK61JKqWqgXiqM7Y2hf7LzEEYpiz4cs7g2LZH0F9zbnAdtDd0cMJ5je84WEiQKXF
UCVtcib7DNBovT+8zXF4oc5H1smWc4/MkNVnxBFY6tKuV/djMvYa3PSHi10EdiFsu9coYmoDJC+Q
zWdaos5AH7acgNVyf6cKtYMsHGE3UHCrk7brsHtv0F0oFCjLf0H202vagoGdXsnaCRPi3t9atP65
TtsaVQssFUcHeZkLxHBZ04CFpF6mC5c5cZLlX6uPkrEGN/QKEyRgwhhybm90SnpSp/15PY7imzuj
6tpyd1hkIqJZAmPAIb7KxNbCfl5btg4vrxuXxB1sZCt7J1qBrwvWKpTbBKr+x/1Ar1WtVTTOhyMu
FS+hdCHxIUMfpYNtSn/C38NOEkxGiHMXyFY/Z0sqUmDrFrDVyQYQlufCEzwbmvkR/SjHGFU6UADE
lorm9EUOIkx1rgDhPakzMsEpb/rjT5elar4lQmq1DdWxobELm2Kd0Lk1r1wyzH5ec0UYt1x7hyJg
kLNo32SUTcxXBMJgxJ0iT+j4Q+BH6mkvfCP7Q27EL7F2A5R22sltMZhsL+QjI7tW1KA9sndV6Gac
R5uYonwMuuqjSY025MBSwf5swjretwqZ4Yo1hyghW3bImBsTTAfbGc5pGAkXewmNexCw+YPsQkgP
tewYQ9SpL5+zMb4yc7fCVumqvD9JNOYTD9JTju1SZmHMfCW95PxhZ/OqYiOmXaPvjVVcgSYBz9hq
bwTeBqHal4Yu3iAE60gXTCtYLG7AwRf6n1w4DNjfQrh4eOUEEWSov8ex3HKyITbyGtn7Zx03Yzej
otz2H/xuCrq66Wy90yJWKqmgdxumi4tK6+NHWEF33XJ6n+Eq2o2lg2DD+4ZxdgZqZpweIuKtxNoL
82CLIkIn5/dWo/ksLfiU3HTKRGuyPjyJLGFUbdEcq4lMm9N1rYigQIO3GJi47o68frpmZZBTNZB3
1FHIg6GoACs2b00HS1o6NN/4Q3lmM1VHdDYfCF4P4n9NRJZs6Hg9h1b89RstP6tvhm2YW/2DWm+O
QUmJotm5MWzndlEbcOIPJJJUMMb91mmCOJ3iwaayO+wO6n1UiFHHyV+ZanipgFigbfS+YgM9YUY4
zgD0eWRNL5tc9oioaPg1Tox+fTsl50DhDZtt1C3QN8uO6HntLDg1ixUwMGz5iQJVRMDQ9NZHMQM5
jRkR8Hv3m5bjLWDfeS2Z5/9c8ez2wpS3ZJE8FKm17UEauX+hupnzUsbCQTrdN52RlObLvrk+ZkSP
csZYaI9lpkpM9tP+4m4w/PEKbY5v+ybRXXudzcBDpL6YVlFjPWxzEohvloPcAzG+JZT2JblMN5vf
FusTW8KCib+ERwduZsT63ih/DA3Ol1r93AlU1mxRRsOwyHQEsUa9w07OBUN8kB0+ujKF2J8zDKsV
9wYfoJ9dJqa4brnqU5udWoRpYuvdaCCtPxiZfOUpajJ0+/LhzikCBuDF5mCgKZE0cgCZVmYWUboU
SAKUVZd2iXuyUooP3W7+QuBoHC3E8ixy+/COyiMGynRCt1RYnYETLRJGk2vbBVMiZxhFnV52wm8p
a8tH7bZZchK7T+wblzlQograHqdF5dK4/B+90Tho4qYh8FpYpONjuiI7XBgaWdMAu2rrYCjBJrih
9TJSgN+BeLfHPk0fqjWG3yg4gfVwzqcraRQiwgYroq5lQ5AbNiUGPycDz/ZpmeqptWnXqjRbVRfV
5ckjSPilxWQgn9/rec64Z8TlRejPdnag5FJEPKy8S95LyZFFlPx/xdzZFeTcB1/wj/KlepuuzPgu
IQTL6BRjv6rMACbqklAB6JVrnSU/66bugc6JkRhke4AVqA59IBcZhB7PF8Kcw7CsdygftfZyfPPB
/Y6zul6W/f74xEGD8B8kBLIJl3z0gpuWdDXOZoihPg2zKYfDiiPGixmUxkTovktUTNo1oRYf8vwg
JQFTQ3eCOY7t6Go4C5eodXbGUZ3fJuw3ARa6zrKSFRp+wyjn0/Ha0oHJXUS8Z7Aa9iC8WTMLu1Ki
gGC/A7BCf1if/5Hh9piKSIsA9zDI0MxI2PhcBYQ9yl1twddl/rj17S7T2c0MTYA4TkjRm3rqe/co
aQn021+NRliyvLj1DJXwa/oAtKLdWX9Q2Zi/TedKqHZZSD+NFpiDvZYoTpZDeCnAzlInbKVdhV9v
fPwEwSc9ZkBTQDusQP59zORQCmFn1vSTLrnv+rOKMFXbDyGR4BdVKDTQfdprT3Hh/5ADy+v/NtI2
RjK199IA0nIOpz+a8LM+/jjfiV76KbgIUYnbdjG5JJmqIFL8/+f1KKZ/v+gXuLhgeGifhksHzTTi
6L74sN8OZyXFoysg4ouhJhXn2g4vCwuLgpD03opL6WtpSfpXLOef0XmBMqFngDSWwytINuqXnawL
0qF5+nPhBoXNAl0101j7YsaqOq0bl5ZrZfYxsZD9RiJrcGrAicUxsIeO+K1XFLsYWimqqWK9hJyI
SOs75Es/2gqP4qH/zSG3O6rhR4ogxeL0frbEloQb3P6EYy52ziHaLa1O43Hi9nruYSVrXlaugma0
MZfmEfSidPlWTm6snp9PwnRRPZDppb9ZIm7mjoNfa1AQY/uzuCisll1XbT502NheAPuUeSgrgkZq
ATXME6wwkyZuB5hYMKLmREnpVHo/9wR+y8aWUxUoDHE6SlZc+QczETeitdJ3Org00g7nZ5OrYTjJ
DCUa6fw9l7unU0nfImzCX1mMDhaELohpJppPfaaKGd/EX+T77i0bLyLlTg6ktTZ6in6+VD9g3i6g
8EAbOdU5kIc0cdj1p6Phv1eLhU56nK3kWgivPZZav5hBZ8vOl8iMK0k7ELlfPOoiRTuIBqokeYME
y/LiyYvg7MitNIIKZEhMYxFZahG6Cs5KKBNZp1gakdmj0v2Ly7dmApbrSsSmTobd6lfP/S0dZqdQ
mSEZ612TY2FpLHXKudFkU6JwU7iSDTjKkQyWF3wXi/1DttypogqQtWR+gRMiAOGQ/pstLYC4c5Ho
DzwBYjJ80EMf2BY+rCpxH4M5ET1jibxBnQLjakkrsacOE2dxRvzHu+O3gTw2NQs6xHVFQNHj1Axt
mMNZ4aY6vQ5n6S6paUJ7lobbCPJHQB4GyQv/uCeSVNE0mN/re2IF6ww9NNARb5dD3IucD1G4XDpQ
+MOQSMEQM/Nq8B29zU7NgC9sYsIkKpIYlKvtOl1ebc/PkdusIftfnhxULNuAYzzoALylxREEDqe4
LrRhhT0XklW/nld2nTzkvVFdDR+HSRzgXAUTWzoKXv2HwgFRxc5zvYyvYPGyCE61YERb1rz8rUxe
9VXFSdUccmqe5z/tZjxdrdhCQb6Ea6QvPog8qsnyX0FZmlCgSS0nAdIS8hROOFqPXRKTHSCnkcnx
41ycAG3a1DqJAjM5tmNSc2ozn0KdfbmK9d1GtAvZeGS6uRrGcUYI6Xguz9++ZZmXUvfLzYNiZYgw
wLkD2AqJrbxdW/8G1IaEhUveFQfQQXajJKlaoBsJQXFyg5/Ig3WruBI1kbPrD06kHwV76eDqTTF0
nzkrDHUIJDuUL3zisjHxDLG1uEy/OMOyUQ3clPI4LLobED4Z8VXiWJuiKtC3KowXN0uE4/Df7wj3
LibM6SwiWPWqtsfscD6HOBo9sqej5P7VrZZIE9Gm5cf5S1XZByz4wice9yREBc4Q7bVD4MtkxUnB
lTwDcJ8bUMj1vFiiIYxqe3QfyOZkqCxUVwOpeVVUZbPoPwRUexeYmr6bvn1yi2za8nhnxdJ1EQQZ
brTal7bgVHXrYKymf5iST95c74yhqZnwESvv+sAB2G1gZ1CdEBDG421R0YeDfzi6laQUR2Wg6L4t
CU3NfS7bbIKZnu++JHSv4AsQFrhQwt5e7jj2HiTqdm+aJa2GgV8Wmv6pk8t2cxMNhvJCUxU5//5S
tbWMefcyKyrpxkJHGDovZLno/8jNL61CVoNvH5mNPgBoE80T5EM1qvjXP0fxZV5UXwgUOMtD5R9d
q9i63H/6hORuNIp1e9Dw1iCdPctgYD5RKiJ5jEmq+OIB40J0d7plq7IwV2kjtJ8LJlXC6pakdNAy
jrH6OIQbdyqZkt18GC07ZeObyr3u8qlFbbPuF66UISii9wEyjMpJ3PW6tABpPjLksRr30Gn+Ra6R
XaNZpPNnCkTgkyRbuPLwLivbgGWcUVE7b1ZZDnKjINLFSs800Mi7WVXuFI8Qvp7bAve3WU+Fq1zl
Rad7+BpkbL9z8p0kr4q42y3esIKMnngJKSZ68QsvifK3VmDtwWEcE4GJdFxCqYtX8F1LUs9djVJD
xCmA3+dRqBAKTyx1IoHlDr1b7GmXWYbxVlW8TQ2Pev/EJnqlgwSqZC+Bf+8OhhAzdN5gCabUr91N
CFfCUzQeqT34vc1HpMbfBgpKsg6SiaRC8vYC18jgJJEOTqVLb4NUhxzwnAC+MhAa2soFLEsxO8qP
vmpkLPx3iFBQL02GsVF/J2JqG52Trds1PI3I20G7hKxbmRqRPRz4XHU/lsNeUocDdKRz6bHi6/8c
BNTvavVRzPgEYq1dPoniScaGMUIt4R0Fs+Zf5B4C7j5hDsH1p4YeN+pDXRriz+KtPn/RZ4uJVZWG
dKr1P3stMIXwlLEpE9crSlYCDhkbF/U02oxMuFey1SDy7ORWH2RrqolvHGRbvpjMYmzyyE1nFznn
2eGvIAWIrn1YMCgpkGQtyy8ZFmCd0MX0hbh8rWeGTGz0egKdJ/Q43lhHVyJ+ekZVhJT8qMSk8etA
/K+Xv02LcvzvQ+p7cZchI2bfzoevUpsmb+h87g+hb/98mgIDCnQJWWjo0SEJU9pvN5gnDLXaAOSB
baZ5NXKIIDuZKaW8pv46v6hDthBdi5DQXg+7Cn5Rn7hJEgFvdRGA+RqPR0fkZu5PilKyfBCuxoua
aDnL+L4O24a2oeNDam0v7cOiX9/EhXsK5x51FLXlpKLvpAaU73OmNmQAiIuL2PMEhxD2JOFHG0kl
Kc3jwypwk2wbWCY9gQrenzNDbl6skVkIc0Q2GBGJqMPK7G2t+PX7BrH3+PMvl3IML18poh2pjnjz
HnfyDyTQiVqQx42bVgcq0BY6A8pIJ1UIFkzNyRBCte2676Ub/ZkK0NxSs7qK0GfhbZyED2AVXrVs
igQGlRNjNuhdD0QQw2ZzQw+rqKF7PfAkgAB1D8d12AbNcYh5WD8n1DvAcUfdyPT7yV6RWoCkSRsh
4G4znEtSdhJiCoIe24Zl6N7GPQO+YoC9H4A4McwOWYNGlQVootfiIT0/wDmdQ9ra0F/EJDc2/3fE
p58aeTt3VRV85M3ygFOFA1b1UEI1Utt90i024wnL7MOFc80JLGXonVUODORQJY8Nln2JJ0B79rSY
EbN3gV717IY6HItc//vIq8MEUmYT8ZYe63mBzqCxRprlz6vGTsWTDbIey8XOkfKDNqDzIie1Zmpy
WCzo7NjvYKFDW+2Sp+qbyBJuzVsRDGrCOanvdAyc/ZyDjWnITj+tZnrMtwVEoybVB/77cE8p2y8e
3TPK4qp+KA1DsZElpdsotELcGeCXzoAGrkTkAls8gQ25Zkya6PMRv0SzUkwV/w75L/DHID2CttUT
fo4+ksPgtmD88RsLRxuRKmN9RbxeKQfX28LbgiqZgi9lBw35Zm+H/zGs7ZAsuI9vgNyiHE7hVf93
Ca249gD3bTLTJPt5b1cVdn4/BO/VeyfSkyFi9DLoKJ9zIkUS+gg4EQa4P/faSKdhCmHy0Ui13SDq
vA/abXqlpBkPiZyLWOhFrdimIWnysfCqaEA/TG9lXTSw88oy9A5sjfncvsXvTzVnH2USAp+hMGWJ
IJRld9lPIWdKMMx+z9Zti+UEggV4BUj2DUVMoI/YaqhyEap2zlt+dVBSTuU2tOK6mnQV+hlbNYoC
yBLIMKdh89wLPe4ACrsAe3kJgnw38tegRP7PoXA7q6yvn25EtSgzEh/2vzFeNXQqm6trzxecdeU4
GkYcu5Nm+xifRuUnhNvrO0vbEq46sirYRcc2E/Hk24JSp3lP7eW5vmHzBmmT3FLRHZsXsPpWN/h+
3KAMycbyn4TI1BGwr9B+6CclDiA8tlrw9znIdyTRdH8Y85SCo+HQ+/RqAPdxfkmNJg8zUFmhda2c
2EdXE7LFPM8cZBhjI2kGx0YPzT4O54PBV5KqgQve2J+jq/EHArVj33WQIBO5sRYmC4DNGCDJ6Qbd
2CFXPuKkTZvIq2FfpMulTDpvcP1iN3bjTgbtRpQcD/7+1aw+n7yatVQMNoEpofEHzqK29/ONy3YU
wsJDY3KPKTSvhsMaetmYpQ4ChB6Q4oeinvcbD+xieKniYUDhZZtuiV9THhOV4ksFKuTyntHVSx5k
dE85IR+ORaQPHKBf/lyr+O3WZvNH9OjyxHtzt8O8ltHObN5yw70LMk5Q5/JSgrk8YJ11mMfWQkG8
hC9nM010otM/qVZurHEizX9VRMVegumK2GdOYC0ho4T3fv+jHJAMlCvmiU6RSLVlqox/lAJGSIG7
p7EdR0XW/NvUs5Mn/RXYzTb8QTWKk6UGTqKegFVZhdSo1+wTU2sRhmSq+XzpPSEmubCw5OPZgzSa
zfJw/LPbSbw2D35xIAadJjbDTxbtsx3YO6KWXZJfPn12PWv93bAmFKiXgpli4Au4sK0p70Dpr9Ty
cTRs78mttQ6/tIYQ8nWJBAFHWKmBl0/rCHHDTiZHcHxUtVLYHb7M3vIZ5LohBo7n27zUmWmuSlKm
r42vUHIMc7HrFc8Ywbhy1+0U3ObA0EzoSIoPFQdComW5DVMHmXm1U921djg5cLuckNXrAuS4Uwwv
FByQqJuy5Ls3UPJqEQ8UcWv5C/LTnY7mJ+X3T/R1B2/3iCWkPE9X0yRLpaJhJTAmEPp3/f88I4XX
S28GPjr5tOgCMdKfQzt24OHDaFRo0XqJKF327VsxL2sdfOq8Yh/2HxQ3FEtDVVl5CdbtjLhLmd/t
QitjLgk3nFPnxl40rcLB3uXaoXCjMvojcxYYaTTnR5YYTsyN+sx2wuxfzN0qB5VjVKw6t7P1SAwf
swU3+y6V7dXhB3BZP72LjGoGbQwBDzMxvxXhfsodwWwqwsnpJByGrFrdy0d5b+3qBisuUWjTxOpv
pr2IUsNHDPt9xvyCMS/KHv3Oz/I82A5iZWo7U4VvmF6IZZMAYmR7XdACwS9DyAZJsLsSU9Lf5r+9
x8xDCIYj+1EudGJyrjiyebbdPUprxv7Xp2rll7dbVh1ioiGRH93hrtxItNCMduc9T1RQP9r7GDwl
ECWVbrjLqMB5NRvW97IYae0ww9uP6o1tIQcoy59IwgXLYR+k22UIEqi+1B51peQz2pbyyjr2lPTq
sYu2XpGgdzYKJFIALIWkmRoI+ArEHrUuE3xxZgD/f6JbjuyeZZy1p2TxhzBs2g5/PCAKTKPXrFEN
NJR/lIR1httAVM7wkh5+BltKskdoxmRekSgpibUBCWhj6xRONjohGi1x5bJcQ913CUnlJF4mW0J9
RMAFOmN+DdLAZVXx5WYTbgUYtFdYR34d9YyPStiaC8w50fJMzfD1XVxCC8/ZL3qQDp1fkh6Mv4sc
tG/8g0DAztgGa4LW9shj0nJrg9vM/b7VMjso9Oy/k0DLZtqxgaI1cVeTQ8HrxXAP4JW/Ubyy9L7B
fNRYTg/2V3+po7IV84ucGmJ8uDdlp627r00RkXFIx83OtufFJ2WVNUekU3qVQJGXXZ+8ySBxXVVG
aCNNxQQ9PwPMp8QwFX90nEWgY3CiODkJ8OlPme13rgKrrOei6Mz/jKDBcpPt5K0rHOmj9Zqs10T2
zvE2tAXCL/tvy7J5VkUi+GFrZtOWZIsro4NGl0Fyqwx+SXJth5d4bUpntjCKFk3qxFSEna81CFnx
K4B08xh/RJIqiCtZFlWVijxhUSFv3G4+1Ey5w+bAgUAng6qimvNSjmAD4o+Ro1VOhhMgRuUtOEF1
xqK3rvyf61k017WkJSN2/QCEYRCcdyVXRgs5w/umvwtBDe0Q+PsLje9uFK4+h4oVt8qe84S3YeUt
Qod6QbBqFDksgTR9qYTHEUnze8OUgixJEve9PrxRqdWLyA6Wefr/Sul8pRUSVqf/sDlGGihn7vJi
ihguw/p/SIUsEpf7izLvxkH8GlffLSbu5guUanhE+cmxQxmKeV6q3dcyCa2DAkrpHJ7OkiB3GajB
90Nzie1N5ULIjmVfBnzqd/VDKUWFunGz8dP5VolCtahaUKNmD4R1PVfL981QKErv4f8mJAP9E3SF
IGElBwxWoH+zaDNffUeeW5CfgotS+BQbVd2dshgw/wmOqQNZatN8ommRqi+G7NweNkcsWofMetaX
gWM5zBQxSNnEDtyO37X2E29qs0nHDzXk3J1y4HzP+LXKlUi4qYjEo+LEgXB15nqpCMu153Hl3Z62
4hvMjhCWHmZqE9QOHgNjLrZbRlYbz1ZMXkcfVcHRmTe/rssiWJcEneO9wGBBaPL93Iep/Alfoz4B
qNU4GrzaorkYw6O6D78suxHoS/0MyNADrM9n3rLQNWRWSdEI/edIWoEAzFVu9Vg7fYsz3er4X25m
ateWmny0GWYlUGSPMGlCeXCaxq8mwj4SYcdjlMNm7Nf38DISx0kbRqj/6EMx0Gaqj9fI/+n875z9
bNg9ewmASf1U0Shyn/DAYacKhcdkVE0JZA2M4l6/91wqK9i0QzTJ3CbY10nGlRjRwly/43evzcbe
Ao9Lho64RMG0yb9UAFy1IiGSjjnh/22e5w+WUtZY+vbLxAVnbaO0yqdCdl0iDf/v+1eBP5Nk4Eml
7zOLB/RZ992/JZMPOhenGwlFJNvfOg8jJK97da3qUobhgn3/4/jkwr1iIkDGlAB2N+if6QIxOyIE
FeXgptqa9P+AWRD7wwwxg9KbB3JvhnXAFDEvd5mdWxr0C5rb6pKlPgQzsVwNQeGK8OpgZzUrqmwY
OntqIG8UiO84c+/EGLPdjMUIt6zM4PjBdfEKyhWF3qMt0/zGxTqFMSfZmuJxEFXrGqtlAYMzN8gJ
n+4CkEKO1lKQJw94xRplpDy5J+sXI5IvUjRfLfOXwfxQstJseq3fismtHKsCXDrrh2kvumLEv2I0
Iv+dX+yrqtD7PwKsJMJ5vnzIS4oxuwfeHy73au7yvyRgzyd1g452t30FuzFKs0egYLpP+mhi9IDN
I5jdTtcF5nhbkQuiAeC53TsJkz3tdAvsvdAlIchtWErDiubD8zsFPrEIEaxzoeD2FBwjZKuEl1lP
htuGR8o7QqsZm+juwRdbNfZZKTy5ymyuD0FwGxpQa2qYjARDym5h/hUWtmxUW5U9KISlYc08QFsZ
Ojxgr9y3KWTerGwTDssfr+ZOeWsPEn4TkQsXOkDL/kz46ByDt4kf8+yWfaR1mx4PO/ny7Em3g+z/
IAhWr1fl6C3TzHPAKNcTLjN7B8YaEjJ6y+5wx9vbNbJxBqq/h7ZkZtH/oQu+D/k23PB1zbZVaR/X
SXHlEgZt22fXyOhzZDHS/7oBmM9iSfibSvMDwcoYrgqZPa1vB/O9XhMR6N1yoJ6NDtGrmUW+umEj
h4I/UYowojMYMmwEDBax/s1eDsbf5h9f8fq6BzqTwBcfKloltMXNO1DDWkbIGip/aQGYm1ec64vC
TN8kmge/wLEt/wbvG8JYRKfjl9wSpKfN38YDDz5MEjnHzJfKFj+YeypknqQi/eo4ZO7A+KfDnA9g
jCrJAvhYV7UAeLqmQfRSYImgrEV329nNQVISowKdrSFL8MLRXtdve6AWUBlzobPyCFyAnCRNE7io
IaGwVwbeMMDuac5gHEedJ4LR3iezqGaxAdqCRHI4QSM5g2OCBkzs6G6Y5b5fjjFu/DqeX7y/5gWJ
D9/OIi3lNcJSdqlrGsO1J8JXjuXInKwYX5PsBHuKy1CaLwhTSmeOGhMsnJ5Gg7M8oigz3pFp/ba/
UmI777jW3vuxQCocGBOR7JTFQN5GpTH3ML9YBldUTXN4i8hB7An8Cwbm7WuymcX1TcdRJtRF6Oyj
pEZNjPyZQ7XemuHAQwtbqiDCiwUM5AnhqUE3YLwkSAKLqpuRocwBvq9KVeOqnwPxQ3qwWxKEkZF1
cxpzQsMKmsjw9A5838WJU5gZK4Uk17nBlbK+WFyJseADuxslpLykryj4k1iWo54yKDDU/u/A+5ie
I8B55pBv14g3hgGhfGYRS/I94sLk5JYsfJ5eQcJ8cObIlCj8JNWrXnHNqFCDqI+AilLdpPQJc7uY
DVNkrrYtjG/Z2jRcrqbbfEn/qrA7iXjO4KyqluNVApK89jWnTHx5KW5H32LiIBCzLjyo+wR7sH9I
69mQ/YC5082kDLgstEpUlB4XE3zy959MnpTaCwf5DCmrCcfO5+3ME6x/3sTV//khtfPeB9y2sdj0
NnCooa7TyNNZdlpZPGz0DbWTB/sKGR2uO0/XjCgQCDdjgIqdYavxW6tR+xL/i4bJvw3iixWgE+tN
DRHQ/1pvRbTSqcoJCktr75xanDuN9uwSQmP/JGy9h6Q1LnfFnT5w3gK1ks0GnWh1uNBLGinnjK4l
PF6oP/ZoDMfSEyg/ZBIbiLsNaoxByz7clJVqbT6k1aPHuh85frxb06wv0rA4S+fqjOhF2/YGss/S
BJ/rEJ3sdb8Xf/ffxi2hgoR5RYj+ye9OtIO8COsyjSlTOePCULH44R+Q6g3Gc64wVdDLzPgKdlif
7y4CLK1EWiIabhwX5i4vazSSxOQ9JWXtMHtwWAobCfhIgQUTK0erMdZ84Sdxc2/h5zExxQGuwIYD
CK2Mlo4mjIhBcBEA7msbEERbNtUfYeKTashpyDlnmr9KtqCyyKc+gxdKlCDrPWzAziFnJNDJSLO5
Ze2f5u8hoCfp7rSMmt2GLBfe/sivdPvYkpcEA1BoiwIsRNPywqLtYhCMybw1bUPkmljyFELCNv+1
3SYdEuqcqjgVfyiZvh28folAhYdc+s/HmHd9IpPLylfViGVXfd8BbQbbVqBtBjJrWh1Be2KWaZHH
eKJZMTjqYh/jqrOVHY5Y8DfUncYytiU1wf2FOJbFlw9TkGBLfXsp6ZdCgiW+2wZiY6ZWdGtA5zL8
1UFlkR0IFKAL/DpBbDeIiP2cwYl0eYD/kYsQazWHq8YhDtoI6tXbZXZ/2eVpVdHcXqp3zjvr/LAx
4lXt5E+71k1FdFowczAjbTzADbohDCNbRi8Oja5VQQx2nfVCWTqhibLZFS3SWnnK0jJk19LcKcoT
nmNNwPoZE/ooQHEH5cY9Yr7732e7nHSWG+8KWzVwU9jRPxqmlUKOI73MmjmmcvK2HEZ2M7SfnJ+B
J8HHfwQZ8+pVtOBHCbBmyx8VzXtemveHPfGVisSq+NJcl2Ow9XskYmfsOOqxni/8zHve/4dUG8pH
Jq6GjTwktyInJCwVbyTvaV+XwZp/itXC+9JyIRtANau4gWb+Sszv/oHpg3o6UVn0xx7d9/ZjT1ft
k4Shjv1uu+I2VKt03PUBa2V/TMsi25gHc1lfCCYHlDRvAtkulBiebl1IAVsll2y6ykZXuw1btOcM
XG/BO0fSRk0BR/Z6jVSK+JIqTi8DmgEDbv8iOoy49pOTntrx6cA7TQi9lieD0BABnIoHA0tklzEu
nyuw27Fu8OAkPikp8wlXGl2z2C7beuM2YsAFe3rI4WWknpqJCngqRVDOVnEZK1TNGtqdeqKkdyfw
a+gDStXknuiyDDX8hQHiMaZcFstj+GrYjP0rNdIwxrv2OE9N3gYMYzgtfFWsFDj+pjtAUG9VLS22
WzKLh+WcOCSCFX+plvtTKOOMdJcyCBNV6D2DTKFtzRuPezEhyRHew042Ra6VRkP9Y/wn86wN5EuG
bqWC9F2Q4h0laJOXCNO9b3XKvmGFNnfqNnt1uCmayKAQZel06oHS5xTCNIYLB82RFTTM9HegK1rC
hwJAKeTDkrh+LpYs+K2K1ZvYa8J4dAwN5JQi7fZJQo5+blvGHLz96HoWNjs6DeVImuhAgdwFCGFC
3wMLM0Ho9sIjA1PilyYRRV871rdqALu26GAQP4u52G3YDIqmaAboCCjCNJFSPVfgqFeDX6VxKkv+
lxCYr5WRIAnIc2L8Kw6SnImUw9mnmZLgZ2UTVb4WB4oo8xUrkMN33iYeq6yJnOsIBtw0k0ru4Iai
4Csy/y210C6ckn1fPFg+0ioUg9DhyAo6Cq/BlWCMvn2XYy5WsE7NHiTbShGOM1OCXhacYwWIdpf8
6/X3xtj3QYhlcT6qEkILLEGLsIZq4aFKTkNgywvoYRKEjy9QklW39cJA5SZ8mc564IGX5F40uSzP
9rqHGXVihl+Jir7gAkt9a6ZdTi4xuT4XyeFaxvQ09ryC3xaU1G/bxIYnWwJn6E+KzOyAkv80SpP3
wOq0hqGfc7N84hLm9jqpT+WyRXwM+11ne8gK6/ViJ9uOvqHxMahqxCUHI5v2WBgw1kqyPnGXbYK0
2Uu3arRpvBfRw3z/2KlBnvhZobZ4NiBRJ5OZ1MNoN7AgiK1fps0+s1DteHVeFt7R7RCWJx01CxCF
H7urgfhoqn6H0x6KdQ2cSAKvW9zCV37isQEd+YjKeY7lqhnL54aNva9NtqAxX9BnVqXtB5PiANmV
HJo3bXKlLdD/zYvss/zhO61T+bnyoeylpf273Ihi0zG857O31Ui6hn7XmKFoSCcLxOepzm6+i/3b
4jI7LMFEJL+ku9LFWKO3P2az8TLlkCKKUxUQ4yyr0Xt3sxcTL0zXW2OTIxDG/Zel1o1OY7QRnB7v
cxAjdvF2XU6/8aFAA6pSJjwNUc9k0OS7If8nbofO9B4Fma+0RhpsMoLumEEALcJn0BBues+sQeLu
22myFZOC+HRC4W1N5tK0aplzn9wpF01BGbdKA7utAL7TzxkPNe3zFzGAPDAlpdHSg3D4goQJzabZ
SJF48RYxjBc8lj0mdhVO7Ihox0RwILs3CwEqgCwgPoumm8BpZOyEOKMF+GY8+GkwNW7fplrumGYW
qp8bb1QNELTSDm4LALgS5SJZd8SApeo6LguyK88OFn6p2sQVuuQsaN4DJnCg0LpQtWE/bLRGJ1Gv
sxg7pC4RZPmKee7Fcs2h7H4CaQQSJtesrlKWuV66XicO2V13x+5ej0oPyU/tXmopyNmG9f6ikOwN
YQLAiX2y7yCslY9gLZ84Nxem6nJO9WzRI5hcNpyl2q8STOVGsBcLlRAzow6u3n95t+GLYVT7JDrU
yE9m3ABPQgo/DFPuWNNMwuQP791QtyRRlgaOH8LtlvzCyz5m+97EK/TsNqC6PU7MZ+5UJ6eMEuxb
leVaEk+hahpHbTBnxQm9uCf9Bp1bLNJ0g2IJUxwLT0i9e97i9OdEyEnqai57Zx2ME2qOR/ZJxadm
av+P+iX2t7z2naC1VKCIZlVwbiytlTbEjOKVo7VQ1l+vSjJx/L4X3LZFqvqNk0ncEoxAX4kOwEcw
PhGga2Pz+BIClZA0LfjAlVrJpsevrndj4R6c4rxid/arVf8JZS2zj9XLtnTBG4IM4HZXkWHgg8nq
1GLqHqKDlRTUr2bLNB5JU0ywTIMfUa17uZOpSq3+cN1yr4bAgju6PJ7b9yKqqLl/fTCVYyZzFe3z
GSrEXCdunEe5bAVWtO3PB1cEXHp6o3rMfTZfliKCIW6rIP8G1kiRi69oc4nwZtSMbYphzEDLylt5
OPy6KS5luliZUFh8uarJJGokVCCgz6mqPuI00AjGMSsrZJ063pe4kByiNdFh43roTDVVZv/sj+gR
yZKaXCDcKXZEVB/vXcid7ERm029/bXeihvNDIJc/DpJrf0/FQzscrswvVYpQm4G0ytNpkxu0TglW
vmvRjZ9Oap08y4Hk8FwjRcl7OYeMQ/paa6Mb8TLYLmzAscVtjeM4jiOF4I5NDlOWzosR4tb/Qd/c
yxpN/ubLyfB3hCWqemO6z24QExkTZE4P2KzBPYSdbcx8fIJKp2UxsVDnXJBVq6R0sedlDpQY6uuM
5bdE/+ENZjYdUqoh2GzNpPSvjGRPTOAugJQ+btp0Ad8HqN8gBo9B9podzG1drQp/+hjj0ex1LHVa
ZMzBw1OI6U9urC7qziHbzLNH99b7gs65a7yyFCYuRDg5z1e3Pl+IEH9biWCacN9r2bMtXCtkuld9
JWXZUpw7g56zke/uuMW28lrqsYK9SSZwBvtEYYCRg7AzwaflHguQZIraPx3HI8y7eHGrECUS98ig
5YzfBWA/GK+ut9Y51EUe0WZYyJPznmLMEpbnZmpTKPb5fcQooxIpnJ7vM+T05tOqWBqzCUJaur00
qa0LS6ijtf2uA+r3PuZdbC2FGOpiKA0OxEgjllEBjQBI8mirBjUmr3pnL2CgoKFUgNdojlqahv8R
6ww6eJLApDvxEsT17bXQspmh+FXwtLFNUANNQcv0EcPdlXKoFmL14FnNE5vapqjvaQPk5B2jRiVP
i5FiRcZpAhmhgXll/Te9siNdG4pSPNWtMlH4DB/CzxZ0tn1bz/zfz0UURAQvJ+1X6pmGERNFKnJF
eIjeR1ZTuXeITlA9TQuMbsRsU6fffqpJHN/xq2HtJoUOxwF2k+hhoc19YS+MUp9r9iRrfeCwB2i6
McWU+nWK/S6EI1IIpVQCL50qTEG5gESRHbdfaJj9Z8KZ4AlbJ6JEsqBUM8/TTWM6gUVSiSPGqXkY
OHI8XRze47jnl4GBZXnyYg3Aqe3UZzIS1EhRaw36mNaspo5G3mRe4JVagpWiRH3UwrgA86TuAG96
8pwU8LguOleCLcOWyhXua0ezp4xGUu92NSWhhJoqwDnZaYqJWWpZBgEiVClNmHYDjChA5jB59yXX
yZvvM9e5sJXR5LKjE+BrdosEicNJAe5QwrrKWEaXjWcFYev1jmw2fPhQvPyM/I50dYNnqOpCm5aw
hG/T4nu+JbhtQwtGADBfSfOyOI3N4s06L5RlnlUKqemZYQekHFg22pLDDT48ahnt2f732QOGtsg2
7rmcuWPIYm3UquxTE2xWzUOZ7Odojp3BMEKlXB1E0PoMWzsat0jTDaDO54XihzhFyfqVj76pmDot
8jyj/ABVnA4CrkcYw2C5jtKGomDNCRcKdL6GGB2lLxqeejU+ED08a8jgi+ghQ8Q9PV3bjGHdOlhq
zQqc01GYPb6lGGXeAo2ho+oZTTM7MSKJ3zrbBsE3cRUez9mS+s5Fkk/Vw/qmii5C8gNmw293FqAT
QS8ZzGu8C/gld2b4DT89DDRCXc/oyfkLRbxIj0hO0y8mriSklHU9VI9UGt0fcKDk59SWDDwlbtnx
MUBQ72WHMSOT02MaRFszLG1zMJQb5YcbAqNEd+KlgNfyOuMDfD/UgKlPOSQg6IsBJjDDS8Wwipys
eOh3shd3gdjqVAtkmt1hzBJVlb9x893zMqPpUtlkD5xmLEDuUNdS0tDYabZUi0+d90/a11RpsPDO
3J4JTTbEbrkXXsGMTwWoAmOTVCwk/RC3xncSYQkOngIk3Ag3XGiZ92K8mDi3NufdkZxi6KmFj5oo
R8YlTMyh1ej72HTWhvp5X9bdLszcaJLWPborxKlHE7yiR7YXeYtfBPG2t1TeHTZNuhxg/3wMhcpS
Aw8x3iD22avDwQlLcLOBvkJTEve8c6aMCDaduT2tY2UZl8soLpYvmL2mU54RKXD+ve5tThbnzpAk
kFNkm4lIF/IPB+1cMUyKL8uWyI2YoYAC0ntvblMpuGshVg0lUsmj0xu7EJGQ+gdfHpHOsnz28OYD
LnPY0kAk9XSxUwVlDzsqGP3e9eqEf5gYgHHvNu6A49P6VK04Ij9pmYLxIA2c4TzAFXMeR++V6Xb4
ndjQ8rSxPI2rWo3/4ieLFN59R54qdkHJ8jyMmj6U6PqMjJkVoL9CFoDcuivEXP7Zg3KtCTwtXWtl
0zlYGLWegspE/rCwq5RzjCsonb5LTmif0q/PBkaheJRv2aaLoEYvxK/YD6XwWoIJzMCMVILlkh7i
Q+8pwcA8WYhuag6FuHgXPHRIXcOxGjZw947lwjdaXuHIJTGHfFbah2J/f0jb4GWtL43Odx+Mqxpj
mfrvsuCgKvb20P3fC40EeEaNbfS68pdIS9SISeRd94uMOh9D46IEVGQv/Y+L5/ClH4m1uA47u78+
FUeLyFkKRwX9IHkx3ayVeEIBFosh8930fJWfUZgvKteJpcBLTjGMeZqqC8dvvHliNGsy4kBpZja0
WxCDoTy9brtXTXMYekp4pOQ4lVZinPHzPY6KY25zdWTy8RxzBBGO0uTJZUvkdzXAihWfMhQTZJMe
Y1opnrmwG9PUUyqBqQxzi0C0KyxAp6XJMw96XXTnHZe2PuravFMmnGJlOJARXULcRh3DjbZiE3Ac
GzDi2LcZ+cb47bRzkRPcJYHSVwz97DzCjY3hEYuIlPzoDiygcQ49tOJmBsbhhLUdjUgOFVyAcQqj
BPiM1P8WfVfAucf2oM5QIGBgx3nIBycmk2R6wFm24bEvmJ/APmY4/svmp0bmgU/jP1pSJnctGYk3
TRnh2eWnvRZD68pRt/VgoY/J7r6lrgj5zwAFTIwm+wvgRRRPFTBa6gTGpPvCT2WlRXx8EkssqH6j
wkY5SJXj5nuFN9JhrNo+UXuaPUSasMEpfhkg8K+hc6Dww5NhDoQ4DI9LCt4gQGYTvleu1MmIqR02
oPwBLnvVYbW5oI3kll7cmxhHVsyV+jo3sjlfUdnU2/92urPaZSOFotdcxcluvgxuwIJofxl4vQxK
NxYVrbpP+R9UBFR6WDkS/zGPyL2/0mAD4hzoo5UIxOMpqrpthsb6bZPv01cYZRChDG1AL3v+WQeZ
C7i0g71OSsbR/ZH6y9bngRnXnuC0VH2f4YEzYoV8p7/ndSK4t69Z4TipE3efGFOryb6fQycBo9vg
aZJGQZMQxWrlbU6FmXs9qHFVvWRbWN75471MnGw5tyceVbbuXAuMbH4aa6PXYFbsdBMVAyMZJvo4
IYxgN5P1Fn4QxkIFA4vbPIZBIM5hBeMeKFtRhrM3Pb+171kqRgrhsN4T83mzzy+kQd3NbrMN8Wcm
+Jn5DhCkZDp44ETeDfa9VmoxeRM7Y4r2LmrGbfHvLDaRaFNcxhHVCCVDWoYDabZBxkMRNEaeee9c
yN8KQxwY3QdrIzrS5YA7IpdSrdyGcCOiaCu4StQJuf0g5yfn0eX7zmnhgkcTokSKmoD85sajkLfk
11RzdHn/0El5lEZtu/3eI8cwdRwoiONMa0AbLLMsKp8G7aWXFOnzw0iOPeS2JL7rOVkuJFJiDres
M0kuaUACl2G8YuK2hPOmQJ2vDRo8Zls0sRFH9M4dFgArTZXoPvE6RQkoqoWKfSwTA729yfyKJPqa
EFLNdJfu4z6kqDwBbIjV+mbcLMLo+gfUL7v2xjYUaabENF79C8nhW0YXuiqJgpA5G15zvLX1Sr19
ImfRu6UaO3kqr/4Pu2RzYO/Fs5czLbYERWJ1lRT8qVhC3SfPJxUfI0PW3OIeiFH0PMiad/whKtE9
SgV/dqwJ8EFOhonNJ6lssbr8qC24C+CsuYtgmfedF+ZFSCBIapE/iJyAVfbSGA32odJbXg/2ZO6p
vLSvAW3YGwutu4KZWTurqqeJMyApp3KsN+D4zNXG9HOCNKtBo+pr4friRgFlvNjNdjhsOLfBSL4i
zTWHHQ5EsMTBLZtRXSighKua4Q/DkXT6WiC1BluATr0TyVfLu+koFkYNuKzQvsf264YFDq+aIT5i
eRD3rHa/waJWZYO4o9CY9snUp65UILa5ATEYP70m8m3VS9zrxF3NS/ox56Y8M1n+WsiBfGLvw1tO
j90qlXomKI/Sh9lx2q55OV0VuHFC1+CqoNpEz98hzohaOoKX4znLUTZZmO0uspE8hwLS662PUkTW
L3eOzNtXTOmkluqrXsZBKGNjU3YKUw/md/ibL/2K5eamzsomRC8FEgdMv4gPrzd9X8ry3RtEGwnC
Iedek8mAFyeXXqdQMgyP3dfDuETsBGyrr9+0h6vsEzBEDHJLiyU69WFeA5ujiBvqEjLUfV/3WZ0E
1RyuDhGPPn5tlrNXJOAV809YD5W70MxcN2PQfen8QPh8FSUkdX6iaXyO0EGbw6w2ORHRqE0sJDvI
fjezEbmnqx5gN1/lRjtmC75lztdoCMA1oM9XbhNdPq/JC45N6jGNUbAkhSk8dPkHIqujx320gyRO
jY7augRu3Wubl400H+AbB71r+QiiTxjMtRneWjYfCzDMZ7/wKsfca2P30F4aZn4pDWoj5IskoRto
Z7f0k6LFpbBFcSUT7MJMR+qgoaYLK3FIOfW80/ndtIvAao91MZSCkXa8XWuOe77HkHOJ1ZNR73H+
TMmOE13MM3V38wOFv7+O3NosBw5DwIKk6IpggnhkyrPkgDBwVMZEz/hPGQIIWBfoPZAuPjc8+/vG
gPRhlDdn8aKEMYsllncp0G0Ko5kwiZ6g7B0kqgzuX87AZiTAzSHUBEYo55sg1Fup6Y8jgLnjQ1AR
LZ2eIWH8VXwSvb5vUBe6+6svVukKJbiNM4AA/VLDVRXrIcx0I7c0quzlScXYlUNFXZzReAz4jUZs
dv3HKu+8WfMtCFYrjhmxrP3fR0pP0w9AbbajfB8Pr6pzpNnaDQR0B2EqSHGO0XB8cC26hwOrPYqz
sFzqcXU9/Z9SIeRyMpiGpnrfZpy1wK/UWE7fZ+L4LjcyH9hsS7aE3PcG4/T/3Va5ujEU7P6D/rUV
z3OI+A1w9+HayajAME5+2oNFJAfM3q+squHxUyrv9mTCwWkZGZaponlaqU3b/zTPV5x/p1YcGuxQ
4sb9fKXLIe1lJoS3yZkapY8xSuHHDbqH7fPNDrY/wTJkIlRculwokKIW9V0em1dHxB8tK39ATXgW
Rr8IXNVfJEqZ7WWJsBJXIN2CvpQ42RYPFdwqbmJaz6RJvVOgXp08WX0YjY2+VYPv9pnZ18yGOYTe
jc46m4I0jCEdULUfT1P//2Qlxt8pkaBUoTaYtBmnI1jiqrEQ50pp9jwPnNuX/VZjKqZfByvxv9/Y
hg8ZFQg4XO6FnCj/vi/hILu//pordqa2DtJwo0yv5uDGj6YIOQXiOIeLJIg+xUK100CcUawNW+um
Ek4waMjzGHLRu7/ZcZy9xiQg25MZwdZB4PzfaMp++PKvjTC5+xRJEw5Up3go5POwo1qiDBqgDuex
xEg8aeyjqowXaOXbeDGqD1m/O2Zp26fzNKEQygbfkUM4+VCLLKxQiZCL5VItD29ITgwcGQpKxPb6
nlueLTWsghCPUtAysA5+nxXBCyM9POz9Bjdjt41mOb3wFrtZhBLhx8PAyoumMxKLko/vFTZXSw5q
mDpEtoKOrOmTvzae8VV5oeNnY0imZc4+eEXpzhVgqQSiAY2sMaRLcDIcz9kXWziDHR3IlsI6UsPa
uGJXTbEB7ltrAZ7iRWtiKtKE83/rFB+OY1JcuecEdJHaIgM4ZFBFMEPnWw+6lqCD5RbO4PbYvRsB
oTJ3YU2qGKB4ZGzFDb9tTlzJwZy/wnKlbE+xHk5oW2CE1mzrilBxjVKnmjfgCJs6IODoDrRkkrL5
iVaz0yFwGIVdPk1cK6yZwDFJf/DSGK4P/ASjRB4WPG+G9vV41bU9i0mL0aVq0ThrjY4AKn5uRPZZ
Hjh64kVUaZWzu9FM7Qz8lkGGYrKQX1wgfNoY+xmuYKD7bChv5S61AP4YE+Ggu9T2FmJiBACJ1sV8
WgQ8dwBZa+mqCH5G13jzGISc6l4ydzy9KW8kKK1yLyLKidMGuxmmnCWSrbwrxSGL09Lp74iAydTj
to80aYrvLQts74324buUkpXGRcG0XakxPewTB13FWJZUoErWwfZIYnil7bicc2Vmce91PnSsZ5RE
NQX0o4tTZ9vnnrk7KGfvaQJbxMfgqh23gnk8RdFmPK2b4HDKn/dvtBS0GsqA1NdPL3iNi17vwxa2
8Yx/NARGEoggv14JKLV43s2W8ZC19kWeHhISsZ1NhlkhqMGWuyGboZCYlGWL0wKAalo5YJfV6mNw
WH/sfAAtMHeob/EQzgmjZd634/hQ4T8r2h67ZVaLj9xgYX1ldhne08Pkx1PuoeM4fGMukStbu8Zk
fBapfzKER3epMoDk28UtKVIXc0mbwDQDVz8Zk9XCCgqVTq1Hgo9yhfjLHMD0K8FWrcu06oA9rxB8
xGOUcNe2epshIxahcxRsBb8tpCuvjWEMxdqtf8SR0Ppt9UP44q3iYJjrL/rg9z61xTZiDyvki/F3
6BXSA3+sWrDhl0H9CMEjhsWslnLV1+d4pLTK+wDdgPojBnu/eOY+I7wKL82yD2Dhadp4pbEnzSG6
dHamty4D5xTJ8mDvwDiNymjKk66p6cfHUd/1D7fbllp9a/rPnwjd9TtG9LkISW+Tm3W5EL02Q2Se
FLH5dqBrp+EfMkHvAqoLmidhR8QNZ7C5AMdVgdTnnVVs8GYhNmQFC2u9NBvrKTWDsAnc0veo3c8R
5MsYNMCOcHizwWsPFzfefrzwHkbLQXzJ2WWeG542HmFeiN7dUckAvz0sRhSYo10Mz57MpTgaWnGN
19CWpsH5Zbz+77sicPnoCURlHh5dTChA0dJcbKD/hOq4IbRlqSeH3XY8m83OGHpvH/cRgknRKlIl
pi5rEE0Ncgmg3WBxpuG/g+XY4lDex/mu8EVwWLZ0gh/KgWD9mDWpCMQ5h674nWZmMIQazq8E7TYV
HwIAcaTcQQLHxeWNDDX7HwGBK1ruRfGdj+XemicRq5t8Qu8Z1U9YMI8HqoMnPU2GggPx3iZDWJHX
WO08ujTIjbkvMG/c7kIGnry5tyFv9kQSjmpkFmCuRoNSjE6jCGpyg1HdZ1OKKCANERf2gqo5272A
PPleS7lYcd4OtjgNJQAIcfv+qQaDP+wY9TR+ZSxt8n+QMUAw0EGkGCeWO8aFTtH3KoVhUaZ/l5t8
E44/VZYFJ/PIGvibPWiyMrXftTGBbJjPLaLTOVJXhSfgc71Mww6t7DZPdyY7TxnCxXEw9hs8gdqU
MXHx6yZVOb4EmR2iJF+MxTp/ipyPRsxA5F7zDhvIgn1yzn74wNzuz19c0UIIlIGjsXWhtMbq9VrJ
OXHnNw5kctRAEH4Io5XnNSWSFDuQYxSnC+SHRQTXHnuI1i2FdQib/vyrpkXTAmDdAIUh0l3hJPR/
R8PFRtX2oDtXjByNGXFoO3/emBp9vIuS4PbLdpizqyEP+rzdgAeeAPxSYvx8NigSOFcG+is7MqQE
zXciYWdqO6U56xgOtXjXYzmga/COtkgs2vwe46QxIuWLwNMT8S2nd0T5DVcSEoOtSrLX0dYIgHuo
iC96l5pkFnL/POvK3NnYvTN5+a47mFoxqHUpgZi07Fkn5pV8XtpCHsa2T4CNAFM+VaK6gAQfOnry
LtlJjJkkOIvKaj5steTynX+57pv1iauzfWEttGjRBoPn0t1+/ihADOLVsvFNjRat0UvhYTMGV4ul
uOiTjXuY8j2JADKbn0CaxgL4CGLRVsz782VTsx1nfYIQBtO6FXgAhsgqY9TM/yH5ZrN+wSLxJj4C
QoEDt7Pn0IPjKNVGLCwLyALCnlUT3+oJCAYXCrxKtYa8iWPM/p954nt3swSdgVBu6afzcztmuL2S
EkT2ydWuJwP3iVAKJJs9fDQUkcB9DO0sJoVZ2fO3kIboyV1lYRAErE/E0LvtVJK2Y/oCUP2h7CuU
xoYwN6NuSdLlnpBZ6U+y7fToU9UX4IITI67zly/6NVi+T//JYB994pOUWr0MF8g9iVTruBvGigta
2H1IGL+umlzLVPyKbrL/EDrWxcuF+inOhMmCR63JwVA8lBogTrVmbteVjJ/TJquHxNbcotFYvEbQ
znJX+OHn7lDIs3bupzqJ4UC49ZmUmJHnbsy6Cw9ovR8/GL9X8fAeUIuR8N9IN0vsbFe/oXJA5OG2
UqMudEHYVh8XuQ/Cm5Nt9O9KlPBjwl8FQwAKDKPIa19CiQDQK8ysG8C6I2ucvGgyk+wzfnCoU6y3
65mqGyL5fgwHpk9/WdRUC2kAkPoEM02j3WNYiPLvpxjSrivRV42hAYTITi/xYRgPkEP96QMmvgCs
6XdhI6IQggCoh59X4dGORA1M7QnNyqofXFycsQ9E81wtUmmaFJSrkbY99NVCdUJ1ru4R/yI6tWQE
rb9TxlpMW0rliGORrmWuK4OwcnIVgHo0J7cSPRiSfOMRfz55InA1ZJvgqkwlQC9nrWa/J2UrAEuT
4ZO6Nv2P4KEidMqt2KCzjMj1NdC6nyIbyviKTwX2IS3HjAdcynrYNYGLDWxSwuBfrTN4dmBDo85G
FKQ9UflXAJj0T+jS/1plM5BmGwKOCTglxloWCIHQ7Bwfdp4H/ulF3tzhk44sVNE/InjYQkFChwFB
enCPq4bqA6WZmlt9SdfAEwIrQ3cqVRPMq0EIJokntrQrvUP496bVoM6NEJMEP0gLm9nyI+fY+XG8
FZY2NdIrWEL4Hm0WyI6bO7ZSUaIFtCq5AUdCceUZ+/WrIka2yi1YvrKhV32Cv5zxDgeqUCVFU2Uc
P98uezrJub6c3MvKpFZ2lpR0slDO2O5iZgBO0BJ2JOzsDU4IbDZ9UQpi4xR/luTK//cb1YgKUBL7
SDqwpWD3sE0FSWaw/bJGG8HCAXClaFUeUj5O/VGgtcV0ya/erilyQeso3L2WUTyCRShkoX1CR/y6
ttT+jWcB/KYnnc3vu9nCNty3PDq9F3sTPhI+9Wpqo9XAzn/rLvts8eMjQCmyuSajenmIxb/DtWb2
mUXOOjy/mKFAGGav9yovLZCxE8rlblvSJ9Uk7AZmRUsCEjItm356/FWiutC95gfSpe1kKu00g3Aq
NoEcFMKgNDh2uYW1OrXTlkUkJwS4t3B8O8pz5qPXXYlwMGr+qZ5cmUD208OPO7+LO55F4NUMjF5d
xCVp9Gxj45uzLuAXGl/0GUdIMttcy1D+2XIig4lhsnwb76iNNYWUtnHWU5PZo0AkjeYuYDi/5h5G
e9cNifjkhHZbJmob2dEFpynt3+OrgNxrGHaA1K0U65W2yGjFTBnJn27OclyUjgG/ENWHCD9fly7o
Fuq6S4uMB+Dc6f5T8A6Z9dZ5qg6Z0y/v5e8HdgFtlT9Ut30bSgI1r1SZR/pbsoGF83auu/bEwtCA
Z310vjL8jdYP5AaGLZZ+NeEIoKGmTafCiCHnaFf8bQVI1q2vVgTkcMUY/hLIkk+/C34/KumFEiKH
sUc8tbufQEtNfQQ/lXo4sOLCTc99iz9ZwPkt47vO8aeEoXgcgki9SMEhVNOz8GfJlxRVDBpIqBhL
DVGrxd0V/DdUh8e3a9fS8sYtvsIeJVyrIbjei0KXAXc/LEg+qq4HC4n8l5z9Mwr4GkZ5Bj/W+8/w
W4nsHSzuGn41L1pSIGLzHFJlJ5wyZYIoE3q7U2LqyxyhjXqScPfnIg76/ZP13mIgegli7vKy3HKB
4w0tvUDVcR981EoWv7EC/05B/7RkEnM2TX7bDGXr1xJ733DqRbUXw5UkVYJ3EgryRhqtAT5mJBey
DhaEvL0u2AuOBt9BrKGZvMhPiGovj2iZzVivR663mOa9ThYurURqDlSNr3y3QBK9VYkmNGBRWl3M
ItxDBR99/dbJRwYuEAV+Z6+0Eb72Dtuk5dkH9ctmOG/rFGDxlTUfVL+Rt08i4IpQEg/Do+ek01lL
swFf1d3BX7gdF2KBLBsVKiwrK3UqisCvTjDKIds+LJ/gnqnrvRsZz3muRbWOqMS2p0iljMcU34wl
MnBtfd+UY6EGWYJwyCGLf7ACRW6UQbZ9YDX/kL/bV5V6jo5KmEQp0LaHGtkYQAzaHgYGv0RQD6rO
zpErRjM33ICQRDte6NShn0FotFRyY2g6Sz3ovZNmk4ugOzHpaDqxHaa+JS0ROZtAOuACM5s2Gm05
VEpsjd+a2RFvu9a5b0QkMsH9CuotG41AAbCupCef2wPlQx7oUFsitnrEkh/F2McdfgAG3sEDCkIN
2PyB/PrXoDZNazG8OjIP0uIUbAIev56N3khrnUt7kKW0driW0TWiDwj5yoGbeS9Zl4rEVnrbU52z
9AJxF4ZmiFA9q1+U7roRWukHMeNTW4R8JcgetS37iQas2/DuxP01jPuYZCDVk9zjBTrEWqgqWyqb
QgClDhPjmuNnTONdgt3DqyXSTw+3b/h3ek8MzGujCVQjQRRitaqWmZtkWgOThnXYqNvvbLKp7oq2
xsSFQmhiLHo354k4/1acVChdJbzVW0uLw0NtooI2YWZEFhumXtMjDRSiodlAy00WiRvoIUgBYXb/
Vgy/DqXSNwla+AREqDOqf0dMqeJ2xrdeuYhdJqAEDOIELJWBLs4meH9mWqFDySxjB3f7s2ghOEjx
HjVTYyBtlat3CVgY6U3HQ7jj2yg2X1LiLN8f6NfwIAmRKKtQAnpo9XoYJ4c/WqBMzLkMKm0R7f8s
++rBtRrdcXatwSth41veERC1wXV880w49FAKUb93xInraiCtBXy//RJ2uvX0CMTltjcY2dmf7SsS
A5o9tvpo7KgFK0W97i16s06mWO3rBFn8ypXU4TfTY0MaKlO4firIgjDmSsAOHk7I8lsTYfzpyDh9
hJ70Kc1MHg1AP+knoN6zYdt5HSlVXU5lTq5FcZasv7yv1YtQlq0hti+dNx8ji2LqlO5jfV3ZqPnf
yRPfl7pkMtyU0b7CgKMFeQbal5XGtxIX1UaMJfdMEMpW85V7wvmyGgX/6nQPVufdI7sHAVAiUtL0
rpZHn3RpCG3KQ6hLaQv2IXqTvZhpr/KjiDEFIoLVVSsQfj5G5sbGoXZ6Ng/fUqnpo88YY51yLbmK
fOa3NG+gw4cqCEMFZx+GXEizQ8yMsimK5svFGutO2763srG1VD8uh77gj1d1UNooJqRLb7PBPUh7
BxtpUMuRr6OCmauIyVaTAUIB8OCawjbEiFKKK4MNEquNsiO5LvCKsTFPjm7X6IPMz7fJ+XzE7tBm
QvUkx7ZOyfZxABwQypEvv+MBmVAvQk3R7YkQDitTbCOfBZJrK8v2FThMblXL/f+yKR6i80983Xyo
t4LSRM7RHp79FKEg/aJFbz76pVOHygmSgeHzt9SOsGe6zG5lVcpuA0KZLMNQbuWKUhcKdC6j9WiV
cApYoxyT7ZqbSI0Nr1yxmZlt6VxqVLPp0xSK6/qIeLJmeoDxER/vBk7vCrOMUeD0y65h+DweVlvz
XjPPv0Y115EjStEblsS8EJtQcH9dEuWYM4ZED7XFbW/ih2mkl99ETgdhB5jEb2I6cGhFKgg4shSY
2ck34wJN9coo2OByWGemKsn/M7V46OeaLi3DbkVuYBDSznPOkPWxYETlsPodDJeE/nlwi3udMwnw
yOZVON/sZUVxG7Qk5CWCLJkc8AnNgj1oejDopPgkPJ4YcMcyYh2txeRRkjIjlBMw0TYiHezA+98q
KAPs01ASzlTOXf0MYHl6rXuLrQweMbMnBT7GMdkrM9lDwl4RmIGX2WmyoDlU9iyMok+LtrcV3oOB
5gRSOZC973MF6Fwc7o/pmuqlCVBa4X4dbcISRPKbePOTbteT6Oe3ZqgLZLNx1jlC8MpkevvKyCGJ
wGs15/9+fVczLt3bRzKpIcMPxi5MHWukDlfMjMwdPPFmSKhEtNKNLcD+4dvmA1ZHLFfhQqYHkyT9
49qIZpQ7FZuPJIgvT2pBntqxXnxj28EJCUJlqV4fsN8gdyyI1kZiNfY/U2lXCbjIXXwQpM2a5ifn
puq5TDdRnaQSNduHdyAH0CYfp2nXRSrY0YPh4Y4p5nJgFBalr1mwltHg0s1u8VysRpwGtA0qh5W4
zA3yqSWU5yYToCkfG/Iyki4Ts4zr32lVqjrQumVBhDO2+7H5BoM0yBZb+07RFcxGAAgLuHtT/JYj
8m5280CArBLAOdeaJkqM0fEtnqrPTz2qygSTJiErNV69URAhR/aUV3zJaTqcysMxW58QQw88kpcV
yaNqZGHH3HUE8opek4w2qVf13bfRXmuMU2pOvaysW0utmV5H8zU5S9rgexLKkzZgwID7v87hCyf3
T97cfq766Xp3WcPI0D1gzNmxSftlhNz41GyRlDaewVIlZcD252xg0JtmlmLE43YNjQ9vqx4km7qh
56ixYfqv7x2mc6fWn6QxreovzVMNHoL6iLr7V0p5S01bWanWSF5J6FVMvMWQT3E9+rc4HiICGt75
WGqPaQTPA97TdBHE9678XsmT6ixrsMQ5AnUQ0WgwtzIDlNZaK7lsVhnzItC+I4a2VtB3qIu/pHEw
m7ufK0TeCMowMnbWQ7k3B4Hv1fLWTKjsGHF9TYbXJ+OlxfRilqNJj9RzjyLGquVDFGvQbAqiAsmr
4X7Aan3+e0tmi1uHBTq1VsY5Pcmi+vh2w2/MA2WQvA/bTHEKoKgkpuBEURVCCJYUBTSshdRCryvU
UGDWfwUffmYOMrJ7OEKcyToU1dy2C+FsdtKKd8VZFavEw+ttyMw/BjUC9xd5b/3KwQJ+pcOBfD7G
W9cgXjgxNGhsB6dQwWfyWs/zP0na7y7NabN0mvjqIGF0AMP6l6r6mwVU2WKFznWxokHKRv2qkOXp
uz61lW1XBxGMv1yEmnK8PaoGkXMVT0DVnm2FzsHd4YDm7NRYzGMkeGWA6O/maFmaqA1LY6V8uHV9
7GLmj5k/KWhYfKk9QNnJYz1/773KpUZJmi2aN7veFY73/XPa7Qo2cM0FoWtzrpKFK3jGmYvkoWYS
9iLR/LGkoi66QjepExI/m731UhcOwWQershdXz+KxvxHytdxR0Jw/EqkU534Xq/EQvifhWmzt8Y9
PWe1yvg8Lk/IL+Zp3gBT39KCbH8TbNZi0dEQ7bpEYNMiqBPVAe6/YiuEkREh30xDF6g/N5DS0jM/
HDepUkKTPzLoXlQ7TvU7S2NH0ah1sxiJljZ1KUzkBNFgR0z+L0CvqEGyHKkJU2bmgSl5/L9gceHL
gks2aBf0nEVk9+82n1qPXbIlf7GHxIspdysdSt81tN5kSDAqhfVYr5iEfUtNlkefxW/sjRvWeT+a
7YLFqhxiOHXnN7XFboeaEgkS9anO0Uzh6t5ndFcEc03H88q46K1S5KZVqmV1QYdbTGy9CR6yi2ii
yyzsqoyS/bjAmMwhv5gF0bW8JXU+QEZU1GgCIA7n2GtjM0e7VFv6+QnNUC5oy4Ud4pmapdBBbac1
F7wcQi6NHS0NBj6vNKJfxrCt1ns/yZ0FaqltGiit+PiNAeAL582tze5IVd7ZpNiis0qbjjBeF2+5
2GnxJ4BzJPDUK/C+aeZJgqhfX0OAXDr5Vidl1GJp7Ma9qSX2SUDk37T1gSMsVXpBYj1A0WSVSv5u
se6rJtEeTtI4h8xa8fK7jRNCYveFBWJpcbMBqCE7tEA+SFhC+UpSwQl8rJFBE2xft8Fda6erixEQ
Sf1UYwP7zWu+rOw/2fW/KziK/vfeVRzb79T0rwqaJHq7pAKA0GUNCZxNxwnRfFMiAp/X2tKrT/zt
2aBC97RpY6Ti3LYRa24tBIitYhyIMk5yO6iZrp0FUMfe2VB+1peaZCxtwipIFwKsjUQsuFk1Dllm
wfbhxd6U/kygh6g+d4B7itV+8J+IFNO/hcdg9Ocp+zFY21QiwxgdG63A9BVF2i3//Oog+l+x9cX5
rJR4bqI9m0GCtwgkHOJT/PAySvSkRHrxgdLtFIjtCeBGyXH+IedJO5AB3l9ohFWY/S6L47rxe5jF
KHsUyY7GPMPlAoB2YJjKBsli38kaTKaFMY6tmIbXxtaiHN6GimGYaVW492j7kd4vz4mQooJ8L6KB
Xzu8g5hFNe5pQjjhooojDrhxJJA6zuf3mZOARULhQXlb4khkN7AR9VGvxh6SZlZGV49WgBwRMP6N
g6CvU2p+wpDiDkY9i0BX0v0/E13+FTAcC97zzPcUwJijAEX2nK7j7WPN108U7sJz7PqeVqcWt1ah
VlgE17KgQXq3XApNH9f3O0jDgOltPE6Xo7ByHKEeQIF7kfags5ZJHHPVcJe160GOpd8fj/QUbaA2
JtO8US6q0TTMs7Um2dL3OL/wdurpCGrgcTR5p2M+ptTeOxsyuVGVX+GpA1NRZI8uD3GHPeJQteX1
3szELoZPo4BTmzcFGTcS8k30H1i8ABQwc2teJDfUO9CC3H71hkafTWFtd4Jb7xVK1n073xonfFsv
F8d5e9WER7LUoYQjTnQ3omTXeGViTqjIzbszbBOUNF/1JjpItQHp0MoByK0DKg1b7BKoQ9SnnBUA
IcxixoAfE1FNlmXUrfBnb5Rv5FAuIAt+4kSnk7P1Y8OYMKgljNVv2cbAKLbt+ik5pDjRyrhf8sNN
pxZL0yZcFvE4ox+Jm5PRn2Jb6TRw3Ut6W39lPlDIE8pfGS5JHtrPG/hziUO8HCm6Wbyt/SoomGhq
5oJrjoo5izRXVPTynVg/tmmkV1XgjYndMGhXOtj5+MMLuWJA06QcBXTb9s9LtQByHNB4lq4j3BYc
K0I9ohEz7/KYdhdztbqIM0dpK6AnJKxWzHo8nTfp0/vsB0lRuyyAR38Gywv96hba0H7IMFgknuXY
YGMHFAQ8daP1CjUhe8UMCPxobjNjjc0N098y1SthdO2B56P0sR56SZU48Fb7I/G98zuizy0FTFKk
wpsEaRBWeDTzHBA7rrEvObmg9Hwx3NU4FnOUPsMU1v0HfsYlS0af3XNGrc5CEiU/6YkPXOsnII2I
s54tikDj+EASPZOy5MlB+GnSIblms0Xc7QbLrSkR670qyTTxCqgbDUuAz/Lex7pRVP5bwpRSYfHN
ekI8D4bOkntK3JGTYBLQUAt05rxozw8kXy5RWGnoXWyVqodpcFECqBdgkyfuexGSuddeuB8fkA6q
CtJHtuWLYmyMqpQJBmaXgN7jzuuaBlastKF+YCSqD36ioQn272JgNoW1Wb6DCJ+5stZr7RlHA0St
LfrHqf6lvv1IsvQbQmG0LXZumnNAcWAqte+2qsmtqS4MLUFzbloE9XFY84zrNQjzD2xL+ghLOASL
h+IXIkD6zOpzXP2Ed45UQ5nA+1NmOWsgLjEI2n5cGfbETne/8dfGfKsARmgCq4criF964kLLpMyG
OUnQNAGIBjlqkDOfBDQ2Rsxz7WnjUsDXyjP3pXbGTSZK1JQJGeolKDM0m7IbIVAPwqipHcB9RaI1
s9VUan9PBHNLS0ehuhmQo73Ox+zi1A6o6iNOgwFl7kw7JTn8a56xPgOdUfzDR/d1yNcTaIxRlJ1N
8eVOVNTALkySRLxrCFbPQFQcYeXDftY7eMbMteG1o/j+rW+8/sOUnmTfOmHJgZEO4m3M3lkG82x/
1UKiXhMJnW9Op4ZTeRN5lp1TSqimgC0rhsB8nTR0Ylr/Y7+MHrll0ReFisl6/FNaVuVt6uMJGsCY
hhSw1fcqu/S/k6t14PaD6SY6l1ajxcy46EfZtekLxUkDmU22sTjp2DrmcrgfJQnJKcIjGqFOZzqR
sAa3z+WWKPpDhYg2A9IzSFgjnY5/VDvwPY3wSqSmA05bkD3i6QcK3T8/3iTAnIYbJpeJ6IRbzL4A
SPh/lFlgT5RkQbSF+Dz/3jnAAp51cXNUcuaYm1QYxDPYUbdaZiql91uFMpX/9UF61sX8JhTDwhb9
sJ6Wg57n4O6Ig5WB9Jkh37v569Xyotc45Nzz7H3tHrulEAGsqt9I9xA4iUkSgnsRkyuSmlbv4yol
3PNM6Krj9tHjXw/a5tEnL/TjaNjXv82yNAr7GFD/9cv7mouxtpsYt9O7PQ+oEQBnYbYxCu7+hz14
kD0fbYTed7ziANFAMGc3sSTwaYenyXLUrN/JOcOI1gqWOg9JDMQ9J6UgY+fZdlMGLpkhbaOjhOKr
2aKjraeIuevw6ZjqsSg7Hf67chWbWJv9dYGrQthYtitFc3R1P/ooS4uxNIYhNxrJDi7yaJ7+c24P
8Yrvf0djT4oNrx0dNinsJBlYzS+IotMM0aIW5zhQWTqcOsvoy+IA4VZCS9gBfUx1BiE26hzzKqOE
HhPNhcsjO1soM7keg8Lp3VLYIxKkzX7u8MrhPqk2Lwc3N0T9GifVG647v/IlLaUoI1uSVlSZJ0Ej
CxrppT8Px6IY7967JWhBHAPOG5QdHPgjBNNwSUy1kz4q1uUBKDjQT7/JSmy3E7V611er9qctlM8s
7FHujaEIazczbuaOlxm+BAdDpWCEa58V/CDE/iWz5byR/XZS+08ugHj7sqxK12DeP9CpX5Ois/0o
xYpM5QIIDE003CRv1kwJ2WevY4TRhRwiLNcI4GdbpSCNHgDqOV6lBkYT8+U0A1L7S1pNQrvEZOhX
tNJ9fNheuHDmHgsnGpQyJ/ibwS7eHR45Qnv7qWvYQl6nTZgq3/BhVBTBO4toBjTEM2Uk+Bci4mET
+61YNlQ0teI+97bWABQoSdgiVsQfp3HHO9L/IlGIPnPREOra4CQJ637Ibi1AtA4ylTYXVvDMaWqK
vietglBBcmkKZ18cp+3LmXgOFeFcI77K01d50TbCBOYNUf1CuCsJZis/5WmBCuhFYHtwQCjiABbH
Ef1ExZqyXkmKd6pH9UNtkzTXSHSXagKkQfj6K5HfSo8MBzHr6bF0PGQhE+faYTYF9sRRUUxxteyw
WVHSPAB1btFWoBhMOQPXHFID/ytjemOXRc+yuygHsO0paisBjY8aGpthG4Xkp3KnBIh5aDYKQH++
DV41sEhHre92m/mzcVD19oluhKJwrKQcRK4xdvONhv2kuVapVGnbgLWuIOT6D8vLRqLJgJhqmyS1
H57SJEAhtZ6nM86hBVhluRg8P11IRoQoRUpSDTXl6g5Pa+psSTaI5HwWt+eBstHdNFBnr7ybRKPF
na+kHbCkbyf/zRAoXWJuIMsvW32z8u9X4Zxeazy64hc5rg7z9sk9ALucj3ynfWwaLhkmRiljQYfE
fbrZobxnXhBj2Vn9bATTpdCefDrDqb+DdEXmZmRsdFyGTC3JRKRUQG9D5gitz37lRch9zyfqQhI2
IUYAjwf97itvvLJDRKESgEiKOsaZoTlBtjIPJ+Dppd3YelWHc9VG7mbVdGi4wmfLsNTMHdWL5BK7
nrIeNYpjnab4eU/vHQQh2GojhoROd8FvUcBckdb8tWwIlP6Y8RF/nBBq1kM+/a+j51l+lKEVKPu3
lgo79w0WHE1bmnV0NVUqyp+I8eKNFv2zW+E4M8n2IUtAgatxRNtGQt5LItYFTPs1b68UL/7lTurN
xDTN0Crbqxw72ZW+US7mAYsxLdB6fmV/emWC9J6To9Tn1QmfyvyZZzOVA4EhTUyeQ61gwqvGz7Q+
MEDVZIcSEve13oSV2fyzfhZwPcm2hl8ClqzC6HrA0brfx25uPDu+om2olWrLJQ8ItE+ZQ3V36x6r
Rxk+55//7ikRqOwRftx+bVH+rWeCzxgH96HJQPuDB3AF0OeFipOZet8T1F5b/jO9R6X+bFhNGU+u
sIQp5zYFN6L4K+q2Y4dkWPG1tlanbVzRO+4QsDvL6ATYpP8EenYq29D40mH9r0uAZtNXO1aIgf/O
hPqUpa2tD3X45S9eo282ksEdpHCrxxVb1l7HtvstjaR281GxKVm3ewzHpy2TmfYhbdhdqGiZREII
jzKXPUN+BWmzVFDS1/ePjPQXKKs8CjmaeneRwf4UUPSjyWPTdRnwGAGy7JzzhOGDY0kaJejrVdSG
s1K39Jk8lPi9a/7nWF8nyTXwq9EfukBPip7JbkGEO4jPLJSocliVX2wk3IErgn2jazPtRCLGOWUR
KJDlyMFICQ8iT07qSEjetBSWsoFado2q7KUjyLUwNeh6M2nlk9zozBzLrQ97W6qkEp/HDnqnqaXU
gHyvlCdhkzLIJ+sUhR0HHlZr64XSxjtI9CA23+Gya1FePnh8IsqWbfE/DNquBQtmm730DmQXZ1UK
5hFJAzdXcBqWSAxRKqOCSaD+cZLsbjaCXSma5jZBPuj8bCeqrGoEhWBHOXWMe0eJ+FiIqhqLzmOd
zMNRuXa1b1TBBxRkqYiph5Ke7wT8bKO3gMZy44ORMnhYITfsGOrVVR3StgucqaM3VgOJo0pZ6kG2
Rny6HJ5GHAEf7Fj55fHylV3Fz+cyhLBlHTC+uVjG/cvAHNZn2JNroCfRB89cR591AP5k6eEw8wRG
v7jOKBFVJVRIgcNgkqrSDTZpAyAMN/ltSVQ9t2zgTtRnYTMsVCt4nB6HmOAtJ3Y48CxOD0SOh6/L
V86yZqiNIuFSinnj07qhzwLVi08B0N5SqeUIxYZ8VbVJ83t351cXJdoRd8nt4oUeTlbJ+3O9dSHH
cvQS9Eppl26j5ZmZZC0tr8hs4kZGKaDA+KNpp+LwtN1WA0IoxoZ9WX5fhEKbnmsSR+pAy9L+CT8A
s6vr7HO0aY/TZwsmrgW+RsSeDTVqZUk3nrc4un0Bt/Tl9dNJHTkAwuoha3HDjtq7xqjnOgQMgOxt
chzTxOg1vR7TrBiF9Dt06cZydmVMQzwnQ7+K0UzWM7ri0ocDILM4C8QPtPKIiOfnrMkXzHdPMiNn
tkgVbtvM0V7SwGy0cONSoXRV/odTRxZMkZU2qn2+jLQmaUbGc78Ccgr1Vtyb1eIDY1e9DPhROak/
xEVHXsK5q3or49bqPVBuy1Y+wrTAy/LczZpeYvCidYNa6nCSKQWnUWMV5PJHAvLM8lHvzRI5cHdY
BriucE95TQIsZh9Tyf+00Hc8189Sa7JLQUOnUambXGezgq7sxNPcxscKjoEhbG+hL+QPIsFyroVW
VS8FsSZJUS5FHif2pzke/lKAtcYbjNdrMuE17Q8HdgCWDmi8FjzDRe1CV5geAovhTqbgvXXJ3DE6
vibsT18RLLx3bhGA37ZltZ5RziP9Pq7DksuCyxSkYeGY172OKKLbv9GRjfNfcS0bbgBkZl3ntOYd
1KXa8yyUuQoWQveJkzpWnuY9tUGc6IGIw9hWrIAoV090S76XOpQ+KHlX826Fp2YnhgtIWNhALPJ3
4rDYFAv9MjkZyekNWZ//WMF6vC8cHURLoDNdM9IYsA4hjaXyz1wzIJq4OVsd2IeDKBGPugbtsTAY
mX90iMVnJePRek2J/vdM2FaR3CLSNpaERckgtYSpAr24D4UrcRd/wKX11teRSZRbR+Q3W1RJBx/+
wntqffPPLezrLmo+xCP38BNXCEHWcF7sFQFn2UcHhoB2qzRHw79cmipECJFAZyFZZIR/QwkJf7ua
F9avQe2eZo98KZcg0TteGaO/NfF/N9DrrYdGCE1Revi4DW3jFqMRxqsskR95kIM9Mf9bf3yx+wi9
tv4SHBBApUi/Ge0FaYL969rkg8gef18m+yog3gZbYN5joQwrRbm/Wl6GkjIsppzr1ITajJgigNWU
XWVRItze6dNJNN3WPZziuQhBXFU9WBHnAklw2oJuouwi0y4pGt3Y2KBOuZhriRx40SI+lgxcG+U8
3mM7ZjsNLn2/X13OIakKdmGOD+XREhoSvcDdTAZFOUVzdkG3dgarLcQs2t4PnM4bgOqvEV5GBFYS
sRr9eiXg9rCxssCuRwHwKPHYwJymzrwxpkCjJltCkkbPnCUh2eOUy00KRQTdNlV3cqROFxj+yqM4
OzuLb1UBA77QKcT9LRL+HpUXeoM7nCA7mEb416n/e0rD0fRGTY2pBmRmPgyo7vcmDW3Uu5VXjD7F
3S85g9WgutVLJMV5qKmaE7JqsN2BEeGiT8ToqK7g1XDGJmYIMAMf0IGlndDTaICt5XwOWAt7s2Tg
at7Sv9H0H7Yv/mwo38WtCLtjo62QJg39kz9teeNoIIPC+HMJL4vKnb//bKKrhfLokPPOlwSRLy7y
rwP781BFBriBm7FOMrv+2H7IOUR4eOAT1gFMyGjmrcCgKIbo5l/ropTfwqlG0jBAzpjm4PZ0McaW
dqk6WB1shzqAEXfE8PYZm7aSLPHAzxDkqCaL+RyBl4v/Fz28XinSrgAr+jun1y1XeWB/ak0WPn6G
cjpajuLq8w+Ei9QXeLrODEjfHrxV8jBTJnTSTsjkUnJqC7agYq58LbDPzHDRajqEIB9zgGOBqo/J
Bw+SPQthdyeLzu//zBQDYjhtReh7jdVpOkLv+HHa2W7Ctz5fObEHxLHsWbSwEuFZshUzAUk93Z55
p0/uirSnSyUJKFM8V3UV3giw75fBEwWzq85kzOFWotLLarKQIQVAzlc1Dw7GhJIAPm1fBldN2vBz
s0ggDSuw9f/L+w5p2jVkxjB7t1fCa9WJ0WskiPSsq9WaNbOGFQB/tYY1uWWZD/05cPjBe7b+a9Gb
LAxh80n3qg5w+sHuc4mYRtZVKTZwVolyrPobpxLbZtK8ZbB2o0CxtzsmeYexaD8SrjaHhoDnJxdf
44IDwpFiLd6F6EIbCo4zWFRRFSRdwvxK+oR7/W/qCgZxNZvw/a66LnxgP1ZTi4ZAe9nvIuRlvx9J
gxzI3tI6ScJ9hGptvL6ytYaIsDeI3diOhaX+7kfFsRlVSxav3Z4eNMDuJ+9xpFV2bP8NPXnGsdpy
NLY04JdLIY+nwOgfUVMwZuzuOtmcrwa1f4ilm5lv6QED4vDXDf63kqR2vzEWiIq/puH9sXImzUat
Id+tsoudPqoHWM9dNSXmnmbUMh1Ras2Sqt8Jymc1y6xSKZFJ4S4vnZmwhKC/QrxdeSu5dZKcXp6u
M9i3nw6dTZbqJUKInulsKBEhsg9NQ2m0vmyED9Ni9B8BtFN7pC82yoTfCcUyA40E1Izl6ZwNWqHU
YX0Su5MWXyqOmb4nwiNyXAMRb/Eo3yMxSbuCvFkAqDcOf9vI+xIyHcsXcAG1NYVagcNl86PhwlDr
M738y3ASvK1YyPBFXUcSFZd3iTebROKMO6LUbmv/uofLrWL32h4zc/kMNXBr2qMlAacJuf0UJxdT
9V/27qE0psLg4yy+IVYvD4dKEREJVsB2nhLyt+Iza3wtw2kRdzJoLNgYpXXSyW9y2IZeY0ltTFYA
vvtqqbwERsQBdbWrZWyCXgRlJKO7J7qe8iQm7rQ+mNDnn+KUCDeGK845yJ88ndDYOy/YW4xZ9V+Z
7gQzxMo8xKblZQ7NEjbMGHxHC9CVK8EtmxglA+pwhP8qDd7CHdh3u4dxJQ+nprfkiUwo7cAH3JUG
HNlJOXJH7Iyd7rFJr420gKQ5r1KQ0YckAHJBoOTxb157FZdX/IZtHScDr3yCPKHZIJVmSCfsVpgc
+AHESMiYM/s+w6QmdShOzNyGVRyGKsajthkrpnPJ70V6W0EMqIQNX2gO8n9pPBFj6EueAymG9YxZ
1zXRrMBeeJxmWrLSs/ht+YC+rxam/BjhZHjGTdmKeOcH5zAhP06Zr4ZrGfQfFYBUV2jJQKKTLN3F
/LQI/yde63GhIQ4+T3jdWQyFhzJgUJwDMiXrHKCBdzL8ACw71WJtnfBxRQvblhgV4wsQmbC4cpM4
YRo6LJV95Kq1gTIlK5b2XANCXRjTR0usBkYmeZZSPET/BfWGgFt+p2ev1E/mfo/d0u3qqj0rIfoL
uDmghFm4Mbzhb4DNIg0oAQKGoQfOgibBdNQzMOFwS//b95211jLedQdOKdRpCU8VL1VbJgdR8YM+
2tsmPy5jn1WKzya+0V55ecXPGTO1HdN4OgsnOwm+y/kfcQuakV3ocMp+FVxwfgvLVp9+nHSHoe68
A6mH9tJDvSEmgpM9ae5hBv02Yua5yV7WO/pKAbDaXVGGxw5Q0yZtapKwKT2i/M/Vxe5tLfcDTNm9
BbyyFyXV1F0bgwc0J5WVUmbsP/XB/E/W5mt/vWEC3qx4WoW7FlybjWlt2EU/LDGCllXuErc/mCC9
/kPgsgcwg2oZkJG9HQ0gkzxlB2+05r5KvfDJRFodit8/ikPYLUpVnKggluii/bBM/5P+ok7heAI0
UctADp6AwwGIxqhlf3UKBULjdLDZIGrBfuZcilWr04oCd4hy+zIMheWoi1LtKsFo3PLV9gVyEBF2
NMdiJeiELml5zGDkNwDtZkUzGQn0XwE5Dbkio2AHGM+I5YD8lEw/XqL6kxHec2byDk8WmETZsv0u
UbbPdG5Fmry6REV4GA9XB8/hpCPcDcyJaLXHEJNkdKjZxGHG8DoeGP1T3LX6v/NHhdHV3EGbiqb9
nw01ZShP08Oacq8i8JhvenaBdbciyWCmf9BZDpsRsFm19g1zW17G2/y3kbLO6LzxA09stvKq90vk
F2ddn+qPj7MDXCofXaZdyN5aRUZoDuqCtYjO+x4XxDJ8V/KMM1FqAnE+ZIziQGJftHjM6PNqGrxn
GFqMTMcsQttxsYMyNrWaJvsVvGyH90xqRsMQsOe58as12ZQdy3vi9mYvNtOEo8p7Kkxa3eCB+hnG
uCQPrWn+r89lA5c44bm+ex0Jax8wm2RGVDb/wyVY546bFjdu3flewDFcSbGG2EgUTcOHPabLarM/
Ocv9dF8gD8ykEXyf+BAwSL9sWcTZUzYbkhODZXZHkMHihIgF7PY6IZtwDTwR1QwzPsBhI5OwMgqz
5k7QePjr0C46BBTa64yOCIbT8WbtHHkLfTgsUstZIGXWjK+paApo0V/qipJlkD6Pw+GZOeWnJaa8
pnGXZlfM1kEwZOdJgAK4He4O69ZGFpj6OmnZjCpSXaG8fTeDyiYV6gj5mlv/OcslcbkbtIF2ky1Z
3T0muXihGnhhgWgQWDwW4oAqwRRssHpT1SVi3j54pVdRBZQHYsYD5vQ/Mo/kYIhyx5x66t5ulWHt
Bt4mlZFANPqIo20SLMuMWxP0QIeOi0Jtz5YO2Fx9H88lkcya7+QfzAIbqrsbH75uEZ8ji2Uajinw
GOWId1H5xRF7jeDVYY4LnQrYB8TWxWKGYVYr/mmzZQ9puPilEwrEAn0/1txIv6QpjFSeGBXtFrB8
Sh9zBV7rAuIOCzzC/4rvaROnlbwuhKqIsboiHKJm6WUlpL2gSGzR7jZKkva8CFe7Fd/GOMvhaARi
Ahw+q+SHng6ZMogQlqW31Lb8N1Z5aoNHrdkjykiIEAOWNcV8BPeBt/tRkXofHsnyA/sPktCEv/QU
CBMeWZFieEOeBKdy+scbQ8u5of7llnH6YA4OCgT7hQdV7o0PH6YLiCQ7N5WXsWs326DRYXXgDNyI
GSR/e0hiJLHEPqZWcgVx3Tay3Vaz4YTgXUzt35NKq0P/Sao3SdwvqAeqtc4BFJof0KjanhYNYPsJ
M8AL7EtwYqjRxgZT44TbCOpzdooUp5rGkRa9ozWNBNa4vgV9qbvhcmOU26RInNQLEMWiSIU+I1kI
AbqWfGgL8g/Kp8c75YQIwXBQj3Nfsm3f405uauh9vNRxzcX5B9YE0oT5ohTjFMHzQ25xwCZJxwY1
ojCiz6t6hXFUrlh5VutcRE/smHQLoJBLk7/CrHND3RdZJgJaZe0SyROn6LtTlMUGUEkJRhvFOeP+
gNXH/d19ADmZ4f+iAK+jxdNsWOKg9TLZhTeZKtLflZfol9ZxabHpNpmi93FdE/n2KgJHioRIGUMZ
ecsPknNHZC/C7NOb6fe2WjGmnzyF2P2NCrFm1JM3ltPi4QfIXignNP2HKoHYPFPSR6jgywgJxS0A
YfkMJLJY7VfdrncnTiliFNUF0/sOVOiZfe6avzy7bPFKrTR19F55vpsV5esh2KqQBqbFhcq2QRpC
dQPvMmVbVr0rw7qboHfMOtUVKL6hN8D2hsIipVIDVjMIt6YFc4PPxl5CO6hvy23E1RTPGUfrM3Oz
hyOKbpyXWOnGWi9bK2sRwcXuPG34jO9Ld+2mTSA04hb8Pwlf3aMM5nt7W5Yit0/d4aN5zpVNIGby
gVBpStrgLh6fKUkgBDaXoMI0IUYLqIW/6LGV3PFqT7IGqpaPOHADvvpFVawYI7XLCGsUFhCJjM2P
7mHL8zBoIwQmCVF4vkT9P1ywyKWJxtIqbiCKAB5+9ipQa2d3UucKqwgBhbmAQCa4iJq7nXjYTs6E
5XXiiWGznqisW1tG9I418kHZPRBhQawebNUY885rgy5/UTuHkTlbBfmLXHXD8m6FfJRkXnTeYzu4
LI35z9tO/2PenL6cr3wh6S4Lrw7QxXpUcoyaPowSUt/cYdmRc1jdMOT3MMikTSmLhiw6qOsxyib3
4re72EvJ3ezqbGnzboQLWKkjBvF5SBxleusZLS3/LaBYfagnMgl6ko1jSm66oL2ofcMV8h/jkihU
+S0phqMxqe+UoKZNzNqhyE7ayao0Vr4Xct4Ze14s6DQMKaYHliaYuVc1x6DEfbs1IBoaeG8kBWiJ
7H6eEh4zIq6YdorsuCAaJZYPVes+Jg+mLfPs8GUWNLkNj/xNIL2afHbSnSZWZKQQJOy7Enp+pNWg
/PtqkoPEDSPFLMossPhBU1o5ql2Hh9bpsjeWisr+D/NrlASpZDLTOaRXFH4BnsSzLlClYaX4pV6z
3yB1Z2a0Y55py5eRgyksE3H2H9UwRrG8T2dHvbjWunMLWAVCHalysVzv7jIlgvhnhKZVakeWHy1l
Qt2BW7VBbcuEmXjdIlb0MRfjj+klOWLGNCzngdGKoCLsmQZQzkey0IH56wXL0T4TWMw7P/uAKP/d
g30OdaxtsZl/wYaOlyb8qkXB9CaynHjXJHYUH+P2Kltwsbr7SglYh8Z0qOcjxo8TiwZyKUOcL9Ci
6pjgxwdX09a4Gz6yudUMCzpKNaB7bG4MtZPPqtOIi7nKx8jVHwo4JWut6qwkvK5xu9Lq3CSq4EnM
C7T2QAF2piG3syhb17eQ4xu4mSKiGYwGhDp4tJxORQETMvG142mTeQ0AUhb6UkIwCMiQScRUEHwf
FFrXWI+IxSwICL7ADoTbli24DCmGzYk3R/Eg9+M3mfYmpMIVWJR7g6Stm8W6FWPvFYeUacwMQU6K
VT7swwB4tbqbJQMnzya9meiysqPx8yF8RqFKzpDyLNN+M7RzA9iqzR2Zytet3/FDW7sxaIjBf2T4
meu4nPyARmS13KO7SqUsd/QTtxgFNN3ddfmKjpWaOGaX7iwRSpyPx0K/ufUT6Dj2/kcoyVHxqgRT
3aXtOEST1wKh0wlIj0/GSJGpfse4RIvDN8uSAuvJAppYsMp+aLAvNKfHMD0ZMB55cnum2lkgvhuO
sLxbd59dx+ClDqk/LNoqErvxTww6Qx08CamfG8vcoqgyrgwHGwK2pLcc9jju2pMnRaSp0U/OHHbV
+sCaobXHYlMbllMrc4IBTKcxFmNOC6P1W1U3JI8soC6m0A/WPFvwxhjBQe0bRY80SbNGnT7fXr5x
9AOXk05cD2JednTqcKHXmX+TJKdZgh9lZl+pi+j4VbBQthy33gBfFUUwqdnFz7KOOih1WmQWFGt5
tvvsR1oA6Qn7XK7pAVU4iBk5ckhxo9+EbDA4eJwUeEFu3B23fKx384InQSsmGqu8qryvNOwWQTkQ
2Dq3EhYRX04/M3ynqbSB/+126Gz3Sd6MWi/s0D1tnI3+bcGQJmYjg1yychLTi9skLeo3UISv0mOr
1HDJxFX73rBZcRlR7rU9DshgFdQWbi/YpDMrfuh54TfsD/dUSjV6ComPSzLSrw8V2x7Hpahk/X/m
vJ5q3xNnIzQJoS4cgC1trWerAJ0MNWa2LvHzxH0NESTNvEHVsbaRMl519iLN82kuVBpSQKjXINJ1
CquVqku+7KGLjpfrPQVCDuR8N1VpV6NY0Wuu2AgW2SxeCM4YzPIDLbX27siQZg6iK2AGO7akEzfC
/5gqqhCzlJCLLTU+kiooo4x13J6CfxyISEr+E3nxu8HU6zRcC/q7IVDWj2jp4VQAqbCZbfDLSSQa
/1aNVu2tE3pXjPCh/JgCW1qmQfAGDFJuNVzkaGcYqvL9B8IVwSHnjHkOEi5VR8+AkzjA/0JXczH1
YH9OBFkNZJ7qgpm0Bx2unL1pOLZC4fKc7oBTqUIYs/JH18D8W6mGdsqsYwZwR0Bo5rmgVqO1wRc8
Bc7HWqNEtlquQ8y8mXfaOhqwJoUQuAfZm0Hj0BhIea3ZtvWSrY+yInTmooeOi29A5a7CmUHf7YUD
DEL0uaZ82YLkJ89Ir7+9+Yl5kX014nWYIqNkSpxmvweD9abueY3UHprR6fdUFDClIVadRcQbv+Xf
nB+wgZjTShR+yYlgJG89H8HyhjK72TKQsgDfSHAlYgGTHQlhfAKu1aIYeiycRoNDLGYWqUTs8Dnr
QXqDd/tpInjjsPZUiSkSeKWdPzv2V79Gf5aRQkvRgNG+hfHc4xHgK4UtsSuoSAn9gsorcpUd+StM
IHSzSEirvrJhhhPDV5ecw32fJenpzAVc7TlUA7Sp3OZLVYQiAHSyLGxw3TkJueoOFAHs6CfwJX2p
GjGKJ1RkxC368NwTUrWVTIgDYRKt9peyVP8ZGuW6ap7L9Ki2sR7k3KX+EpagHpHA6Bq7UbiiFexa
vePG0pyv5BFu0+hxfdKRDDosvQthm+rK22YYua5bGWjV3DNuD3TTij3zL/ixSSRGUXKS705sssi1
VKBEZwzspGrgg6sbm9O6rqi9DhmO3dpzZxXwsV+zylVcsy4wOfaj7beUT2Nobvlgi7wD5ARgQLNB
HahmRWczed3kr0Jl1J8YE5YPjDmWgQ9JYwb35XYlFf3zDu+16Emp/fj6tS8DhA7QgI13q++uh2hs
n5gJrd/qIsQ2kGhN1fj7JRaVPeP7jadc+yyq1PneYXOprnfxr/516X/6W8ESVVPXK56JjentDMwF
06qcKWNV8N4yb+skTB48GebqNNc2hSxsmWM9kZykAGN2sTc4ovy0JsShTKbs8rEOz6CTWicRT2ir
RJx3NEN8x4GKX1o7+LqA4DTNIP1A3C5sst1NxrK/xXOiBNp0jH8CY7U1zNF+yo1IFmhtr8aqOeJo
rqGL9nZs9oi/OhfQO3yDe+gCeaP/+qmZlUEUOpEKSSKZ7KQRQ03sC2/kVglaS9M07LMItWUaMvCr
uRkHGwgPayxQ66zlQW3dQGp0lflF9z5iXRx5kuLQJOwirjryZtB/1GjHePvVBq2T73TzkGMjnlT7
JbYLJe92wt+q9nKCqESOJtApTOE9VqEkRsxgxJXqvnJyf3u/7O8pUoNjyGRP6YffN1Sczu/RLfNG
endCEVe8aPqvcjxWArPZzNo8B0ZBD035Zfk60EznD/nLUEUR4TBhWMsm1kXIOlqLGyKLOMzjOOSw
dW4NBIA4RzsqR82lNHIzHDEJYJUm5LPdYpOfoaB6YPkIcRy+yScVaemNnGVmMi1pAILXDmSpFXJD
1H4S6eVkh3F9XScIf9MfX9dNRdDTNOo6Yl1eOGHylVYbc9hB0rWKtsLOCuIvL1qQ0iwZBSMrB6yV
Ka3hNcgGjC4h3PEELBptfnD1E8N28YIvhNT0odxxttpRvf3/2QBJNDfo3CH1BC1phNvl64+kqcVG
JmCvcDGO9cZrfvc1iqBcNQgESt0BqzWbvdJ3v97oDkauhOyfD628hOF2Db8VXXfaLZ03FC7NrTJh
C87zN9e4E5zkkUZuzilEYyquHsIMmRmUiH9yHKJ3/DzUtBUHI0g6VZuyBNldgBAgNKVSp06c/ZwC
qY5cp4IsmSyl80N8eVyDOf8Nn4FZ0s7GgkBQJt38n/jdOCeXVAcQEYaaqspPz0vDYncN8F4pemMY
mH7QKUrZmL6FEwe+lrt4VZsaDhzpk2XGsgRM8t/rHnFjAMBZqFYOi/TFNQgMDbuJIwJXaZxneG0f
6eZ1GNLhNxhTtcWA2alkKV+11BfFCluhg7C/XVglkJ1Ph3aKe6B4Srdl8nsfRr96t4PKO7UfNUo9
WlEz95Wa9uF0jURLNdkHCJ4MyZFoGI1H80xyfL1R58sOtmiDDlWWF4/er89clKcDU5VPvEEQaqwA
4dhDQvabAKQsRF0m94ht3PmCWFTnb+s9GLK9qs1WGQONq0kM6Hn2Nwfx3iJPoDv5avLnW92sPcEQ
i6Bid/HIYuzwCFiGfMTzLpmjZgjgST045erLvXeU+E0GwzwdeyI0WZ17d2wxGis3l2PbfKvf8KH0
DGIIo+CWDxa4YH1yaxklN6+eJF+hQAE4QW2fpfSgM5sEm/1gNArgG9LJxx36gTDOvvZi4LOkes9/
2bG4pR8v+DxCx/MTf2uPMXWIBgAeYUiOUZwh2RdDQSbUKeZNWlDgnnuJb9jgDxcuDi86We2DFKS8
ynDjRcEcyQbyKEYWMmx25UhlgGFD423mrVeJshCZLK9ur7s9m7Jcg3aQpI62eV9pr1ncMYbAxNb3
0KS6TdYjE2GISfhDPKWzLHDpLoysBldrm5vJTsKRNSLhCoQsj99Waljrn7wKPY8As2RWjY6sE042
3RQvDGppknQ20hQsQy/Y8E8gYkLw2PP3MQQ7h3blx8DaOzqY53e+6V3DRjd2UKMSJ7uG86sS4hb8
tkSen/6z4oVNLvp0KH2HWInGT/83x+n7OPXFC92+aERQ7/IawlaTCENk2ab8ciYtmcI4cDpKuF2I
eIcyWH8ry3sJfiXsJA0mJv0CGRYbs4PVsBDRyL2CY0SlsaTaOhaRVCuVFWo8GWULX0m9Wtty+OU3
2AaKxNSG8+P+C9hgXGyxkvJ8yec9/6rKn/kNTxSwd04hulg329YKeUMZJajp4CiM9XReHghtQw6W
9AqlHw8YeY5w/k4vls8UxIR+FERlFZWw7B+UweFaJ88GpV/xRbvDa9xnkXJQV7ZKP2HWwtW7akGF
7/w05moeA70OmIqSHbwvNaS+0rrjW6Kc2hvakTIoDxpEGnrh+Cv8g9+t08ZlINR0ZF8jUZfWfwoI
yTse7kbuk0vCU58XyiOT+r8owUmcdaaz5ceJyV3b8hZmN85jV2D3RWKUABZ1yP/VeeBFCrVZ/Mh8
RvDQWchSI1ui2EibNYs+jukIGUFIl8Q3L4YQXz+44krW620VGdw/aaN6MBw0+FZunbqVIQWbPRfB
9qwH9IGyrpAkvKUBHoYV1/MDKnK2uDEczC2LZhRkhU0t+Ls93fCg53gIpYgeRSbURh7X6n+7O2/v
knavn2joZNHs1vSUsApmaQm0GcRstSc4XespDs90H22d2msBv3uhUAJBZYUlxS3wljlr11Mw5h5D
hcI+vZrRaJkE0uyJu/Im+yLnTkTQsXUU4eZvBGmD5isPedkC1eWGOjhE4AHS89GmgbnLsePGBV7D
ZnXmPIaS6vO4z4C1kzHZMW/nI5PTw9WySAua7kq6ol4EHceYw3d3r2FIaaXaZcFBHgw8V2HNZ86C
UFEY5Arh0YvPjnO3flkD8FdtOmndzxTyZoxtqlsDtGgTM9ZSjx9c+grHYa9c7vraMRjraoQ9tC6o
sfZhNm/5Za2Rx2rhOSOibHqSrplW4Qw2ohe8im8h/C9+M76iABfBNY+dkXYCKqXRMiJjr/lvx6pD
F2vlkX+OGzt9zLvRmcPPtSZB6LouVHc8mlmxo2RqQX7mHO2nv0PHFfQ9/bwRJBlXPYtDp2Xk5qLg
3LNi1G7r1fx2IbkIlXToKrZkMSNwCK1AfbuQXlEiz68RDyB7GTgfC/pCAoGg6ZO88H3HXw2BxQ88
kL5yCSvfZOSIKhwHrtW1O4rj0t859XE56C3XXPyyVx2F98ChKxLU17pXqG7rr5lrj3+tVxaZrFE5
dS0+fOe3+uswQC3xk9fxSJB2v1yh+2Pxbxew6jUVo0iSSJLw0Zf6xufYUfu8fvyajQUk1HnhFeUt
Y2CPu48wjjeTBu7Q/4QG0YimkJjc/C6nQOWaUdB1sq6+0+jmNsafLJtXQsRiCPJSRNopINeDt4y9
zrb6XNa9NLz9BTE0zCFOIZALMz+zvOeO1e8UYWNNuZWPbMpnKBdIFwjNFLJDvJenOLZIqmOma1AZ
jgq93N3Ju9ZjBU4N6VKC1D5Wcgsw/Ot+OA2uD/YEac2+2eaiufq9zqUcl2NOeOGxcLYONQfS3ITR
ju9EyCZYzNFQco9+Lxqn0fywknFOK64DOwTpAcAR9xu2Pnbt4nck9LowCOBmj0aowZX/JiBJQRCW
1LsC+IJO+FM8DVf8u24OfBtLryEcpSio23NK8+D2JsD5v4ih8nAOicJRL3m8boIYMw5iLFviyLhw
ew0xdV3yGiXJAQF4pBkzuohVE0mFWi2W5xHeO5sQg6M3jp2YzLCzKE4RFlXIlvJ8OkL/y/b8FIFM
0seetA61wcRMfTN3pacEjB9YvmHlIcpuDd/QzpHaMov5k3vZpsHbv1s5sqApmuld7/KZzJhqr0nN
QZnf0EqkAcBFv2oyYPbD+OKN5A/Fq7XuA+JLEYQCtdDVdpAdqVJWto1KiPSdCNK35uXPGpMo/hr3
eE6ZMe3QXNDvE37tOnKxx8nx0rT4XQtyW0Q6sL+r9JgRJ7Ya8qfiOGZacVtVWDBrQktnylDHDg5q
geNk2XKAhO0JN+0PP3lPuxhbKmQ9EHxXsdL9dDhYo6U8bHDYobX/IPOmQvrruh9yCYquLUeIgCxC
pLmWh9wsVAcYbRlTdzyKAtWXtfZyoUj6RTsC9tzrzLZdny2+rTBeKCwxwKWiPIrkB7FTCjsZLp1V
qlU1et/C7fGrqopp7v+cBV/OSezP79Wart8cRv9c/P/uBV/zPyqlp7vNVqTQLUd2t2h8DMjBavth
50ntfl1Bfle41T+/YmRPhQLOA1ikML5tl5IgULuTmnWfziTUeXffpIccOUDDRcE6Rl4K9UandVHM
cVZ4GAMBdXUk1Fy5nStbn8MXzsAAUf1JDSrvb4SrZmczFnCoCZqc2gzIvouD0BG+IaDiJ1+hn27H
/judXs4HU4rBduiYB47+YCAmkulRxVqR/SoU3+m9NFoOWhe/AYPXFGGS1ZJzXCvMdNzNOtYEdwCe
f2FQKcaoToA4IvMuvv2pgPnynRuahq7CS87NUICT54ScAty7gR9j/qBYtOLKrdFcLf2VPO6NfBHI
/THkXVLYVdAdsiNvD3yQQJ5/98EbuPZShDDG9qgsWLaNisgmFasWeAyZqXhXOHrsbC4odpTTbFql
5qYoMyGdYt2IifZc7CFKmJvTm0ia0RN5G8hstSoKucugIlTGlrjvRDNzEH/8DZ71cCsJUo+qGCmi
JOYYkM9YIqk6k06qfZgB/VplQFb8ihfegfnQ0avJkHtxxLog7Hq6dX76zo0wC0PWsAPH3+tid6VR
lYLYZf8StL5vfxFxbAskF8jO67C+InJE0Q3zsISu5lI3Oy8I6SNlTKNknOlGAiwpxBqg4uEcdN4E
/Eri6LEAXkqqVJY7R4xkBdu9/RWN9ZAs1p0s4Nr1uA7SL9hC7pUmvPG58skAc4Uy75Gs5pu2d/+J
3kq2BJM6H/2Wbj1bn5RAD3alhwMAabsR1f8Y+bnAM4pl/qBTAiykd8+hlWH7QI/0w+Ta33uZytz9
/kQVE4F4Haz9+/XgF/0UbR+Vc+gCE4SRzLRHqO01mZfrV3Cwe+cKT9bnuVWdWsphwwwFekjWhCSm
VBjzXSop8TKbEgoZc1AiHaFaiDfg9Bk8FoAqaHg+4leBt7lU5SX6g8IFKI7oCxADVlzO4oU1hwf+
91p1tDySvsy8RcATfxOLlUJBlur03In9beuN62dgd8qNe5tzMlGB7s4vtyYTMOA1ZiN+xe9jcoCq
yWUQQNsqigTkRgfGLLRWoMbILWmg/2DXLbm4aOvVbDL4rJNBhBd36JJQcq1MEOk6mOB6dXSGWLW0
Nb+pZdT7/ng9l92WddIsfjRC3y4LKylym9vOC7F8eCaFbGF03BDAxjnwrJeZY4f+4CU6c5lLLa7p
Jy8HVWDpFIFVFoWUhhDRlURBkM717tXxfaLxadLoibrfC9G7ZQBIjcZzcCMRuiNjU2YZVvK84Fsx
B1SVhoESr2t3bXVYOlwf1cGpZMxJQJDAj/wVZDqvQs62MJN70PfykIWzHklwhkb4/cL9pFfYx2hJ
6vZG5dhvrOmxeyknu+agEgtgzR7btuPqbHaWHfriIHxTLc9GQekt8ynt7VWORMtJHKPqWGLadm1g
imtwi0iEzMR1wgaVQZhdmUHyQrsaOxGxrT91uPDmaP4iYmtS9BXO5cERbJmSU7vf1sQRf7d030Eb
UKTBo7AVCRlFsfNCpTsaN/EKQYzI93FMUzkiqzdZPl3SjUuQTVik6KDLOtX2HjyiBwVcqkHXrdDW
+HCbl2n9RAYw/BNaIy0QhmHgeQOMS8TIyqIQ1ONmzeNK5pIh+mGmVUasd6/vanQEBwxVWBW7gqzC
c3Q4AFmXZVWg3s0tCyYwsoaY0feywP605iOuin+kRGi6UPu2oBj75XE7CYVGVFk1jj4S5FYwie+a
8WzZAXaKvvRiqMLZquWwF3RIR7XrF7bitj8wVdZa76ZOTKpVaDFpLcnp97mbVrGvTDFcy2Cdhzkk
8uK+gm1bQJ7+oXTWYHifl6e4hZpARFyLR0KTjuiMmO9yYNQASos7NxxWFvHQKicP2No4QcJ824p2
qC6BQWXHSeGAjPvJIPInkV2w+nK5tEAgoQTpxwtQYPGpFDHJprSN2ypvdnAgkmEXFe9Aqs/xWwLb
MTFHPqgsO3aB3d2sxGyz+3+m66JXnBGvWX06Cu7uqr1R+dzUCLURaq8+2MzJc/686XIrG+AnDuBJ
MKvYpvKMEm5FX1pz/YNiThrpaEXeAJeWULHpo1SU3DePL5VzEwHEiO+dKVaNsFIcExTf2wsgi7Yy
LuSz1+YFEVjJt2faBqxXRpyN5MgG3rJEs6WHGCAMYJ3E1A0sQBDoG6Az65R0VPkkJPLhxgVoeYnw
T5avbpSYVaP0VNutji8reCfOPb460PGtulCIJd/nZrwqaDoHOZ37sW1zqi4OWPAHmfW/ocqexYoL
76GF6isTyiPVwmF3z5J5W6GfpdR7KV6+fN/8DVF60/153PLf6LodT4wPmADV/dqRTc39wtGTDqIm
Zm7potCgcPRKJt1zyDnKzmxHkH0hJwXY1ytPtFnwWTPbVj8HMS1fHiRIv4W17BC/ihalrgwcplWm
uDiFYIhGFqfTpgS5OVAG+1GH1k2DQmY5RZNgFGOEN+1v7ys7ht0F1FZaKRM2HsC5VgA6OZbP0whE
qlcc2GlRW8S+Nb4G0yeB/jqmhR1c6Z/Xy9smlTtSOoC1+F36+LR2iAFqvB5p08sEloi8FMPtMSRh
Hbgimu1LH9nrRAyWqCubXZ5WGk8v11lSF2xMJIrEdGCPRC/M9LBES2QJv/frgt3OeJ+HVGjt5Mss
wDH9yyhyYA8utDfHtl5aDQgK45MF0gjjp3mh8OtXj03+1PUyu0d0nHlKswP3r/T5sOWdUYcYSWXq
BY04xy4o99ZWP94IZROSaGkNVP4ojGI+5IE1KrFL5B1dfpC8fRLDbKJEZ9tfBj+Jx6DHXn45agFi
RUzeprGJ4A9wpV1zQsiyAlvH6gQqDklxhNJRUE0GE/lGJ06MWaeQjt53kSKUU7Z0LFdNcdUBwpVk
tJ5CU5SK1uIIOl4EgzIMyPDVQ7aZ4McptVRl80oocXK1NGxEXMuLAOyTn3IqR/aTI7I60y8Q4U82
lfdSjJpnG6azWg/ATWwYEGTqBmgFIHOKU422v3ymb4Mq22GsLrfnLsfK6Ho9RmkLr/pkIfMkF60x
X3WfYnAr9oqqPtZNtiStJtDqkKsKgz1DjSgShMnM/1XcIkK0mpYmAdC7/YBSFGRSfUKVnqgnx6/r
w1FAdr/mxsnBUo7yjcB+Z8dAaJN/O47zNCys8JnTUUG9VjUqYSUj5/L5QOfzs5erSdhuDifijrSp
n4FuStIGXUtCsh+8YV18nMM1qYjN94z6KBkAjvyag9xGfH/nQoeHo/cINDOOA6+Alj1/txLc8RN7
9q2I1qa1hXf5WYQmCX7yxcezoJzaHTOqg6xUr8DuRqGjMregqlASORuGbShfPtW4TGnMsCYUJwEV
PVoD2/aQU9gTTj153NvCuiXKaOkCkJu/yc1+ZHjbNd/WistvFMrRhEtVF6eVBFlpMD8sReeG6XkA
vMq+QbR677qt7FXF94tp/Hkx8H7MSX7hjVjwb3+qHx7YjkqjmiehGNq74jgN4XM+wlboCvfUVVNi
vbPPUlD/5EJGmysGSinLdbrzMQB5dslDYRZZbhOlMo/4pDoLtrqVaP3d4eoCR4dacNMb0EUTg4xH
ANBcamIuhWhxklFPCLkbCeVLAD/Tol234pIJQPkmUcyULvodkiIyffyRRegOmZhsrN6nfOCOcgPu
705dB5ZpjnSkDKaUanXgNBfbxrRMd3TPVqDN65XGg5SlbQkQ+7wupQoPN/AT1pYw7V+12sTW1Uky
s7kPSVh1z3iG0JHHp/dTZ1mKuDC1N1XlfvX4rwXECXQn9DNKnXFCgKHVtTWTXnRHtfvgPCqnwpqc
MzWr/kPUUHEpjn0mxznTCVBNq2zHMhsWqgDverqH0XFgfB/4kn1MIxwMQZZKSo5II8RNq7G4TCZa
GHU4thhQF6qstQD5PO70IxBHJVmYRdmZJSeo4bWGMTr599wKo6CqgZV5Ls/yNO0LOOHctoQiuIj5
EZ/+X93+60b2KK3uPpVtJq+D9Ner2jMnLQmAXfurYyHwlDDXsHH7QRXDB1S9AmxSPstWe0mA7Wrz
ZHJ8iCZ0NX3k5Spy/eWX8wcUfcE1I/wQ3B0xkDVXmF560OpiypetSmnWlj4DRz8ETxhG5xNQQe0N
N+tQsczsd1h9avvqgeW1uGRfo7ik6nh2HFAO4HedIJi3axrow6Pe+le17GRKJXbccyUIV40U3ehE
EtvYaMmoB6yUCMYpSNSNUkkY0oWoTIpkK7LGjigbzUjP2K9soFwW7WlWuH5SCNv7yZYED87N3hKh
MEPRIqWoPNVaZWvOwWtEoWsF1OKlvbJRv8cpqRlb99X7QWWbq00oG04Y18t0wl3iyjdv1NVphVXA
dZTIWx+38+DxO7UpntfOWm3kWGaO/DCRQLdCgZJFGMCxfMlfuqyRPCIHgfOTRPS99IGs6LOmBQoO
bmtWDAOto5su0qxHkDnc2Zic86LslfOfAbFhX2XPlJpuftkwGpGBSiLo6bhgbfdJYNW7geGxIdl6
jYqvHD0y4DeOd/etJ0jMRud/q4yXPedItPqITSR6C1LE10fWI+02+7rDBqBxCW2u6JtsLwuSZKvF
plvyFFDTQpF4lFGqrOmBHpYXNUwpVtF/MOgyAyQxLmw5hpeoQRvUbO/7wzkK94FTlE26pK7eW/yF
+vTbYCeVeMZTPFkErkSeywQX+dEW17iBRTij7E9EjVOwyxyuTPqbnnqMnIpiv6BJi2FPL338IiTF
TfZ2tSD42G3rh8PvGoPE2VxbHrnqKmgcGjr4QBrCDxuZuEH/Dz17CZK8zv3iaiDbBeH4O/CP2UNE
3jUSwTV//dp8yOWgCfb62DKbltMuZa/HwG9ROXGPCoC0buf9WetSKKCAqr0M96lduiwaQUBYfmpc
jGofvH9YxxLerFs1ViMcXqWR+lZbU5W4+nGK4LyX8N/HGl4mcciNgebxSSaFz9ZZ5NDVZjAAjUwP
8mRE0YCqibMiQli4BTaki9OoIK5jif2lS7QsEnxB8MeZvNdfBHITMNPGVkdS9sH7q2+y3cLSBKhT
kR63lYidP33d6OONUKVbnEOgS9Qi0/8m5wUfdWKS6JbGd6brSFt5ixLXMintdy+N0Ues9HI0b6t2
HLKOtGKTYy4Y/hjXxm5xJA5UG2NAxnQ0z0WuQ18xoevVi9h9egERBkACkod/87u5BIB9wntKOCkx
d9jEqeE5q/SIX/szKCM/bakKCoW+ckPIqytEQ2O6ruMiwCAFueB0YoXUc9Rl8wh1i7OPonlWaYgM
P4aW87lh1Jx+gQ9j2e99TLhzxLGuVZcB6D1GfUEkVAfHGdyxdlB4oEHYVZkfoqzhBY1j86MMWt0N
eBNWiTbS8zbShRZiiS/t24omCauuVjy+WQ2Vrw5iuQr9uuAqz2hbuVjZJWBLyAqJvfIs/zYV5eW5
ZirHFQTAIIfWfOlIoI1fwKWpysgz6XGGZW5Q512El57OJi162YIe6f6kQDJYzA84ydxNzARNNfY4
vpZIg8naxajvuu7a+PFhz4YtZ5UuE3LPMsAP/MshsxJGtmQWmf6/in3ZAYiDF+qZLkMb6pnOnyZu
EicPs/5iurahNzK+/g8+9oCI45aIiw/5F7vtIwSWX1Gv96sI0O1bY8Y2qGv4oT1QoQtqC9lxhpn5
0kTOaMkF7s3XKnz1aATDoPDt3lsGnP8+uwflcVRrgizj8ffK9tylWhFIYdiBOL9y1iMoYsHHPVON
pLzO7MeX1fvMRyv3w9PmR0mkmUG7Q+fYz57LZ6Amr4pP3rImeNux6CvK2SLlD2rxk3XRjrAdV9eP
5itU80KWKEuxRwvEvpI/EKKct4I+YiI44eK1gcyBWU+dg4ukI8FyTSTi1fvUv6j2ap2kuDon1wa7
wXaPZhHBm9nRzEspe6iwOGSj0TrY62hXCOZgzMf7fyEnLjs8RTVvC67Oj2tu44fo1JJqczBO2QjJ
ZUJg1smwz2Nqrc3BOMgqBpeBtgWzicAR+plAQq68EJgbpzF7Gk6VCaoL3xXKzSffDxCoOOHufoEJ
jcOsE/mTlj5Bs9czpMO+qGrP/F6nE0P4PuIf3sDuZ/ejG5Ht8A3HF3qQmy7uFPWKycuYjPguamjo
yJ5Nh/kYAyo3f+XmCXo9mjlucKCmSzArHr5zeYpJF40hCHrItEP1Hu4hZRTxukuABl7nmt/5Hwsd
Ri5sHjwaENyoeB1nDZ5lM+J0/oOtLJr5GDq7x2CVLPnFhrW0FkfOVL//PXDUMu1Ffwd2ZqAZZP8z
cv0fZwrwwCTVapahry2TurdQxOLfMo/UD63g2CWRp51j8xtzBumRqJcHQqmp8bvO/kn6ImlqvXXS
OoMzJ8P1Q9B1Lj64bz976VD/jLAkWYScwMyYPzZ6XDcq8hrxelXkMV3WOIp0jiC8p89KeGp3/jYC
aqEOaTPNU/nLDa+y2ODj+6t7QHJryHHVQSts94pAvzyTo5c4yG7Hj7DLfiynUzSBA2npy++LzX2e
lHFXkF71W7Clk2Wk/xP7/ZRHVQjiRl4pvYl4hd6as2XH2MtKcY/vcVy9mcDK2DRzp1YOFxsnr+2P
GsXfFiSbnhewCmbC3d79nksTlHZegFAjQCIv6S5Mx6A/6JXnqe38q24VTqZtowrVGWzS08snpWMr
zDSOYoFnKpl/xxIrd/zFfEEeAUGyMK5fe5hsfnWqF/jEPrE0ex29BQfGDs2i4pBS9QcsqW+ELyul
4jmgv0h+JGvS2ss+/34JDRgQjurQlQgyC0DpMNMdUrJzoiOZfo4ka78qDWXEIqT+dgVEOHy+3FmL
d+3yUkTx8CxGT4IwrdKEGl/uXTLqsml6JKyPef11p/fyYvB6uGLTnqS/ifDtBRfFU/feHmXzW9N8
4M0t8PJJFywT1rg/trNIcdKHaW8wfFoo/zMFgcjvnPy3DxGd9eFpoEyovQkjP2ujL2ToHHSwXJ7R
4L2qX8E7I5ZGjJ6ZNXHC88M4BMsRDI19/62u8NmnqzN2cXot423PRP0IZtSRSIO55vzqJbFkchfn
vRaarHwnIZlDyDiev6Qx4svcCNXKNrIyyUJwDGgVvT16/2Se8N599F3JSXfp4WpunWfMN+A8cRs5
cg9ssOKeAG4xzK0YtDI/tsmFBtMX0HQZKa0nyiF4I5pM7TQcvTMEbYxoMnRnKUZk7ADyDvgBhu1c
8LSYMPbXIdXxxbVelToaUMjysjVnZAt57IbWWqANr0wFBIocJq0XTEIK9fLdqOcrJgmkSKmxO4pD
YdUit6mN820rORE9qOslUB5xi0hyabxcpn9qFDCt6g/lsthY3+c6DZC3z5YZiPHTxNfEjuoSlCt0
XWhg8SoYZom3GNt3naybab18YPS1+lj915TaSGNpnaQjhqKw+Pupl7H/hux9BNNU2dZSKQhh6Dyk
ZlMImQQAeLMzyjst3y4OOTRVbZW6zfgpO38w0zGywwc+V0saZ0ERfrJY9oUejFmngeX5HZ1MgMfm
VsLkOf2TCQphVU8SVLh6CsULjO9zC93YXgguLXB2TVJqJLHy0D73fN5XL9KpcmGwOt3RAquvFd00
pQtWpRTyFYbLFMoGH8C7VxPgPYyTts5znDWZ2siTtz+aq1K537ALF5FHttxigjA9kc4g6AvCZ2fX
/wljPOssOB5aHusKKqa6rz1wqAM8UShOC1uOayEWhxP8jxHkOulQIfAl06hyR7SJBytI35e3qeXM
MALphjYL/KDja2JrYHfjY7YUBRBlLl+nwRvlxB72niE2tkAqrwVjeWU9i+/XK3pi5lLYEKU4ZaRB
y+6cJ4Ry6Qqas2dDN6WJoVYLXWwZN8BZg1G4view8/3PsMtlnZO5+d1X2cIpTdvrYOoK0QXsHh3k
OlrVs7LvNRqRDTrL5OGsUoDlx4R7ymAjHjWW79KefhzU1i6PH9SbL6b+CeGFdR+dxm5bCj0du81a
nxL3KX7GXLMd2eHfV2NwTdeZ01UaiGia+llyD9gFN5pYQv/etZfXfrTgtyiWI4XdqoRyzZne31yD
YdZ1ErtRqs2s8sCkLES7CvvYhBgY2QPvGJPcKfcyUyQVYr/Qe/CEwGRHfSH3FzZFs1lR9QDEus3E
QryJ5kp8foS4+RhSsXXdEI4tYaqe4eXBeJhvZEy8RSTAXDfw/A6sRrD1rRCRWzU5eELc/ubMO+cI
rr79nlq3c1IrG0dF6OrsXJAfwW+eup2Fu5vhxTV7FXyX3frWGvD19LplpnhbSzgPSNrb+CYjnQaP
zYxMGW0JL0gYgbNudlltR46M5M90e0KkJ/lS+K1DW596z/pHXwEBUliIWpFFmAvfvAOv9MWjVZYh
1AZ3446Liwh016ih5PWLYUXCjTp13m3H1v7XKuBPhnlhFDCCOoHVm4Frg+ASMuqdx/weIDtOJE3w
MOBirGQVJcLFg1MdAT4Q9RrZTL0eUjR1TzyE8U6P1tIo2Xd/560th0H374zRuWJ7orA1Y0mHg0N9
o3S41f9XrmixyNlLBibcOeHhonz5tRjdd9br1LU3EMvu2LWDbLRLXz3wHWXOWHMPa/5AhOAyhcBb
Vrj8Ypn0tddeN5idm7XXTPkx/jRkEpCL+oBmHESPqOae3rBNz5uqQu+dD8eygr+grnKKLHxDNkdT
meQXHzD5MqZHhktIT4INRAzX1yqKjyn0j0z9iOkqj7IEpnu0zhhFnQIfAexV23zvq2mktUGSM6U+
pAsPu//Kcnm8dQns3BOTR79N17i80YsuH1xLlCvBxTpq4O2utbspgaAAUYB+jaYH6+3CyOYWGuVk
wAWeswnDxsl+SVV+AfW3BF9iU999Hcq/VNk5GHZStO1GFzoZHMNpU9+HIX5zPAAEACZhRl//dUS4
4rf143nuMx9m6NuCrBa55QYusjXsfA3brvstdxQAfRBfTZOqg4TUhj73f+p0wPSKCMCsAXLzHEZc
CccBRyQhJKU7la+feKzdQpu7cIR5mmI6147xA9cM6AnfR90lrK3ECqe093OPnfrVqJ6O9JIyvZk2
GIK7GEfFdvWihui/bkpqztYCp7dLXUnDmjGi5ixsvLdj4I32wx79Z7Ex+tOwc8S5ZWR4brEysbfR
M40OqCQeuSa/j+JG77m7i9fSfknNaJPl3RQJMVeL0ECv6TCitJ2xN8AWZa/xY3B9ndjM1I8Fb76w
Hfk485RRevmvLuagfHf72n+GM2Z1eo0629KokYBbYOquZWf1LoX3aEfWr3IxQNAVyXFmU7T0fG8r
U36phq2TX3oHRuVTWTrdVx8nPKZGed8+DGlmYfrtYY2YYbtthUSjWBSmr3ewQAzckJUYP76IFqlx
PtgU+3VbOmKbDFZzQQk7DhrkdKpbXJbRfMfh5TVIBsnXX/oQW6VZj8sET9sJD6rCnP17Z0qVEF84
zAqlkcU5BdfCbYAiyW1uvUSNp5QwftFclbXtoasAk0fAvrbzGY0xksOhSN7etBnTsZ2VzMV9pInz
g52pYHmXfxrdwzUMTzx3s5itRthERuM3B4bzNbEFhT2bEoIoy04UAM/euv7G2K0GQ3PUO/yvQGzv
l7+jIQThAWxewWWdUkY8/sYI1Vvzh1MNPCOVDKMyewo5bbyWjzGbFZkHPsUEp79ySZ32nknMjoyQ
uxJ2gO6A27udzu7q720keCQ2za7VP/kyUDUPQZbGy/FrX1sKEhWusEB+C+B+kEc5LyFOhk4Lq0aM
fWG88eaP3VXlHI1kcMWs3Gkgc4emgHxR6Is5VQGU+/s8Gktb8SxpV9c5/NGQY4tdeze6ArjVxbj1
6tDarD/m9D6E9rg1KMVzd6WGEH1I9A6BS3v+/SY3DL+sYdlGSvixWCu2u+Bq9EZ40a8MkFagrJiP
JFmBLbj9dsrDAYIz9CNAMONrXmNc7NrgrgQeJrXz3CP8dqO02Qi28ctQoB8ZLIrJf6P+wseKkFVc
qxDYgjiOCVskwu/W5i+MO1FM5ma/pPDkprLmjIuZhTtVlDikb00cEW7Xl6nirOF+CJspk3Y8XGvg
cwn7bF6uWV/1XklSYG60Ai4W9PA9YE7M4IPfTyrmIdsAjjJ/OFLKYl4IQWCyNcFW5/7MwsK6aDha
3mYugznu1uxlFcH7sP9mbNBfBJs2Zy3JUN6g8CyDXs1+6xpnkjzzia1F1EfvUuBHYJkHNvQM2b8T
pt1eMdLiGZGNHaYOVlycNvjlmpoBsRcnyqOFwfb2Ox72xezEnu80pxoD8JvaHLNvMQagqoFR6b0u
CgOgeWBSMyNCvSn/n1JD0vrsTCjZW7X6+BSD0oNWrKInOuc2EB2XRD0vNYJ782IUfNilHJ6wIfaN
NjyYYC4wefFu/22B/qmWDix/WRNxcd8mBo6m3DTamEnPUlgp/S6XpbGkw36lRTWBUxOPh3d3Juls
3/neqkC+qheCyLR2jksbDgN7nQB5hIFSoeodIuTlSaSEDfqhghTv4i5ZfkkNkZ2LpTuVDCZnqlBZ
+l5RPSWz815lcQMXdxmL0P+2igdHROX+dZULJ+3NOL0FtwovHyjO45DM6KqF8B3eSp5dQnNncfU5
ly0KtChshD7yXXbvJOKw/S1LKoaN503ke3SP+QeDsnaGqUTIjhFsH1dVWHG+mesWAuCMsX0NqxZg
XorPeqpnCJcPJBeUXzGDwHGXUhDXI/cQ1fLNfDCJg/iRWEFXzlEnAsDm8ocJCh1tWmEeLsOl0oKf
mTp93RZiSx5OOaiVMLeapsYw4T6v9RcljM8ncsg5aYLB9wEPfpiG6w28x+fqO7WlEIJXX8iGbhX7
AvSU1XMp/qx5rWxm3EOfggLMNJZXM3aD7N2/OkG0mw8+0OORtCFlPStF/DwRHR0eUf4E1QGyDXlW
XZu5Lc4K7rZSzGIYgiYbXvshsooql19698nmc4qFh2KFsTNHWjRuK2fAdg7gMTs1WpHS89dtJ7ei
CIe9dUBzX5w33RkjLbLlymui+iy5hpgyTwdqN/YCRe+AW7/qZGDLyjVW48RDtjzvAa/x0OvBgoiu
JQJ9yaWBoxKokOHjFmYFx9ov9jcnqkxyeqk1/5QeWRBxCZszvbFETPeEyHRrbFUN7+ml29oRzWNb
vSw/D5AfU0JGTibSNY6BY2B5vkKaMpUFCTCzxM1VcaRZebocNg8RnKY9NfR2Xudn64DwBrDD7xUm
K4SJW457hovS6B9HvXJwg7ZGXnkKln+ruQV0ZT3gtSy8gGeQag7v19PgKltbME9IcmC2nOAlpmB6
M22ouS62hW3JvUl5z6qG+ZJRUqZxeXW+4zzweQJPErJ67KAczofiyWcPAtCM0s74xSQSIj5ztVwO
cw1JBD1IwcY2lDztvmS/gyPyP/LkAKxxN85hIkicZZUeRzWLIxGinmyFtsFiDEPNwqK8x2ZY2Q/6
K0XQa9YxFPWOB72qs/RVIUURLaAkdFY/lKFmMWzJKkBM2DWcHaZMyUyNsjJ4BD910EBMOUVEPWrg
a4WcYkHrm0CtMmHsT9OnOwBCqVNbqIDhixODmzaTS4kuhkWZPjkR/JQTAxA6j6OuPNw5uXvJTC3z
y7ag116nAob0yiJ4E7YfgjZ3DtZVVyphCIrJ68KCra0Q0ZvNLG9h5E3zHv426QBwYt6emIJcFtYt
NEKhOoYc/dXxdhlE4P56UJCrhFSzF3O8LY/PNEUg/ZIaDDxIQa66R87k7GKf5WftgmvmX4Fkm9vj
6O39wYtrlujC7CdR5Pv13Kbyktu8DnSsYd3fqnvpMqHtBBvnsw0YXlPagsdOeZX7q1fxlkQngD62
CxUEMc+QPs/4cJfCcE0QLm5B6iPpqQgz7ck5Bddp6ZedUam8I6Z+27EN/hmhZ677I5bZT+6HVU+S
8grwgcXqsmgQKz0/QxFjzw9dvDpDqnxX0wAzcGRUpYoUs9eR6g2de4iI2n+CKpjV2dZfweRu+Ouy
9ojAuO24cl3V+WF8T2TECBTr4kDkqwMLX2F0UoOboaY/0kYj+MldAOL6iatum9W+5llW/f1JrWD0
QmzVAvTeoRsOENnncBqcHHjBkcq96wsl3YNXi4PWMJJbKeUgaLMWblZHn4hPpvzxQy9MOflRQ0od
AZlMGew//EOcr5yiZ9X6r/2sgOWF1UsQ06evMujmL9QBmWKkFly0ZaI8iIxQ6hKVOhp0244G7Rgq
prd/NZxEHdng7nlZW3IPPtlb1NxjAtUs6O+PuDFZIC5tm1KkzDMrvhsMzz3yHzxSvB1YIhFdKjvl
8IO8UiNdh2K4APk6MRZdnyNifpy+tyEmC0JFfycNXtH0a5ab85cTlhG7axAiKRZsutSO38OBrJCD
hB22C6qeO4BzA3rhw2oy3q65ke4GhaQG7zwCMc8VffaeJMpJrALwERXa+QHFkxC1fKDiKink4vuR
DoCSvO50EkAhL9QxyyXvsD3kFHbzgRBsx0ANKkK6X21mOYKlIHNLFsUvm2S+hW/D9w9PIGr4f+st
PS6i86f3L7QQu+/Z1CH7AoxYK1OpsM0lIsAWfeJsP8DkQBxPfob5DfxGMD2DPS7vlWXmP7u6XP0h
ZuAc8JB0jDCGcDK7CKDl8BAZG9ZVYbE7dZDPWQbQfBfD1ymBsBi5IlT2YiHmkbk5xdlr5bjHoxNa
oaRS36ajC0FOp9YXhCMu0cXkUbfp4fYhPyWjM/Jjf34ZnU5jPHs7WuWBye9LhX9tlXm5qeB1ZJdo
6yNRaz1XFkiBPLKQMQ7E8xKcQDKyXmnLfs1BGk0EyqMz3BFl85Fm3qsfYf8QzJ7xu+Xw1t0uMZbJ
bOU51BFzb03a+k0OsF1Mwd+bjgX9M4Pj203ugKpjeeCfJS51LE9sPbgYkkBideb2c0KJDYFT+mTA
qpfGp0FWsnZ6zBnZgpYD9MaF/jWpa4COrvk2cQzx1y7ifjfUCbdjfamftgpaY6PK8H7KGy5HS/l2
BGxIfvqG9FLToFAdmNkMIbC9A+fx34/+iS+0RhQ4GY166Sw9QBKd8n0taE2YN+yDNJKG+XqmvzBh
nnb02GeioWsu97ZrHsQzAktdJ3k5lr6+0/eD1OYjQjSUKHKnS+RQfsKmzTTikyyP4+/cJy5p73Y5
2qfNO18VrjEpUY3cgITLABZoL1fHMgv8MjctblPDr8UlgzDPIrIRvXuIx/vj6qwnDFAsSBek6+Y4
C6ZytZJuyMH8ocnDnAgLttZ3ccacqKY4SOUj4/GEA9ETbL3IwEywzm12TWjCD3UXDdTnfSYtAVOL
cv3QnJeA8QVnUby6SR66rEtzxGbLpK0UdmEgvABftWi0E6bj4UL96Hl4eVJ+WrvNuHzKv+YcVpxL
5CC7CisP4KXzNu8svSsBJ/ldTHZqH1Btc2bsZV9WQX4D/rmFg019H7zu69vuDb7LKbkYXw/pasWX
93FVLPcDaSZTNJDByAz3BFNKpNkWKNVT+4Hag89P8RPTskqX+sqICcUSZ6vh+WLnwAg8475LgQkf
VdsKqKPP5HU8Ixam/e2vFweMJ0xZz+wTW+fu0+eb+pmZkBiEJiFXpv5k60i0cm5JifPZ89+xWqGn
SVUs5wlaiT6gHAJFLsf9D3a+mocQ5oLmpccQ99C8lA1DhIHu+uRMkLjzS2RevaViQTT/ldUioslM
woASGRjn4Wyq20K9l1DoHe3p1Ggj0Rq4hnzHyyprlcdKwbHoWAvmAJdts4WB4bWFLE1D/S1107lF
ZRxs+NuYmYH76CSnVvGWb7Jju1jjuEdAi4YvrxxtZmAP8D1r5GzWcBpdf4fBJ1t15XDhoJDIMQ/0
zqoGDPih1wtBH6Z5ZykZD7i+65BPm7SVUT2m5buU6v+BvYryaz+sBzytq/3eba8TaWqp1zF+OQWe
j2mIEcYrZ5at1Sjp1hEzl+1+KUeG1imxNZ8xtmSdVc4Ew3mQrHVCVymxujGnDp0OC2Aa7Ge2fd19
kK0M9QutaPSq4r/TTgzYe5c5Y/WkHyTD7Wjjz47FhET56lQW+rPld1j4JpugJGuO7bJd+0Takjn9
tvIHLSb+FNYT6OInu+lXnRqNom+JTr9LXuYGmhqBQgyzL47DtiX77/jqnVjymSX1FiM1GKIZ3iGb
E762bquV7Jq2NiLV4SPtGW1vDhjujv+p2z1h8MkRr37BPfsa/FnrGbP2B8xa54mzoexDtjdjIzOw
xu2KkKfpm6VdsqOzwQiXTsHnh1/JL55PbbkookdFbz9Ql8xPoV2ohLVTm3exK3nc4Uvt92lpNFzi
bwQlGKuvIc+b+uQOTuJThgcCufgns+/hRhxBUbliIg+ZHwxu2Sy3jgIaH4TgFGSlYlxAREhi2DXw
E+HpDwKVE7lqlosTBLE1vOef08cWnSAH5FzGg02PPU+kkxjtjeQS/BA4fpy2PQm6LmtVLtXdKlJ4
BsYUhQwfOiWjLf2+xhKGDsONqXzp52KqDqqzVXjCq31wcnboXQDQ+rODNkP1zbBele23tr1wLyvv
UegV2zqJrHoERrUxckwnnSo1n16F/snTaqQV7TRmlGcfdG/4PkRkHc/mSMHpTg1oI0WZJeTwZth5
gXGsfPEX5LIIDbpkdAOSl3bQMin1J+h3Onjd9C3JzB5c/YP8vAH4Ig4JFOA3SyAECMRLPpc4IH7V
Cw3RMJk3cPURB1ua5WaAls6c0lG05apWNdchzJtJJc8gL80DAmrEv6TaNhyeSnbqYpmU+kccBDK5
TxWEc4dyR3/3f57CGzPaMVlQJGyPFUi5GWcfRPORU/5eJTlS9RDUGXkv/RHYnPpmzmZr99Dt0a4Q
5nagHKRdGSYJ5GMxTJg+a1DE61YMEekt4T4pA9LytUsocTrKwk30j5RiaQ7wNNzgO59KSjEPoQpe
ssdE01+DgTJ1tTAAti9XzDoBqjFen2DSMfgGAco8qKp+8QpmyAlb5VvVqeZ7c4r8OhiHMHxEK0n3
s+G7Lk39skmdwFgxaIkQn9h1dsMhqUtcuR7FIU1AlO33RSx6aY4+Sc1wTP+PAh8W1x4f33cUTojq
yof0ukZ+S+wSdFnO2x8I7JEez63t5mcKUE6gKE+AWubD/SJ72Bu/c2Eq9wuFwDqUa6bg6Qe1zHDJ
Le4w0JT869N4bdnWNjS4rPWZEO+FcUMNXAc3sU6gF5ZOnvmMu9G3lZ5+y0c/C+TonNxn3WZ2X3Du
wJA3ikEQI7LFAwukJcrG6lBw+Q7VvTl92etNQMKOCWmwo5xOdmwK+RvAXaNtt0GuBZCRU++g12YA
e4bfaJT6qyDBygR4YAe6q2jzK3VWolG1ImniheAVXoL7stka0xJxRzmQyBhbg19gwbKxpWPxjhiC
0E5eEt1vxn+p+PQIST2KGUXLLaBzEvldjE98UzVWp0goQMr3/hekN/kvjKs00jpcsJbE6JVdRzKe
gDLguqu1T93be3thg3QkHyF+Tbb+LNqX2MwQ0w1XnSrWVYZO27ZYdxig4A7aPbDpQN7DHNDlnNgi
gKw6iY3Us+F/2AOrSQ47IliCEQt4KFJiejCGnrZsXCN/NEgZ9VdSkQn+re3b4HxaQzEs5KYWp6KF
9pKhWK9+BXXqk3gC0uGmy5Il+Vp6hYoUtEl4DiaCoR+VUj+Vityy7Flt9V6pzrmflv14ZDqMQoa2
yyed5AonyLrjI8qHZxhlanHh6HYsJAiqEAf9tzgl+vgR2W/xZZ8xekQjGfjTmP6fAWIP9fnI+UkL
Y0GjkyMVmKVNiSPc3VVvxlmGumHQUui71dK78JMn/z2sRhGNTlwCwS8o0BCVrmUcR5BgFw4E5lu+
3GbpXwLpJqlW8+2qPkxzdMNL1+yJ9eR89ounUNANpfj02//9pHxg3MwmzI0rjlUsYz+59WpgvCjM
GacO9LDCX1V06kwPNRZtCor2MkyKri8+MizK1jpzDD1QMMxmXt2PZ3+jvLoTMwJr/K9ObkICr8zP
KQMX8tHTMq3pCVG6hrArPTuUnGJ0A5NrBiQs8XfzomjB27sKQakfA1mhpU3URMeB520RLkvdPGSj
og3VIyyki+QPXgSyW3bIQVUBROchgBSpAadzYmDnv4S6YKfi8UFSOKbirg2eGL+LXmy6ScDeaE6D
xHcx6VHpoj+wfSO1mSMQ5AKghRyrcM3QD8hVTtSCOF8mJuLeOHl6xzRLRkse7c+y9UcDzOgIcJsh
FeiCF9kx7+UQPIKFNeGvp++UVHvSKATHDQqiHyUO89Bi65qAlM5rA/GWwWftbTo4AdKrL/+OeSYk
93hdrn5E3qXEpYGncKsXCJXqpuiqcs1bBMC0tTw8ys1HggpBCdmbEoWZDJPwuf5KAAs8k0ThIMmJ
4qH5NUYwovJQlz+YCv+kKjhelG/+YS2q6aA+Zol2diK9XulvDSW/BfNvW9g3kCSPM2jMwqTfePgz
qtfQ57SRFmnmpRWfzipOoIP+lrdB3q1idB2y6lYhwB72mWN4tDekQzJFEtfxUfDE/fDmFhyf8e2e
1Ga1s3v+HWK6wTjuHnW0n1rteqP1h6fEFTUsGWdMinShMw6bfBr37ZWOMczwvXU5elMZ1pm/tXZj
4cdW+zWVQGrnWza4rvG4O7Ts7GdpobOgQs6Y7UUv75XZ6qPnPH+GtNdNqOXDM7BibT9fLSjWdoiE
paAC2BdqdKKxgItsEBC5XKgkJOrdh8rn/liv/oPzziDjaSRA9b9MTGI1YT4t+wOtdqo4C4ZFOPog
3BRY6Nt1GEC5PKAy4SIHcuNgCdLorrCpy4yUJX/xtHRKe0AyaJpRUjndX/gaGyBPzbqlEpW+gAv5
AVHQc1AHrBd6XINnAS8Qc8+mwI0+1s0pQZXhlungVgiXd2bhDwavzNAo0bhn/Q+ouTli9iONyHgg
cttFRyWJgEULtZfDAXjcGIfNf2uY5pVUOzPl3kYpziO7misPtt/6QgKEh3n8WblkP2W1jHA2XEAo
ThzwR9lOkVJl4aVOWj6VuMCSG5x+N9/fJWLX/6lKq6bPVb5U+0s/NDyRUYMMtdzsg1BP0mBasIn3
7c+CrVaA9Yi/MLcYjhxZuDieGKuhcBZTnHpQ3PefLxP/EI2E6vkR7abeQs3d69cS9AxToQvMuO+z
iNv68f8d92mrCKTX/3+P9diyQBIhV056j5Z3KeyBMRBZZM7dX7CKeQQh8EhuAR6ldRqMUEa3jR0/
yEjoIX3Eeo7nBETPgWLIrMX8u6TF2Q7mXz+sguGg0JYj6ppwn7Dn33J2t3toekxQJ7kpi/5hXJ+f
FRQTHNzDQpkdfpEbxYJ/7GjAPEDbFFWaV/rlmbgCzdqiuA0YMKPMYeHT4s2T29sUQsdFWuVCOif4
KSv3bCkz3NeP8XUgrUDDMTxu8YdnyqlJjjJv6a0KCnuVXXeHPwlHnC05NvDc1/4yIdT3wHJB20Xa
lbem5MV/NPzu8YQRc8dr0vRIq5PRkchZJL22gEbRrJemsKYpAxKJZ5jNRA4bXrxIUQkkVVoi4ewe
wn7thTOaMmpSFL1FCCzMwETPKiGRfmCn4BKVmpZSgsJEMcR5H2GM4KJwPXplq109r32/kPqndqjz
RIrA+chdc2dR0McdV3s+TF32jFuWwK+IwY2HCLkhkKnn1ffGrhs/J0tvmoxu7SyvRFcaoctkCbAn
mziUoWMrj/qhNhCfCyRidQ6qTmn/JzR9+ObUf6UhxI07SG779ZagCtbqEPDejet1gd2WSTN4UACz
3F99viBYSjxR9nXZJP2aSlIdsLjLaL+pGcNnbJm2+ZG+3VxAAOnCKWHyeo3y+LYY3A6kuasCXkEG
i7ZcBMAoDYGbzMbcvzKZUEdnN8LWXtA6skaFks8NPFAbn8z6+kt+3Wdsm3S79Y9cxeydgvGM+P9O
OdTDQd9Z2/IbYCS50Oi4hfz/T81vHPOzjOmJRIWXngGLv+PulCT29WqVnOlhOfJvZ5tvSQz48uB8
Vu2YwU/0lcXl8T0cCibY0MQO/yJKpaXEqXj7omttEo4kNcNitSAmr4k58jQAdwyAnDWLNMQdrRLm
G7qYR5hvamCi5rY6SovSrYLJaO2KeZ+JwYqJX45H79FsPJwXV9Mxt1/NvuK3cCilzah7W6lGlmgV
0f9NqFgLHeMEXMglFQqRYR37PtWb8YXglMGAyZE6ZgyGWcDlLIjBbCfumt8JS+0+C46s2j72tK/L
UM0m2va7aq6feIujL2pOxvnTn+v8ksnug3XBZJpSI8WMBE/iFUHA6XF7brSY7X3yIc8L9wIIlfL3
U0l55sBKJIu8MBJHR5P3IZQtVQR09HtiiE58JaFdsp42dWBWkz5S2rIbpo3t4DVAWuy6f2eRodmA
FbepoSisT853DEn6nSXSU+E2ihWzZrJxIKvDb+OFyvLIJ89uri5Va6+au7to96R5bvsJAo+1K/8m
e9fdEEqQCicRQw7PIw+2Z71iIhrBNHBgvdeMJSlI0bAjjJTGpFznkRQvKoNmSmuPnZnUiNs/NnTT
1mOkSRydJpRLtfLS/kl7YnCGzEaT7y28PYU6ZjXeav0heKl9iKsTcZgB3dCDpw+FJwlktRK1ubC8
nldzZPoM9whDwMdlLUCiGO+Xln+l4FZO55WZRnwrLAoVBvjaxvKGYd/rriNny32yu7HGRyAS0g9p
eqhQafVv3ZGQxxtU0v9Sa+GFJX0l1OFha7XqOsgIu7hp7nlWbFAXIP3Csn1ecmiHNADlEjZ+fMWs
Uus5nsl67AP7pkO7IymUItQVBRpAedifQ2U3Isvyb+ibxm1bjtkwfrdBM71lKuuekGzwHysss7rY
IGn6dxKprJhaUgEOXVVQowRQF2frfHuol5nAeoFiuC4WOIUwgGhLsQK6uGDn2ePLeMOXEhOCeoi8
Ad21dTN/eUwW0r2iMXwFaVnex5dCxVi3QjmFVJRyeHdonQzsgeZgksumSnL9H03J45jQAZvhGSXP
QYN56PFSCSUwKI6+e3N0ow4ZqCddjCwCgcQuk51Y52TcgOMyXZA0iYYjLxQNqxSUD/4yz6cKsrLR
q6QS0FgAu0W5NhDNAcHCoLf1lk3GSY92uaLl0LzDKWxXCaczaI4WrRhbZEmc9YfUMKDbUOQ8oL6l
3U1X8XYOkMYoXZ0Gtw5JUOAkYSQLISRwuwvtoMs7aGps2LgkCuHhIXJeyzW4rgb8v/2I1xtS9qtr
hBLHTom4AfeyNhzflEIjDz1/zV7aXHSYlCac6v1Tu8qKaZBeUSaAAzFDDbwYIk2hkNa+lGoPXz4d
4w0FEv+RuI+WuStN7cBJmT7w35AJzJxekjUMGHIC1Cfk6xESo4Xl8poyv2MPcOmv4S6XgIIHBISB
+oNP1k8J05Fn0iSZK7Xpr6ERpcqdruNI8gghxCoLrBqDA3diF5L/IKnnmjG6ga+95GRdAJkZFizC
j366Ivy5v1YiVbRTtsixCDPF4yHnGpPK0DB6ptSUXKF6mXsal58CM4Wgmp7IMRHOn3ZbpNC80VZ/
V2RQYCJvnQGri7PVfPiPo1gOPajfiNbPfKu1tyf4KNOeYAl0MLFTSV04cPvOUPQAnjj7TT63uA6Z
E1Lt1yOktgVDN6ANDB0KKvM9BzFt8XAQ9Mw/atyV4N6CTO4IocxuBpQAl5b6/EYqivq0k9M88kNf
SxXtHw7/LFJx4kFFmh7ye1qGKvdhF4fmIf60YkVrCwf76CbektWckm9qCfk81vYoTHCjcRTL6W2Y
1hVjLpHF3LZ0nq91o3hwXaVr9Xsvy8mIdjljCZ8p+eTxFoiaJ1Z6PkVfXh5SoqEZauMYjotNZ9zk
MI0uQoxxyfpHX13XLlo7jAB1lWSDS795T+KCfGo4sZ8jbwQseAcrFZHVjTYQ/3Kjotzh3k8m6iRQ
jlHsHvIoIlCJ7PwtpDlm4deTT7HVd9wirpk0nHIIhnkkcegFkPT+g5j10fsmj4e16rciyx+7kl5x
ft1lpaqQ8PUsgavri+I9aaugNZr1Xw32ZsgSOLcSIYVnsRoNL4yLAYU5b4bIRALCPBKPAaQOxu0T
rycQqU0FpaisGAjuoET38mx/UF8Ak/c5KdVx+I7dAFXW8AL+UaRx0v7qqcmbTwpUbaSL0PcipyZt
Jn8GYoCcOzmrvjVbNGj9BXrGVI3jEiRP9gTJ472VCZ6g5EifWzic94pqnOERC8hngFJECEhm1g+v
mWUuQGTX2B4iSzQwWtFlLVFbyHRkEHafSBihJ7qoSqmdI71GCQr4rWPplO4TlDeRjehgAeNldnv0
TqSGNtv45nuKuilm/VdGdK+KEUdkvILRBh3FcHjcanMwUZa5zzt0H5WSSvoT463ZfhyezE76Rcgj
dB2HCN645MhsxIV59b0yZWd4yFIvJiLCvqCCClZkfx6nuuKA381VbPXbp3DtGdYo1m4J1fQmfOUK
zgvwIDSKc/KkN/AZ46redA7ju06PHGVaHt9jdGlrmr606ykCL7z4xNZWMVtDKuh0zE1d7Xk/hfZ4
TrZla3PN/ZdeVBN7wFezCsOTkcQEa7wY/uIfJzsMJPNIgT07HG1w9eKuHa0k7QrJB0M7gOg8R2B2
HjHGrYQtpMCMiH601ljSjzds/uw/PoJlvFca+vQMZvWRjMDoynNWXC1U5bJlHtonFn26VGbexHeE
kzD8FNUF7UciH16d42rjiNRirIy95ITR9kAb5VND5zwGuKw96CwMZH7AhQd2a2u381BBydFDSvIi
ElsP/Rj1HtXIW310Bzm+pLVAo4Gfd9Sm0Siz5ozbosJI3/qBebJLeDloaic+JfoXSlmoYdrpUQg/
Rzy1VM2MyR/VJkojgZfIvj1Jle//Ptn66muPj1LoX5hlsY07Iluq33yOqV4nkbn9bB5IAihegDOL
W16+U5o/VFdqV3pCXCcZ72WQSj7NYR/xtY04/qQ1j/dfISRP9qNBfIhms0gPiHDcEPQS0L4shO5I
kgK6JkAZneie1GrcOGpocnZiIW71m3XFUidMTu9Lqxr+hXq+wvzcQyeWw0e6OXBBezKWbyRd0eej
CzrO7pmkmQUrLW1Xm/0TVzg7jOPDy2B2rkocBAev/OZzcD4GYKmAYl1rQNVHNUI9yFkSXULvoSi5
IB/cFH/lSpaCDQWFuQjMjBghuwqiks2mI3SAv5aG9eMzzYI+n6BaIxMXgL7Psnlx5epQ3y6O8bld
4YngtkTlHUkYgAWmN9MlI/BhK2vrIJie4OYVun+XKfSmU5JKEfukYHTDDoXrJlufIBh1tPOFmbUq
Bc9u3a9bOpzkrdzkoyRQ9qzfzRplak5pty20PBCAfwGpRr6pTqX7wdHL7dy2TWazjd6AxwML3dSV
TwLCSwsWic11u7jdgvADKMNYu9W4YHv1W7OnAH0xTQQWbA8lKnd1jLMzB80wAIHn0g+yIIoswf4/
PTX6vZbDKH0LQQTEddT/kp+Y0P0uslu6qA2C7hxLIhbu1gpZkBpvczR/NpN+S+x08+UIP5Z65OL1
jc6IjEVZVT9ZJti/HUPMYSPsE6AjchNLBijDZ3pGgI418BIca7o0BXEo/sPZNalfUZyCbZA8Nvet
eOlWRZ2aNbebBF6QfhOhrBoQhnvbWZ9fFJzh0YETmYg03BorobHUF7aXw3laRcr580ncrxxjfiBS
pSk6A/Vq0Jp2iFafn+WRhPIlLlVzZJ84GGSKbjGg59f2zp3Dbt1qvBc+wlaA9D0fHKxTUNBQyCyN
71OOzo/KUp+T+zc/tiAHwPm3szo6Mk3vBESMgki8dmo89lMF53YQUjuVN/HFwB+QsuGhTVW0g97Q
d/7hBJPoHW386ygck/srtza0BRMRgCX7a8TW32F9skWtnD0Etr0WZl5LOb3L1214oLLDhHXnflpl
6gppsnym3TakXPDDG43Tzrz6XJuPAFffKnazpMsd0c64FJUnSqUZIiKOEXf5F2O9O8cfA0JNEtdk
lSys5jwkIJtL3CKRjHXq9b2ju9qHeZgsYB16XSlsncskOTuEWGkoautprgY6M2uy/DWBHe12zNye
hKLbuP3zsjGyZKdl+/ddSH56SX4t9bTrsyoznSTgNNixyIFTFUqRLUouwri3jypwd+8rtVlSO66w
vaIEbBK2t4dihapsE9X6t5/tBA6ZBR4cM/JiLSf65jDulG2hPsOLHteDob/yZ7ld8jenKJndKp/y
xg0a3HSJA4Kzc+T4YWeTZ3eShD4V1h+PWH1afhtlbbBCY5wCst/0zwD18/0klitJeI8K/bI2NwN+
7Ecwg6mN9wDG/eXuk//vNNlukQKXQrqmDW2ZO2k/gsTzCr+Jq5QdvA1gC2u7C6qKl3X5cDBimbH8
dPXXq5WXvSo4JR9qKqaefajwbq/f6Twz/I8vAhre+IXSMbOoCrQRA7txWBtwjsu6rSTwMInCBHwR
bmsoTrwg2GfZaKgEo5Fz1TWGX9sxjs4DbQh3dOw5DVbES+yiOL7jvH4Q07kEd9KPK41XQS0tL8fI
PnABb3igP5H0SLIc2BUJ6pxbMuW4usudQmgUsAKsJN89JVeCi1SASyvfp1syKn/pZElg95t6YeMZ
4SwplDs8aBZFr/iPE/2g0ld0nl4phCCTeArOgiubKOIPhQQ/vWzz8IkKXaXGywpHowM2tIMGsryq
vW67dW2gG+l57hEAkl+Sfjuez4aTnTvGP863KWdJF7o7vtOTx3pPWGpmEtXOPO5OH1jyrYXWkaYq
0SeOAzwkcOKXhDidDNGoqiHkwGI4ZYy48ltYtrFWFzOSzThrjdh0iB/E28v2fpDeCq4OtOdLJ/cD
7BMjfmcZMzrkbh21ttJe7bN6QYlpB9xR5BdtQa1cFX16B026R0js+jP5W7hVSY9Tdm6NhAFvOn8U
a4VKb4tNIbcfxoq/zjE+RmxhU36IPFzVxdw+XPpP7zx8gn2HZyK4c1tqTigvExtaELfy6Jkp4plK
e86INZUkJtis+dcTn3bRVfKqASbfPdCGn8YGRz7KzH+4F673mOQg01g7hKqiSPdz8PA5r2Brx4yl
bj35k5ITruYLRJH4AxAewRfbeWmr7w8cKq/IRxOMgf/3Ounp3PVintTl+DT+1oGeYSa9tFDANRvF
rSK+aJtrPw78ZEAB+ABFuMqFeHmgXN80RX1yVaNpiLWv7I5S1evfCAp2UASSM8BMM6Rs/8j4V2hM
BizondBwP6SMnsmkrtEHiV8CuE1qFQ5qCihSAIp1ylAJ1LtmR+DFuCFngiO5Z+2G9yQltX2ZP+kG
vQRRCj36Ofy1qvAyiDmoKnee7Kd4sMxoTg2jAvtRb6IHA7hso2npswxElI1KVTIdCkhItXScDNqX
dDK9ytY7GUByKD5GsvoxegdgBYjuEbH2XZIFG5hetaS1ZZf4kwgd0fdveO/2yXwQ3nDRYEw5qOn0
6pqOzWsbHTf0sMBLH139fM1Hkf04WnkqjRFwg+16zO/MzJXcLcUDsodT+joQ8e7BXpcfHjQiLTH/
tr4yjOjPgzg4WCpl3SZHhl7m018nqmx3DSJ70q3i/JVXzmKCmYBghwFqGZYskMIKCzxjqbr0jgO5
+bV/J41Uv3Hl5SOiG71qr6WanczWrMQtvHYRayjlFXAHk24B628sXQpZrP8DGCGjdioBQqwu8VSg
fdPD5c5f6WfnedwiaNDe08hiyOJO7jkqWWOfo70/q3ipE54glC9aVHyB+RCXZPejkcr1ZSKs0n+8
wWA3x3+saxDSvDYeSjCtU/dAGBAOHA4QMRMnbVIVCuA6t/zPZ9EKPPUZBvwH4eed++3reQvCaDhi
jWdFe1HpWC9g2yCO+MTPEyJ8gy9FOFlzwT1LiNOAvot44jcqwAyNaTL43Rd1abRVz9p/QzFbwRsg
YleD+8ZI203XA9xa8dxh2qJTgzFzDWjYA5Lo7b7imyBPea3YjCNJ+Amuzj1m+6UV/yravfFPakPN
EaT7AfBrDAOo75HuZpZEQ5ijgAM5U4W1FLN+2zAjwDVBxIQynvANsvwsxCYRWSNAyO1x3c/y39RM
Usf3Ud7bdHXczk6Id64XiUnuv9XxsKzBikzN0cBMQDr+8jqZorJAkVZkMRljWvhmCgyCssnmWcKm
8zql0my+1zN2zRC4BbUexwGLmnRZZM/VRi3+2S6G0XlghauXX7iQZiuh7nv5rWbythqOQ+GDAZ88
XPhdD+9gzC2rnp1hp65mYV+ZCp/U8OlgDW/9LYUCReqNSqgMgj9Bqu3Ua2Yv2d1RVW5lrEU2cw/s
udW+HWq3HIKeUi8vqNDt+27iHXtVcBquCjvHQ6MSvlvnyauKv/2bbhU85dGt9PJGxtcuoR2PcgmY
bghGhsRPHvbJ6elSzj79PzMqIXzHFQdXbPhVbGHtajgAVL7/DUmZdszcUZ4yW96/bL5HvEAhqSwo
nh43Wo/r71mglrs/9J5+CGoph1+66hMSqtBCvU5o3zjfCa84HL1kB/wDg5TUUhByVWgfFWu/z3H/
MZeWNSEx8jcGtMIbNgzIH1AdjAmZ8ETx0R6BEC8GWLpsU/tJNUn1rS1KxIHl7EqYhVw9MBaZ5Cns
DXymzyFwoqhuPTwYAFPidJGMP9gzF7u1dF1a0LYjvIQxqrOf1kihSTbA5+Y4Vgy+PRRMzFIUa0o9
FMTEeqHOVWqse6XCzIhuVIoeoRy6rseChpviDb4NK5Dosqib5BXMohgsne6uQy1S8VdUX03F+b7C
J6jd76K7Qrhc7qSIWO3cIEjAM8XpTzq8cgYAHT+yTZp1FknoI1FiwmKgN51PuCxkoR0D8xrGocqb
kdkUQDMHv2R4Vxlql4ouBmGMdlJ3ZwD0iMqF0AuVovAT48bsWOXEP5WxEkf7lgBvU/v4BGzvh9Wu
32oOhI4JGdHuZRazDsvQTdzh1f4YxO4+cxl/91/E8Ql58aNwfX09xxK9tXCY+mXy9zcdAMOtwmZu
LxxJ3SIImtr8N2wbAFydlJDOzAL5DUmOIHGFv0drZnFCXImh/BpwceAFScvbruMZh8M9i6+AFE2V
57GQHFinouRS1CZVcZGxGm5z3ti6FE4NLq1qSaeKV/kjMUeiQrcpZnyHPBuVGIpPqYzxDE0sbqla
sToVsK4JAB9NgcbS1sRWl0Oc1GL/K8F6Q8GrWSCc6CaB7Geb3Gft0CYkjXClytTxMmIJkWuIOqlV
h14Dgt+HZ0YnD0PS6m+ceovIcSfw5aO+jbduPNe77Fu7vQs8eeJ9JeJIqJtSuWedzcFvFJREBqmh
3UWZ5Utb65I2XCMc3lz8nnNMONBjQzdWWFvZm4yzHOhy9ZZ47VxIt8xSjNZj3zrq8YAOkp4U/qIO
D5/SGXCMiXcR3vANYx9Cle2THBg9uQHBEo74Ct37HJHTBZtr11YcPrqpZRxeMAAAHzMpo1mwBZcS
sJ5yEXkmYMacj3EzmtJyT4cPhCZPsc4rTSzGrXa9GeCJRNvmSdOyCaCPW094LOgidbd61wnjiTAj
MJuE9tRYI6HEgs/sOm5oGcj8/7Q6mMvanHUjSRKunFnIKYa+xyH7/ffyHxoAY48t+eMZYMjNXOna
dFn5DD+EggcgkZGwCVfpgNI+Zsy5i7551m4SvqIn7ZrnJA1SGk5PK2C7XiCWyGGf3ispg3xGsEr+
r1QNVBliDDsauiMfkz6YuXl6OyddtU6XdPK4BBeqK9ucp58SqGci2tAoysoyfKcev6ngq7+srly0
UrAPFIERbH660fks0fhJ7lZsrZGcsC0O9GmyIPWSrPe6vv4A5jmyQw5U4IN2bjHLlXjlSq0+DmzE
dUlTaLSJt21+/tOkEwlVaVgDPN425mKKh/qieLvMhidI+qb901ip9q5czWHynNit/2ToFLwRWavb
2tUkYS8KYKOkHU5/TQLOxXKNoTZYhFNsY9FKqEttUVCQ/1I7cJapth649FBEVxY0BcU0nNOyeWbG
2rFN7yk9Q4padm5iGT/lidazGUaAi9YX5EJ82nLQCr11f3+1yTk9spTapySaZgPuwzvMRf2+GA3k
pPVPW20h/lI/FHhVcvKZ3f4UKHkJWj33AnHftz2aQW3DbRROolrckDqP9CXjEmjQt8ZpnS8gOmaZ
fPTCpk4Lmf+h0+be9urvfuLFaLvfcXg+Rn3cQNWLvfCsasT87S+5wGqULtE9qSJUx0bgYXnBH2cg
ycS/uhiXNeQxjBmMY59msAhs3CBMn/f7YQ8BRP8ehYJfP7oC2MrRTFinOIMCvps61/CB8uCyv3Hc
Sq5V1J1KFinZbfb4qLG0RP5iZQhyMSRTbNDLwVf5nGf+REmKZG27uQ3MrmWGRRfCJ5LoMmEIXROb
QAcup9pMpVhTq2TthHJ8s2ikAtWjPA0jgWZ4H7uiJow7fS+iSy5GwYC2kBIslhNJRQ9XeiEft3RE
kCMVYyPm9Qx328vz1xaQiA9HWGysCM7R2GFH/l7fioRzgj7unlu6WzdeARCFDEB68GKgjDm0Ah3p
YDGDBgRpNM9k/KlHobEDuADLiaRUQ4OT1qWKJxh2ZJiDqa6yvDbgrOpZWjoCpVAa1EF+W+bOWZDP
DNXITajBVMT3WkUeKSLK01cI0FKNyl2wS95aAiukyv30bjKDRwv/ax1ITjhsE6XY+djkxHq52cQq
GIgacOPXv0SVgj1tdL2W1Rds6teoRQLTgSRZhm/XY25ceUH1SZBlKOeb10zAhM7U/hmqfINacbkN
W/dCT5nDVA/y2DWpMYL1N8/83T3FOD/sRVspMMRlOzEjjpYajaaVNWH5vOC8DxYN5U5v0ikDQk8u
YcYc7IqgIDbIDWHD4EHLjVjJV66OPp/S5RDtfUrT11PL2BRvjklxs3kcVDSC4xil2/B3LsJRPrAg
uf7PD87Nemw0ux/1OixCcZf0wg+HHkdeTtt5eKELKvctY8H4yh2C0XSn4aseI5dF8020eebsR0Et
NiCocrRcDkqNVip3kGbjjGfjKSvt5OkrYgA9Uxvs9NkwQTpXc2GalotBiOApjoKk2gO98HEv/ldF
Np5OQPmuirVEGPEqUwjMUb5xBqVRvbhFf7YZyLRcFw/E2CHn8TQLC49iHMfjeOtxbKWPVsKQVcdB
lAndQQ8G+WTtN2NFl/VV2fjMfUV5P3l5WfMlq8aSstCA3KxskVuBEi/o+iwIcKAU8xjdtIm2Q12H
wxpTkLUtDWUuG8XZADOWt3R6kzVYXhThP0eCBAnpu/4w0yN02rbqt6OpVg+j/T+84ZyIudcxkd78
8sxgnrGqD6aYolbMikNeeS5upMGuGuYqIbhHqgIjH2Dck77QMA3813d9k+LG6CTvEVV05rPtiGLT
5wzoleKTRS1LMj8Mp/o3Zkt4WuCTTiBs/G74hQC2NmSHNPirLsXL6wRm4fuz66JMsgvPweDiL9B5
ICjyeeQT3/oZN60VuRPYAGG4lfRJ3DpVvQ0KpZpGC8fWM8WlcjlyUu/X9CbwsL/KIXrI+XI6Uf0F
4F5RYEFjGWY1Xy07fcLeARfDs8LgSjSuCZUCQ/TxVFtH/DuV26+ePmCO59ICUF6xvWrmj80Nlszv
UC+4z1BpFI2PkMhs5LVFRFTaQN11QjMUD0mD18BYJuKmHZ/B1c8+DIMtyHx9cRUIbZMwGm0H36iP
T7mMLoFLJRdojFFuwCKjQ2unGexPrOWPWH/7wQ7owsx9QvJYn1rQ+CQXMuz8EI7im1MMwZjjM+Jt
AMQZpa+1aXuJ0bgZgDa+IMbx8G7Hz0Pl+zv0fUo2f91Q0M8PIwMbqKeIhA+04wUdSXSy3Z+b0va4
YGFBvqQ1iDwBAJsDIQr5cchqrPBYEZ8nb26cUpaszUlopHcuenliGcpkqpQgwoycNKbU9N+UCZFG
qKyEsjCCBqYeCIA5VqciFsRpMARXJZ+3JlBKw8sRE0I5sTVaokIxRdDsRgTEriQ9dIqgHgPw+5o4
2uq3czGKppklg30BhcW6C+EVITggv9KLkjs3syFS8zCuOwVDTRE4D+Aroq9kMeMkl5E/8bA4YsKH
a2bEpOyNGazYeTV2UbafLRSB+fIRruQuhVPnfqfZusRaXqi622/7H3Ul1RSLT6mhZJavZONbCfvg
8t+u3yFTM/Eod8rHRF7e6CALdYTLim0kzsVOtW0NKMLxrznJiB/RZQQ0CakdmvYgQBGh7tSiUpft
LHvRYEYPp465Rm1P8dhhWwfiBs6+Ya0Na/+yPRuYYgFVd2ZT3Y4zL6lERnjy8HNoM41omr4vcqId
P/mVG/SRz+mVVZUlXIY/Mu80JaRUE2oXSkY82fGIj4qJCaGElTi+75sDJ5n47Mbe24S1Umg6v16/
MY4cvBvE7ThXtHWy7ECLtcBtEVM/TeGOK4x8/EWxLbycbWlf5ELf9NZtSAACQD2OJzX1lmEX+Bcg
TXnZ3EfaiTyTbiUBsk31UZ83EELYu3Z8f36ZiEauu8Fk7grbyQf1MKdo5p6loWCU/dfoYBNpozJI
QlA1X39vpM7tZd6BMfVmm3c283noSe6mpIrvwPhZet1XcpVPLAoQzfVRQsFyHVV637Q2CWN1ImIr
aMNauOCNEN3x1kPPwt8/JxFK90cbW8+bDFbnkGZpHeuiH5QJBzQs4mq+ZwAXiHmYpbzeIgPtShf8
Cn201daYYTUBzDeRt5/LQwl9tXiDmW/nVtQw8eHXOCClNYD/dy7IAc9LsxvZn2wIJtjLhGWMV7ZQ
JnZhZmWsbSheoa8Y+ubQHVP1ayGMU/GznFAH2kJdc650698rxkEvAmo0t9TFgpwHlYuZ0cOl1vK5
177KJ2CY+vUANNvyGKjJqbwi3gyTvsIj2SkCiaNASxkK+UjXXRj3TPsp/1VkN8XTxHGt9JPtsZQC
TaS39YTpoeUFiyUyJZOUQUg1v7TPh7uIUK6yxHnx2lECHHKNVRhjigFXjs5mk/od9JtnhAw9iaO+
aVOpXUSVRodMQstysfOFdXez2MDDnl/FBauVNHW0mfvi/BytecHIxNcjXnUVHFMngKafrVFacRFr
V0/xrEMRzAs3ON1r4UN0T6BsDVtKqtWXQ9HkyBLxr6W6RtYN2TCVXVdr8BfwEdkDaQbWk6FyJmOb
TuL5l7SaoG/ARroBUZF3kFlOCG3dnSY6XTxw5cn495KoQExqHjRGVa56/flqk2ruipD1OS11QvVh
hclLTtzf6GmEp0ug1rCnma9cbKF+wKQYjF0IvmHPUiQqFYcMC7gCmxE4ZdMX6gGy++DPoOl9rw9o
EDvcWeGRAw8SOrwdw6iotdZimSqBTZjQt4bbawU/75e7TM88tXkt16lhGGCDlwsFQ2bmpwQS8Q+n
2TWWdqhJRQ5K+hbJBfFAX8wSN5fflM4PUOeZX/cNt7v+2eQT1524lxtZ9ZLkACd0SrSjIR5KvIJi
TeernAFZDTH4k6mmncgbskBDprIcMyNHf1x1AJ8zxuj/bFXgKBF8UbAYrKAtsWfeF9xmaaWf6RlO
wae4izompcexNRbeC7BZzuQM1X3u8XiminCQ5xUZiK1rQQuXvXp3rx3HNBF/tzcYfmAQUJcdeJeY
OKxqc0UXJDm8pwNFX44NVtqjRrv7qP4hQN4fiQ8mXu6jL9hwwswgz2glAzGdWeVWE+dImsfoshjm
f0gxNHGoJhALWktAffI6fdRKXOvgYgl+qwk8uyQqqj0p+2BYyw2UsYxisvum0w+vpOIL1sdkvsiG
XjK6ewEXDO/Qia0XURGCqxATGcOOJ3+8LZe/7RVqWEgOpjiUp/k6E4VokZ7VqJj4GYG47biofPc3
tsTq5MWG3+MrxxfAS5bHxTe5L0ZeUztDC54wlIP7Q0e4/jyhJAgpSuqx2JV0Tw6bP6R5BZvW63CH
PPr4wVf6cez5WaiC9c9MFA4ZBRGZe5vD+pOv8JO8pQz0ACd/ZMRymUGMzy1fOuiKbzDYJQ9FDNnh
89KG6w1ZPKzq40yNEWqK1Xrfmt5swTISZoBIqc38zI8WbUB714rM6CDdSINyoZLzaveIGASZnP3z
8Xj3l27vi54b4TgGiGNocXn0akQ0Pz2rHLlU9RSV2vuWn8hMqeeb6eozRrv5nL6crpDwUf1I+OIY
kkF6OcQZFaI8cbh+i/patr3gf2JFCrvwEMdyekwvqrBmOFnOV+od9kddkFZvhQywOxPGJK4mqjtb
+Gfn13gzPFX1Y0oUNQFU+uoJw5SwdobK2EIuOsgwnV5B7UArV7MMdMDPLQpXKiHutFPwC3ha+jRe
aCbeB0GwS//OAycOUHbpm7hAWpoOjoFBlrmH4n1K+z5xixqBzcUfa8FqH20RtHdxpzAkGxOdy9S9
tN5Z/1DeykLQgJkQTx5xP8RDN/mo0FHDNeE8LC1CGMpAqlergFGWiQP63Is1dZyHUKDMoviSs+m9
3ipL8xoT3JciUZqtCjSbFj8brD4/XEoPFZZ+upPu6Adsaf6Jd9N3yeYSOrbD9O5vK+yNlRRJRoV3
UCDyotHR1eCYj4C+rfUluJrU7tUeilgGxrvnWh7g1PGUzedftXLsSDjzZz71R5CEBYFaO19t/ycm
rM1lBLD2jwebkgyP4+K9PVHMHj1DsPMKQwUAIxWvqpUjAUHFQewTv7KTbFf4qxZl09XanDmcY/qk
Oe7GvRPByDJZcNPhv7jdvkY+1pUfGWXnGPI3kiV6sstMqtLZtytOM5EJAtCQrFF4x98BhGazlyrS
eYpKWMAQGEUcFGBFPgsWbvhs5D4tgFf2n/werHRzievX65ygX5oZuG62kOaKGR+sHB2+ZjcsoySx
0sv5IQOyQ8u7D/MERlO7SQaPCPGfyOpV9mT8af8M0ytSgtyFYH4pyuEpI7Or+9k35yki8z19Q4QD
CTQjECiu6xrue1HyXSeAmQDk3NJJZAVFE5b874KPGz9/VxsVjDLTcZcwTULWsLmlsY+OpdVbCoIs
n6mn6Ufqk6eJrw+9jQloZSGzJ3y/dIQ2+6j0tX32q4LXY85KzhuKhaQ/1yeChO/GB6IuX9UtdmFI
mtZ6OwmsyQqO61WIa+JKwh5C34WtaijI6tDwfwNrq2Of1hL6eLG9RldzwnuTPwTf3KgPZSH606at
Xuv2quLga2Lqh0rZYOYeWH4/KQEMrxMIZ3x4vcqIhwaVyiJpP5DqW6WFhWzDof8SS3XDw++2oagE
moCTy96WU71IGLrk3ZIq7iOGUkdn+5R1m4hFojjRsiz0PKX3GjfoomWwPajLkvaUDpPg/TTbc3DG
8W06s11ZWl2W0A06WA6aNh47WiZPsR0O/f8iZVUdMXY4NlA3HgPi1uZIUo5RAHVEd0xFt4DhLYxM
6fWuDodA4eHPf0VJHpuESanUIQMzNtfclBwmiH2SgVkGBnvzT9q1M0+Pt2VeituT6tZJnroOuta3
9JnspsTGgU/xr3dAwwUoMsdqnG9Kym2vklRVwYH8FON45TvPPEtwnRxy4shBOLYuAQpnvKuo8nIl
TCCt3Fh1gi+xZULA3K0rBikQLzbUO8zMuMChaHgpOr8cP7jcpEMkJ3hCCQwJrYBZ1UOzJou4H+A0
iJgH66OJb1OnGABGLL/pNV6JcsLlDbqYcLIUf+FmTeuL6tf1Lol4buzK1aMWPbAIeqdQtEXM1QZA
OOz/DSinOxUyqgaot7KwhUXKAd1XwINgySKJOdoLX5umJSjvfixWdN6Wt8XwH30K+l+OxkOKEzi+
LRwfg2isxW/EHW9+qU4LeWBth1VPyh3+yZUAyRwBJG2X2jGUw1NUGxirc/l8LMvQr0eoFh2xHklt
Fx2tuB35lWormemSQkOq/ORIr07tsDIGo4xzYBunr3QWwCrU4OZVYKrNi9DHqQwyRzaYSeSgwNWE
iJLwwK3UaxINahAoopeqNlTifinyE1KNOiYZlstBJ6AySKEoIcfZ40BRbv5HT0/zkw1SimWElD8p
21PX+DSJl5IdE/kbRmwz858bWAdfL3Li4AdQ5Zv/W7SFEo39BkY9X/PAcU9NHmsdrbPMEaw5hwwd
QY5qlb/EJ5HV1XPJjIYC63I+mfem1wthzPPWTz503cMbg8mxFM4Bf5F3Xb2oyg12m/ScMn43W+wJ
kq9jr2jnuRizTBiTUuYtpG0/a7eZOZmN1GRhUUZbrbV8gWnEIhW5qHLPpHJ8199TyMBt265+pAns
/UUiThMC0Pf3scNmtKl6qrtmVVYf7MamltCFFAz6zcalDg7PndbqkACSoNAQg89JsxcACBVt5XMQ
BwgA/i2dTMBwZo6TuTIzRMpIZCAlV7elAG3MMFFf1qdAQTroIZhEBTtYCYZoTR4F57cJvZ7r4Lcr
cJFP+RGe8jCFxk036xmRrgCWUJ/IVkP5o6S67unzZHRK+liteAr58B1H50bwIGd5l+7tb9zMF/z0
RXpQf3KwDxh9HP7WVl8TOrWywM2qtSpMtbqXUFQZxqlP9EUgeHSF4FpAPoGTs/fHqyA6DNe0srlK
HMyIpzNOIyzAIyaMyLPB8hZoAy1w/v793sznthfrTwH4c3qYeRsw2q+uTbC+Z5ZiF4izJFqBsRG5
LX0/Fep5PdX/Dv7Y73DgS8hgXA5r3hkPyNM5HPBR0bz1gLzANmy9ZCFJ+LRoO5o4LRZf1prElNY3
Eb31di79X/g12yMMBLXQb3UNaTxkZumIVH6/DbYJcB9kn6L3+wq3PSRlLgytrVOkwqjwyx04ctT7
lQmsU6H0J6me7fX8nyeOfFSClClSocP0rZWuHtkPTfIYfLmmAkB9RjWXZERLN2QV/nuMTCrakKJC
2Rx42mjY4+EvO2uaA1dTztTdKWBTFmawSxl+2YGLwFyLMvR8x2oMOe/8lJk6UHHyCTYhGKEMjvRH
LdAocw7OZ4s93zRYolnZNTdphhcSebLkJfg3ALmBMtdGObTjrAUZ4TsGbPmmHb5x+qIg0a+RAmwj
c+hhrkVIQsS9LHyA7KGDD/oM0l+y7483mMWy06AQyh6sOHMm8CHlo7v/YzDitE53Ra+jzJP7PbYz
c94o3qrXJ3JOExRmbvVtQpAFBXbWmSfCeJOlsn9w2pQaRWQzA7qAH34dFPd+KoY2XZeGmUaCw/+t
1dmuhG82H3aqLIJL0w9F4n4Qy9IxN0RQBkdFkJgd+cXF5rN+QZtV7ReowlIGinTOvXeDVw/JtfTu
7FbZDDMycn5MzZbom6idi+h0J9VPBVA6hHOd+86AI0g7MP2ClwB1SjL0mPqZPGI9d56+9kWeOv8y
/Oo03gEdu3iMbAckPkcN85p9Qdso5DnEcFENpQsSroendh6T1Qs531Vdp4XLHYICJYirXDxp9boy
FfK41TSAIsUv6/IhkqJ8gd4mG49DAzjGo2AlrzxC66MSiHjJ1i7IyzWoUhb7FDp9sUlYcYx4PbF+
XN/xxb9uabQ6UeyFR+gNjCSj+kdDYcfoDecQRgAiufY=
`protect end_protected
