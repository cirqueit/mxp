`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17056)
`protect data_block
HC2IEycByGBtCQVSGQ0iss4OhT2vAhDr9pt/crRWFGUEyZR/4Hx+KtDZRB6XUIPiFMF2pepc/k3W
iQktpDjSUrCZ5j5G2jziCsebk+2mgLJHYfNe73XwX0aB2lt7gYpElQHBoje4Cqr4JtuJtFvrVi8i
FVqzycvfz0tGs7NrxhSKeOZTU0JdKnBHVDstoY+nyvG2Vy+rRXG1/8poLTvdcXOGTm9pa7cnGwCl
hENFHt2NfDVjfEKmLO48yG4Z0FazjJPHNOFyw3iMXwfBXiQYv4uwH8W0OQ6f7nzGjgNHo5ig17Vy
wwLVgL0AKsNGKXVClmahOpKGKNJ9k84BkGSJpY77gXrroS/K1wbr4N3NGVfPRlVi6fEpFWnxcqd0
8Dy9DU8+nYjFOL7OEgIFhZt45mM+y5etxY32G01K/d4HNa6jZdIAFVoecIRBEBPmFrHaeP6to0k5
pHFsj8e3AoIpst77FQrJwSk/kDrFnHZUSq0QrPO584KgCMYXNA5RRJ6/xsvi/zRLtgDRBxONHBzX
xJvNcCd0eXeQlTolADY0u+cmMOFJdT/8EiXuG08fXccvGsugHAsD0sOTF9cVr/Vu6ck/mvalo0UA
tUkd3VPCMywSudMCuuixogHeJKqXIAg9elE1jRpguf2fvqszlnIvBzSedU0yZERw2Nw+KiPJ60oc
oSFvOWX3MBkHMr9FdRS45TH2zIujxBVC0ur7tIebbSPl1UqHGJuKvO+nIDV2zknlabIPdq4Rt+So
9Ohy52o9F1FhyPGpiZpF7i4fYsh2tc3324a824lsg2e7KR77HUYeFHqUxC7wstVLjhrQDixgPF4M
qWZwMwuaJD3ODocSoSG4vZLYKeEigetNb9lvcEGRBAlCX1z/cvAthWc5D0evOraoSjmDwC6ksvwQ
eNLaEtT7sX1TI6xQkpRInYoZNNWFo/jRFXdMKwXgb6w38PAO8iFV8ikDsSLTFv7lWbmWRM7gXn2s
gOrUi+5uB3SS0U8KggLoQYun3r2nmPTOwqex56T7OFHFa5PTSTc/EEyiE/DQNRqtNnIDmXeaoLID
KOIIu26dGCyWSbpzAgovc8PUFzxtaQCgZIHBWANrJBNR/Dcc1SDabkqsV/XRd3PA+WJDxR+POsK1
tI6vLLiDErNchR4UfBPsT+x6amGFXQ1URnX/Lovb39mFlaIWgQO7MDy+1VmCLhfQU0XhkEqSymfE
NRDLy2G7SdivdUTjqv+rPVQk3o3wBP2Q402F1UtNY7Hryr2yamJiY1gC5he8+m/WPWOonB/KrNdW
qkh6opYKsEJAOli6nyHE170LGlXQ4iQ6Ah7fmZcQwPmCSmwULdNZvdIp39nY/j6r1xBOUlD0jaiB
pj4wqLZjlJnMafGObh5kv0rthYzKdt5fl+NsP2FMZMk0t5xd67gkT4pxw4Dp/YGYNbHb7+aquPtb
u/OG5DHRxWtn3b/O/Xb1vWmGV/2tUw/4Sw+DsQDmep7sYRkc9scxJe+8/rjJVyn3hudQB8E7G+Tc
1VK4hSZ/qYDP6TfoLUGIZgKS3nN6i0Qa8JwGHkzNv8FOzFfegFbUWnbCuQrkvOoT+3BZRYmxgvA2
JpO4ABCjOC43tCBMKYov1FNuo54lcw7WsDyG/GaQLlpAodljya6ugy6aDTT8WWIsPz7xyAGyTOBq
wtpP+KkKJN+Xc0TxDEJMnDtcH3YABhpVNusgEv8MXislIToD1I/t/UE9FN4dqxVTJREVqpAPX8mv
JTlaxSnbFsVm3EzQdW+gDL4OyNsjTkvaRJssbYG/qFHBFdu5O3cx4id6h2Li5eYS+NWlgJGX/d9n
NOAuPt94DMWXCJlbPZ1VRO2PCtjeY0i1DC79hnIE6nEp9QRWGSEDmltmCime6HraKhTO52ZA91eI
WEGRJeQkPAudQALmjKzUHRuzKx1ZCWva6y0Zgh6RTXimBTiq/SLIcb491eGadrZtpweaSleNI+4y
UDjxGUtft/nMkRBmhmzreOPYkSBkzgrmkL9u1EM/5q3n+IklIteCsEu9HvX/LPMoSl08UwueZTGO
0LUoS676/NhsjUyAvFFzz1FIqpbW0Zk2e3zGn7kBewLGIaSo7mAkQ0mEEfFPhR4oIW+9SN2y76+7
T6v6QPjSItLRtlrJTOY21fV7Wnlnol1iiPGWyMnnlrRHZ6HumV4F3Y07eP+s7j17H9ZRNVdbtZoP
LmMYZBOHPtFA+J1L22kDYLL1QrVkw+DFa0HoyC7u70OaD8lGgxtwvCDr6NtB2F6e+bSKyCbgZs9R
jlGz2/Y4IfpKsI2vunpY6lrsVCVsX9+jPsE7icPGv0Mr8Y28XASuKBfUL13D9OHrib2xGjSokcpl
Yxh0wkauKu/ZqvlYi/SzbGImT85bxpLu5+PTpWjV4I9feC9TcIrRrG+iAZCtRa2oMY2va+NufJOg
vk85FSdOjXxh2cC9Rpa3sU5nHuXfhX4FkVtv7UoxJECdFk2HXTHftYwMsyZ2PIS9nQUjS8gAU1hD
TLB5mOiXEeqmcLkyn2k4yrp2KtM98a7CJwbOQe+FpvdAP30no0xFNEamR0rldRGtaA4lRNX+yRda
dght7dg8NKkQS0I2ux68iX1lCdeNI0bJh2W5WDzINWQL74vvTLlCrPHT2YiJpIHO92jkiYdCyGcq
F2unJSB2oGCPIGz4XTR1aiVUInTOsabqXLhqUqdQqGnPXlchzZXocwk9JVnJYUn/Izy3Iv8eR5bj
TVkrbW7Bph+pnDriE6PtQCxbS5TfAiwtZWyQV74U8hHfZaRZVyLO/D80+oF5iV1NKFfTbcAp4sry
QDs3tDE9tjv87zPe9+6979mRcsbNA47MmiNCk0T1ZXpRwFzQNfhD8uEhxvFQ4Bq7YB5aHgExll9C
khkzqMtGYFClP3f2gf0MytOLU9vFRfn+Ft4TiwliUxvp90yArrZTXT8lWDqOrCc3s66v2sZvSw7m
TIjIODWHmOi36Y63nRITbL1HcK8zw3VlzNowfQaKUdO9HqjFU6VN43KoV3myJ/QpTW0L8rVHVNZO
5gDJ23kAaW5d0rIxOhFhl2qMKYYiOknLv6L1bP1J4boiOcgQ+eOjzZiHVDca7VsRJMobWt8eBhyB
dHxL9c8KogoDo1+0XPfx5x6uXpN78Gnmaxpmm60qKrhZUe0upLU3FvYqpIXb1fBNGZ6PpGnAv0Nf
+5mzqjdGV2TVJDYhNvctLt3dEIodbOEdQEY5vWKgVAscH1quVblDW+/NfnSbVHJeLUNS9MSpV3ou
LmWRrDs64PfJ/yIJWsGftq5pjsZ/5LrYZDgslJ+ewqHefSqRo0n9J7vUnTWdnDDGUy5WVdMz8iZO
4WrvN9+8+zHxh3skB41/uNNZL148gMmyXy5rWvv4Xxt4u3w7IZyZgqQ4JmomQf6Vl+Lkg97iq/2L
RHEB8AlXHMRAfQTUkgZCFDihGtaa0HsoxOOrfGkvB+bu6fk4eAVt8tvcjYxjGPVuUEMmZ30km+xq
BrRKfVj53eAIxL9ekRbcYeJY6ek5O4WsVkPFpdnJW3CdsVcqjOos5iK04vdQkvOq68lDXnwzMEwi
miaH1bKD/cEg12vckN/+bou/pqZmbdbzyYryJ1+VaJrtf+sT3RT3xjrvcRlTQygKeJu0Sct96HB2
EdHl/92pJfd4qo7ogmLYkNtA5EAd/5rGMJKftpp7xjkWrPL8I7NN5uSWDY2vP2LZ7V1Rg07YJyf/
+qYhUrZo28kZVffuUXrG1Cic/fQfyklxHQZR+Lw0w4zUw5cIhPMveR7ftnoXR0hD0v60l3iorX0W
+COQH+gwwNuaPUb3afSVmhgwCzbM9BgDnAJlVcVlb2T/zFtSFbiUErh6W6F9cXA2+j2qg0akF0vF
4qaHei57fMNxbGQ3w9j9MlhXO8LNdLH5VNaLJlRkUR/5MbaPiAarREu3VR6U10cZbaSaSxamuqSp
WuS0S1NgMSnjYARSUmBGkQbntiZH3UUDDs+WM8jD7Bu3x5vbSrP/eZOGAW/aYFGPX8NAsXn14ntX
IB3IdcnvEFvfUGfet/1X/qyLrVJ2Me/3AFO0PWRMfDiqwuEV/bdefJRsnkmZMLlp5acq6sPag3Xh
D3S9NdA42lwt9C1AZzwZlL69CkMIHzrHut2VbHnlbJriOlAltIkT2XIeQdd4pafytYw3tbCUvtAU
fvxLAFdj8gLoqoFzXMpucIaMrQbBsBCllDcJZf8CoeXG0qTPPR5EGr5VFwDjZ28Tq/6ZjKN2QCa2
/NuU2uKTaVmdJ+OTJC9PTqwYEKM5CqOL36LwD+ue9IF8xOgmjD1iJF75tHB836dikIFobmW5OA22
AxRFppHu8iwNQ3y6rE5m8SVijalmu8i4I2yQxYUjLjCh1s3+hojDOdY/SVcwkbYhNy4y43dH+AyL
87/lt1oWBewO7Vq6O+S5LRqRBX6U2LVAwfxtA+wDU3R5fUfQrarmsNfYyCluPrKJV0REXOzsdAYu
weMDUJCLD+bqsv1TuMKckY/PZLjbgZm0PH49kcvlVqJKuez8y1cVp3tWbyLr6AeNivgW5icb1Jct
SdKSxlwDkI3b31snROq+YCELOWqNbyGrPThmGUr1+glfe8bMOY9ja6caMGpTzuaLHBGpsLBjqAWS
vu6uP8xRz3l/O2PVMYtjkeAphZDbgam4kmlEGFBBf4+tlRrPPuMZ7rEG3FMCBpHTp6X0UT9NT5c/
S5DwiBjbbXcm4c7jPJ76IlIQlHekPZdGiaJNmT7p1CdKcFQcPyJsD4V6jLtRFXiwZ5yQ/bpTaIQ8
i1ImwB2hE4JiX+KSMy4LnY1MUf+s4qMAnu3vuvrsODfHbTvrUdQddKeZRm9Yvvmb8Ik7Hv8Ekp08
7j3ESGTvpkfy5sBOQCyzbD585rxk8Y2jL4Gk56AnpmURXmt7ktU5S8Xuaj8lZJXX4JahEGXRWLac
1lXnrq+dZ6/BJww0KAJcFOhg2nk/nfosIj4Qur19gzJgG1jik6b8cpGWGp24H7SYF3Fp/cTypLpY
/vPd55NfdDgH+un/Ke/KpWFBlPHTSYqRO7GkxDoJGDHxeaVVtmZX+TQsZ/1edVlQQ92bbIPSJORa
tm3wu/WvwQfBHtRRe31JYtySCBE4ofx8tCvioD3xFPKXiqE2ib9XTcPk6drvgf9o+u6TXPT4nlFF
SrFNHhHlu/p5w5Dnc4YCHfmksGhq483CTI+6oYDR/7dyp1PMfAe7RFT8JUbxwahe+6z86m0ntVlN
68EtkEU1oD546UZwpLwDh5NVaSrUTyqKljurib6HgwEWBPXkCh9/835DZgoQMf2/fz4wKyDXVzF8
3wz05yHJMBnF8khEWZopxbzERiTBPzY/pkqpaE1oyiOOW7vBjlOr8jImJU9wBiSgD+Tkrs7XTMvu
KNRQ3SHptsGO6QYsavRgdJdh2fKJt+9Pn8wzUftmft8fze62gwdQhz+FSALKH/HMVoVIjOM4OYgt
ZT1lf4LIMYs+FOtGesw6pZtwHpHudTgazXkG3k3Zj/50Dr/u6RjS+zYf+rqbMm19FpFWLJsCnyZO
ZJum67RgqRf7QvghrHni//vnKPY4hfQcVOJ4XPoWTZLnoNdZUI0np0LJgfOo9QPxvo/Ja30Ak8Mn
iusy743ris++Pbfmmcvv6OzjauudPv3WPQ9bFmCu4d0xFvcKYln/mFIg7GMnVVv7pNVL7bICoBhg
HsqH86lVxQALbMZ/phMRlqd5WhaHH3GAxu/QXnaXUFTTwkR9lKqZ7VBc41gc9kz7Mpy917k52NU3
Lr8YakWfYgyvsVxQbn085U08l6Z0iB4ua6qQUal9ccVhqnYjZtTid+kVNY7s0bhz9xvwz3uUc/p1
MD2VMdNZSWOTOBTaW4XA855/Aw8RbdBG3gsUuMWpw9m/F5jaEGB6W4qGJ8l04GZJ/6uvoIl+a28T
tnRangs7zhKNWsO/n62pysx/L0E35CGxsNWXHCqfwVgy8ZS7Klcr+wLmUTVsmtC+51QH1LZpq09Y
bK+IRAm8kO0opB3L/S3tl89rsQwF0ZYhaFYqxOb/Jy6vykk9PczJaV+u/gw4TJpG/cxqFaxHyMVy
sAydA4GVe6fx76jQog+ZBf4dezW6Nu1tuSNUvkowFcWXnYMKo5x1xqf4L9HOsESuJxP0ZmbTDWfJ
6CctMlnbvQggKc4ESTlCUa+1474D7arvFejW4ayjmG/F5hCsJSipzzABsXu5aF6ttx/NGfM66uAY
2wTJ7J7mDb9SW9U4/uTGgiCop3nnByFKE8AanFrzF6mKu8Ruk/yI0eiSu80Hcjp3RTw/4WAfzxPp
hNH9y7ovN2CD9P+Tk4haUqMvM/bk7CnvEktMoxj1peSQZz1ldABAF2qq0ZlHADAOWntqcGF/4Q/n
1rvb12KUlWeDDaL/ZmefqnAzN1vteSxcS/7rU0L89LW3HyZ13/MXF2gEhfLvBJXuT2mU7MYpL5ZU
JbudDFk0kOQUuCYopluM07Ko5jfav2FpMhBOQVQWvJNqLumS4djtTmZ1+sTZvSLKrs5Lpr4BMSvW
VNffhJd0fV8LjG30bnopWOAbg38Vx1kIj1bT4oeDqpTIski/vToA9SwgFOPHEUoQBO4J2samj9YP
7deBX0xWm/yQjfQdG9C+yArXp9Q21OrkBr4oDgmpi9i6BY7nyAEXeQ/Lyv6EUGPKbpaTdL5kLCPk
OIOfmiTtCDY/KaiGg0KoZz36s8xItGkXZje7tfEpIpwuiMzXKfCVxpiElJAWL664Vp9h4pRs90+b
WIEGbT4T5VC0MWtcI0opyEyf7oM599wgKz/SsDqcduviY3T00xvxGkyX1y60YxVocg8LL5z9QIHL
sRKv5It6ixzckj1eVX9SwKlZfoWtvQeCu8eWvXyJvC48MR7+ov6VhU2P++71yB6CmKDBdXf7ifKF
H5jb/7CXNifSykTLxRtRE1zbg6ugUTR+w+Upq0jTpstB5urDzo60BSbzGROFi8ECcn4++bK8bpQW
oqw2RyCCyAp9Vlo3oB57RhMyM2dHy+OV/Pk4eGm/fFOEkkA6f4w4EIGboKrXxxLrkgtY4X1Qs7mW
E6wOSKX1G1Q33kHlvUT27GhQeJ/5Lu2El4Bc4hHk6EEivWt6YrqGaKKMij+ZGZrTzobV9TbH+Cgj
tFwEtR6c1ukoAzTVfS04dalIh/ebTk5GBD0PVE9S3+rfAe9m+LynPK34A3FTiQExmzKniaCoNZ7L
F5LltisEMLr4CcUDhgvYygXOdttdvMCnGPRt00AUFAwZajo5IwrcsK9iruG5oG/M0P7EFjHyoWH6
yE71WH29304Op6+n7Y7XN0AQe8vUKr3Qr7/B1T+FTUj1/gpWjvPMC6h7p9XTLhsyhMDNroAZLGFd
IxTz1mY46CpI7wKlDH8w40iz1OafOc+ahBessBfavv+y2dZngih8/X49nbpM/cH+6r0cSctHh7so
zT/H0SWmObSu7DGw0ZdbGrwk6qwtC1TVElfcEhgWnnf39Sojkm/c+OJJfWBIwR8MMxJATmXz/LsI
0x5fxuaDpjUEdB4/Tl6SsVRGNuX6i+Z+LYAm/tzDP1ED+Uyvz8WchGEt7U98jg16x+HEWV0h+xsf
cwOFIrn7cRuqUWxD5eDV5i15lcJngb+C8HB6lKkJpYth6YpM3o2mbx5NSxONsf7FP4JSUK895G+T
Xu00rx21WMcSloJaQcKh3kI2rEj3cM47vF4l8HYba6kzkLjU2AR5vhATC3Yk1HkPNiqkSj06/JX+
LvDnFvdzrN2cFLx7UTCJv7SXpvSnpT0yZjs55N49IKtPWrdgqmsxCzH1GwApb5RX3m99L/B9Bpr2
+pMdCH5NtybaupT6AEA0rbiw4P3F5/Q6yDgcl4kORMJ2Npj8PqGhNZLTw1aGGIanc+TJqBHh1slE
xCfdSjKPo7agOWIqmYXdDIfYP3Rr1VjVQSAKM7HMFdymKKveCt8QP48MYD85lVpSm4Cdo4YgzOCR
gVCKbMnzWEOGRnS4AJrF5HsTHd56q4tGq8W7HpgduqJVQ7U3QX5kA6sKVO+GyMc1d2PxByYH9CFY
GrIPzG9sdyCDxhAq+RNaf7exUjEzNM8b6T8Ubng4s1Yxjt0edkoN0W4CvFpDxT7lMqwYaVEVOSGA
LI4ZVp1sWyLsai2iy4VHGOLCQhrRHZA9UdgV9gcPR8QsDtWpvRvc2rQOSMYh4S4Z/P8WMplaaxgA
75wKj4DJXZg0OHVCWBQgMhy0HsHUOsKGwybz9Hp8TggXGXvrQ0MP0LNXFKE3V4U3CRBdcMrHiGWa
X2FNc3ZyQn/oeDyoaPOfOn35VvQkyQP8759jXR6KB2kFRmI11M+QWheyJ6pz4SjsEyDWS7XMBABB
3RLUtcoznNLhp9Dx695IFN+vrzjbwO4FngnAo1lNsYhq1FoeSpbnt7umtFdtI0UJaf3MNhE96f/P
wmgjkJyCsc599VcmXmopNHOom/E9Nnrz9nKey7RBFu6w8PbO+fqB8lAA4871VR8ywbA3wm0LDmlQ
x3edQ4ZsTYQZoN9rbMy8qYcTTJW2/HlmLPjN/gL/uArRUTv5VSXr68YLqlsSn2K6x7sZblNNY8ji
gXg8o/NEhwZ/xMsGwsxZhIDPYJLeH3ktli2F2L1gPPi3/HBpePQYh+UETFX3tsQ27DxJxoMIDuvX
z+8EhLsZI1aJ46ggJhMiIGhGNY2UIcccyD6y5NIwkBxxFCCR54J7FjLK7xnrOQwKSjSZO3DJoa2a
KqDd5bjiwP4m3/Y2Ii4irUNJZV2b4NU3Nmwb6t+eH6p8oSC1g1LxGPazM0nVCRI6EhNTa4FRSztl
16yVM4z1qZlRPf/HQIHCsCdwr7WVER6LXL2OmfUSj6eajQ55XcrjImMAf017z1t0I8k7xg2ohCq3
wEfb2MfruGTqO0lBl44nLwrneIqmLmZAebBkK+h32EiHka/t8g+dCRbYy+sQ8kZ8qwIzoErTmH27
hDrXboHbdIIvWRsHUAp1SXzG99QTSWHgAvsvxdzfpZDgXoicRzFC0e8atNUp2H9VyQir2rGUKr6w
A0InxzH8Fg4CJsvfX9ArqOjEVdNApCQIHhOmC58z9lGciY7JR68RUqsigStfLrzswDtVFoo8Gix8
IaDj4tqDIlXPPOBzpqaftbMmUZdOwZvdSabrmUiWI7LQogv1fP6SRjcASXEPDH9iTaRgc79iSo5S
ad2B9KR0RI4Kzl9ebj2i4SvdclD8faLeXaVLInYtIuzZktcefVVMOlgi3ZqvwYFy6yg+FeZLrVvq
HsSoWl1TkmT8yQ4fOvynbNbMxWztVXIiAmJwwiycYXznpC76sn2gRL1w3s4P8PwUmqovey/h2Uw4
2v3gTWMTpXwzDIwCf7E48GOTHvQ9uVAzXhlG6nym7y0YIW7JvsDTyj5grAs+BSB8Zx4/j8Yrl8iD
HRpYOn20R4l9uEA1GSPsGsT4DHL1h2Eo2ayKZxb81hHsF7/B4LLJXPBm60gZS1WsKHQN0bL/ezSA
0aNBkHdUGrxsx+ie6WpZDDPBZqPiw+guo+CBNSdvKlvdgBOxDMuxPXg70tUIVCRG1IFZKhrpbBR/
zhr/qEJdGDn2oHDD6dVyGITTHsCtnrW/hFV0aw1BDWXnDyQxUSJJ8lU4hT37dsOu8b8kSIJ4EKF+
CZvjJKtQEfAR+DgV6c3I9kl73LF2Lhi0MmUVyVLK1OQgX6uzIWSo04chvJpyR9c7PmCDUPN+1oyo
7xlV10PVtWeWv1MlQCNNz/UCBlUwBo0BN39m5YaUc90bpBv8RIY903t1OyBlWvrEOW96wKphffsO
jjT21A7jO+AiHBqZVYVsQE8OiHfe1Yq03L9b0Dy2fXsKR3JI21veCZHm5D8W3PtUWw72fESmwgjC
gYJe8vMs4OxuYwRVt7YArjvZDv5NB9FU/z/Uiyf8lm2BIBmKH+P4BSw/byJ3SDoy1wi+FG0mAyD9
t+NYhFuSsCMT+ABCO87fHbpf8KrfbRNLjhhwzq7lGWwIEGpvW8SZ9B0Nquidc0s98mna9poOTQ7J
HiaMHRAPT2pxUDk/JBia10qOYWQ7f78deCU5MARKl3C1/q1UxwmwhKd9O2UqA3D8uJ0PK0YyjYfE
9EabM+Zr0+VXP/MqFEXXyN2UbjjoVsEsgs/vRMgUccWimFmF2olDfLPLL3zcLOz5NOCkunLm3W02
A51T6/0HM+UQfP3S3tcBeq4is2PqmY72t7xVaqphj74LDb6KB4T5kqb8q2kYETfoVOkKAT3RXYhO
rTuQrMCHoGJYhkBr8w4PaYWP2zqUcXhD0Vw8b1xr+8+dW1adF6qwtyH6gFE780PC7QiaUSPBEpk5
VT9J4CKx5K0w+pnnQcr78FHzsa+jUFQ99sujYGe90xf7S1lJsxhFLuo9Sshca+uY4JgbdBlcWv8I
EU2FrRXkktbZEZBQ9dMUaOkxoE9V+gJtomBd9fJGr9cGX+V6L1TQP28zzscvVwh9dOhXlBb1Atrm
ZCimMddukQdIOVKTsuPfvhetl0k+zbH6vsoI10uHbMiSH8EGo/DYIj3YvMrMzY4ut+IzWPXW6i+U
qsHv4Ji0oHwxbKlrj9OdlvSH9FLu72AQuTcM3Nx0LilsFZbguVplGKm6Op3viHpJBOsSBTRXz+JQ
P8guDTQcBcGxvMNUabWNJN7P+UmRnjOat5y5VmUrB8FTb8EZStxuvsXEkZKTCi8xySdMdapTW801
9APswBS0VF1DNoxaIntpEhpyi+NCCDQpsW1evokq7O7nM3Y0dx4u61glsEWwb39fOFBc97EPDQt1
tHd6X9dk7lq7UywUpop/XBsgct5XvwnXEXoL2od9y3NBs8Uztdd/UPFFAKrndWkWWHVOb2ia/hWy
DSlGZ8GvXgK0Vvx8X5jeBpv5lvXWYGeKJrXLyhsD352Ueqkh2ntBzJLMOhTcsc0uIKjogA13nK7t
5bzzc3Znplm7aCTBP+He0Ll+i2VY2RbAh4schocemaVFBfk7mAzyMaxErcb/mQqrzzBa6sT4PL57
2eRHBqeAb6qyeYNM/rFreE/tH+DrF8Z/yksSEQ2V4zvZjQdXHyQu+ePvBSf4O9BCZDjzTo8kiQCq
4H/KdfBc4AXD97n0p0iA2TvnlgTfKaUHPOPlqRWB4clacxG8K26FQAqfCr1MVYjL+Y+Tmt/urpYq
ehsI4t27dJfuIlhN1CgRbMwe9AIoK4eDFv/kRW7BtJZk4FiIoaVcZgjbn/Tv6nRF+ko/c+RtOlrl
l5Kaxm4krtqIb/Eyoq5ejd6xJvBWX7j9pMPYIvMxd9RY2PQijwa/L2HbYomnM8T4uAcAquwb6rSw
0oMmSyFa5mTeywWqrhIX6BoWuADKnv66dqTdJjKP8EvjmqX87BFxT/V31S0PmNQLAWBJnLesxFBo
QU8miUjeo/1EAcuuSLVd5AvogUpv9Wb4cZ4Zgm0RLQZcwBOuIEiBzRyVV5ds41/J9yCVYZ3w1oUC
pZ8mtRcJJJClyvKdRz7mp+ByGjlQkLCO5OYRnO/TJcajXSbpFqw+ABQlxaNaMuMhMvwQABxmSb3l
obpDZpMhT9dqHqSX6PF55ViZb+8Bgimm/CoMZwpRRB/QOkTpZf7JkkSOZnDF0ZEkKC25JvXxN+5i
yXNKZfBBEFbOV446RElBkSMp4D+2FT/ZpC3ldaUD2qcnEO4JBHOz172tOZ6GAMQST92rbKtQpsmp
u6c2du+U7aRtmHYnTtbpHWp5EZpl9bLQg7bm02FU9Zec4si1yYTPOIzZKoSLtgj+XRj05cRtLQy5
HDTeJWL7IRACP4XM9GhqZyIRhfZ8s6NrNNsOzEDGT027l49nfCaKKgA8n5KebZOR29uooWKHN77s
LRltz8HLuFe971qigxB9/Jc8hfK1XwigV6E8JrbFYjFKFj/puDEo1pAPndFH7goFxOqsLJsbdTC5
0q8QAtmbEymu5IZPM4RVtQdCYLAiLJqTdy8F067U66/VuCvTQs0dWep+nPyxHIqAefuqWi5fMPox
UKBJY0FOXRSc7qhgjlxuA+dnF1zfNvvSuaa3TO/STFAOdKfvhK/sMakfOdO2z/4OqhIm6nqouQjK
1WseoUY+ZejsJE+/ORBz4YW9dtEwbmVkcpAv6BIL2mCc6GZhFLPbrmftbkXhh3XwKB1EuzP3kZg5
+GpuoqSY4uf/DpMT2oe2tkz5/D8b/jFUepy4o+CwudhIWOtRjeQRc4Eu4gR6ewjuUxuyv1b3abBq
9qTwPKlFGJtcrviqAqBwg2p5zqdbt/rYk06wW36SKUxVhJWjgzl7h9eDhWfok8XRoXe/kFCzkb1k
XsHncKRoaUj77Qb66qawhL7o2gn50wpuYHi5SNF2TDXOjcZlTG4+gSQHF0GaiHmZNVVxFsV2ZLqy
Uj4lEyWVJXM4iexHEUYOUUb4wt2vDUlSTZHiM6SfTcwX96UulSSE6yP7qWWmSVHtsRV2Hj/jR6nb
Uudqoa4mYqYj9koU940O7NdTivn2urzu3NM3kcNRxVgLRwpWJ5mtLs1z2EQht8EOGfaS3BJ57X4G
HZBkK9NyFunFkwik5uCPT0WHiVJoLM7lbx7URM+CokWXIFnPKFtBmYz9yTaKmdZNMI48B9iK9gEr
Or2KEXqkzkaQP6bJurIrLwrIlC1Yf8RD9mwYHQhcl1wIp8iVkYCxORWf38NLid7fa6VnP0NmPqaf
cKYc4qA7bAYt2fweXTQkxlM/pVFvksk9pR5gL5QhnzmSvpEt/BuWDadhU8hy7mvkbpUU0O4BtBhA
E93KTNEL+d53+Jx66nriq5/n8qC0JIJmyinu1eFbg0B4eKHeff4rE+9dMdq1iGVQeSeDBDSeDnka
dNXINF0f/UFh9aMqx6LpjbQngQ3FvYdYrUMQ95acCPdNzVDU1+v6y4ENnAhqMy1rHfey9R6yovot
8J4HBH6Cg08jQMeC6NBlwSI0C1pgxSaC+1Bdm7zxr5RdIkAMvuPJ+RiWHknkweKakJTv/c7WK80g
AMjLQ15rfNYTw6edQ6lRJgEC/ZIcpQFmXofbD/aqFYcG9UiiMu8rodoOALp3Z21tACPvBtM4rh5b
3F/hQl6KyAvuwIYWbOn1FFXwuCT0r9ADVRQgk6jx0qyLqwolEVYH0YF75kxhDx5DGdwxu1ogMrCn
qUlOEMTM9kcmtWaWsfDkgOQ8kKDWNDkTjkoei/PjmRSV5N1kjWQpLtabD5g6Fx2UyAc2a/wt89zK
p0TZiTaF0/dhIC5RCqslYQyN0ilLitX5FzJfLSKXcCrd2DDhZ2pcmVap7sf1f8ERyVhLsy393Bn4
+IHCVQZAlXQasxw4QSZyMKiCL93uxezn6hoNE07+NHAsHXwZZhcKyMYjRHio6FlaQ/kwyqkvFg1h
SkiA4m8doHNbUEXB3L7vYG2kT85nGJAS3RcNBSspEjDy5l9Sjc6yWw89+itdS3/U7vrHZuqK+mr+
hrh9MkTUTYIM18KdWy0FYISID7Ou95pQ5Por3xlALkvGpT8PWUrRprVB5btzbpE3vbPA8epoypb6
sRox6Oi6zJMIfuAZlT4bjlBFNCO/O2nlAA7fS6IBouSvkjZwMQyhBp6pG1xOPnpUbc0Ypc9rvH6b
luCVYn33Cw1UwbFY2CPCjXaXRo9h4QXv/S+YlqgZpL0DeqIIvX46Hfyzla3WtJvNbKnc4R8p/llo
a4zkh4g/n0aTGQxY/0CXREGKoHkZGVhLbNNhuipajSlk0X4nCPykzbM1Qlz2aeiLYnPuGYhldtfS
7nuix+mIYNdbxLQ/wzznbX09ZRWItzL4C2PBYPCXF/7dxV8ECBTp6ik5z1tmMKp4zcbXSM1YCBXj
/QI70vgrA3V8iCu94xIPlrMNST15RTKaI/tzkHLqJ3MmKXFIwx9yDCzwtKBaCKZ5SrzzR5SIKQP+
UZvcT6OzkoKbl3cRDMzorvVQAZn1JPRkCVM91hP0dF9VO2T5AYXgpj0b7hn0HO9/6+JaqHxUNSCn
mm7XY+zqU8PeDtzm3l2rYRrrBvMTiqSeBwHh3tP0h0sn7TN3dbnFMUWiOOmbDyHAieVqNAqGb1Du
yAroLaqwuN2BkqfJ1V4dXVMgM6Er15+g39JSjgUsRDLVeZBby80aN6rZoLEKDpND//7lEe5wlNz4
xvluUbVQtW0ujMcBH45cqS/kuNv5I2bmdoSOi7p7DE04riW2X76kM274lCdiJjTx3K3eQH5QzKcd
hr0JxgmI10U4Cu9I/6uc7mqqs7nWiG5FA42CsfPi2moCeQE4WTAqYzTTwT9M4rvyvV4Lj01BKS0V
Ogg0dB7JdsRvcK67ZjcQwdAZwxBA9JbqUpZznHe6QdZ+0sX81szCceE/Ogq4mwitupaMZX5K4FDO
bJs+g4958DWQNmb1kazJuxXs5KjAGuy7oElUfE0LXoJd7KZPNCiooM+u6ZQht9ajmAFtrsNsPNux
wJN0lmsWMqoeoqNcZ6s7Lwg7xoxh4mXT0Rln4LrdL27XJpxhAxyM4os5n+D2pQ4rYizh4PakFDJ8
OpimlR6wQDctN/Uy3Cq8RUas3R4FLoKIndda75mzXSiMWCOembG5WMJEd5ckghfA0Wgd6LnB9iwo
qosZkmrrHWW/b9tbwhpgQMmF+CZtl+3WEToukqdfFxj/Oe4UwFMxk5vqYlbtn0Z5CSjUnoC1cQ8c
SH2JWR7PUx+P5Vqs9yd+CqPIf+MCtGLFKrXY8ebwznVUhvMuiA0bPXrC2vhf6dvgQfy6ecXufhYa
WDVm+ebB3v3BpD01ewmrLzRQhBQ3AVM3eeBnKQb+ujvJrxT/TPxsik/VYx8qq823T5LVxkOmLk9I
wNAIhFBiMcTBERPdHgbzGwTDdDTZTuScoAnjfPe3fjjCzmE0L+6mqaxqCbUmnpngdT6aMQ3TmUJb
tfpEzD3Tvrd5SxV2UaURdSAGWdR/ANzZnr8mRdtM7zapXB/iBndmuyz76mEMX5GEARToVXW0Xwvf
GliG0K3WLk/y5S/D1tniLLFWh5qTyfaWGPoWfPkkYCg4ZKYij3AJuVIk/Br+xc6S3wCApZzD652r
WkuRPEW84uWXaKCtjRlmjZNqV/s9V5PJg+ZOdJDIojufog25N4ochORgYILjG0piNWAyiZa1s5px
Mbzsicp7uQ5jRF7Jwr6v+dw1H+Batl+Ao+p+YKkFhXne2rWkNTdKq1X9u9TqgtN10BvQfOk6OW0+
aoGILVZohOkoe4nl9nfRLTRK4nMkjN2/7N2OappnH1Ad3QGK063J3W5MPUdezw++xnWXamUN8Gth
CUMrvC/Whu8RDj/jeeO6MHNur7X3WJ6afRaiVigcGgK4/+4cLJH4k4f/oL6+mdGFL3mt7bAPMqoh
wtiCi2n//mVkDm/65b/Eu50sk+j3+KkvmEqMW863OV0n8rjgWfSO0ShLodVRyexryRNnnE6KIAKi
aqB2YthE48pptAK6n1tZKcIind55isWW4RXqEomBHbXqB6msKPurz3Dj524xt/ysacRDlgu3oF4A
/+DqDj2Su8eqfQMAim8EJ2qVvqFf3Ilcv/2UA49iyVnD5pBV407JarkzwfkZr+zAfPKpQWEXmCYM
nQ+q6pKv2SNUCygOPi9LApaOC3YVhr31fKYp6xPDKMxLPc5yKwT+7e9TtzwGlQOm/tH/QzIn4Mn0
Kw2gJ2V4q/qcy5Vot6iUGJOSKkgjfQkkOWhrM/uo7ETfXgCf8x5s0J9KA5n1H4jZFXZAeNNHSG6o
wFo5A8ZA/I9qPeG3XppzT+ebgtkNyMvws+TX/w98xMaL6yz2tPdrS6hQfe0o8ZNGEhUzUNVm4ErB
V/ifeOr74eqialnups31apnGosv6EB7kEKmB65KrxgRKJtK/0LzeyeHOn3IFXHlT/vyv/XAbxeA1
PsVsjCziCyPPGI2Jm45QJK2NPEb4Y8PGuRp0pMOAhN93dldU6H58h2oLCvkE3Yv+qYAouC1/0CBX
rxh27NDGfDOslJlxyhJBBIgXpqpb5EIdFCph8pZ6pba1BzKZiGEIZMQIvr+5wvSVCCW9r3LYmxKH
Alx/W48eksohC3ozTgebamhxVjjMEqT66bBFMvkMaG7vhjjqHikukJfS3U0LL8YqQJqj74p2J5wj
Iq8EdPbQIsZ1ev9JuOQT7tQySuDEF1ceWBg2tpwAfJVZEayfGtliP8u3RkJ5837GIZkjVZoF0/Rl
+LKDtEAmyVcY0aAP3S8SCJVGRViHQJtdUUWkdvkHSXzKIgHUDuDX7EWKOdsWOx+g622Le2o1M+rF
VhM6hTzXTYWNWO4IFSp7uzebobjEatXvDB3B/iadhiO6QCtrcIgYlRHl2r7QU2NPcsTt8Yuw2q0v
fmr2md/m8bc5qxVB+zA/sRYRZb/Vy3Z9IYp9JDN7s4II2P6O2pNcQ3473Sn+0Ik/pd3mhwl8fnv0
V4K3RFRDbw4aYY+dk4B8kMl08YITSGdqIGn4M4Q1nA9uC5gICq9Vr9/M54lN7YfmA26sdC1c9ikS
HB1evKFMZNGT1SEAESq9D0nSvmbLOKTCIPBFwbvv8w8tjMH7eX1FkCg0h6k+ymbRD5L6IG7rkwbD
kK1DbGlJtEXXOBMia9U188L9gw/ALQkUwEGjK+ebznkGdp7DjQTOrYHo1DXHZZS9nMZ/jnUQyiYC
GpYpCDwX0swttCYodxeTCmMMpspLs86f0z1jY9EVqKQriv0RiJ9wPWZjPKxxDUtkVPK0bIvMgXi7
hsr/muAVpnO2Z9bhcBQs426hlMUVADH9+SnvLeqOAdxjVmZaWSum1zJNNTcxv0ROHTUmPFI2LjYX
a8in5x0itJySiF4PzKFw2KpOH7buPDLYPxk/fL1N9Vla2oidtungpMLBclyev3kyQppF05+Z1MJh
S50m3NBYOlMAicpFGcsVqDb5A/MAupOi1apZ2oll6Cmzr2WTRtOelC/0wAcINCkPRCWJVQpjEzOa
L/bRhhPp6YO3RNwx+IweTvjO+nwoYHbhHqJB5XSPXVhxDZVE3JEsoIRXL4W9qEdQz1qwG9zwo3+n
NljoRVpv/SpdBALmoL/OqKx/Y2dh4sPa3bV3XROm3/ErryuFpiQ+7DgY6/0fZEoZ6it9HpccPADj
ZS/Wx+AhYkaWMAF0KoX7GxEfguwhpVDAa3Jp0kE4BHsHU6YpI2bUMafIkqZayuag/QTJrcjFmuiV
m68S6gng0kpkNdKc9k+hW9i9MquLFXWJXvFOubkK3YcUqajaBxp9NSuKKCubc6iFmdUIXNbaxr/6
ifMKyjPK0EO0lBRvD38NoAR2QgIsxIg16BS0FmuUCU+pVWGvJiusTdIn99uhPnNWoeMn1vzNRmQQ
a++V3s/qRYp6Usty2sXT9GfX7Pw3Q2d95r+HawfuIvjqefljF4+kL8CvO2rNm9vcL9hzjPTWeVNt
bWihelY6jNLo1Z2jl33JB5L8pte4Nfvhwoyc/kzx0U7dnL20mnmnesKttwFANiyCrsXmEhbG4ax/
xi4tEiC9vRIQIgNH6KzDbIB8qGYMthstrlu1A8p6SyGDtXLZWEewPsaBdXijfPGpu9PKkEvURVdb
+ro7Nzy6SThIM+m/Ma3F4qZ8h3Ag1ACOyrrmo9fwV9GcPDij9ZgLIS/+9+LTEE/7dlUWXL0oVrNS
0KovTaL4rCWUFvdADV7lwmEEVJ3hmQ5WcMtPQ2N28/jdtDJ/+LBuEidI7gNaAc9/cvYcwR8PNPh9
Hsy5hbjMYL7e9wZckyzuV0FLfZN9Bx+jN2j9oTOtsEANm9EWLSarHRz/ddE/37B9Uc1W/FLuMQO0
h3vg5KhcPZu6kZpCufz3R28+XfqnOqXGC4J+0SmlwuK03RvN/sa4FD0Jce/nZNE0b9ZP3IVGr9ob
gN4iJRHl94xxX9+Q6dSHgwSM6GUN9x89eUvThc69TqVHgqhSRXCDfpyUT0YqjvOvqXc0XHiP87M3
cnCCsNufASy0Yf2HB6WEGZIJUBjIZyXkR6xanWJGJLHw5B2AZqOj5HHMkAzoVw1sVS4EFfqSHdw5
k1IJdS74u2niqylP4CroLy3AzvDAQMAeYRTJJam1ghnMdEebSEVyKq1BmTbWku4Doiwntrf2n5Zr
lczO9xJaSqi0rCOMSZ7ylfpKVEIPF8TNUeHrjY1bg5TlBrDvWhtLBQVxWLP86aeG+jbJ3NGItOa1
IUMctSs+x140FXko176h9G8ksMJKzaig9wdGj6Pjmd+cfbLB1k6SvPfb/uHX4YsYdvp7RS+FFiGM
ZqhWckw57I+CJx9vVvoBvSk6Dj7HAxLV3Ml7z1y7y3Q8df/AvbxlH9PEddgHkvlrkADiMzNHkJuN
9WZFjsK7EhzLZlmnWRVSUZ1eL4jlWLuj7wALkW/oKcCGZHDjQ+hzsIq2ux5JDjwIIyIv3A760dBI
vEG64u0GwHf05kfDOxwgOVLLW1kogIbM8u7WDZkofei0MrcgMGuZ56MH6jP7stnimT1tRWdHatGp
9seEhA2UhPXDZNMbFepafXGvWuCr6cgz8N/cPPgqltP40xhvKkWx0YM7JMDD/qZnDExe8QkX+ual
wTNd5nO74R0GmbaYyuQHMsTm0yTUMkPHNyGrm+fFu0MvEijzGSqrLxS44fEzJaaBJhOjFza1If3t
5+rkAEIyqmGfty04TJX5/4RhigMcoJOJ67jdz4Rph0Av2xDfL69f1h2odeMlufKjkskPvBNsmfII
7Z23Fnm/ewJlVnxPSiahm+Rdfh2gN+Lpg6K7X+wbIA89OSQcztH106TidbtheS6fzVP/E9aRs+gX
38Ihat/+XZr34BhBClnPViBChVm4EiARTh+oGJCH6MI6j+kiS+Yrlt7QvNProDsQq4aLH/LCZP/n
078nhErLEA8aCP6LqkFYj3iuDjxwKr0cgz6DRNp2P3oZtP0cDdBanAvPPgmyxgDzieWMFOOri+0T
l/QPaz+q8M7r1a7ncyIRLcJZcar1fAK9TpIBNjxiucTWtc+sfkIZI0u4NWFn0xm163OOmFSKdsFi
cuhBa+rELvqm79UXJHFig/guZ3oY6J2FtmJcNBC+wyfu+Zp0dknkNnFhInxw2DxCBM5/UL6rtV4G
XK+AVoPLY6QjxmvwaFbsKmBQpiLpWikRQxAbBkT2JM48gF2GgeNvOv9VX9EAt8UBUnv/J6Cyg9JR
HybCV0Ghg1zTxpwpHlVQdcWa6Fjf1bscTfrhtSFdiAy14eDtUfjDzC8rN0BqT2Yrw9XqoL89bIRL
ZC3jGIaUS3VSB7DvQxgwRJF6+Sj6Lfc8qC2onTg4cBMr1ARb4fMwDN51PS59sHESqrjKBn5kJMFe
IM4qEZDWP8+EUEmOIFeC38li0SZMlKkbOUpCxnQuAgrgpf/UXVlJZlLypHm+ikiqPezqq+48p+Kr
/MT6VqatbmxALA6XoBANzuKkf+9p4Z7YwquE6+rk6xXLpPdroPSVC9p2M138JqdwyqO1HnNC/uvy
5WutvwZbqdgXQyej8HHOFdxrltuUuVCTldcrfXuoWSMpf7O+6dEvAzTY8T1M7zxoEUnNda053F8D
SyKK/q84kueQ3ctk4kP8AUFCiHl8Ze8nhue5cYJlzHTY684Z6dkqg+m9/Ej3fZ4/Lqps7yghLIok
79SUn3HpCixrMlmDdzh1TQxsf+d846oVDP3CI450/MuKC8AlLQhDpeGjtbwyX78TuipYL866jhzq
2hyPl6Zzt9lkJx2sHkYNoFfH3jwjuFxi3BwcVWI4VFsjrrJpjWMN8WXpHs4lDrOk2eXRYNKl3Kzl
XRjxN2+DAx65AW4rCf+sb+jFupfurYq6BFfNDQIeQO+j8kUKE37ELz9LmiqEZ8Z6FIqNRod7rztA
TaB/i8viK1oRRvbB2qz9LORLT8AZq5f66o6tj5KwFyxdCmfU5802pvSLuQ0qeZlVdjDdAhyv9j3h
y2AOccMKv+MoU1rUopkvfZXzrlYyR8sju7iT9L3hRxCzNZXAJiJbBhaZojkXV/IyxKBcILhZdGKg
Mcn3fbP186hNwxRYKcPNp6L5+zrVcPVRsi+EivJ1fhCr/ZOB7KuuN6Oj/PrbayHwrkHpfd9fUvLK
Dgr1pMe5thu8LbBD4/WDrJD1PqSxBTHm9Q+Vfp8K38ZHgG8YA2spis2eV6URom9CLqtlYvY71EQi
xGUZy+P68tsrgHeGJgmBOkVSSIbx2I43uX9pBI+srObnnTNv8ANSLdOGJvRX+ezfiJsmoWGlw/jm
dfHFes6QGwhWpJpKq/gXaWe242OHElzQda0AO80LlMWF2j4NbJVtH9LV2LbkjcbDMs4kNg8D8bik
N4abyjhTtqvvTPcNtSEOPXAUpvN4oSqM/ZeF3V3pYHWAQShKmXJx9ctVDdBHRKvPVki68q3AWkNK
0Pl9S8pcztJjTCyX3a8LQrtiHeqVBBhk0vyYyF8LX7Rn4/CxEzy+m6uMvbCjPHB+WQ5N1AT91GP9
qKTzXnZ7NyCkVGd//6nYg7xMZtV2pZ0WL2sQTwuAiSZlYaQba3UxB+AMULnDukHXc3zdBUouYyy5
B9u/jQU38j6n6YB4frn55+siX6jNQs5TAEOepINanA/HTl/QorXKg8vO6g2fn32OsoiHE+hAKD0h
nHb8vkbXDrHcv9legvA7Y3f4QXIR7+7qdg/QkJiON4kYhuHGrrlXX36zmEsCMqj5ausWsWQcNm3e
NJ95PRZAB40fYLSglWqA4XsT03K6lpKv2rRfeWSQPCH1G5r7zctSm+zzNpzSEgkahWQSs2NCa7rl
PA6NZRRNarfeuI/MezJc4y9VAnAHtMHBBXUOy1+dY0UFRta4BQXJIxm1JnLo2THvFFcd74ysMxDB
gvQoGuIH97eQ/k0Tqj6P+6PDnOUUEtIIF+tmnEgTKczdGBGvBvEOG82d1kx2xirHfKLRMq0QJKAC
X7xix//JEjgDbYTir1RXCBeEtGbckrfEm8XtgE/jDvt9QxdESlO5yj1VW17g5COd/vlqmIjcC8sT
Xd3Gn0900WKnmDPuYnKzzAw5LP3me8tz2cRiSaxfXvj6yV6im2ESAZqeZF8k8XXV4QNrYpR2+9z/
1dIwJvPWLMF0hHMChfd3RO1c7/yRf2E9YhS75CdywLgCha6Gcr6pTanjayVICjHzY0yiYxWPvdJJ
ofYSusA84ipMQ/VZV7JFMwXM3RTGm5DzgFOD7DR5Yya6pU5t+JzyiKozuhyW2WRwJno1OqaTA136
CyA6ybg89OZY+2ysn6tATO6VDO+Lz1f3Pt4X6g/wJW40pXLHi8+swwQm1d2AHRiaEVt/vcMYPo5V
dnF7QZCadkALwxGIfhZJfYGdTJZn+SDFX+09XbKc2hepQZnuluIxgpejsjVLJkrQMvJqSHhvojQC
yJvCn3oh+6SWB45LyUPh7326OMql3k01Do7cob1icVmWE4fphhd8wOJAfZ69RhNa+HzWwvTjDNBi
ekado3Ur9q1oyd2GTw5NSYM4D4qDi2IsqSQ8kAFeSCh4ZMy2fU5DhS+EGiMg6ptOqWm+8S0QC6Q1
kr92htQLthZCWygOJ6/9CjRf8S7guj4FfIRFIAQj4REmiammMJMdBmxgNrXZSKEI2ejeXdqgv5o5
YX1MJTYA+1t/cqQZ+twirQc+cJEXuBys7oFmEwbRQyDmkRMCPk/5h0oAMjM7z12SDUZOQ9gJR24S
WucPvkzXtcsEjvU40QAiGAFcyFy00IdqWnTEZcxS8eRH5EijBYFc09+VHKk5TWQeodgO/AUDFMLN
UMR8Fjz48TZeVbxP5/KcoJl4gnlmrKJbAcRGQNAiXjcZIUm7QHYiGwSbUtkkct+4QXbl7ghsfyjT
at9yFZqZaH1j0/oh3waTUqCUaAw4K6EzPzM8V7rOC31X5qdfSkqtk2OXwDWe428Agybi0jt9jLer
okeFRtMQ3e4Hf/w+17Tm3yldHBadgbxbEWCpRHQxE1pnQXmA+ekY52dlPP8NIOQ3AKLmsPE/D+g3
ZVfG5mz6eOLUqevVJs/EgseWhH2OjAZ/qWzaND39F5bo6Yunb0duHqkS2iOAlgl70wbkS6uiWlpr
uzJIQWV4xTf7zIrNJStyC/zNhVaox3VIL+Fhc1TLY9/DUbI7+fKwgnRMnOwq27K83ZIQMue4c68q
rqgKYcGySX57nfd8ikhzDZ4b9aslyTPRyuSyd+7XlsBwLZN9yP6TJ8zHvNrY1RkylugNZ5R8c+9I
sgNzULCkBWHT3cN4uUcHJxbKxtzCyKZRNedYWuwmLnER7DhTMEwysQVNaxriFd3BkYtSlt2kEJ2E
m1lP9M19YUvvcQClJKCRVc/qURnNy26m9ZqG02OgJwFXwNrMlGMjHLSVflVXehLz8l4ZSJtx5l2R
vrECDQ+QfXV3fMoMo1oZRWyirv0jTQABUFtQ+LADr0mwUOEy0QCugZKmAkLGh9gF3ApXAHWPAC0G
hqhSXVmK4TkF5BU8oK+NsQUJyIjhuzKDb56izqkUM+19Sa3lTUSc7QBlV3Q8drnaSsv/WGJbql03
MLb1TUhx5Ux4HVBplIg/A6FQqvlAEpFoYMEPQtXDIq6hVhIWZKuXzvKmrQZFoezsTYcmFukYbcuV
Ks1p+HXAZ76OCD096H5lW5U1LRatm03Br7NTmaefAIBrcsK4nQIkHK6ynfJSLmiVL+Hbje6IRzTj
MG1k2SEz/rMfVdQR+Ecbbsusj/kQvwkst/dPlLTAfmmH24kJ4KLIwwA3R/mKr5BjoxxLYN4+7YHi
Xzg8XnyBOwQBs7AA1Q==
`protect end_protected
