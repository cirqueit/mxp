XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����`+�6�cw�ɉp�i�7�VFYlg��b���G�|@A��ҔiC;��cz#�$<��^|��B�DD�bH�U�����fM�m0r��]�;�����Ǩ.�b�9$ؚ�:��O��� ��Q��4�$>r;ʀN���"�b�Q#�º��v\�1w�޷���-ΗYk�*9=4ǐ�썄g}$��]c��M�a�qiשּׂ(֚�inދh��_�,yt][�J�S�t�x�Ý/ ��&����Po��ɭ(�GH]D�Y�;�U��)��=�Pr��S��
=f�����J��;�;�>�p�~�t����|�m��6�C��W1� �o��i��Vȏ���h��\��/�ns.�23�� ,�C�>��.D��V8�0,0�4I�]����%i�Os��m�zտ/�7�(q١��cB��G���S���<�:�};"�c�Xo#~� n���"���(�k��>)\�6���K��4�=���k%ǉ��5�7=b-!���+R$�l��?ɷ�#,��脐���Ku��=���%vÕ59����6��fQ��d�2�n�-K�E��9'.���ܯgE���x��P;h���>Q���i�F����M����ܑ	C���X�S@.�.�
0#ia�sz�������MM���%�
{��0�7���h:���+*t
[zl	V�^���S"�Y��q�s̺L�|�\�D�i� ����迣�^y��!QPm �������%H�XY���ۀC��K���XlxVHYEB     400     240D�͙ʶ���8�#�8�rkF\�=q[>8O	�x@,�X)y�EPwϻ�<>{��V�˶_rM��t�3dL�Ȕ�申itO�N�nTsj���� �F��H|É+�Q�7!�m��mN�t�8��aMƔ+I�`�g:�B��C1���=�bC'���WQ4�%?����e3֛�>=������Hv��Ѝ�Qn��U��y�n=��7���r�;��y���!��	��M�W�����ù��:��;L։�9 �r5���i��[��RD���yN M9�b\�ɑ50aD��-8�fIx^0�F�%,�,.d>.h�I�5fܥ�aP�_A�#g���%��UP�$�m���`e�BU��nyZ����mR8����5oo|]'dN���$�4�3n�i��V��sK��)��,�}�X�f�qAhY
�~�n��/p��P$?��
��DI�T�nl)���) j��/ Č�4ޜ\)Po��ҋ���^_�R63ʄ6,�)vZX8P��ŘaR�`E#Ӎ�K�(㟠��]kTi��`��y<�BҾ���?;]9���%�H=�SXlxVHYEB     400     210���o��+�'
.�6�̇^�(\�O:�Pv�@)=��"P�����s�/�}��� c�	$H̀��]��f�o��S��ʤQl���7(����A��Xu��Q��S��MD��:��҂;6h��*l����a��[���<w򽌖<����l2^��>b� �����9�5��㸬�Vw/��<�k�ZT���<A�% $7[wthj�4·ӕ!�l���������$����i���_�)��o�(2�|����n\#��d��ӹ�e�Ⱥ3��{T�	_�cMR_�q=���z>{��GK-:A�uU �����Ye�(��	RR?�H���2h6����&�H�:!��˜���A�qr�: ą�K/��z�2���t|	���o�W�������N���Ey̌�W�4q{��#��1�� H�`�3 1�v;�}�t�vEh|3Qs4B2�,�*���SچrA'wʽD�Š;?Y�U�b5"�,�B�~ND_�$��d�?�}��r��ۦU������3���4XlxVHYEB     400     1f03ݘ"*��a��B�;�"\A�#���.�Pc[��񬑌:Cq����6
������M��e/�b`!�_:���mw����e���M�=���~�����l~%�:on��O#�̅��\<7�CO�1Dc,VpD�S>�Nƶ�RJq������o�U0��S��f�*�s �]/mD�U�C��M�D��
��.M2H��j���E�hH�k��/��,������9�M�u�	�p���./���u/+�p �3	��b�DcҌ`:��惚�[�c��ŀ��Ů���Q�p��0W�9�֌�� ���t�����p.>��]��v�[��A"]���!{d��s�</�&G�	q�Ppc�L:� �H
`*�L�|*����ty
a�=/���PL�1.�&�d�#�Τ��V+�`�$4�i�o�~(lǃ�Z�aX�F�v�����`���QE�y�z�Np*��7V
'my����c5v���p�?�e�oXlxVHYEB     400     1c0o������ëv����C�y�����槊c�x�<�Ɛj�~��D��?r肣�Ɏ�/!�"��.ؼg�R^9)#Pm9����!�Yi���Y��<��̈́pB��T9wÂ��n�����Y����φ��n*c��F����1M��K����H�;�~���2m�'�����M^�r�7pP��Tr!�$��|��Q[�}V�y����gb�g�����0�C��I��['UdkR���gy�UM|Y,<�.ϳ��9o�~�4���x[�	a����c�.Kd��\ߪO�c�u���[D�QAH�!�B�펰�Y�A�1y�ky^����CE��kH93���0�vr�B ,��ZFj@N��hL�Ejw�#]��c a����U��P�<�zwS~�HR�yi�Ý��NΪ�8!&�8�wB���(�!����vC,I҃�x�����XlxVHYEB     400     200-|,v�Qs�ρN�'��ғ�&�����FB}��F)� ��w��`'���	_��v�]������ѩz��ϺopK���)���+!�*ϰ&�xi�� �g�p|���� �	��`my��6���E��e�Zj�zi����t�r�Ʉ��Ø��Q�yB�����\�3o�U~SR��Y3;�+-t�VWzڈ�YƁ���lvн�Iz��Ĵ���=�{������ͿL8JVf�����0c�A@ooF��5��$bN��^i������˩�$�sHPF)�T��v[�
����5���>)�孁����&o�<���N��}���c��m���$����
�s��&5sV�};z�8	ѥV4\ ϟ�:QG�<���@G7ߣ)B[�l���g9]�\��3w�&^�ςh̙B�l;}]��)������k�3��c��	�zTO��ݮ����J���%�3�
�2<��{Bޑ�D�^/�?N��s�"	n��?�m9���;mXlxVHYEB     400     120��n�H�ҋ�m���ǁ9p��W�߶Y~&�Ui6Ex��Dw���,J�_��./$�Q�����'�g��FB����g��:6��+����n�?PE�:��4�f�2�U�l)wh�}�gE'�(hXC�f"��p�z���+�Buf�ÝDw���an���������xyХ����~A�{e= ��ߡ���N� w�·eki�E�kM�T��xck!�@�4(�>�R'$�a�*�T���L����B�l��c�.�7Rab>Fxjq=�sƿ��DF_!w+�F�XlxVHYEB     400     1a0A��Ԕ#��aE����y}��EK��\!�tn��^3􇦁���0���x	�F�TWz���>J��{x�:&c8���nZ��[n_�<������`I�	9ê�Z�^�K����d�+�6U�I����E-+yP�6�m���`��+���P���"o��r��r���R��ܓ�Bc",�p�A�Q�����#���%���N�����K�l� Ʊ'I#a�Ԛ�����?'��2%Γi6複����Q�R萿e��o ��!�]�Ö��8�O�0Ĩ���>P�KA���be�`_Ђ�����?�K��ܔs��fM!��萘ЎV#�^�І��j�w�b,/
wh�F����o�z"���l���
;vb�m��0P�����ٳ���M�wL(R���/�.\��)�3�V��p�XlxVHYEB     400     110�C���
4A���.��n�=����/��i��/�V��(�٢T����9upOZ���fUI�)뇁�5<�@K��j	����t�ҧ�,97��gx���(s���f������Ѵd�Ȱ�"�S�ə���1g��;8�� ^k�+@7��N��r���8���b���p �W���r%�nj�����֚w�_L6�~�G��{ᨦ�+��%�� ��(���"	����⚲.�:�8���x�!v�����A�%�f��I�R��H#�I�]E��~p���XlxVHYEB     400      f0#���ſ�۴r���͗&
����L��P> #�����c���Sتg[���X�_HZ�D¥��*�Q	_�:���h��<�+��_��翋�wR��tfQkd����Ab���Ԥ��'�W�0�6���f��=��Fr`��g0�{�j�E������x�ښ���`>C�>�{�hZ^�]���^�E_Z2��و4u 6�f�q�I���)��a}�����!�$ �L���.*ᓭ�����XlxVHYEB     400     130G[`��n�o*�LCP#��E�+���i{�^��"U�^�"3��h��Y�x�\���ʹ:F(r F��Fy���RvR$ߩ����r�XwA���o��],9����1�Ͳɷ����ooG����2Gpe����Ne��������p�b�2BqO��=���韭���U�Mx�/S�\="��>�Ǡ�Z1����C�����>ǫ��p��gf��~{�6�w� Z�JI.�kh����K:���k\�+i�=NLQ�1�yJ���x�B���b���ʑDET��U{�ԭP<�QN�+�#fE��QXlxVHYEB     400     130U�}��ziUML�6kٵ\��y����胷��B�)�M`���Ջ��"3*���0��9�fA���K�X�����M	�f�˃�͑�J�R{MgF�q.�1�+:R�?��$*���H|��d�;�g���7	����� �#�0�if���#+��+j^��wQ=W)�9�Q�OmҶx�A�H�h-�.=�XT.���Z�`h9f�yەOԪC:F6�Y����A]��	Y�&�ϲ<�i��	���f����£(��6'�!ho����P���X��h� ��DxoA��]�J��CN�	XlxVHYEB     400     130!"���@@��;������!0�,����������(�Wϒ	�9�JIh��
\�Қ�LR�]/[$��ߜ�������RG'כ?7J3�%�:��Cwa�a�CZN�*���i���e��演��7qLU��W�SI��+�$���O�;MI�w�1�?c�é�G�K�d�l�T�F��5r�i=�����r�g �:pVD��R@`+ S�3%��t(8別^�{Nd�O�(��:�9�g՝&�7	g�h��h����~�bT�)|�`w[C�ڂٰ�ܡ�vpeլD�#?HѴ�Y���XlxVHYEB     400     190I�@i�� x̄�2 Hy�%�s��@���o�n@�g^R����{,oY+Q�S��TJ��9H��J`TNS�����|^w�﯃����ݦ���Q�݁��&@��`�+���$���g�󆧤�`m��N��#��[=�y(�;1�m�r�B� �r�2�	$�|ۡr��~���*$��|�����J�P����"o6Nh �1X
(�_J��D6�r�f�s�t`��6��(����3��+�	 �ySE��.Z�Wh��72;� H���w-����T��-�߮�$��~�<��xc"���N ��o3&@�����3O*���?��F������.��E�CYs��o�W�d���1���3';�}�B:��M�Oa��OHI��bm��NC��
�%�w�XlxVHYEB     400     110vr��w��g';�G;q�S�����-��Mkf:�C*�VPhN��( x�fO��Y�ȍP�p�p��d�)^U�%�q{U�qq�L���z֛O�A�����]pU��Q��N�F������~3�C�#�{���C���Ks��P���M�M��b������,s7{��;O���/B���.&��n�ڠKv0���t�������=�n�^l8��b"�;.�v�T߁9T�ev���a1	D�<�Xx=��|/��v��[����J@��l| ��Dtt3�YuXlxVHYEB     400     1b0\S"�����$.���:���ae3��3\�B�Nj��H�D�	� :u�̐�1�x��b����/��r]>a�)##�dO����`g�|�2�%G��Q�,�Lh�dM��W��|sC��fP~O�-_���|�5�I'Hd�M�
��j�n�G ��x�f��1��͔�y��o1�{���*iJ�\����E�T\
��`��=�+�����u��eW���0�X@SZ#|GdR�� ��hC�RpQL�$�&��5yY���QIbP��S�<7J��Q%"W��#�Z3D�� �R��l1�4z���|�M�s��U�O ��R��e���وQ�n��H��s���X�����O�`�n]&'8*�����|F�]x)����Xp��m2eId@�Y��s��ȉo�|��A�"���q�����XlxVHYEB     400     190nvG�m��$�$��A���%��t�A��	z����c,��92�} ^~�A,߁�����̞�b�^��%�͸�#�>

����*��$E�O�v�Ɏ�hGѣ�gm��x.�Q���6\�]��w��QQ=(&�to��^2��QI|�_���\�������,���5uԤ���qf�"����K�A�����p�{e�u�d��v�_�̆�=�"Gw�_V�� E�w�ڴ�M�%C���N�3��&��%��@��8XoQ���OE���_f�n5.X�H.�h'�W<��5�28n{°�	� �`f�$iU������؃�9�l *�.���bY�ꞤTh��Z�,</bډ�T�5)k�Ό%Н�
ɧ���S��8#aR��0>�)[��gu���XlxVHYEB     400     1202}H�"gc�fD��=C�Xz�X���:lN��TOn唴����S��a���w\Z�*ɧV!���04���(Tx\��!��y5�b�R���o��e�0��D(^Z	a~i�|V��/�C.)�)>�S(U�śd��n������.�(�7A�^K�i�&qpӯYh0(��o#�w�L�PTH/�~Z�m���f+�9�BWg�>�+G��̝��&:�t��i�^)F�c��d� u���O]b.Ď����3�L,���w�b�#�=�B�2 (�e9�b��JXlxVHYEB     400     120�R�6�f>��M��I��W�92,����+��4��{R��*]��#��r	�q�b�2|$z�~��vc5�(��Lt�Y�Uz�h Y����N���=�+����̻���D��9�O�Fp�����9���~wW=ͧ���w����z8�)B:�l�lyw��_
P<���y���ON0&;��HR�}30�Ȱ���?`R�-Q�l�C��i�䀘��2�˥`<����L]ZiVeW�<Rh�������'o��w�S��=�e�uh�q�BH����-XlxVHYEB     400     160���Fk98���:3ꊘ���6VR�d�
jy��_����HcLeǃ�����p��M(� z:n�I�Ŧl�Z�S��A���&��90�tƆ�2����&u�ް��ٚ���D�D;��UE���A�s����1 �Հv�z݉L���ϯcK:��Z�� ��y_�Nl#L�E�^=	ClP�)�H��p��BxQ�=V!\т��bFP��3H��'M�D���Hy�6e-�m��a{=Z`B�o\���,�e�m�qw	��Vf�g�Q�zցrOΙ֏9V���F�C/1��BԷ ��Y�E�̴�d�V�:�us/�K�ԍ%yG����?)#=�)e_&��D1j�����i!��XlxVHYEB     400     150�Z���ų�p_���׆`ќ�N�+�����
B��6��8D,�d�����^楻'�7S�(6�u���\ ({��7N��G�\��q�D�m�VH9�2@��Q��t�Ƚ������P�������p��b�&�wX�>�W_��*�p�� 9�eذ����[�Eu؄�����8AF�V�3��.���B`��q$N�%�cL=�٧4�jS�k3t��{�g�c�]Ҧ��ks��93�V�K�r*���� �7�o��m�'��z'��z������_j��h�R���i�7��|'������V��Sp�<�L[Z~�٥��f�1׼����ςm`*XlxVHYEB     400      e0��v��䩷b,�zyzu����sfe�v��xtU�բĳD���&@�N��˓,C�_b4���ƹ6���o�B�fW�E�!n��Ud��9��J3��m^.8������o7b��8��S"��*�/x��>ц媌�5��G�Jwpn�>�p�Bce�	����8��O"5��;�rk�T���X�H����3�����0TR��ۆ�9��<�)}饸^�XlxVHYEB     400     130uq���d��G��|R�R,��7V(z��]�_d��,|��>�xh�,P��k	(ա7��2~2v���/!�_
����j�� �Aذ>�V�tTd};����
���d�L&i�ɫ׫?&�,]������?�Y��\��9���3��E�(�l�l�i}S&B�Y��n/�a�Q��ڈ�t��R|$k���7�5!�:n}.����$��7�S$�؇���K���?����& ^��j>0ܜ�SG֣��B�o���d��	�� ��Bcs�:�kܘ�S�ӫ��wH���y��(;Yv�M�
d��,�XlxVHYEB     400     140C9�#�-�;twVнO�2��:)��Q"���s�����t�-Uh�n�Lw�:"w`�U�t�ʽaM�bq���Nد��RT�&%a��c�4Բ#w�a�������}�4�	O!�e�`;��w��xy����7�2^���֕7�@&��^-�����,���gޟ�I}�
�:lB���E��ͅ�'fԅCw9�=���o�j�k�8�IU�U���z���[���6��Sz�0Ѻa�	-��)̞PC4s�a�һ�y��f,���A��B�H�{���,�wf�|�����j��x�a�!n�p1������XlxVHYEB     400     150�G���[�?���E�Ŋc���b�y�a0(���쥜%�1vt�dDX�ē3��?})��V9
�V��w��$��٨b��[�4�"��$��O\q��H���]��H_I[5Q"~�@|yP��zK��y�@�<�6_���bF��4��[m4���S�=���f�:�3�yտ�A��c�4�\#jV|�W7N?3ΗNY_���>.3B��?�������0�@�7
2�ŵ쵅���f&����f`�k v/�% 4�W��\YLѭ���;���� !jPؗ�;��3q�w0μ ]�4 F�r y��������wTr)��P����@�Il[��XlxVHYEB     400     150��N����Ǻ���j,}��{oѢ�e����J�
�Gx{���_�):���a2�E�Em~��9❒��a&��%)s%��S�<�*PK� ��gt`J���+��O{��x9_��
�5۩��I��IxE��pnw�t���̜���Њ[��A)��;I��z��bah��r����U({k�n�H�p�ۼ�@��Yνj)�BI��H�Jg��&�d
��C���A	��V(��;���W�$\�JKۧ
F޼�����X8�md�Ij������<	�╾ɑ��Xf���F��:���5$tHda� ҏ[��3|4�l�Y�p��C��XlxVHYEB     400     120ӏ�A;�؉�HƇ5��t�x�z~g(�<2,Pp���q�*@�6y��T'�;֐�����ϩ)�G��Ou����A�zlں�׊��d*b(?��g�dA��Dj�B.òJN�������:S��Q�ޜ���4+�\d�P?x��מr��1_�y�h�#���D�E�E���	�/��'���2:���UQ�BHSt��ӊa\fO!� ���Љ��!}LNIyn�������&��H
�fջ����'EۨD�\7B����{hc{Ҹm|�T�X[f�!�;DXlxVHYEB     400     130�\7���3tٞ��2%�%��At|�.� )��HQG�:��e��R�3	�0�����-��]�xՊ�� �\OF(��F���/)�N�JVb�w�R�C����s��Ð��jWQ8_P�#,)�Bwǝ���fA��J�g.s~�(��ü�����S���nxm�^Y��2��-�j�0�hG�e��8�llC�b�?��Qa������)\Ҥ�:x�e.�X�r ��]$|�b\[�lb�U�Y�m�P�.*i}�Q��Z��F�52��1z�:u�B�*D� ���H�ZL��q9"NXlxVHYEB     400     140�^k�0�����#z:7�:х�/��z�D��.�����&�Y�dBBJͅ�Q�ޫ=�w� ��G����ÎI�
��U>Dz\W�d�MѢh
�f14��c����ԑ�vvy���㮙Pe*0��!�� �ME�h�k�g�QY��=��ݐ����d*ה�m5��������,=}
8;|U��)�L(�}{|IPγ0�v���Fc�B�*����	��i��m$����Q����N?M7s���f��X�,Dfm��2��e5���b��|f�F�^�aZz�]���	?�#�w`@�'k_M��XlxVHYEB     400     120H���z�jx]�����u���P{����f��v�v���UP����f�5�N��Pn$������K6�,@�aC�g��72N@�Q���]�ƽ0�痮d[6����P��[хnd.���a��B.�um���.����eEt�f�-��Jf2�A���������ZR��	��|u!~j�:i�ɢZ�h!�}��L�Ra���{�"_%�8.��&J�KM�c��H�(z�K���@�M_h�����;�ҿ����j*���?RRv(�=�{�3L)�H!���.�XlxVHYEB     400     150M?FAC"n��K�H!�:e>y�Ozu4'�: 	ԖƜۚVl)(��h����ƾ��?!�h���L�� k�&X�Vx[���]�m�������n�iB�+��4����qb_�(��IoKB���N��.;��˷�4���z�t�X�v��5�B�:�X'p��9 s��~Q�t�%<}`Hi����O��'+O7\�U��7#C>ٵ�d2'wnh	��ݖ�Yg�������5W"eB�2di:B����ҡ4A�Z�7,-�����fx@k�iX3�����mP������lJ?J���/�!'�m�d�J��@���w{���\v)�w�e����XlxVHYEB     400     1509�@lx�ڻd��5�K�&L��e�箔���ś��R�����|R�ɵ"�5�����v���%�C鐎h���e/�`l�I\��|�ZZOi�e=9J��{���:	%�<�N��L��/�6�[�ۥ�)��@�b[/��Ctf�"�2mތ�M=�ӿ#`�����6���)�i�������tX��I��4h�vmW4:E{nJ �$�d���S3OH��c.m�����.�zvp��Fe�{�1U7�H2&;�a.jF2v���9ن���G�Z6������FX'��8�d���oq*\��8N�WS���������"�Tz���G�L��ao�i�/VXlxVHYEB     400      c01�	[�h^)}:����J/ �GҔ��� �a�4AC>�Pri^]�T�1���v��z�\�����H[ ��g僡��P����d���b�o�˹C��׈dw.H�L(W�2_uu�i������&=�9���+���0n:����O�V 02�B�r1`Զ�8���+�}�����qШ
�b_XlxVHYEB     400      c0nmӜ>M��b�ֹ1ti8MoCR�<׫��wI�~�c���:)�U�UZl5�oZK�a�9Ř�X�yʜ��*�N&����&GQ|8�G�e\C�KC�r/����׹4��cqVP'֩`U�H���Ӣ����eR�QjS�%*>��`�<���is+�R���xt:.�&h-O) �7����D4kXlxVHYEB     400     130�����t��~�U���4R����>��)�d���x_�]2@��ٱ�S�Fx-�D��}'ɮT�����r9@�+~��i�͝�b�݁p�
�_�TT:�yZ5:	��b"�z=y�jo���
}�^_��������c��rM��p<�G!�:,����}A^^pÆMiGWG}���һ=�P����+��\N%� :4 ��S>����$��؂���G�Q��ַ/�轀 NVWС�(ŉ	�c�8�M��/�� ��w� ��{l��~�hT�Y��!�<�f�%~���_�=��XlxVHYEB     400     120�r䏰I|��2u�m!���዆6��`�G?�-'*.�����`<����N��\��o���zz����%럂]�k�,h�+~�g'?�^�)z������6Ŧ\��<��f8�rN�k��3η�q¨wv�&Q�!�w�w;lT�Ϟ�5����n�jUi�r�ie�{�1��s���%��H����;��`��L�'c�Ե)���7q#�W�	�*�iQ#.0,�/-|3K_H\;�"�vh�'�\OגU}}�᣺s&"3.�7�3��4"�5�lF�XlxVHYEB     400     100��ۥ���ḑ4���H���#ϡ<�
������T,0ID��#�!�^h���}3�+٘��h�V����h+�N+�d�%��KZ�=�[O�������Ni��T�"9=<��U��+���:�9gB«t��1�h���1����,��Ȋ'9��.B���(hFE�3�{'�pR��ò�]K�j�U=_c��iT{)rL����I60O�'�JQ(3�n۸��n!(�i�8AB��j~m�N���#qİ	�kӼ�a3XlxVHYEB     400     160�xU��uV���g��E]��mΈ���$@`t�%-oea�Rv&|(Ԟ!�3(?�~�F;�}��m�}!A��j\�ٵ��YrY�n~Sȓ����G��R�����0(��αF*kaR����C ��g��1������O�}�+�B"��A<G��p�Cd����u�s��f~�v��p�����%����W4c]Ih`�N����i�8�@�F��Nϩ3���T��|���-�j�Jי����+���Tzk�a���<X��A�bu�.U�R���� |wp �8��LQ<@�7�2gs�nA�<�ãli�� DǛk��+%� ��J�b�F<T�J:����N�8�f�XlxVHYEB     400     1c0��^T��I32w���/�|Fh1��Gw��\^cns&�Q�YR�=�����1wS���[��L(���H�P�����$��w=�����	�.�L��u�#m���D�&���\��P�3��Q۬��UZ��|>�,���E1!�-@��f�3��Y(,6��CeZDJ�/�We;)���>���|a���.�@%������>.�*������ǻ6'@Qj�c�t�������zj9��ѫ<H��G�)�P[_�G�r;������2����A�k�t��:2l=��j�>K]H�].T����O[��# ^���%^N=�7Y\��Ѷ1�b �t��JW6�/)	p�S��t��M�rI0�@�b�k�V������6P����$��K6`=
�=��B-�\uĵ��?J��NT��N�0����H���=O/���/XlxVHYEB     400     1d0W4~���3�=��I��!'���^!���^�܂L{3�Ţ�l��,g�p���6z��f"�2
�r۾%^� ;�w���	�}+��*�ӯ�K�E��l�^%v�ɡHr��3�-���GK2�@6�Y��'U�R�h�������-Bاq|��>��^pV��:�;�|�DG����������U��\j�R81���xųb:X������&"c�d�A�+}�Cm���.��~�Ms�B�n_wn�4�
3�E�H����֖��Ë-Ù�٭�熶{�?�=L��&�C,�͠����(��}�D2f�A۸����U���A࠼n4���d8�ke��6j��!H$�=Q���̿wJ�2pf���u9� ���?�w�P�"p�AX�����U�e-=�)���P]e�l`&N!L�L�:CV�z�w�
5sB�ܥ��Վ�v ��DM�xVL�@���1XlxVHYEB     400     1b0���%��!�˼�|7�6���a^�D��[q�<���O�������--���� 3޺lF����<i ޒ�x}b�p��Ht�	��9U�CaW'G8�%<i��Q|go��n���o�y�ࢠ�.2k��]_���9U7��(gh<�p.�ҳp̝�S& �]셭:I/U �
��E��
��QE>�t=P֔�)����^�Vl��u��+�`�!(V����MF��{N���c�/o�۪2˼� ��آ�ݧ���nG��K�۟�{�L���AZ�E6mTJ������4k��RE��J�ve�U��dқ0B���{��2/��1�k����5����^�J�����t:�]�����HE�p�@�ѷi1E�-{ Ul������J$|�!�TAp�y&�i.�E�t�N�;B
�6:XlxVHYEB     400     1a0�۔
�5��A�:�^��U6�Ɨ�[k��ӹX �������O�o� u���UL�$R�{��( ט�,�5tu,�K�QDNeD�?�>Bb���jG��U��uaF�5�H�Ci�&h��v�����ča��~2�ANq���8��F9ͤ���?Q
��i�q�_�V�ß�� �4�n �/Kh�!�?H�{�Nbԁ��5nE'�� ��h�&`�p4k`�h�\�w��d_���ܐ����}�QO>P�~�t�/e�-��5���;}��n���UX�,R/^�|�$;a����E�Z/f�w�r�d��E�(�0_��E��B�PC0���;A���K c��&����N�l愅��<������APK����#�H�v7H_q{���Vڻ�R����lOe�\V�r����B_Ƒ��XlxVHYEB     400     160�Dr
M��t`i�n�\����k���qZW�������آ\=����K=͑�d�I���'j�zr(�B�n��-��̇ 6%5���e|Iu�8���'Hd��� W�N~|2ҹ���yA&aѽ+t�#�� �e�U��H�A�*�K�P�|��M�1���Ԣ�Z�<f��R�V�i��)ה�y1������A����bz .���\P)�y?9�]pF{���M����o:71O�"R��Wϯ��}]���O^:b�GRI��y��n�����@蠏,�/vP��?�u���A_�8n����8s�A�>���5/��w��\9�O�A����֝�!��pl��?�tƻ�opCXlxVHYEB     400     160��wGb����=]3!9^��,�F���e�� ��x%lz�R�v��4�5�{��$U�s%�w�c���+5��3�%��0*�kí�$`�}�m�f���a��TV��h��|������7q8L2G��)�����yNۉf��ʩ����|�����C�3̤��\��&��G�B�~����v)�.K
�Qvtq�];&#��~�8&9~�o�}�,0�w����>����ٓ� ���u�Ҹ��|
j�O���K*3�KZ�/�&<�<�h�(��G0t��t1�~l�����Y�`��Ŵ��0e�$i� Qm�v;��4�g��C�U�*t����j)�u�����gyXlxVHYEB     400     180�j��N?Ъ�5��6�9�D��Єvʉ�1b��+����AG�1,i�@�oTZ�q౾9�Uγ� M��E���e-	>�P��#8�_��d����" D�]P����h�r�����>/������J(��*ަvF�V���k�X��!J|D�&H�&/*�ZQ�@8�q�v2pP��]Ⱥ�3�ݞ,l����Ǜܻ1��\�`�ߨA~�����F��TZ16R��zYm;]2( �!�����u[���M9�H��w�x$�- F�4eZ����{���Z�c&���y�� U��k5��c�-:�T	ք��gM����Fb�.��l�<��V��rs�F4����[��"�D���
�N�E���UJr^K�p}5j�F�q)b1XlxVHYEB     2ed     130T�;��H�;$�'�*7��!ɬo|�5�qr( ��^�28��l�?ܸ��O&ڵ�s���_��*����(ت$�p���ڤP��n]&b�`�J�(Sؐ#��;qD�2�w9ԥu�+^�&	[�7�����J���ȇs�⭸����i��{�@�Q����"Ӻ�$_����H�����ѕ��b;�i>��g��X���z�0�p�̉6���߼q��8�����P��y�o[_q�j�B�6E�w�G��p��]��^��M��4ڹdƃ�L>;��~~�rG�F�L'��m����~��!#���z��c