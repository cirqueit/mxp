XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w�X�}f7�-��S)��Q�b>q;n�b���z��¹�(�[��uܱ��q����Yr{���E�]rab�H<y��������<��M<���l6�柟��)�)G�cr��i$��6v��� y3��l�.��T��qd#��������+o{���� ��M��Ϙ
�]��c?U!Ds<M�_c�ONz�ۖ�+��x����{�q�B24��kn�w�ɗ�ۡވ�Џn^�d��䄚�Ts�)� �(;��tHr�s������KJNN�<�6Z)"�ڎ�=�\�N7�{���[Ն�d�W��(��7�Y��tk�ժ�9��_?�.�csk�1�H�f��VkD���5K7�p%ꘐ$k���N�$�9�V�6,��P��oK��W�ѿ��+�WH57v������?�3�ytT�]P�;���ZCB�$s�����	_��^�����4�z����!��64�$���Qn1�����%[�A7޴�$���Lxxq��ن���_��IN~�ɑR�)�s�s���pe�N�7}aw��zpJaȔ3��k%7glz���gR�*�o��E��p�n�9�<	*6B ��G��e���s��NǨx�nT�;	P�"v{xX��ɞx�SX��Z�� �{
��j�YhyA��_��ݠY���A��_?��r\�Keڊ�eP���u�}�KM߻\W̠���F��`y �1��3�zW��y�s���_ e.3fU߅���u;QU�2	�����a��"�XlxVHYEB     400     190���EQ�k���C�b��ދm�:�@�ŝ{�U�0ȹ�����>a��7S��:�T�K�?<���3����7����U�aw�{��{��@O��E5{Z���T�%c�|��c,��"X���F�Qw����3��N*����T*G����Jr3"�0j�@ I)C�J����C_I��lq9aj86@�YkdhrE��kNOC [�L�M���Q�O��6�:b�k��d{�����fb�DIvE���&*I�K��X-P�IF�p�Q�H�H���*�7���r4ɯ���e,�܊[�9�o�8R`�֩4�V��PM��`|�`B��jj;PY�}�����~��	�ޥ�K#yC��X_d06Vvd��tF&��6P�Im��xٮVk~`�;�XlxVHYEB      3f      50k~���a~����ܸj��pP�)H H��_���-��L�����C�Yн8;ĄשN.h	�3;��}.�	"��"���Q�zz6�