XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8;v��p��1F"�%��+M��!��=�_�;I�g��5R�UeH~7�6Н_A��i\ �A���xL���م�!�ߚ���u�� �<z�M�47gk���t�������˅��<��=,w#C^� V�e%�R��ec���/�`8�g�A�>Y� �)��i|vU1�lv�ςrʪH�Y��h�j����&Ǹ
]�#�����Ԥ#<_�d��F;���!8bPc��B�=ټ"
'�a���su4�Ki:IG����N6�*�z�sZ�R�^x���J�	=as�X2"�/˾@nm�nN^����sP��5a�0b*����xE���v������|J.j����j ;��� ���F ��?{��ACl�$L�s�s�"��D���N?���ɬ�0�� NT3�s�"004�cu���k�j�b�G��'�=�2z��*��\�$�%�`5񠞊I\MI����'���������K��8ȅ�F�]y�ͷ��u��Ѝ{�v��o�|#Z�����ђP�щ��\wp�ȍƦ�x���oG"ݭ������ב��(���ֳV��cvc�K+f,J37�ՄK�{����Y�.����Dg��u���j
	��-�yנ|MhW�~��P�F~<��#>E���D ׎n-odu�!�C!��b��-��GO�a�)嫂~-�r�tj�Gst���a�p�sW�Rb��Vw��v^*Bk�kSgnp �ęL E�[�>�2������utVR�7�Y_�K�ˊ�Z��W�;Ø�]�>��ش'jN�XlxVHYEB     400     190h@S�?��<�/�`�KnP�V|�rRHY;qH[t�i�x�H��'�(��e�zށ��}$j�=����K��~��L�<m��;!�ܘ���{��D�`PZ����L��
�l�OHm�Ry��?����!���d�dc�>i��%1h�>8����2��}� �K����CC�B�LlҰy�~w��xm>9��Awp��2����BH�l�َ{h�>�8�1��xsֈ���Đ��/�N�{��s�f��7���r ˅�J�B�v��q�|̰P�"�+@��ْպwy�"�Rv�x��x-��:	��^Ʀ�\i�3Lj�}�>�BTF�*�>X?p��ɫ#o�m\bd��n5�x����u�ddn)J*�ig(8q-M$��?~���HNXlxVHYEB      3f      50L�`/��_��E4��I�L���p/����YS������r�[�D���"�H�� 4��&�{ϗZ:���}�mCy�