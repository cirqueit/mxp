`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9152)
`protect data_block
EmvOZQT6a5gKkDc8PhfBsJ0GLrw0aiFC75yUZaVoMVhh+YXfn/hiQ/IKAUxG2sPsmO5jTimjUlbR
ClldoZDn00xLQ/JDOWbwlKDt/XST5b/ryryKIa6OwqYrTXWTYMrorCwdgeZgBVuiV5qBNSbQ8Vi0
moa5DlqzOuZ8HK704kbJBDQUBJiS34hVeptYZrrDKszfrxsxTPz94IW/jVJU3rQCruTvp+N05IbX
GI1QprEJ6DEmXNLvWL8Fkm6rQKV+9yCkqeHL1WFGfdkQO2yA95QmmQICEQka8USxChYYWGmFX/C0
dfjC/0UTg6Oxr2pQoBWRaYXbFFZEPuWYa98fF9mFqEb2C8t1k5BmX0s+3S30kKU4V5V7iSj5eEgO
6W3vhaONmnVrPBhoIa6y4wzB0PBRRbsXbtW5bFAlVA/io9JHNPDmNntZIWl4HW6YVBIKrB7WHveM
n1vGvVyqMJ0JSESnd+9s7kxHTKDDAUh4RQyLdfrv4nwTKaDxXyh4xZzctmmmu6zkUASJ1tAANdyh
05A6WzKVsZDAIiXW3VpJsIRAXh7k9akVzaoaEf+CEvH+O9Y0m5u4Xsi2juq9wvjKMrCHOk9YsfNc
OAShR2fy+JcZtyUSb5fo6tDhBx5NkyT5qE3YGYjHkheMpDgAuMHKv64B6J65gy6w0CqjgHlpTMWj
fm44Xsb/ALJLhRVK4bxbVguxzzswKyxDXG0T+V3euQzgOob/LDuVYK4A5yfGrJb47Gm/XS75HQCB
ZQ7TC8jNRXpcJgTlIG4BmzSIevILRGXs2qWhPxGeaMseHLywt8LFIQGriyP9fBnxMo8bbvz8TUL7
hNdDOFqwOBnHruwNFDYf6CsVFNHRnmV3SPSuOkoCQPUW4lu8hziUPxZhrXjXR6wrymSVKG4UOjto
yufQwQQg9yM/BBijnVocKKsECxow5iWm/ciaPMP8pIHWMur3Ye145tagVpBiGCUyy2uOnh0nocsT
bAs4k2W6ohLCzBqausUnZpPCjNxMYxQKW3ckEbgkojTgXa4YPd9sluQedGH+v4OH+LAQ9ue4z1u3
mW+7lBjSdICUXznJQIjSaIewvJttBj0U33KKL0poXxEijVVTyHsPFbKZ5PxRlXUoO5xJ+cAA8gHd
9mi9yplJawqq+s9i8g+3NlHl/UfwAfNT6I4cWma2EuLYdtD6/QPUlVIwH8DjHqmaw6cBxKUByQ5L
PHxmlUHHs/RZebtayIQJPX/cHkiOfcGMHdh6tTPf2MJaZahAoGLuvAOTP4KAMyroiR3Q5eJpqCx+
QPR/X2bl0EweGiryt6UBubl61n4JLNXoVe2SNV61hGwF8czaEb6SgiuJvwdD6hTagp6PP4SolM02
ltSDQZ1cewrWWlgG+pzR6VdIy72P3ROsdE/CfyVdUJmltd9dyJVtz+xE8H7dPh3w968Xk3bvJfpc
OYEdxYqr95sfOrtxdHDY1VcwXJh623/IwaFMYUxayNrEqLBsF+Wbrwtu2R8IU9sWTKwJYdnkSAM6
J6iMPNAZvd9saX0dodJHfEL/SK42ERjW7wlbZqIJr3Ev4lgimgieEUF9exWgpG0dXze9RqeRdZaD
mcXYHwamnZ6Bk+BEIQDukiSNi4ac/apntYRBsWLuKQ4cnkAiuAFQHeO3YgSkFhlkIuqEgO6vC5uQ
wwQDNu5hZG/FOxx0l9aD6OjbhsLIqFNLOVZMqzL8EoTZDgmLqbgs8xGYlUg/1fPJGBJNiAgB/CTT
IPgJR4UOXDCWgLqyi0XdPgM0nZz2U7evInlL0qKPQlyJnBniSC0gQzZ8OztnbNBey+CZqB5Dq3YH
xpxU4llv7VgGemjrgKa1qwx05GDgEi9zRmOQLN116w9muFBtPqIscoErQL3kDx2PmYCjbBeGhj4/
kkZIIQvnD4+bY6nZs4HolhQ0eWwQHD0PJv5152wLWDs/SWSHT4eXoFuKXx7GKm09aM1GIXjCShfo
aRtRJtEk1IxMWgqcrLy+g8d1fTS4reDmSBWRdeQi8sBhMeHULjGPfmiHm+YeA0Df8mjBk/HJn9+Y
V96potx/Rj3NWg0LemkO1FmIoJTbsR0WiEFt4+HkUK73jF1v7+mxOsN6p/3fxMQouEufniJN+w9s
hoL9bQNfMAbZgmNdvMOLUA2KUvnWsMAlbzWC0ObTMyjbQM5QMA+cJ0Lfwv4xwBF1z+odVouvF/HT
WQQABIa6edwDnpYtr3kf7cfnGJWv6W42q3nOmpBpLRU96E56x11/FKody/Co/tvyUorGrn1l8SIq
zWjZzyZMwr5c0uBY8PPNTdqv4YurzlVjqAKdkNHV9Eqz/Mm2mygDU7r33IbrcZi2NLxV8ElVHbU5
vA5VthlxEqLFmj6OWN+pDo5I2XUKwACa4iNwP2Rffkx/GGqpB7aq0jSxaNMMhhZ2XNOKRfEdbWoV
crYck1dwzNZ5pm3vHGFDmP9XJQTnwGMVZ0l69I4+7TAFDwrKq/QCcprvE+FI3FvZ/zAzMu306NAk
iceimg4mp0U1bAmSwrf7BlfhaoTBjycmAualQzVKJIcRQcJp4iOyt58O+H8S9SAtcwaC0r6Cmd7Q
UsePbPPiyQbKa1+sTht3lwKvEygwKoa7FI+1j0uqbc6bL7R8sWUoDeAcObUC4R8jSg1cD8C2CO75
qmuKbPdWniVuYRuOkoMNzJnFKIL/yU3B/CCxkne3mJIgPYT3bo4DiXJxNEv6VrNW/4Y0/VV24ZSE
BUs+hKKcqf56A7KQSST7yn/d7Fuog824u3wsxcYmSJkXReGawR76Pd/gnjELXIN3tH85IXUw59Mm
jLz9Diy66ueExKsAyMlvlKz0njE0Y3BY0MxBtghSJ0GxbRu5asLXGG4pXbBf0hg/ktINGlk5mq/1
P/qWdCTVX8lzXnuzjuhBGcrNrX/yrcCXswbEvZr+bqkiYa+/tnZqSnp174SdPjrVYdFmwdTfRFqw
kc9Ex+6+jil8bg61h+EEZ7HG0BGeD6Yk8kf4RStFXsnPaPXfBU4udRmRJimS9nIkT/qiL7kBo32h
YxvoC7akv/61aNu9AzX4dODMdLCEDYAwisH5fprotdxsocFzn92DmU9YRWQktSDA5MPyNe+IhbJH
BMo4mK8/Dor+BV0jUF63rs5yZwnUP7p76ZWj+t27VAWDznnQzgGdxaNjt45Xuzff+PL6wy8wPNfk
lqyJUemkgHCYCvPsE7pKpfkYtQ96t/g6HyALoaV5EWpB+lbtjrFsIbmFjpT+Mi0JGRmsGxj1Lzsb
wie9w5dKul0Br2uEjF8eVVWvMZNr2rkHsWg40EUfY2PJE7Ge24J9K7ZxekkQ1AGaZCLIPrAP+bJB
BFdH3Fga+1sUo44QqYDgZv8CqHt1ZhIpjJ97VQf0fU4DDINsdVG58/HH8vptMVNpMJ5+iGeoR90a
blgfhJ6ozNnTwys30vniCYipCoDLArkWj4vszw7oAybHrotrp41tJ8qnd0a+4o70b4OdfjcypKLI
rAaoDg+twIGdmEy4lsHaCXby5HYiBaTnSVRg1z92cQO+cMGn5302QKAwTC2EJRTI5K+BCGrP9TI6
0IeHfLidn4FTLIVbYbntu2RY7fNAiU2PkYHDuijaVe5vMylNRjAu1MVtuURB7M/Rd6p26Nv3BnZH
Q3rvAgXz/dEfgndjXZ0l8iv3fgJNaeh3XQqXeGkR18DGo2k5PhiBSIMcBJhGMTdlxkXs/R02o2g6
7Uz/H7SahUc78T9tqIAwGVcgv5/OcrWrYvULE0ZO2jORYXPMMiKzTn6gXeFwpCQTvmpSdpCNsCNq
JXqpbyVv5cFLxPQ4YsFxIgHcxbPGGI4uomvDDuj9Ajw0TUvUOrqiao+a84rd49Gz3pjyt8nOyb3b
kqkNUA1EwIMqT69MSBGmzR4T/EScg8PODL4JGGQBFVY2JArIp2JmmqeQF+SfQx49YlV1T4ufwpQ0
49HKCmaQp5Xk7XmoynTLysob3RgIFV9M/sMfaQn86Oqn0HrHw2exk+CfFqueC0FV35xNsWlIWgCo
nxmnCRat6J+sAzqPLnSvjB2zwuS9G7RPT+C2Ff0K2oU5yFhp7XXefGHEJApBA0Cj33Cs3WQCoFD9
UWzPnHlsPS7cqYfozrXOyzUHW4mCicB+gR6L83hAzFeXbht3QhdqS/nsrRQCpgjbedsudhl00eSI
7Agx4pbIQ2OC6MoQn30U0b50cxuC1njAYWRJvdEVqXzoeFOfvg8wm6WwPajexoYtU3fo4XbXW5wp
bAmGwBcrEKeYQ5RUB7aEFfolvxUx6m42QvpTPt0/3sgkj8lOEifgnwfsUhTHdbnFtuPtH+CQGdGd
5iyGJ1xu/lJPgSd5qMDwYXT5AjLe6i9+THDQtvINBHbUUpXeLWImTXUnV/mgPxvUJ4AGEkhQrWs9
FCIVCMV9S2RfnK7Dc9HAQx9N4WMXWa3jKFFTk/1+40LVe9u3qkXWCcAaLQWVxaR0KJvEPgYX+RfM
+n3I6AhQcDdIqEplwpqA21Ewmum54srFFXJlEYlP0oEkJOqPlG9dn6tKTMg7R3lzRolR8RL93eVW
Yxpjed24aj8pLR2ZsXuk4PfXZ9I7EYb07Cb0MTxSXeOjJzrVZDXHfE+r12Of/Cb//MpzZr2kLiou
+kTq2bvZG47YnjJ65wjouinFNxEdchexJ8OPUsYrmxTdxcr+UKIGxnY0mTA9NNtgRUOTgzL+ZgqT
cJxy0DlkWdznqTQnVrj9tRLjAPtGsjZkzTwbR6Xkd9g8Q2jfRKlka81p4VvUUWcPEhliy0zN1Ehz
zJGPJrYFs0ZXnTZZnroRfBqjToRwUKixEAzfTO/45js9dtAtrhX0afV20/OAeZJx/Jd2ydJKlwra
BNsezPodMgESfU++yJrQ7yijklZNqeThs/IJJBHE2T4dMleTX0PMGEftCRkGhDjCXlFZ5dh+u4Me
GF/51NnD6bFZX9DnopKn2FynHRlZ1dfpqFHEtPcKgNu8hzkW9i0xP7//OgJl2QtiDzYIQ1m+7I9T
BwUxHHCqZgWCeRe5CMYOuM8u+PMaquz7jFLO4uqgSqGozNZyGNuOVilPpo7lc5zpKG/lDP82QhqU
l3ijBS6jpLsQVjUZM8DODgmGeDh6S9Yd9mzMAO1H+TNtb79rGUdG8QdfJKdAPVKKi5NA3bmDR7QV
dszQHOfWf5Pnd7cwXgwW0rqQ9CXmOzmrzCckjOncNvxmfbPeipRVUSyso0gB9S1ogxBh0rAXpA6R
56onamjmAbfqYdGgns0Kie3o3QiRuhNxMFUk26QBhGqWpgE8RVwQT3CmAIDBIYSDyScDIPu4ZNIG
zVHZMo2Lf7F0RQBl67NttrS7jgic7P/rdEqfGai8nASrXqH0VUOWt1pLpcoYJa2lBt7PtShyQFIO
o2w8bjL2vJk4uazmf1XCk/Doi916LSQD3yaeyEPsk2xvOD8Yu/F16O33VR2dplCoVGCx9GpwZhVe
+j37NGwNgeIsKjugbm4aq0EevNuwR3MwSMvN0AHTTx4wWMK0fgrIxFBdwl7QswGiP64z2nhKhvQy
VCzX+VKtnkmWrICycECFXw4WOhcQFEL+LZMvGxmefZACwx3EkQAza2Q/wK5jsjNfza9I4BFyynLk
9a/webn6XYvGgZOBXBrsswmVoJbfEoC7Ad9Ey4hg0KOVkD2X+rPLc05Hv2i3dnCRAfYaZil8kXdC
rkxd1WLMc+N5r474L3LudOrCRgAxmpOKNDmrERSrzzYM/QbhUdSVBREDs05udJQ7Vqwgt+jtU+La
8FOowcTtYMd31bClDlX0HEDhp8rbftrcfqxORKVh0wbdWE7QUFrYpQhQSTOyPXSQ9LDLiaEU7m+P
oh78FTUfyLL6hRQXlPUD6cJdXvHQwRdoOZEhXPbcoCCZsKVd/2vtdHYdx6wOThNB/vQpV9j4JipR
WX7PN/fbWZjT1VZg+f7WnR+3mI+erFnJQhcAvodYEgxfIjw2UxY9PsBqTsSWdxucUL8Jl5RZQkK9
mJLC98J0laL46SSiaF5GAl9xzznOjQPxbtqruO5Vkr8iDD/1emkHXTXFaWm3uzPrW335M/Q9Ce/q
JeMrj2MexMBlhFIK4p470ysC8qo/tBZ69BwXLHKlAYdrm5Xv4ltKelkpZlPzgNng6L4zvYcnPo6P
V8jC1831/O05l7BCr6MWis4IHlZycFdSk8Pw8w51g2H1FkFYAGJk11PfeKD0lUMvuK2na1k3zxYB
3MCoMING5nKUs1YggGSd7oaAtaD8xPBPCmnMxWJn5n7wWD1nYoy6/HhJQSGBe5bZjsKHW/8NwCbG
1Fl3w8igdiAz4SIRmpsSGQKGjd7FC4rZrcXEtyViCRkvnJdabHwBIAW7E1S/4OzaUfdf2WdFHPC0
iGwdKwXsWyk/s02u9l3dlLayJ7Axqg8z07NG5HuU+Gsajp1AskvNih1tPfoXCxNvDvYvT3hu051W
9RiADezeAruCAszMRt8wOa9wgt0dAEQsCF2A4K3rdTYUDtuWKLvPPOAS32EDMV1Kma5drZLVdB8F
5JouNXdmGmjYuCZThqewE37iQw0EUuZ1M+IEQIwYwIQTJ9naEphyCN17rsJ2QGUyseYoNWq9hHqG
bwUDErgpADBWZ7avADirQdnWaZ6xp3Z7AyPOxKfdwtXO9aLeoL6/KNE+Xc1ZgGCXWyecr3yWfh7w
whELckjW0xcxIz+OWbvQhmxE7vqXYSDyv5YL/kyC5tvrXsqKzbRNB8tDUUnYMz77auvF7JJjueq4
unSjZ8gdP7jCvM3hq5z2oz0bzOJv2W3+1obWiIVGoriIWOiSZ2nnDj///T3A3owKxaqTXgS19FGJ
ostoRRQ3HHuYRp8g01+4T5PPsEXzQfpVCsQKmb2mTJcNp26/wRtRuaVBsYd1G+20UQGHNM8ho59x
HaaDCJ5yVE8SGlj1+Q564zwkqaM9Dah4ZCj+JjR5KC5X5tp+65vUxfBEattsmD1iN4ET/KvN7gHo
Yj6pkVSW7P34B50eDg8ZLVnEAOKo3rTIFHPqlas1JkYwffoBOQ8bb32e7Q1JSP79ybnaLFk6u1ip
jah0zYyse4uilSm/QUfe7EO6fuwvqca9eeRgKJUcyFUKO6CEXsJcy1P0KhBt21UTdkWsjXCJ/iVc
iqo7MHDXWmht27xYBbrGhcrD9uIXFTJUiC2a9SuPP9tNWy9Wi9uk1bEkt3troCHm+azP4fD+Hl6H
n6n/jn5dYrU+CNPxgJkVpsA8s9RObFG/2Sgn5QmU1J8u5f+/bS8SbYVXeKpYgOxP25K1y87RU0b7
GOj8HHyZ4uoWl/qiRxtYXz+PVmCJtvh2ZJfLcbkZv6Jo1N1kxly2RUT/sOyMLcG59xtXrPchFqxg
1DpHJ0r/2N6wvk7sOQd1Db/pili8j+KJ8YvosWG4B9hGkB/fNBY6CvDPwlDThfKYCYgwP0ruO4Q6
+BaI4vOuFTWp0l6WnLjBUtyjdsyOIV+bahhn1B4bPeJLflhwmL+mGsNcU07lb4oXfNKKFcRfm4Vk
wDVZ4Kd6ELVjtjbGwHOhACpoysCKxskvpxpmzB0qL+Z4phjjRz8Fhty8p2CTc10juclMyLL4VuJg
ifZePdWo78BzZkpenS8ONCAzLhNMrV99riB30yfDG46b+v1MHZNgDcR+7n/Lh0ZejCl3iTlIoPNq
NK0u8AcLbsQFU+56OcpGpkT3KZHh6icXdhOK1JHrXwqyti5w3gcoc/ecapgaMN5Tn/HIJ1eBswCV
gUtgrLgxMswGmFdrpVYadgxKkcnBCM47HEpMnOuX7ILMNC8ce/X/pI3rH0B2kbynIWmwKk1I1+kp
/sZU6b2eIdJRYP4B6InVTOqcG3XUNH9KXnFINnPOh4NvFmCl4IukhxVtsik/Z6kM8lzzXoB2d5Rd
qSZ5lypSkM1Pco5aflhZgv9wEFjD+PP06F3okEpL5E9QLi9zI/BwlMd6QhwenR2Huw0VqXKVOg0Q
g9cAkUHL5XdGx3Pl//eRcl8f9A6ye62mtorvFCTcAo7I6Xdnzse7jCMPn+Eo9OoyXJzi7nrXLSW+
4PAcKrmw1KpOmJTr2n/SYXJDy9byLU0TrewT7awfPyS3EVG/jgwwIbxT10p2PQw7PIFi8SoWTVsz
yJrB5Dx6awkTw0NYpRsHeaNWhVWM+gszGrFS3EqQ+oAQGpvtxck6DJfZRxF7OVfIwHCjI9RHhpos
qOMefRmSFi/SuR3HoOfW/pQ25WKjSOq5DIXFOmIq6qgeauF3V4661YRUuW44QzTBzi5jW28UHIx5
eF/7eN2dS2zxNeXbn5cKvmoKmmjxIyv4YS/XH0fSWEcffxNKUSVetPULCTHsDRyXRxBsD6VwR/p+
iVn3VMCo4wsRN0x8w86b0IwFxjDdwQBxoL0Gya5/2EIg7MlzaEqeQJ+/pPcbm+FuwklYc2iQJx/M
JO+TsQFIeYfVvfWcosC7BLsuZ6GJERU0j6pdEEldQ/DulOybgf8qZzRvxrEzJ1x5zo3tK14tvcTE
gkMPAO+Y5r3ND8q8xwafn/mb8XTvURA6zqdT/MpnzSQkIGABKqUbX5XgCwjwokAjucFWoY1tghWV
wuOGvUd4VjQhaUdB7hpUWm2OKGvt3piRGCI+L04CPVTX4Q09YM7G2w1paJ+15LQb3NZKvaKiLyQd
64fOWnJ5S8nCdMmeTOefbMxywzWJG4av/f4HRxMWSUoCBPn4eQ7rzKfU6PZyCBxMxb6OK56K2g0W
39bIcLVubrL47PsQleHDXmSSPohmdVa0ncUrf3WwT4LdqwYPLARwyb39ZM9ngqGDOwPmVgqZVOrr
Ybk4ExzIyiytPhWRZ3NAPlxBiuTHBxpISvW1TE8ICDUXB4kjGeDSrANRGZ0XalobTpVisHkdoNJY
E4EbpQ+LOPpKjgQZNmVd7J1Cxh303FpDaVFpCaWNxSCGfV7JmSPj+RuokyrVDwRXf+zhGgiqw5vl
CSZiae5+zKvtcWNLaIQ5VCJLHxPGhzGsxhkU7TShRl6HYqRPwxO+YvV+gBq/+90HpS42SQzaTt0f
NFNAHcTSFukcdBJvDlFESDNDEgA8zfSZYQEiuWRmZkxkwpXNbfGTUzuJcsLz/1D5vxDKYuuXF4sd
Os7yNB4w+ZTecUXMv2tMfWL5YPoh2n5Lk56kV+jLlQmIu2kIT2vZTPC53JlZsEmuk0RlclApCgT1
Lz66EvBcPybti0Z37ARLhCvk5ts9W0pbzSKTknXW+yihZi32B4b6qrtR8STSxGNBpn3EtubUQp3o
AymnKJOckJcL+DZqs6Sh6mCjpWkMaC1X5OmcpWeVqxfPk4dzKmm+YxXk+tCsXrJOoKrV61153TSq
5fYVtKy2VhBl8VDg7UkZ/uiv/y60c1FwCcRziRQttQdqXTm7Mkv1vPDOzXMV+hh2EulD9sV2JjIB
m+NoOjRGGQm7ZQQp+ojjI5rgTwbNDKNDILkc0+wCLrdkNqFDzfJEpDSkIOYyNBaTXjcR1qOEZ+mt
EGM8L3ISsQMC5jQ8dHsd/fWu13SnBLyUurI7U3iO6EEtqJpbnb/PY/mHtUKAIz1C32pzqHuGH0jj
WzXsRd0I8yQPjWhZBVJmGaAxo6F/6vNQ2mjGe/550l8oSKrN63k4bnN40lSS5NlKAHzAUb139tVf
DsS5TWibz+qDfnHnNcdlvjIMH59l+q5YA+NF+7lMElUjEEdINFD6mgulEIT8nYyRj/UQxFBvoKHR
z0XemFQQ19+LGkoDMIheQQtG7ozbNXuU+6puvFWCbmYoZH+4UL7XXxxstX/5z/hDr5QW8FdjDmJU
dtPqP8dCCl74WB3PZapsnihb27J/zIbKnBCK1y39EP9beKsK0/XDKDVu12UhDdl2WisLFcZ4dcrt
FF/0t9/EbJ6NB7CphNZI4sCDD4kZbuyOVbh2YzL0tF8Rpj6A6R9LJo8MwopnCPNYzuk5z7I8DTTy
ufqpDy5lVrPkjWrl7FaDIFWA39o8R35Re6DIhamt/ARGs96B4/VrBoaKI/TOVXdpi0qkECtDRruI
zr7p/c5QfWWzbbMsZtZ0uhj61kilxelpFEKmmxGbHhwrHAWYGEFhr9iSIj87d8pY4iKyp7nUS2ZY
EDUSd6euIBohV8C/hTgcWeokEaM6sok6jNchpV12Zxk4NaSDS291wAnSkD9aH/SLNN+N311cUQAq
+vRvl6OdNMyyBRWPsK7qWd89TokIscAkkQt89KO6ERxbXfGvRo4Qn+ZYAkddXAN0yzBnaxe3I5PU
QfHUtBExDMYaIfwKH8FcgWlnFKB4aaq5dKehwCXYAhYSl8STYmYyW9NWQ6R8uHK/iJrcryLgCCDV
a/yS5hp2CJPTvKUR/UBj5XFB7Hs5sijmJKlkW+NQsAK3oyjcm7I8CV5qmy1bovtkylmoyU+OtLYC
nlmcmwnsvg5peVCsHd77+GhbB8V1nYXKnsngcpydiQf8cAXRdThHZ4GHYz2QHSwJEG9xAssDF72S
tosN5+wUamG77TEEZfd5acKR+UmCnkoAszOO5L+G3CcaOeDh1jfHIRWUQhosapoBfZlNxCv3JGkE
Lwtzn6TzSBOqqw1K8Kzh94pbb37ekklk9Q3Gb0g5PRV/lDeoba2ziUewUsVVZdfv0KLd+jUQyaFB
dT0168ejQwK5N39Zf1UqXOz+X4vTsLWe2x4psMxoRYj3Z32FOcPSca8PCEyQT5krU0p1IbbCQXJM
YelOhB0ZQTNbkjme9zUexduGDalCjHEc1Ofv+EszIQLm6kvRMeCYkrELUDCN+o7V71JfXIR2ns15
iEbN76SehTu6qTyTwVWbRjpcDPNQiqffPJ3XZSdev39eN942YGB88zfsAkzkZ1/P4dJ4n02otfDB
im8ZWsLF+pFty0pJ3P+IEqzWiP91KTfnZc8N3tdpIJcjUGeNYlrsKkr7aq06hzEFphfFqcQT6wgU
DLYQzsBDyqUyJLljPeKicdOz9LcIOHt3gaTfflzHHRHdB0M2RLLr7UhCrYi/4eEdECh1ycVLdgWM
vcheMMHV5+u9GGNXNNazKvS5BY39lm7lhKPlQkphgbwZnzA6drtdXRMUd1sjgj8wxm1+JlE8eKmL
sc7CZbF9fH8rmo5PpawnOiK5cEw8Lsyw6XrdLJIaQgKw1adz5JROgGQcxRMBdWMnwO6hp2kMu0Ib
N3/xtSMKc2JJPNFiVli5IMy9vmcqDaBOcSfYyOdgDAkIKdQLwdPzfbMTiIjC8KCnrzo2zTjZeqPe
xt6RZpghQOS8tnoLen6qdYKdWtlY84dvUvEaeudjGIvHing1GagOn8tQcvdBcWadsaLkTFOoS4Mv
/2kk5br9fpzH+E8568Nz9uVVPvVBHLmNoQHYO1BDsO2UzXDcQ7DI8Mf+L6IHqsnusurI2pmFitp4
NAgFDjE/oKMAG/gNBAhO7dSimL8dL8LEi2hmgMYYspIVH4WHgifR9n0SiHxEAoSrqN4WAmlawc1R
S1PrwjcOSqZs4l0wCAEoYKgHhU4CO1mEQfpAdj8YDK1Nc/Rd1vrvNbVSZ7bvJ30AJZdC4VKWlp53
nfQnNSb9oXY7VocBpf63iJqovvO+p/wdkR4iY3cMXStvSWhM1AeEJhzkNZ3yEhFnKkBkyc4ErJdm
R5cG7zBuZOOmPJ7c+Bx4n6e0sG2uLLwwm4knjiM7AmecWBmlobtLhtjVART3hK0ucyUUiEKclOSm
pZLA/YAS0pA4Q73nrjn8Dq8u4kXKW10A6CmSXEfiVEHn6aSkxQJFRrowA/yM0VFV/jXAbRjMlRya
2PM1M4KWy3U675k1Eut03uTpJN77IxIS9hC/DdZ35kmxJaEDHVJKSBMzjByx+popbILN9oXDKve2
RHhgsyLx2m7NPVLaLrnCS+r3FCLuU0vfYF2zO+r4+DGy8Dj737eGn3EQ64d7RtEqglTBmxGg7fMJ
ZsLHoazP3UfjiNWQHjPHcRH7pMapRWnYxc0RMkECQpscNQ1gbgTxRLSUpLgG267R17cYxjXBMpw0
ZsWbOkbHT+G1lrmuHfsjoq4yi+fkm7TMx0yKYQ4LS8Xx5nPdaBtCskh/2bgzkyv3k+GsSriagBO/
luEFKltd8nFo+quX5OAMmmisV4JDhHi/ABQUKR8phHgJbAAdX8vtjikodAXdTwJ1+BNgEQaT29Bv
zEpkuQ7ZiJJAOGxypcSbEJh9zUsnIp8VCd6tE3CeTDY=
`protect end_protected
