`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11824)
`protect data_block
dcJu1fnBMt4+zoJv73f66AxObnlVujYlSI67EPWhTL9sZCfdTJuKbIq7SQ/RCZpOLOLXWrc8T9hf
D7CEWl2m4IJ+90JzVLyTUfpwmahUga2ftwzYZQGJuovezty97TfWqpCUeAyNNWIf6tIoGbCEWq9Q
r++JgVutQTRlGaWpxX4reKossvZdYMblB1cuc59JfzyZPRYpor3KM2xnF1c0oF+4O22bBc2hAdPD
oqrXajFmad43TtjuM5hjrkqJeh04qf/m904hhdwsPCBgCIbMEjOgy7JFoFtlJRQEeNy+ltPRKi0P
Siqmc/p2cVmtHGxKiz/wpw1vFWX8D4YzDO4eaYY3D+Z2UlZTpZ3BSDyb5Wi8AkhsGWgRIay7Wb6j
9DcKsyeqgCpXol6pw0/M249fo9GJI3Aq13MvYFh2a8d9nCNQ2wT3KFT65Kvp8eMMDB42rX+pcFm8
QfxhJlsPhCDtus/vEVN5FFakMtMtPic9Kmih+0pHk8r+sV9wozpAeEyaN+HmglQuxJbX0KipSkgr
/QcvcQn3P40gJJ+aTw3L2JjZr4CoFJeMSPhTbi6fkPxzQrCh0Yf3gMD7jb0mmHe+IqL4Imsk68xB
Uux1h2TZ27mf0pm5MnZ29bPW19R1Hb42mMcf+BeRtAYdzOFB4H1QcnPAw3Uq6i1SA4ONMF81PMN1
k/oid1q0MEEj/kXs4Al01eVdLU6SL+uyeAXqUyxkVTXX+ptTTTANA84LNGVp/DzX+CVKQsxRp5JY
XLTtLFWKzzvm4hmkwYIMFx72JpuEoEZIEozhuDAwS9LXhy2xdcqZHUD/oujK9FdZ9RTB0BkNQIm2
Kj936NCLSFZAv8js6QoP6NBg1aD62d3JbvgM4X/g6Af1O2YCKGkzDRLZAiPm2KAhCOxQ5y7+5Mcq
zLSvXzNJ4gDwLsHttJYPQKkHiQi7bVbMEj9FJaeLkcNjgozsyWNrhALhJSHswuv68qaXo+9UokQI
liyMwTYwRsUMVZ9Rrm7xnuKNijphiyCbYexQOVTKmQHw0DIT5JlvWGOG6e6l4xmxlJTCtiOuR4M0
dQY7mvs1xi1848Ok47Fy/4Qg3+FHd+fDNzxRGe6n0H+5Q1YDa5DEDyDfC1xSImQST97ZxGSs5chB
9TOk66MEEVMOzAHKCVjrWPNuSbxjjiLMwYVTHGAwxZEJE7M7DoEMRCiHKXFYy4wAhFR/9L9Gsydm
X18sgdr9r9Fa90GUW1di77ryZpSUCQtYt4JAa31Rwf3asIMO1F/sCg6Ck0PHywo62fnzhSA/wM75
eZLPV3IiszOcc519JGJ8IaET9h0mSPoGtLhIXTa58H1XsLHEomwZq1SKHk3vZZTIiYHVioceKtdn
F0yv3T+bNSv23/0MK1uR0HZHSHT7A7/4a3QVJJltvywO7shw0Opn/+441XqmB1VFrv7J1z+xEy2h
QvF5z+8955ykhVidaYxts88Pfcvc4oIk/3pBLYWzrFH5/BNVpVq+Q9ll7hYkzLyCRcTLGdOtSdlr
rDhUPS6shYKVJ8aSGHSD+0+D794L4L2P6fvkO281WB61aglAY8HUSnjdiRklMHOoYm4RDVzhFNK7
CHq30LfeXgVtVbjGG06PAOaRoMqwiFZ5esiNoNIbCDLkyZpIIe8pq2VYlaGmg7zwwB+2UIvLLHBA
mWvytH0zwiH+ergIM+wAZ7gCquTWfzouStH7Bvvw+ay1mV46TGJu4fUR6d9r/yCOV8l6aodpt5cX
k2UYm9VzOX6Yr033Cr7jZviiJZoVlxCtSNHkEcu0j0RHeHWMT+oOkmu4xXwQqsvsjqbFwVpYFxbw
cyK7KQdwco4mByku0lMXKAMZNkvsF/5l4YU+wz2xU/79LdCfpGE1SaGzaN27u+QO75zNQW4IPiZC
3KrlIFQGeZZ5ABClqK9F0dmFo814xgvJ1ViD5RqZiKTE6E2AZJVVgzyunpCTrH0Gt+oJncDKpxHJ
W2YVqQIVkLoS47h9GlLjXQ7rsEfj3S0tFeZZKnxaesYc1NGu0DPj17cuv/gtiDOyRhM7HyYLDgRs
3HIbMI7afpG1krM1QqIkpIr3rDdg4YS0093SMf+5EYvB5oPJASyzdK02fLdGkOZyTd+ox1IHWWZ3
SJmCwzR3BZjkwK8MYynJu/hVLM2jn3jsXmrccSVyS4I0bUU41fK4+uXbdZJPM7GVTjbvmfHHKohc
SSJ2J6eExZ82gUU8QEc4SI6lGeE/gz4HKqo84k3Bau6E6SEoZdnzSzsVLcuovjwpuHFcTJUu+BBx
7nBXiUbpum2MghYxbnK7VcqEa+5FEBg6KzUZ+GOxiWbXG/Jz2g63jVLCyvRPwW01NS7nFic4jTIo
BXV3fRGq7UFIYaa9Q45eJFI2vq9JjsZuCBn8lp1c4PsDK4r8ldxTnZ6nne1K/z/As6xOpBWBUiAl
aT3+q9Jug4JZD74m+ZbNRHqlL8TXTzVXzIFz/veQWBEzHe9nsWBXlvBikA2VQYrBl3dytsmtrfY2
9acTCn4916/ZiMKacyTmOaqwqkwRQb/Utl5Sv4bIs+HzIfrKZHaCOFc3k2NyE6p1v4qak2EO6K61
d5WKKsrMgWA/COAn1vP5MXzHQ5Bqn2KUWTytElRFB9Y9Y7+ypiFhPXV1gM/C/Owg2OMWYQXLHLH2
nmwCi46vDkppYyAxwaNkGPy9SF33styW3VUKiyMJ9NpsA+pSe1vu5NmzSXNZmCpuitN4blaqiAbs
XwYpvd0DjjJtngASsk3kBQkJhOsnoVzs8zGqF7zkU/hcNLgXDo2h3RuaAYtuTaoRfW+wxOHwoNCI
DUKESwx4n0n881TWPf0DAn3t4vEWVwyydiyKrEr5LTLx3UWSXGQT/ByepYiWd2BajJxJQLPMWQKL
/o6zYpHQXPsR0fZA84NfrHGEGrDWjhkBOyxZWWye3eVNyeXsdhinDsSffeH9VBrwY3LlZKd5K/V5
ESJgllkbA6Id7CAeg+5GMpzFk5yuJW68qCb4TogmEmI0N9c3pQkh9TRHZZ01wKFTlvvMMaUeYdSX
TgWWfcp5l21vKrjR2NoeAYaybR7nnPAbvmv7ODTQ5GPTddZR0Pj2ixwcEz45pNYgKZAFzuRGhHvV
+d6dQU5kXfp7kvicu096EaZ977PJSx8uqbIhtP4geEk127JxZ0dOjEARZ6l4quZMJarVJi9SizLk
4uHU+iBRq7lsCLonvScvjGQOQPDNf/oFJAwIlqaBXUIJDFWwT+KMfOcjh26CfAWC6PwvrXAJSRhH
HTReNGLKI6z+z/OEeGKJPAX85G5E8GMSDAWStnQkmrR/ZchS9tXoEXQYv2j9yXGhJxK+TA4WhVKZ
s3EQHsx1A9dgJNG8v6uEUX8pBnOrh0V0rg3mWarZD6S8Vr8YSEagqQTkYOrUCS/MENcUar9iWI49
wDwqstGti0P3Qd6yKvbumKejGcI+1Z9MVQ9uVuT9929I5+134tLPh3OhgCY6qTdToKywEBkBVsPn
3dDL00rBdyxOK26qkvRk0T71IoCVrpcrXjQuCxeFywpV0lXZylgKusAgE2cpgQjeM1BfHBz9VIcJ
JOSCSnEQEedWrCMX1qttqb7ms53K73aBbI7jEl4KK+70pkQFlaiRWZqEksZDHwLcyWFN4NJczE4X
Bqhgf/WRUF2B8CNqriRWnIxwwRoHW12B5sj+BvZeEk1ABBvL0rcTsFkfXor+GHCi0DY6HdFsv//+
vcV7atk3fvHzlEOCpYk3yD7PE3s7z0tvC9qLr+igjaZLjogv8MZDzx/R5d0vvI8/ABhlZOz/EKB/
kCZ3imae5wGA9TD4GX8THErP+Yga5lRuxo2cDnRrBpFZ1N6EgT0seSYhQg1eH3UHDBuWB41+uj03
crUbZd3PraVHKT5pcviRhJTykrlVSluwNmtYKo/x1KoQblYYZNoE6uTOzuV87lOXOzZE4gN4MDHh
gaXCPeHkK3TPbWeRG+Z6eyA6tKQlCzwrEoAqkGwmrw2psIz6PmLRA26QlElnxwUyP/i2SB18t8Ce
+AHMnkgHS5MjpOG4j//hETfSseZAhlbnEgxigAu0sKUczkoXXWyv9t/yo33uRSBMj7Zw4YW9nsaA
rQYbvySk1hDpFOFxVQnmsfwOgq9FaSOANFURIfgTuu5EypFbYxEkOTc122z3rBalBvQp30cEMgw6
SFhawYIhhkHK9rlorZNsqw8weJHDHuDVEctcmarUCkSTcRUmlBh18cW/wy2FNlgxKI3lCWB6/TXF
oIa7BYxJvxRG3y5+/a7bhRdiypZ646luTmTKmcT/eGpqcfEbklmTbNxK3VCUbpkWIVOkyYuJ87qt
/QvK/VYSBMmGHec6HLoCAK4zTr4xNc6/7hN7w6VQy6SoEquoyYV55jQXAfGp4R9XqzmKp9DeBxFI
f44Ig9UJN94DMW4NEdQGZmIXoDsviX7BGBpxn137LTnl63vxPAIRVsl2coPUrf7nXTFXlcFETxJ5
UfR8Thh22uKdgxufmM3IuZV/Ulwu0/ymwUH5H9xLAt/sULwEC9Bs3DsBUf8iK0vS1VqNAGujNeb4
1nNKZ87BkvpZaC/2abPEKn08DIAz7zIJeDSgSnDT83ouLcgtQkQk3HzDF5EiadYKYyEOQwlsAAxr
+T3kxMGRznI7u4SsZG+OroLfZgQvz+/cR6fK4HWcCBL0wyyBd96Lcu2n4erfJllwd5+P5EGrL080
QJOqXbAn15YARUQ4K1Kd5ZVerwku80cEOQ7c7F+zW5X4Y0PmZlpdvB/p456xtI2/O6fWEN8m5aXO
zsCqkPYHASIgFaqKJLNfC0k8kpQ/qtytlDfyMfFRCmgkRoa/capeFYFSFsU/syDTcjZVktD7yP1K
/DGbnnFqDboALb3LvcMu42Pxhg506FqVTwVEsd63mI4yXpkg6GVdksIPW5evbQ7OMRq0dXYPrOTX
/2fHkjbge1ibT+BxEJek/4mFQOjjlYSwIwso5LlUQulcgMAsbNab0rWG2IwycMN688ktDavsPFJS
0ZApVsCh/eKTPIYySYyGSxHVN1PNEEjevn2mCltizHQQDc6PqqbEQ5fSa8UdzBJ4/gErmOwwz0jS
+shusgO0WiAJ3J5HQyZv4+G18bTv1ZwIxanFIeBv2w/TQyDf0NvC9GcME3hYZ4KKjr9wORoCXGG4
dL5W4so9QdZOjGNeQDFCtkJ6KQPwzP3+spV4fn17cvriDKqwLrj3/+9yDRFw+h4s1O2zTvcNG2gX
Wme0aHZo4BSJDFJnX376e1qTBFGAFfX8KAonKFs3bXXbdUCYUKlEa8HHbDhiB70Sy4dzTqFB+mOF
NyN/+NbSIn7j3rfnS1uvqi6r//asDpYKL3aOfnS20I+O6+a8JoMG20I54Hr1R6IbSNx3d32z70c4
Vcl6NC+SH44AZLUAoCc6TudegOm0Gr4Z52KP0ERZS+TURNdZPP9Z/ffFM1k9H1KoEfMCj/L9q5xo
RV4yIl9zM//TZdL1JX0A4OOw3rrRbLMdAOPzm7lMv9oM9KhNic6T/WVhjwegOhV2l51nBd21Zz0F
SjICmkTVjfiRRSWQ1Sw8xtO8d+oclLb1ohgKdgROWF1DAs++hCa6VdTCzQGjvi2E+kppKnMtb0Y4
wZRxx4DmNZOba3TduhyANpcR8okiqMCTqDM0kiHAiYCLE5k/kAknqRTK9E6Cis8qwYflqtnAtGko
JTBikE3QuOGKgG0I7XJSYlRpoQ77fz2G+ITvxTq3wOCfcNBE+aKgAr4c6siZ72QPz1Jf+6E5Zfia
ej2bj4YaXAJ3J2/J9AHtxWkZ2xrKS8Dm2cIpaa3HtTOEfKtT1U+iGa+UxUK9E04o7NLLd7C92u97
N376c4iNrN707koI22GLo/mi438DI6DdawtbE9x1kDeBWO5xAJFunUrDjSQGuvzoZSJn/GCpmESA
ChCvHCC+pTJtZ6pRHR8YSGnEiONfWC1ajhbO9k5kHJk7oMpbwNviAECCR8t+iAzWTKIW/+yEi755
PB/QPIRuIBopPLkCly7rSGWtiQRWAZze5W+RDfvM1MGv+fsChn1KbE4qyXfF4+WfiiPjVP+03B6s
PnlGVgdJWekKKpqQC+SOUsgLP7BK0z64wikKipEr0CNvI7179pSnNRwcimAFB/IBiET7A7tP1G6X
CQQC/AI5zWl0mQJXBcxqcIKE9T9aUkw/y0sH8B/J6vNgVOi9GlpHVX7FPQ4CSPEC4ARzpOtUCQQL
2Dz9cJMnGZn4fYq3rssQBYJTv11PgYDSzAyASvz+rUZbWK/td4GWRRMEcY89llZ49x7zOBU1WWLr
/7UQIfJeZjYxwedrCjf77j7Iqtq+rWVksBoujmr0isNmO5BZ0lcj1IYC3jiFtWCXqcrcCYLMM7ev
Jl3FIgm+zZ25WRPBS3KwHxuH2zDFadS5bzgIvQz9a1oz1/FjnZj51+a2C0Z/3MqZTaYd85KRZZN5
DMUuyxOo7j3OZBEVcZj+x0s1oSqT5/2e97TflKz6q/jqAHxKoFo7ufuOZwO6/avO1fqprow7Afs2
KgT5kyEpNc2rRlfiTjOzWWxKoSMEskWQelBW4i8KlElOnayyowEgG6fymTMQEU9/R5uQx/NVLPRS
l+rvINHIZfWi39IfRs+vLnFqQa80Pte2wnxF7VA6hENnntuEaPCsGwRL1gtaMPTplj3JK0Dv2wR1
UL23qgk2C2Xs/kym7e1cSn0Ao0wP63nd483QBDPoxoNknSg+ZILIgKDbriALrGfdUJn5Vb3J+6S3
+4wPARR3PpJ3DnlU+IZr6U3TOAMT6O6ImqQclFDfpUAXtKyTsYSGl55MNsJWh+RhMpUrvSblpvZ/
pdGAo1xFfWeL5RK7zwWd9RdG5Mcm/Rrd/bzDV2xCW8OQdG3+QxUTNoIopHRCcATLsh8s75K2T0lP
TT4aoG/JcG9ITj8wYUi0zKz5Nlx+/Ibvui5cHbf4EXwoUCdDFjCDlCqe2qO0LgjBeM77/0fpAMqz
rzvPFNkhS/NZw/hnEJFlbkwLvwcLQwbpkhjPU9iPT/1WVDe2GS8YKRFR3fyM3v4Ir5xsKt57n+m7
32v4CChsEGw0A9rNfDrg2dgpPv+ApSEz+1ccV1LhXAtZNOczAoNIpvzP6YcZO5bVqJc43NPHJKq5
rOFUyTfNm4NaZW6O7hKgXRVr4q3k6fjnzsVmsZ+tLEdQy9t1JkbFZkjVGrqR1QDDAfy8EFphXn6b
yrrYMHRXKgCMVlbWSPuNRhVkYR6RqpgvTW2LaLGDMmGdMPXBXohKfEWhOaWD9FnDCGraVO6KlPGA
MY+NbFCr0Lb5jB2FQ8IWGLTHC1RoGEH5K6BnaqLLfir4wp6RWeSADf3cjoejePDp+tuk8vnZawhM
WQRFY59sYcS1r1VMN7LHwe2VzkG7uKOtzLX14sEoeAjO8qizRTjKCWe8TgTGUcuVCIwykHhCQf+c
ejGvC3H+1qI3h5ALalTCsQ7vId7qulHY5+R3DC4MA8+5d8o23CrV+GJZuE5Qa4eTHPw4nOgL6ITy
+rfwB1wKcBppKsM8k7hhx8yCzg6T2+LULlehY71fwDl0utXyqpXfJpRvxkYs5CVIQ6AVYHnJczIe
uMLK1bkGeP0x3J2jdYPer/cKmckT03ttEFrc8/pXcmIQf4/qGRtifznKPqUmPR8wS6EbhjtHA9Oe
Ec3e+jCxGP5BUiOM98oEVU+bKgvJQ3CJULXMgR+6yq07MXacckWzjJmwxTjdJEN2IFFjv24vgFts
K7cWfDlQU9elMweodbjvTzXH2VYeh3AFdlixAq9XOPNkfE95Nn8YOhkUQ7b8myrPWgojJgg77guh
d//u0OZVnncgvpTxaW19VBgX55CImmod+vXJKt45tY0y/mxfwPAIboMSu5ULO7ZH5wTdk/r7P3Oo
u3/u6bZ0vLd8q+LmRBvH8NsewcAAzKfK9C96Yu9YICA206h6UyVzcgkKu4E+zFmhiROiw+Z/uV7G
xGb/AnmqeimCbWksniFbxGpDyOY6Rfq1tihsyB4T+e733BLlVTmV1Q1XRFDOKAorsDKkQuXqOg5U
O9A3ZSN6/uYB8JFBC85mVk9PovTK9mvWLrS5nbKpBglegCfXWuXmMvWGImUdfmx5lBrkjkBwjiR1
Va9JM+Z8AiokHHq9YYuDC+BVt3fJ6SIGHOWnyXmID5oCcQ/DmHW46SgMeoRhZfzUUHoOwj2ANtSH
MYsFBrgfYS+kIn7aroIjl+DQmAhbPBJsb4CPmdTks/nwhZNBHonHoBZdUAbqjJ2aNnw2OQhaKFm2
GfR8S50TrpiDg3FQ5X7raP64JdBdbHH0WVYKuB1a7Xi5EpeHyQoBaaJJ4ug0SkC5TpnszCaVzIZA
gt2kcPyEX+Rf2i6MR0AEUqkLMjaIIe6nJYcXO5P45yQLqjWxypzjsqDsreGEuY+IRut8y9ZSV1RZ
4JPuWCouJ5E3vtQ4lg4zw/w2wmGp0ubPiNMWZD2/j8YScZbrhMcKFd1vf1BmbaNUmE8ljWIilm15
n/aGnFjYklkGPwGum6Q+YBkVeeMQvzjtF34Ftg7iU5p+4hFi/8Uzq/IDMH+FB3lTvpUG/XPV4AG8
kTORI+i9zgFYr6emPHEwJqO3+rlfTMrMP4GEZq+7RUgW8ckkvwDMuorqkRhrddQ7upbCSwp9LCB5
qebHSxcX8rkOE4J3C7l5RJBKijP0bUFiixpEu3hXDRZrYxp0ZkHK+QvqQ8oB+tvpJGOOR6G4YYD1
ffomC6Nn0C+ynsEYYuPSRIu3C5OM1VIlEvP41EmpXmkZFKCQoD0OMfeAMTmqUfsZfg4sVZfU11dT
yqqDt4aYqEECyY9EP2ljnuC507qgZSHA5WuntVpCiyFN6MX3y8eZl41tkFufuU8nH2Fibdh3y0rX
H1FpXsBlNib/BwU89/dYzCY7rxwDcXuuzfj196n/OE4iZcNCwUlU/jJ0dD2N4feSb9GUd/qJUOc0
SRhbQB4gqPfmly2cTb88HOsmu2pY2/U1tBXUStcbyyyFM5x4+uE9KtkDyZf8Ufdq1LVNLONC80Nc
zdBvJNf5SiANQeRvO8WbK2PvOgUZpcnIz2B7p1eYXWz7mlMAc7fM8L0xd0ehbR+sPbJ786aKNmB6
rosrW5vTTJDsKjKSC3c/FkwCuRrjPTPIvMeJICMJlo5PUDiIRS+L6shfj+EYRM/lqxTFKcJ/jZfc
TXC92Y8OucXCiPJLfJ05GxteA5BkThEFVNScQRNPXYgeEOedqH7CBByrjnO9fg4aeeORvogp9UQK
n4Bv8fVX5d6LkpPmETX3I8Ks1TypU5QWnA3/7tkMo/50bmpfLkGW2RRmvjrc0DfMLRRNpKGAKp/N
AaLRaDMSLBllcoYjg4kYJ1GEoySOEitjayqtPYCPX+8xm5PNilG27KoS8HjWz/5iVYLVJf8K5/F5
gfsK2MUV52IxCufqRpwRudUcPacSg67kNMnm3Cw2VYzYCmsWqz5jn713mdIcs6NzpAuseJgRrlTf
YudN2WOvhZxQxoWP/wIj66AT6wXY+beS8YppccsxLNIxi+zSYZA+NMtxWzdeLj0XwM8nQYBtfm9d
PCI+9/B6n6zpxfFoj63k4Xk0ejs7V7hPSIGW5G34Xj0vLOUcUvuz97z09X9bDx1ecINlbwI2wDLl
kYpT9XtGV3v/mNvWGaouJ6mxgivfnUoiSQ8WEqyDdjDaOjZsABtmuv2g6uf7jIQNyMeHDZF1irA9
PoiCQ7M7ujkwU/5jJZgv1+36cyDhiR/RQ3Xb8HWvwiNLzVrEhpJFEP/x/ucQc9sV/SCtc9qxngj6
A5qCNddZ0o0ZcezSfHIC2TOz9bfLRdkX213L8g90I/nlgKCY820eJ83jfF0vg86j8pqwQkHmoVSu
7436cPtolz0iaIHPLG1HiQi8bwzPR/UT7gZbHa2Vq25KFA9HRKISYL0w74v47m/Z9ou4zhQoKbBC
nLXetI0/oxTjGEn4yYOJng+LhmoU43YgchQlAagZ1I1UMqUeedG5PfyZLmukGmMkiyKFkC6Ir4Zu
kLMMF4R2YO0p8qTtHJ2hZkDK28lAZkXpr+WVCm/LQ94AIFdu+4dB1Ho+ennxQZwrzLBXG3D8Kcvy
UyCr5wnC0UsYZUb13VZE0/DMFFM4rldKAO2u6jS9aldR767YD3HSwBFwJesNBOeBeD8KD07Y88FX
j3UKvcJBn1mEeKPT3Zn0Aa8XwVh1UL3TZxl2hu3G9TqBN7pGmiCvgqXrRTKzooWAON6vYZZeMgM0
DH+IfRMwy2v5/ZjnyIQwS/Z9CArcuZ3VpK3daGqX+MXafrQqICB4o6u7hSGIXUoLGhka56mBO+YS
DTucXDuE/Dwv6pvFw9R0t8/7iGPYbFLJw8MD+7eOEs71utiC9z8H1HDXIV9aPLDaNGd9wOLYuHFo
XlVqBultDObEnz/37htvg8OOFKR0Cnql8FAXvLnYpIMBYTMKMha7B8LBRuiUoE8Q1bFrNeu0I53v
VaexL+u3U5l9pgRfJNm3xwhdfopUv4Vl3L2kDUUBtnu2UjCfEwxzCBaeNfqQJMr+vByfd8ZePTNI
T0cPRWsz20GHK+wJz52pg5/Qxy3W+Hd/sv2sewroknMvaWoM24rbzGPwGbuCZXFNGTp81hlnM07p
krg93rPl9XLbVpzj3GCHGhWkXMdsoHPDnfn0K9Ult+U1Ww+690/xnHYTUo9lAUVgzVyUfFfr9O0h
RgQ+cE9Qq7pDdBUyO63ojOGcrr4CZAaX1PkSKh/NJ8asGOPMzxzfm2FtDACAHZV6LWBs52E21i3X
ofGYWbhssF91pJE0SjG2beVsdLI2jG9Py7MfXbBoSq5i8GGU25DGy8hcGMbtGC46yOsdGyoR+RMY
cXdOtRc46hEYNGWxHpel2ktng39oBP1r+7qxINpo8TpyhDTuMYH8VzkqZ3zAzyBQQADZkETBjcT6
RRokDr+xwEELSET/9lpX4PwzVjcxZsAyBdetnexeZWf041mv11hXcE0l+lpcIkS/MjheGRaToSCp
JDfo09cnWl16WojK7ZjxSQVuQd9bEDGpTZNTok+qlBGbKN9rLe9+vD4kyQa51D0nGbdbYYXd6BVx
Qqhkda2PVDDArBi3NGkhK8oK2HYmisYfWbbKZVDanVUP0W/lBC1spVn45c0ym0RkZImFXOogOXgy
DX+yuAlfVCleatCVeCsF/Y5gAFn544dq9VlWhy/3+Hf3/jRwBQulmYwqFVwePiDsC1XJWsjKISOy
GjmvO9CScupjOTZcqXN7WqDpX0PEIw0pkelTmO2wGoMQpHfu+8csjtwH4lbKVe+I9SCYJRKQvJo7
RQBlJ+W5bfofOPmXIY+qlSM7QgJN0zNvOYUwxpPVRvIS9a8CP0FRuNDdff8OOxz2w2OqrInQVLKf
2HgM2qQV9hF5xFOzcRrnOKvPJw9NRts133IJiD4iCoAHPVbSqY2sI3BIWTglUiADqSTjiFggeVZv
GafmF2v7bAf8aJF3cdDa7Iu56weheR21QqKIuPKx7ZtanY+g+sKkjCC6KffROhx4tLCzzn/UlItv
W8RN4DrvzRUF80xVqZZWPU6pUiIfv+KEHOLQhJTUjf8HkWGMTb7cYqCqyzY42/zJu5hj1xAwVtgc
I7BzTbiBFAbeBA4YRg26ULZ9QGgFWUsMgIYMPnmXLb+KHdZIefbdjND39ItuWofC+PxwRIWB2D2j
R6LMxq0i1GAU02VZcT/Pp8+NdePYB/fRw3MYaxNo3Y8eKuiwRGw2IrIbWptXPuJy4qyQdcuL+KNb
+9jVWy0vRihQNXcndXePPApFeYlbYLpjNj30rPknWUIChuDo1h/6gyBz8CdY7mtyOULr4AxIcQQO
oFJ8+s49TmOxdUmjjBI+Ac9WYzITL+NDoN2hg2jE8RBD5Jlwxez2Ez6PAKQ+I0bhyik3R479v89E
FfQtIoOTmIHkxTg02bx8CSrLsUutFKOdLZc+EEmfNB22SEky++Ej2dNZt3r35dFHPsGpjZnEAKwj
k/oxXv2+/jeCMvSZngHNpE7qTk4EFWHLLyg/zNsfvuz4j7QjleCw90z2Qc3i1SN7iD3QfJoEFymR
WJaM73sS0PdyUja6Uh18OjVw397TP/Xo/OXioqTKrBwpvppsbQv6+0xMU0VEVDb/M1Awjv7UUNKV
NiJIUt8DajB86Qp1wNw2gXM3Arh2641UdnXW+xseChce7Z9AQtVCokCgftSABd89p2Fl+tGO4bkC
uL+kVh4o2LpzEBJSs4yHJvyovbLQ2U21OVo8QKNC7hMIgtsVqVlX1kIuJMKRKcZw4HEYiA7gf6BC
nOPyts8Job2gGgRqB/1fJ4+o6BjuBL1sCMRiOtmRBGv1FNPivopoDAfrBsxSMeFJ+yNBUV+N5vXx
TxsGQIF+m3dAYUojYkd52RIzxAnLj+JUhXkVtzHqq0GbLLpPX994iGs/wTqjIUBcuen6UnjEDDue
sSAsiqWKEtgMrxYX/HecQ/WYh9Ho4xQlTIeuOj4ADE3gH0rYcOASZP4Rj4wEfobVPIcY6/pykRSG
hWtIix6EslUeHV+CJLQZQnfckUuuMo8TZ0meQqbXQW2cpfogZdW3SXUG7r8J581PUjRhy/pv9eAS
Noq9nDf4fplU2Y9Z1PY9smUu2rZ1pmY/WMXHdBK6mCTab6O4wygYFKJn3vMXdEarOElMbvJMCqKT
AjK54gfon/bYlIZLD1d2NSB8GJkboGkeQKEwbL4+l1ld2VVA71KxCVS50OR/pHgj+dTkZUiTtyjs
xOYncXlGKgT3LbZ9HNnYhCt0jMW4a9m5V18HqYl7yklL0zSix4r/fxnxSdJ4l4lVB4FSl1iGflDP
fnW/kBrk6Xhr8TJi6ILUY+Xlm16Cj23EsTmcbENgeTAnHBCeCD+T2/WVFb5RWDKMgXne+5Dwc4ET
8aIqpLh9U2HvyfPvuTJxN+NHx5OhqTBKbgxQ6ZL892dRaSRq1a12REZUDw3LPLUEonZFrphcyWT3
H0YIDUb5dxtISwCt3271YOIJybwtfQQrJDkxYL5Hevatz4ZJRvRqYbWyhln7yszfdW/+wQNJZZOx
yRFkUBe/LGx14g8+jzsGHsbf5cy/3HEIFerwFyYcMm9Yng40P1kSjLVfrBqHqCQJDSnzwTtvtSeU
9x4+TKjQFIjL7lMjovnEB96AYX16+fDy9eMgIVYY4ok4JOOTP8vOSSh9KipKJPss/tJW3PYKCnZU
iB/7VuIbgbHBBX4AmExNU00bXtMKR5kag0mB6CZApBgjyvzmzD99nk3dtg7CYal79KAKmccNAvQC
JmN48HtH1F5O8tWTorLNJCYvccnJ1twU7/VCeDr3ZTwmMeg9WX9pljMt+6J0Q7lVtXwlVAS/8N1R
u5u6PMG7MNkM3LvHrGNxznuGiz9PaDY+UA5IUkg7iLM4m05pCKrpQ5t/eHqHZXCNQ7yDjSmAysaN
+Obq4eVXUQYWDx62QfNJcWleFL7rPYhzZxIpperG2OsI8jz7jRf6Fx/w0gyWDPYaEOpVVsn7b2Xn
+6kka8AAWNXJu/xdSFR3Gmv7F4S+L+BeGkiYarsE/Vw52zFL2jDzbTvp757kjq6i+qBXh/n2GY58
L9Wl5HW3za+aILp/YX2c1nGKaVttJoSuTR8TnfiNNXp5mK2fA/V1LgbA4Y15KrvrPryqII6eLkuI
8WYIMZ8UqCY332sf4AOtqiD1vW5fFTOmmhQdrwmtWJjsm8qU37vzpS5FI3XLqHKGxKDp+rReMkXu
MIwFzKQpScNU0FUSD3IvJYnp+fny+26auOY+hyo3OXk+CtylbXBatm5ngwttcD58l62KR+ErnQ0J
8b+x5gNNE8st7eFVs583EnMvpT/9RIq7Yi7H/G6FHcRKToP+nTrwm6M29zrkN0cC7ySr3FMqPp7e
EygJVVUug2+FSGUlfOJPvaUFfnYcDiURhV+kIF+lJihjw6Zr+QBEx7ldQIV0jYxoV+Ta8MKkO0uH
xBoeoxFyWVitrSUwMmzi2H7UXf6cs16WgeNBUgFEJojHVowQKWOiuIWSMJRD5+lCqxfqX1xXFMOV
2T3RiC+GWym0hgW43nlY7Igol9mxHHshTaV32k/vYtrMObrqixb/q6G+lyc7tczAcV8gRvWmcMYg
1CqqzHL9/j2dx70k+cJKQeuY2MPPtytj51GjkitWZ8rFHd5GpwcFHdN0A/MkiCVSQo84PwSH6/VA
XI6u35LwxhQw9tqgrOFmSHfM4Tawyd/X9Es7Wgqih+NfbcleRB+Vv3gUPQ10YoI3YKw4PxgLJt9Z
AhWi9xfjMVSihsUPtmPtsgo22W6UDZ6zDed8FV31SVnUgMbo5pUq0eGB9z5927ygRHudbyq7Dk7E
sNCK+WPmrJqZzqUiGKY+TyZEOKrr2+RVsCmQpM20zrsJzFkfj7qndYmg/WpAFfoMrIEtmu7S//Hg
SlOG3GgOCkKSAhCwNgIwjBbnJXUOWOdWVO/kZxxIGv53sEkiuCUtczp4lKXjCkJLHY+ZxHdC/UfQ
Fys7ofSWOQYrpPsgGFIYogV19TmM7/5Oc5eB3ntfSWH3j/fscFDpxQpdl2rdNPcMV2XPdRtvlE2e
HL1i2NwaAHeLfLz8rvAzoJnVH0fyxdAT0JFELfVRbXBaVgvZvEOvG0dL5GkUIic87Cg7cCzA1xWD
r40XT7b0c5HWwvc9d84o1QS/vVt0fpUAcW4MMzZIcrvd1uCzaoogP+GCBnF39ORluL+MsRa6gdWB
jY/UWizDVeWtLEZD12GsjJgnhg/DHAhavLPY3KI50Q+eXN3mmZ7UYQR7DSy6tsaHIyFSYfEQo+kt
aSasEjwZzNgxVdiHQWuSVd7VZvVha/5ej1Rfn5kgO5hyjfRC0dD5rU+yUEwBe84cLe5gxRHSU6Wz
+5nbXBEmZJYOfY2KrZ4sJWXRj21YV97V/C1zYobFjCsC9zOPERHIrYEP8rayL+MxI330lP3XytJE
Qce+d1LIqyaTNMwc859aIWg2Sab+pT01CxfEFb1yJXmbr6ir+UQ/lE9ZP5fTak056NbUmFcI+JwK
P9Ss8aQCpD1Q3EWgsU/ins+uwtWcFoqGnViyvFtcTImRujSoAIF2Kbjc6iJg7V1e9xsOabhJgcCt
O/Q7hfozfTx9lcndwp/PhWQzCeJU68FQyisdXiLR/xwBr38g/616Qyp5SpcrWCsvJwiykqnsA22k
VZomuabdd2sb57LfCOSiip1P2YA3SY7I1xrWv1Bg6255A/qsKmz3fYh3NbN7sHBb/i01NidRs1qL
0Ib62mg5qqr6tpchUWD7bsQWwH9jBEICsomy3pxzanRXL+d6Kxlbvy71EeCsrYhLx1UyNI0upq6G
IjWhx8oPAdeEmqzF6DijyJ2ho5TVsCdI4hQAI9ORQ3V5O3f6eKXGh7OLjaDtrjYnSKQitW1lRV0n
fNchcgyDQVjqiAxWkiHetixWGZJV9TQAzv81QorQHj9b4xcuZAw7gWbtoTAeOaMK8XsDrw4w1gwz
9I2x9HshiS9pulN0NJQ4nE/NTnpLRFV1zaAwciXmu/HyhYY9fSE6+xq92Zz9MeokLzVEJ2BreNQd
BBmhPJBX5QDl7YjojVpDzTRR+uwr1rXIdb55ZiAq0tLCWM3/LRLkEc9bmcQrsgfeO8Bw8tFBhxyK
McNL3K1ONAU6JYWCbb/4mzNxLHfIXMI2mMfOGLizXG3YBM2mX6VKNYC4Q3GcOcZaOf5xLL/cV9Dy
j2xOHokUZ+1LxNHsNjUR2cnXXpXhOEvO0g==
`protect end_protected
