`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`protect data_block
Nzex0BHfEXL7qKQiiyLQ02s4j1Pty9PyBj7EkeaUhkw4wntQBqazH0Y4xfUBPhcgsojLky2mB2lG
Nq4I8nZOVjJr8dYCKTqXtNx7+m5bz4uBY8Fg9yaIgzP1eWhveWs/jZtZYMCKqTmP581DdEscEIAw
FLBG4WDQRMw1T1+ZtfAcIsvv4IjS61q/BihT5NyS1BZgS1qv37RKcWa9Gm0bBu32YXgkokARKxy6
JTu+SOm5EYCwH6dzT1hDbqS0UlgrxtFUjiS0cZflYpb6Z4q0rmF216/VtNfe3PrMCFA/narJWKdy
bbiTOj+IhMHuYhMrHMUxImJI18MTtIIFkXHhT8Ynb/lfGxhFQZFcbGm8AIDNAnS73vGIcoiRDDrf
W8uLrkO1m4QQtzM+4eIuUX2ThVYfwYfwsxbp4ZgP+ZujchWPS/JicjFIP2Qa0uKfz/u0192FN3nT
PbTQ6VJRe6KSvWgv8RhiKW/zbBEkrp2UXhDLQKXR71OjTpVunPPB/20zVVVZ8QpurkWl+moTKWDm
4uHf+bgqkyKooPQoaZOi8AuQ7553KpfP023LhRsFGFlIOXGKaRIy33NRR3DFnxZjiDAfdgX19mSz
DGoGU4oOKOKs+4oJdb3/PxJ3weQCjleTh7K7kG8Io1CjCThmtB1icvg/zd4511ou/FN8By6nqS6C
8Se4euurMexxcgWqF23zWHjGFHQ8hSCHgRlPM74YuNE4hxi/bdJ+QvkcnUCEohcTEFmZ/W9pjAhJ
Ko5mlIh2Ni/I/ZgGcO+xKWN4yadLj45IXT/bWeGjiiWE4nFVwVSb2lUq7/Dzh36tWpOLI+dwHvjT
URhc9WW0Gwa7ZIuPmzJwmueAmyuC3azq7plMcH7LlDDNj9b5LNpwJdpjRx0qTFDZGR3VeCn1PTpX
BOcp7DIMh856B7oWzeu/5RmACKlLhb83CLcIb28b/GEurSMgc5rDPbT10NzvZ8x1dSmEASNjMddj
7grqD51OVnuHW4FYPq7TYXJRLrxrCt/c7H6rPA2fqsIuBB4LysQ/DsAmeqmOiat6EJqu8YPHY+NB
RJw5c/7mOuF9lMrHwaYWDSWisxywJmOraqv1WLQ5HdOz1BTmxJ0yNJoAAJxCUiRPc8oFc0HYHqwY
x6PB2XBZ+E3Gm+6yy8ZeRxt/1wxZivvr/N7H9NHmMa27il+pqmefrL/gljBIx+kfkX2z7Hc9mPam
hXf0eIIgIKJVvj9AD76K5GkFaYeokwwRtBF5Sbk3jY5tIIIYFTbtL7hZS4E5Chj1GXNTHie0jELj
5LAegKc2CL1pm8RNh4u5NLmHry7VQLvfIbwD6ZK/Uqd+gQmyy+naTx01gK+E5JgluqudvPBGo+3J
XvP8fuN3cZ6SVokNMCUS02yyLhxIiO6fjhFv5Oroh9G4TvibFA4RqL5Ebu1NDXGng6CI8Y/9BkWe
kqwAfpqyYOcSwHG19aE0wRM7xtEfI8rtYzMT/hRNYImW9WZrfWb/JXt5LQ5cUAs/bplUr0RGM9z/
3f+gyJAZ7YarzFexjD8K3CdXKJKa+YrAqhwMv9QuFiRkTH2qexDiclXtj+G0XwxKuH4dU1clUJjE
4L/0IgapWEH5FbeyZK8icUajhdzms7eLhi6PFvqRAwJYMPEGpKLD3z1ug4hV1v9UBVWx0Rvc6r4q
xJo2NRBrtw5oUZAh35XpYIMO8br3pf+NJ1Xp0kpK8Ze7RaNRN4+GKG35Q2K6lrkM8FDKJfWiGger
ajc1k49OqoSjGJhsEog6eugDPoyrTKuBuPgfyT3NOjes1+4QhVB3aGz5clWjrQ3QrpV+lGY9ehh3
Cqk5ly6/2RnKtoVTNie3jQWyeT9Ev47wcEXcRfT3umrsozUzxo9p++R3d7+NOlDmxuGGGftM1SeI
SJ2b+NBqu96sNASOi66K3kz1GS7j6M1ZlqItZTMEbZTpZLgxnpXPRKufkTem2Y5tmQnkGtzdN0Rg
31wdKtHu2p8soOV3rsiBWoE4p9KnQ8lNsB1KwFbNCmX3V49WFEGrQxs9wPH4yoIPBjjFv0Nu1P+U
OH+TqniyYyyImBAVPzCmqKE7eDlHX/mibaYo8KY/jNjdE/1SuUaYsGafF/zk
`protect end_protected
