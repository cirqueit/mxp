`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17472)
`protect data_block
xDWz53Aiv4YPVl5bfVA672qB8dX/cYmelHo9PaUbQiRDQROUvJ7v9oVF0VpYccWyeUAsd53+h/yo
/OUFhgbcZPeIFEuF417MMTZECt5PGuKFdDHm41Y9jByOv3IPDd9p8IpvNRRABqukRQNTmLQCUu01
fWwu2pSMJOVBmmgOeHNcDim4I1nj6Qr26KtN9uVsGePEZ7rPbqyqvidvM0DTRMthEj81OJGACfrr
WC15njCDP206ErGtb1N1v7G9Hn4OqBs2dWl6+Z68f6MmDBhZgVXH89kptle0v60gSemq6SlBZeJJ
xNwxpitEKDRvejeErNkhSXD6gjVS8abzgvIcKbbIcA7vRVKhHHNjzfnB4zAaWS/kLfVMWUd8Nsn9
E11DQUEfQif6YF3kXVs1Z2vfi6LtITixpouM2/3fByuia4MXpXufEYXnx8pvxJMfrtpu+1TP0SNK
/3rrOsy386AgKYhpoTUWmi07UKFUf3S1r9mt9koLUVsXQHRnlWZ12drOIQ8Pb4Iv5x0n2NwA4QtP
VGN0ESSsRpY6i3U2vopcT2gw4srdYehWpxaX/U4kh2T4yThmLOZpqNrvbdZVGtf/N1sBofeVG8IZ
EZ/IlMYyGoOKihhJ84jdMJruJh7hYJuxqPHeyMCXygyUGua02ztlA3qWJ39LGCI0MRrH3eL/WSxe
XEi1grr/TfonDAUPFU1RLP205I0yN7pkAtMFPjck5d3rmc67jKLfkSvDg3SIT0afn+6iWVko7wvo
5YY8qaKRAx02Zjz+6CD+r4dJEP14GAr/kcqx4scyr0+8UecST4EN4qikKg8CuGvs8BYaVLZBOLbf
OOzfliYNomNlXhu8ACUjVZDHsk8loz1wtG1ILGgMuFLnV39fsxfMHMnyvw+ztQeT2nptM+85veg4
vKKqdR6EaNvy3UPFORdCTPRC05+u7fteKdKuIsf/H1OU4b6+g+dLXsZf+YYLtdGgF8UzdHTPJdME
wzxy9O/mje203l/jjickuhYo/xbAwjfO8Z1KiCg1i9Dk2F9Q2zv6SjH0fcHhCzVc8b12nO44PtYD
Qt+dMxOLz7fSXZFq5NTQJyVIBLMLuWu+Plz7DzLqhs1q/cyeN77hlD4GYFHTRaRax0q26vccitYu
Vmsmdhd/0ojUKygdnTelQBI3uyIAdY2icx0C/XGCKxZq5SFcozxj992pD3gxhW6eyp8fiKkh714k
65GinKFBO9noazAe6Zlesg6rS4JyKXHdnVp9dC5875YFkfsdbyRo+kgJQSVNSU3BAurjj4M4GJgW
bu199mMGzAMIXaEUlGaJJLfJIOXb1hyZ8IS0as/8PzAAWCugK6R21RFvu07Mlqe6s4jbJla9wCKD
zavHj257SF3YV+JxuFKMMGRHD4Ajok0gBoCRltKzo7TQ28aJi48gsLq7vZ2ZUhosFqTZ4+i4RoMg
XcQCW7UV/cI0weKGf/pLdBZjjVA1eCu45PayEhAT37wzsOvEF+I0K/dnQRaA0ywzpdOwbi6XWi+E
yntPLaYfPPhZvrjlsXBfJ7H7BOczkYaz6YsELCMWKXaba16v1asKwOEIt3H5P8gxXR7NVyqnr4AE
27IcHm5TX4Z78p6p+XvLLoeiAlNw80Ff48hxICVx8UC1w0vcQKLqHCpClPzw3F6tvf4ndmK+YRYI
IwICi3tIu5HB2R/PEyesDmTserFuoIYfxsElP47xcOOOg/rKBqaYOZ6bnGAWyFDOHonNaxbYfKFx
j4JjYYkpjOt0aFA+XJ2PWlvLNSYv4l2eFL/IEZBHf13vE5yc4nIG2Gfc2z7iKKDdvR/Q/w8Zi+rs
A9xakmJIrP9D88MsrzI+/pneSDHadKFtG8OIVaACZCVGUK1D4sD7HczU8swcLS2h+qYSM//pbF+p
lss5tYg2Uo6Yo9WcmSns7fY9KGe98W4gqcGoMsvCmjtYm1uqro7YZB04kJV7TczU57thT943P20Q
grkid4ua+rKnG4ZWR8nInWwvkjQu2sNzZSvUGW1/dRTV3WeJ3yUh8GA/VopgsEsgBuVd7RLvLr2A
VA1B9BcWp74YRgTwpEmni2Q21/OYd1SE4T1TAfYd8SHsofklTVVdl2B1dS0gKCoCLezwUp3kJZml
o9P8sGDf2B3ziKwMkob/bcd3LupnpkSeJpLFYuHh75Olr2BOne8GgZulP6TsPnFPgal31ir4HNbk
IGfY1xkBfay4W9bAE/aQ6iL9ZbFyfbDj8VMp+DsbSLCbLUKtBfx160Q2rN1JaG7LZ868ciK7rF6H
GiXRKkXrSS8Exj+GwwmQRFB50Z78I8sDciUjy6J747HAt+A6cXv7ILWBYa/SexoR2EAhc83/bqmq
jqGqv0o19WA8+mBoa6+YXN8APQct5ZSLJW42uVOJcfelhKN0SjsUkT8U5nUc51lMkvNqIu93QyvM
E8eiO9DOpXB1CocYgkosTflYiV8yHKsEiJ5wOZa0EpLJdnnxw2RUcmFBvL9MqJiy/yDw3GBSyeNN
AfiEbTociW1zy+j3MBkgznkiJOy9kYA6XvJ/TO6p1FYFQsVCLPQEFM2qsBPAxMu0QdFLUNseDDFz
2y8QlMN8kjx2uUsrRYoRRoPrp40lnbrFCTfKRb50EgT4dfxq6rpw/deLg/4HyXixGzgBG2e2saWX
CXI5tFY/miLpFpSyHu4Dx8px9FpJuGqNv8aT6Jsshrxau8edQ7NRsy2C9YEla3H0ZV6pHOpJ/FCk
3T+9PvWppjrBlCg58mObGxpFmlmK7HkJ33JBcoukluhp24j3T9bW9BaO6CyycDgIgxq56ZszlJ2R
whlBIwDYPjG6asV7Q+5SiCBMZFBLDo+TmjjrYg2Dcfhz8VAhBh/tmW6W3P34EKt6UWsTfp/Qr0QC
8F1+Z524bNMPZEEd3VrOlRDW6wr1igT0PAQYjVVghsSS3s7/JkareENYoDNv9qUqAn+xrrMB3cSu
VqA1RMu3FXV9I2p0N66lWZOMSku/usd7aW+te5fhqcpFl5kYn3xIA+b2PLgxpVQcc0HZrTVny/bU
mBe60cce3aTAlkfx7XJQf/dfI7YbmYudUFYESSOvkObUFkpt7V7/F4QQxSYZd42f+UNytxR3iLIJ
rwZMFsJMT3z1PMa0HhU8ThctMfX1ndieUJ6VbvQxS0gcLwFYEhll7/rWFwDKaY2Xlw++EVSKYSCv
s5hzSCcXz7Xkf+nelbcB7MwJS99XSfuT2YCsy4KxKSHdsJlEE3P3JhAWs/IaMa/ZyaWavj+apUjy
2OfZ3u8qT7f6MGzchSQAM1Q/oeGo+7DVdgkpkpv6kB6DxPWwLIWZhTC+bg+ENxVyZekO4RzdbCW/
Obpxl4DIsDUX+n24XH8l8M/rMo3qYKtTh1nBfqRRCQXc2Sl8vciQ2jHv26EV4Jkhq0iGnGvS7/zH
2MM+rmTjvU+IKx6mzjea1kZu61I6KZzsgiBLULCH2nmGrRrjTI+JmrvVMbq2TtJFk6Wi5IhytYEg
ti+9LFGyAuBET+SWMuc5ELuG1MIKhgqJdU93h/lGAPiiYZpiozazConGVwdlbR92wfl+I4xEZrCL
H12QFS+tvjdi+Q/OiIFziFCy81XZY6EdzbXDUrnCr+vPTXGfskVvN6jty6RtXCrbJ1kDT2zS0R8C
fU9GM2Qx0RdOrh1YqMU9qGmbspg7+UnU24zsFCpAYtBeRNQA4d/Sd9axWHeMv5b5R0TkHA2b/AGp
1alVVHS7ga+xY6b3HRRIJYQ1Dxh+Tc9jK+51wZmhw/k2YuyLi9hrogWoIuOXciw3FR8WPAiPKrsf
Lfk+MStn6TGKNLqy6MhsOVh1CJ7GuG9UOkx4m7oJo57ipIWLEZqffGHG7yS6sg+liMUpP5Lm7s2Z
8xPYU4z8M6dp74MvBpnvwSq24/0/TpPTC++bgg4m4eXDngme2Iq0ENL3okz+pLN0zA12xGTaZLtm
vO8FwfolHO1aert9fLqb1cF+xZ1JN8qlDy7Q+xeXd3/bcrri6pjtP3pW5516nIh0Lj0+rYOI5nr+
sm32bOu/Y/3rb9xa1PISxrCuyfHUqJjyXS8heBGo9mKCqdzM5BBfGHeUNWpGVFIu/BTXOsfcqQXt
VsD7ndi5EFwFGFFSYigy1IT9FjKb6pSBgBQ14SbqKiIyZW3fuE7DTBJelPHnjKHyqpxtNZNHHu2A
SkmZEsTUfCbxXqW0DolbIx7f34szYo0RdfSKXch14Grupkki2upHRqI/UdHjzdXQfV7bFpYnMvnn
RCJsNMgPXeIx8+LIS06aog8BZw5rLFJ1Hh5D1V9yjbzEd+iGZMVH5dQ2jmPpbbaipONyfPsBEy5q
N2oPC62j44OsPnRtW8gEz8zl1c8tM8kHXzJNvrgQLYcomxFZf+b/fZfDkYtYhmQ7p+MH0IenTM+W
+cihpACD4mmIFC/OPs4cVm4UtdrCPATSy8h5gwa7EuBtnkhb3LhqM6U6jRGnpWst0c1quEipiPSK
g6Md8hRjN1mIOGP6yN/mRASyx5edrCBIPgrTnisNe1zBwqgB5Sezvbj1q6m2FL9ennaw6u9hyUUm
y2O8sU/THy3iLtNfrSKN5hQ+ttx+OZiqszR+84agS/AUERjDPqzi6VHjG/eXTc9jPmukmPpYbPy7
4XZp9Mlpe+/YvLPvnF4g+ZMOrkaVGb6a4UfDiO4BqLKH36GhNYW9uFgCKjU0QMZZRmwpJr3HlU9O
1jNl34zeDdsjZyOE1ZloLevjmhusHQxj/wecp0J404BHv1TUUL0DYgAS3A15eLXG99d4GX+sTWHN
Sdyp9wSL4AsmRzGqqg+GaI252ABEzUulPRBiRS431MDjM2lhSA9xKVTWc+ty3sTSbxxX8LSqoLhu
HfGvLgcNaFIvBXTiwSG9oa84mazpV+mrtKn08GTrTprxpFLjjwUJ1q/zFk0RDe8PRYGfJI45dHTK
9Al0T7okHRVitZiAXSm5vF8SiFHxNXSdFCF6Svo7uQ2kkbzGTUFcBhydX+ZU4SwSqfpjHLI5RpJC
FfUrv+QXWmtwtmcCZrZkVgQTFF+tztXBba0dujw5GS/2r1VEUWa85OmI8HvxC0utOz9GegSt9G50
7AVHGJiW0zXwuee3OMIdKEnOruT2NnxEr5t8ZGMxjL8RyOTXTPFA/cc4gk53cDBX2AxptO8GOecY
a8QbSpoEi2S0VA8wNQFrFjZq9gscETcMHSQjws4wgYhg4Ps8lVrEytZbsRBjCFLapCfMbW9V7gxP
eeT3+CIRQBvPvzHzDDSK/NOFhjIsfwf9551Ve2iX2apgVx3VaaAGyjOGA/aauP1fxvQsHar+XCCy
0rdAqutCizREted208fW2N3rBXZgjFcwTWV3pQ67EZ70u3AT54uzuCUjAZ4WOUzWFrLewFNZ0RrT
OBPumiPoWwCHd3tj9PJRB7Gm+soJRaf1JqWA36oOIejdNO1AlugB7+U1A9y5rxt2exu0qqVUI/xQ
jwny8p38i6pg0tOTLPhltr9WD9NaGArQQfPpwbnXJq5VwkSvvYeFR/2JhwNJKPiBJ+j1GNSqWHbq
FZ0XZ0WNhXi3ZL8lb8uHgXScTrQGdv0rgXDyMhpBz9st3B3QjkWLenItuo17R2Qf8WB7f5PXukVj
Bv1d5b0txjnP0iuPb3cyYY9HzJyZgSTv0zUGtRWdgu0GCKewVLEC0K3e1pw4OU7uWYZBzGrBSj2s
QBxprMkIWXK3Fpd9yx+hAOvEwBWRPOCDjdD9s41RSx4Hue+joAqfKmszcYrE2QlRwBAgPv/sncSU
JNhungta2fi/bQK6/Y7YKtplzoAd3FjV63C7+ABLqRUBHrEwU7bGIOOum1f4dUPaiPmyvwMeJ8LJ
0v40aWJFSUTycXx/Sreko7ElrHs/3VDGsoXr9ky99SJYk3CwJZYI2N/a7mnbaUMS0FV2ou6Cp2+7
ScONiY4Fetj/QMwnzYxF6WOoEGRbnwXpjAI+OH5Ct0uQ+Wq/hq1v5inFBTElG9xaVG6qEd/JAnFA
oUJWaBBHvF/LVfBhLCtVvNlmsofnHVF8XNFFfI9Q/xn4lMnW3A51IxEU60iKT7gXAFS4xLHecaZS
G5PCXdFruTdeR7n/X4100VWyZlNZo1QNfItrQw/wPiPpS1vB8D2ehiW7RubI88yBGPUxI2k3SpZG
Wo0OGW3H0raJL5hjKJvZU0qS/Bz1lS9NueXPl5ZjEK89XoHmG/8HT5YyUaaXtVW2NCtRUOp+QKwn
bevr3/53B55yyaYiwkx9u9XW4EZgLfXsLnvQ5ny5Imo1TsnUIMkkJFjeCcDyJWZ3Gni39LZwS6g7
ogmnIpP7BpHHjBqwkFKRM0pKBlzk46j2ZomE2l6x8OebHqLcWea2VPo8mDQKbiFkveTExagFaVLQ
6vcYaB5x/HTUl4D26zMwKG1WwwnWzIEfVlgCIxC5cr9Ojt0av+kKeXPCV4fJMwyPgi0vHAuDiYtP
DFdngmuHMN7SmobPTcipUaV/2tFknJdWCbCjnBhxrrYZ5AXqmzE1TBj09586NntTI/zEYdNNRbMW
s/Mf3JbR7STLG1bxWtDatyPFelrN6Y19gmW1uZC7VeIfogXMbTAeb78rf4LyY0MqfVJpFTOiz9Rl
iamQmXF+nMOaAL8eLpC6KpJYCiiQ4pVHQ+vrYMI43zdSVVL7H0McrwYQvynv89694muk3I+F6qFr
Oo5Kk0gNsP4yspltR9c3QbseyTmiwl8VNI3FCw13VTeOho4T9ldTLFpLUxygFOVEqMLB2+0P1m0v
DQVdBMZM0ei5VjFNmt0qtkQ6Jn35sQOW+f3pQfdEkluYTepsx/gd1CoYbmclpeJhU6LfFqYYYlu0
fvnVY54VWmKoqiDzNDlgOwFERt1Mtnnm4rniQzJvxOSbKneDQACLtH/G5/BUJD9rr70EmuvFQxNK
5FJFWzmXlj0kLbCUN68x5purQCrU9lDrwNWfk1yNYUfqtUjA2b8/JPRdzBtJXlX6QRY41nyuNxbc
OlQWYsGUWyN+BpXenlH+/3JDpvsRbJJxD71+pkR4SpivDhb7ABwVxfdyzFQZAqn6aG9wnAcwvQtO
Eiaz6G9RAF2TruFRFZ3nJ1ldasMPy3POjWbdCumwBsBJRHI7o3jWcTtfS7lhTAuO5C53tfifWoZH
FBFhyLvujmk7MI7biEMAd1KWnGwLwl2k3lgR+ZuoMrYSLTE6I0rrSJAy8V2qEA9QSr7fljwuCogs
SNQcZjwGSWDqOCFHX2i0KgLlnq/U3AKTAPHXkRHEOsI4xt9CmYnrB4AiJXhHta33iymj7LnuMjII
q6Q41Fp36JhYCIuTHUtZuSQbVVEm5++cwyF/JGu45TFk6s6+8X+Eh3m2hAe0KOExhp24MjFISxNL
EQd2uPz6FUQqjklhemcWAbA/d6I4Io1tudkqcJhLUBaWPDm8KOvNEC/HfuS+4utK+UCLWSaLf3wg
U2vWBytGx0P8aiGx1CWIOXN48YrP+BnL5LqkKksGdEmC95GJumJzu2OqUi3mG7bARVK5XVM4C5jc
2wFX9eOTpOczyWG7oCUegILjwEDTUuQDvLrHTzuNP8e74tw44ltCVu4eiQ6LckCxTEwMnf044BEf
o/TRXdLx9ZQTtZtF4FGD84dzGvl1EcSdACCgcBDDqIhLfOCB8eQ/TNkjPR56DOvu8RtRW1Aknmag
d3rnlGJJtxqVjvaAIA+xGQ0r/w7qVaxQTb61y4zv2emQNAC6bcWg4Ypn5PaJ92WA0mdr2H3K5s3X
bl8gxqYBfbsUdxUmN8rV8lZbnHftN1c9WpE368JgD6y7D2slCd84P/uRoliJtt7QnTXYlqGCWDPu
UncsyOxHPUlD9IcXS7czwCEDtm1fbSql2PSSzADIPuIaxnKMlpbaLXrV8qaqFKMwtULosAWjFe0p
oR4A/Ahckpw+WWWQI+Bu4XO0zbwlKbwdi9HYV5z9jRgFVYN+YDmk3AGL71mBUw3bA5m4TyosWR/N
0SacL500tjweUABeUHgh737FHSG26TujvcOPvIz7G0pxeRLB1gIrOoBYGg5nm+Q7Bcj++9WtHSyD
pOL8/Alxt0Oy70eI2Spg7DJiWcvU8jqL1eB+9ZLKl2yRSHb/sixHx/f9JsX5n84UzRLOqXXc9vVr
/eVnKSY1dJoJGjI0PV4MuvTYqRgU7J6Q9WIjjTT593qI3wQkJYaW0N6f9gC5GaJAcfxTmrY6MRIM
FhbUUk6uKtpGChEH2W89ccw5O8DiTZIahuc3oRdbvjBivO/mqEnAm/nAz+VxHPnASCmqv+kysvQG
cDKh4w8V7KkA2lxKWGOUDPueGgDdbwJWDItaWuYNAhw9RVsWLxIyugrUCrPm8nL6sLPWeygbNGAD
bXETU8A026S4LYb/l6mJYNoQkq2f+HGm31dkDemDkIcl1i6WyPShrBlTc9/CR+AFvsD3sOq20kOz
Um7XIdcUN+LmL8PYhu6nBSKYA5DloNOtqlhCrFH/e6C5jDY4iMBzf7LNDA2bUbeoB/rOGWy2mzPy
lJm/EpmXshGKZUkx21zxN5P6xSF85liGIpi1GGGG1wuEy16I1MQALvMxNW6YU2qHeLVy0SbjRFv/
wfUwz3KyKTH4kpq9BQB1ELBY+jsoHnfP9AjX6nB1fhQKRDWaKeJ5Gbt7m8aYHej7ZGVqmMp0HadY
0ZLxjKwDD+eh9R0QpVqK6iXW4Ee7Q01W1D4hhdkrPWcrqYOaqzOtVZDsfpf/+It2xOJRdedJXy+g
1JPmwW8oI86Zs6KrRmJytW3ZTUkEHRXLDD8UeSZqVjDUYU6CaYiNnNrxZU3Q732NLZIcrozHj8j6
Gzird//B6zbGzAGL2yATXBB8P9nY3W5TAdOH+W3pknB2Jnj6LTnB9axWJoIc0rFf054tWiHs/CNp
Zv9clNK9ock3vUt24S0JvfhT2vF4URzIkuVpxoGLawu0ntvMIwrU+eE+or6Og1cW+YO4+lFKgk2y
KGtXyhNJ6yv2v6/ItESJMYK+EFdBbktMNVecIcdi1Qqj7h28rrsdtVosCe/goerwzKeNkzrTm1ud
50qhBA+QJnUSWzdQyWeJvJx5XDYSoJb5IZbJjRCsgr9wmpL7lgmnKzr2eIWdXvs8ieGdGkqiaRa6
D1xVAL51LpP3lCHKp5NluliDaDpzdRaiAdPFqcwcVWaTVJV1DeYZ2r1qCysjMEXQKJkda8Jayz5X
m2X2/dslSWDjBCPdB8TZe+n2aOB0MTM9ligxMrvwzY3OCIDvh2iAkZzSTwRYwKwXF6NjyUcMJVJ1
DII/Hzy2oz5u0VFJqnjoNnuqV4oo50GcI1OJbiAeDQedNe3Z+JKkajYHyGEexEIBZ8/5RX2izwYw
bS7x6p93NJDBNlgXXAqO9wCvuZQRhffdYZ7DGkECPv8uFii96a5t3W4Vj2zG51pmNp/vSSEV/RG3
RdYp2WKdx1n4kWsJCLc5t9Hf+6EbsDZGmjtuD+OyPqjXdNctpO2z/27Maviu2QiN7iRwSqGc8/zl
nx74CsLc90vRFLlJseI7pkIa+pWvAsPVNvsSAH5yZYiHY1rbsX/Y8E2GIkNyRfjtq3rGdEc5qbpk
Pq0/yL1b5sJe32nWxqx9y3t8DE8uxopYnR5ILQUnVjso6iMgb3wFcg2/Jece1yXRd18BUQRWc3IS
FR1QWjXOHALgbDkprpCdzc7DMHZTtvoZVxszhSkZL7tAWqVyjSdPaG6r66usztKXVoMEbp4qBCcW
T1jV9GH9KFyGKbHi1GmWWps7bHbCa9xpoKC0GxdnjcY1OfY49NdtEVBPs0pkjqN67wF1PYlewLyT
App4QpVmaKq2UnG54GpmKA9VlwUZEbwu0Yo/JcKMPEBQgSiqnsDG0cOQJR/+w5LJ3Sm+ZbFZ9gIe
H2IX9Lm9/nrJi0gYsMPDqPpcxjP55U6iZcLtxwCUPH4l0cx0fMgzs66Ygc5MxAthBLSrpXm7GXcS
UQ51IcJaP7z01fQTFqz3ntBdniLa76awi+jCS2ac7y4vqoBLNTcgRxZuEdvTImgIUddq1cD77RXW
R6MUAiFBwoSZ9FBb1oJpGL5VEnbxEBaLmdiLTPd4wmSELGKaKgnMJIpEBhiBSpaCqlw8CExGhyoK
BwDrRUBRNTSHVQH3zKQPNx78sG/R66EwP0l7fWdNpWlu6T/K9Vap+9y9gOoUeRSzS+jLbNVH6U9V
Le/j59gktaOVqo0UiguiJMcolkXX7509zriYaUhUp9N0i09fimkrladITJQto7f2KFE4dMOkbCwW
VSsIQDPVJmO1Odc7D4gclcb+tqFzxJ23+MLR/BonNAgeUTwj36iBx9P4AOyBZXvkMt0eiriLR3qp
W7gkYUQ6qGQJpsu00dDlrvc+xcuBn8Te/1ZyWPg8sjwzRcn5JWLwFZjByktz4mJ6rBBuX1j6UOKx
A/wsnJblZC1BtZP+RGcGQkaadx5rGcw4LZc1eGCwTEQTJv2So2qzVULIyN9Knro2u702iYGPwdyQ
ApcQQSDCHj6kbnzXju2g3g6VawzmDjto2uNEgfDjrliXMoxyux+fmtSVafclUDs4bkcNPWF3YeRX
HHI0AVWPDa3glduuSeY01yR54UxS4ATFL/AS1keAoOVq6Wiict0H5YDL8gSFvWgx9EvJl8XOS+/O
bF2y51FIAq/LSF/OcrMI2XYPHMBgUjnCgmM9Etelxx/TQVgaT98pAliqCI0zHuKMcmjy9kOm1eYL
zAHsK7QzyWj4xvsi21KuUcLsEn2tnSVowQe7Rk6YwAx4eKeZxIWjLhnoFvqIHQcwl3uvQsipGTzX
PyDFmKVlUlpAV+sIG2LZ2ZnK4s9Op7uq5feBvodoTpyDLctSKxyQR37zJDTCAzvLlHm8zbhHtJqz
13Xa1TUPCBX863UAMVomnjGT45u6GOffXamDULR7CWKT53IAR+Tl65KPc9496igjQLwCqVKb0ion
YfrRmvPa2MIaG/Duxj8yXLPwzCdZ5Caw9cS2SKiD203aRYbqdxdzO6GhzP0Z165/Rc0ekjiZ3L7T
dV9+yOLPDwL1zHsZcrhnkJ4kERziyeg95MesagS1dmmLZYZc4chbsO1v+HrmXzDvAm92jbrD6YFG
JD8JkmuauPzlNdcj2F+LiP5EeuUwboaGTg+reQRc4lYfyJYGmzMbAUdfvVwSIjhvRsxQyHffcwIq
64Ycm2jlUvqr1ICOYYK8MD5pg1436fkQFAR+6S6rDeHJu17qmOnlq90ZsYTHIqqdsxwxyxsTQsKV
9JHWxBJeZUx8i8LJsxZzPum/9jcTP2tp35y6opKgascG2HasJMf+hYNavvztqXqPBqgLbd4DIjGK
dUzcnBc0yQRBaEy8zc3ZKPacC4/zY2MsTUvYXRFDY3PgmxnYVvOK7q5WRD6P6ughyhvVM+veX8t/
9NNGtyh2YYaXW5Whcw2NjklVUze+dhIDdRAp4k3K36vHsv+hKzaBa1FTk3XPgjf8JgUrtkdpAzGE
bUawLb4Rab29n8OriXUUMfxU2iERRxYf6E/W/h8BYIr0UBO/ESn7naQ40F7IFGbZyu+d1drwg8Q6
b464flAFMlUP1f62z1hEn6qRlTsQr5OibENUgr5+uVhiWs4k3AiebX2uUZWdTHunDvg/sSaVnYUP
x1uSCCZ2LTVMcugO2E5PiTYNYJec1bMonrBKyGRuDj3N+SIFeWttnEaFqFj6OSzjj5pzCZlpvA23
ScCcqN/MbZZwdVl/gAWo6XG/PYgbjOOWmdgJS7HWeqNY0UYBpDBXXbCiSjB9fXV8+5W/JUFLZU6x
p7+yJYce/Joncc52CcPmOpHf0GGWejjjG/nqUav83S2tMU4aPGkfhY8R+53+iV5HiGtyIxqawBzo
825X15FcnC4kNRqTE1uPPK3jqtwAYxlzE5CDnbrfxkswzzI741KNSMotweffN3KI0EhHk9I3U+y0
wf02fYta58RBlJUtiT5gdq2G2q4LrqlBPBatl/stqSCFyTFalXo7aHWYnVwT7iOo/tizd6sbJ/PR
L3tzpk0WjxRZQ4N13x4dj/MDzJloRVqVrvOGhd4Kg5bUICipqz2Dc53+oB6zxsFD/oRLAj/fhYj7
2u6/GLkHBg1bHNSBKI+8vAMRUxE81shH4Hjy1WJxEUouZMR8NLXyAX97ay1pGchvbTBJysQPmOpo
p2VLFkLYeP3lGKrdF8MM7Ec9yq7A3ZljPMQGwoQmP6zKSKIO9/rU1++7okxdYngRSar4hRMAj9QS
0xzAihn6TKoTwTj1NbDH6HCjfL7Wu/4YRXRfDcF+0QuJzhSmuJeGwu3cJOD6CKR+F9f2F0LQO8v/
0oFt0nnpxupH57XuKjyetRpJ3gHsEigi8O12kmvXuWHf04rOgnObxqBx9rNGlRXs8Dotf/2UESHI
BSG+qR+mGfT6m9bRt36/itjaEcGw3B9Tz3ENcOQMq1zAC6t/u+GHX5sbVoScw/Fkc1G70FCncYTM
21EFuLY7zgVJuNFnkCPaOTp4BqJvGPu0VNttWuOyq3Y9xs6N4/9Pc+eaj/LE/EOIIUT3hNvG76HD
Epke7vsuPjvOkZIhIe0+xNe3udjpmHxoSNj9DE09WlTXU61Q7fGtF+jxG/tcpthaIkhWPuXvRcEN
SiK9c6NS6iuYjGYgQDA8XaeULytSTQxQ19D9RXASbF+KBTkTMKqXz0lEy3rHsiNPgZ8JSxLMxMv6
Qd3ApUT8xrvFD8SqgaCHAe/dn7nv0+xTn4G8iK++8m8RskpoT8xRFtU2K/tvBDe9xiVqmp6Izdqi
uw+fFpUGvvVPiNef2ZlaGENO8JXDLdlqUbe+jOJekph0dfM6GHNZmxJLVnj9H/zuHUxDZ/Aye1qK
W2t/5QSgc3B0llBD/w6mR2+dO0f/M+QZkD3qaCbaPkYiP1qqwlcXUHMZMuMB+6iSJb06s3KtQ0Oo
RLKHrVnKVqx1nRq5b7T60N4IpDORwutsm5a7TGwi/VO/nnhOrKfcZSt8w0KuWgpSqGhdNjMkYiSI
Iyqw+IxFUPN2Kv91kSVX0ugOYUih0qtkwz3IUr65a348r4P5euWOF5foZefY890tnEL7gcMuEUTy
+v9SSKnkwOUQOByC3ZoANiySaLAdGtvIJsWrrXPSG5nEOmi+dqgAxgazV49SJUDhNE5n8I8gRwaU
26iCtjdWjk3n4kghTTtWFKJNKusILdG+nvb+UU+wlmCgnBlj3r5k2Pvurugel+B9bi5gqkagii+E
WvWow9J/mJ1jU6NlBkXNT1N/JPybk5F5CUueQWpH/7cV4W8NP+BYWYR3cospMBCPzgrcPFf2J7Ps
tKzFrO7mJW/y7FwGJiBXoloc8XKDQ0nzSyAsi0LB+b1AbOk4o+vDUzthr6v8Dc0+qWbJbVgtn7xF
zJGbHeMlZIqFzSsnC4RPzj3FdOuZsFJzw073PMRruj0pb0FxbdTfcWY5BggtwxL+0ypHXSniA2u6
ipM5Y3lHa3U0H1+2Bccni4rdP6tTQ6py8WVfjVWwB1Sxt56IlMVOOuMKPO6+yLHP5sayRF9lz17A
IOw7lgsiU+kFTrZrK2uvCoRhLEtIFWigkoV0lhO96W5gKLjVhYBs57HXIK5g57pg4D6sYfy9L1Jn
nY5vfVf9rZCzJjrSnt9gdzYEtX3TY4tn1FOm0jIlxH+lOYMMNKti20c6cdtCEP9kK8wCDcUpMkWx
ElhaAFa5/dAQ9Sn0xahA+wMn55WJjM4zyuZcx6RTSzLocPRqnw/j+0opLyfaP7jSg647k13V/e4b
AkNwdmzDeYJFiKl//3Cm9y9PeKDMfEjgpC09T0Osbzt4Jd22DGG/MG9KO2vb8W4+664duNcy5Yl3
HaHLVmy4NrUHt1486ltY0WERJk238eS1h89JqPOt6jwiEUpedwTr8bApTRuBUk6Ro36S6b7JOxPV
H0LJxgrVri4lRQuk42dor5aDACO/I8qoMhSz539Fx+d3FJsYKJu/XCD4Q6Hs6DHitRemmX8B8wSx
4dnpaoJQjgBMCXEy+gdFi74dH9K4RReAsYv6tRn5Hhe8k1koTptLnXkDLqxsIB45QZkhiD5PtYm2
0qOxOgJLnw+P4VcKWIBNycv0war/TnRX+Tfjryp/MJbH8Zwi1ljffIoDckn4iBjrj26+cMprFj5W
DaCN4Lh3sQ360vNTOHkJtpYXXStl+PLmmKCqCnHN0pqR0qh9m0YpNrYT6B5BTPpPaItZJ/7wbANp
ffKm9B7Ivw25lDA6pz4fkqUxnKUEFfFLvL9n99DsGhCuUhfZunFL8v0gz1vjzpg4kxcMf8A5h4sQ
LV7m5UG/ZbytLXxGTAg4ZzhXiqhcnBqhV2PgdWFiSw/ACx5b77WpGwKEU5cfSA5I+T7hqsqxD+q5
TDtncvmMjvC1X/cmzCAkTU6htMKpT7uZDgk28+mf/JijEglfzQNx0caUi/XeqVPI4d1QKwnD7g6P
TYJfd7KOL28Z64BXUxNg6n5PaEbHg6VfMM3jVWWAh2rETaaAzfPCLHXhq9p97+WYswUm2vU7QExR
19qyMOuouxd5WTX1XoQdxPUHMbj3p/UvXov0iMZPoZ4k205DAqrVdVZzlzfzeWO3gXgcil4D6g9d
/7W0rNOIsBwsan/vhLiGcarxgB5mjen4lYrKwOdtincFDviqDZR2rMleBNtrcTUJCQw0gmzcqfsX
Vfhi5uYoIsEC0Pls0AK6rnWrBLtpdlo+ufFH4VuRuQnbShEvfp0iVS+pKJ30Z/ZBhn44T7ZsqUvT
vJV+5choBFP2s2TY0qZ26KauHujr1talEzqnCy7o7FACVauZO9OcwEWWhjfqBnQ17GVNhffoNsTH
lx4i3kp9OldKcEsDFmVhDQpaddFdOZBlTEELXtexHRpx/QlOod0ThXTQvsCdPagbfrrZMiotuE7/
V3NmSm7Sdh5VVs3LI7IGEilS7awxB/M800psd/si+6i0Kw4jKTrzQA8JZynJxNvXOpYbDrEi5T+Z
gdFEMETugTJUo6bks7YdOtWx92E6q1lLgb3JyvdeXEEhGMhbb4S6UqNiRo+1VdD9ubjWT1t0GCik
nTqrY4/nlS2pbBMRVot6C6suF6W7BSsmRiX0LoXc74i9l7lI+cUqrrZNEoN2LyXs6QTEeya/Vl33
1hLL4HAXgKv/3IB2fJIY7QGh1I6wM6sVxO0aYkViJYnBJSJ7N/PDpROCdViiilXVXlG9RoBNYuG1
fisDxcsi9EWW2sIOXP43wmYbcbNv3BrDtHho2xodUubILdg9pt0vRZhZphjdZvv3zuwYf4EMWJVG
T5KKw1HDR0NSNWuJQrf7Bj70mWMyiApQLpGVjw71uWHtWFdkotf9XzfWjbMcGUovpctVNTVUizgJ
4uH8Cub+UpivEu4dNGg/JbC02Eh/xKT6tAU851+awQL2nxPbdm2jM+y5syqQ7yT+aZZhdAkPILnf
Sw0FjYYnS2wZ3f2LTYlHi8nTsu0lGu//iRt1cmkQsSWNHviHj7QtviajMgItG1wO2BUi+tJR8ZW9
rQO+fRDI3F5MIj9e999X1iCzbrF9gS1HAxQ7iwBUrza55pYJOF1OWoUdnuYe1nIkLovnEM0DDEOg
EOmqnNqCHW9+ZhEO2QtIQpCjuK9BR5mn+nwvC0bIMiDDDK5Hz6tEIb4esIg0GaBwAYvxXv1vdcBw
wuGk29RTPpVemnHMt8XP61zsQsdgpcByQsKutmJCsot4z/DeSyTRTzXIgC5FgtHXHjdWI/SxyEv9
PaTshVLbUi0KHEifRSkMdmBI/D2Lywg3iViXcUrAvPK2MAiMEDNxOtpHC0E1a6Lb90DVVgc4j7U4
+1FdrN4E+pxleeHZzwFGODjohHnVEq7W/B/u1CN5yjhfUdSv069pgN8yJ18dWitbaZ4wbts+uCKs
vmxOPLP6U+bTXRIGtZPvPHr4fM7dsQXReyv1UcfMNhIUfZ10ifaV6Y/c0sWl12oyI4Slwcs8GPeH
vqkEybaXdy7WfYj12Del10n/efhmB3yEuNaOyu8CBYRlmdAgU4eh4/9dk2GYzN+fjbHMlWacwRns
IGK+UyUbxtsssNjYEOE6jRawdaGf+h1co1HFKbnR5CxEkl600F3q+lZ0kefKQOsZa1aeshU7beiv
V9SS/DcShz+9stsQo/PrmbjxoUrY3QOtsU30ynRu7xHxoDTsHjcN88/dg2NdmX2lngJ8IlqTo3hu
Yg1Vb/cdSdaSKRKkaOVizSDXaP9LXmhmnpDp9sZn3cwpdBU2DCzWJKEsX2P/WclTpcprhAPoADgH
ekw//qrVINvYiDMQDgkrNSGhO6G28A0HG2vy5SVkPfAG8QCIl3wDuypzN8AXVYlWN9pwGWIm7Q82
pOQu1hiXH7ZPSTSbn+xWdd6pytl/iBYDjnw4l11b+hT91zyoiju0XU6PVRI0RrCJCmlI2rZBxtMD
+HUb7xiSnW8PEC8kxQRQkF24J28soZfsrqLS3/IgawHyqwRsVrTdIBPM2eOzYOjvkIYaf5gs8z/K
hhGBTsoSwl0o0vMD2L0lfw3kEOoZi93ZT9f2o9MJ0W9qAEPepNLAcX56wQYirpTUkeC8gaZoNOSc
6RHSnPULoYjlJLB3ypq7PMdTnu8bXR/sA2LoUqDSJFEdRb9m7IBYVIfTe0PjbTquh4u8RBEBnqHv
p9euMB3u97dvt3TaZ7+P+I2KDMNgO6aBYYmd9UdlTiHMS6fuYLt4DG74McBSmWl32yL9H7I81Qyu
njEYcX8A1mLRKnUG9cN0TdZsY4WAJdODpd86rA4R/3WoDL4+IPNaY4yYjPRM/yBYXEjY0JpFpcI4
45CaeI9vbnZ8+6ALkHx6I07o5VXVz+yBXku4zPANv9gdflhxElna5zop9xm9efs/3OtsONwlAqlJ
s/oE5SaKKu8mW/487QWzbgZC9/hh7/2JmCvwNXoSs3Rqp9DrEaeC3EvOzYI1vHdiHn4jN9NzZEor
ybYIWb3ka/sdEtRMRguGlygJkIxQOLsvPpTMKJ4YDWpAhlRii0DoS9KZOY4aQMzBOrHymazeN9CI
O6Hqswdo9JtForeiRkNpaGGzWB3GUiRriotaOHZse/YRt48M0VA2dOxDEA9Ca+x3QkarVFUY0+yx
rY1CUrog+XCFZl9ZePQhxZPcizDNg+9yFZnaOz7YC0rH/2AnFbxa6/gAGgnGe7WkeQiEhlDx8DpB
BR/yrgTUp0NUt96pHeU/ximwBs/n3giKTLqv5IZo3LiBi62YKB2HaKO80sjmS1TlGv9ePDxbFeZO
3yz6kIvp54B7jjwTKnGFnUW8J48aiHLb77aBBvpNDkbaeg9tw91oZxYykEDYUfFVZLPPwcQRAUst
x0jQZyoh1fLEIeJ5a7awaBq7l2GABGG9SwPaQ73jgM+RsAIYWILHgk6iwq0j38NJMOUA7p6QT3j9
DHSiqvJhaL1D6Y0NnYuTwlP3ztAut0GEawH4lYP16d7B/6YUnbZe3gw/twsjw2vcG/64pNXiWNeP
HSZ0xnTpvBs0KsETJFNTuotFlNe3U6okbSFtvxePHbNrmxAV7rT259x0jbOoEjsPHNQjqblOYu89
qFfLvCYn8jrAQWveUK1aXfoRGqDPgzKLf7bB4LvgBOrzFagxebmfX+Lbk2W/+V1yr9XRlbLd8yk+
eHVpvQbg1fOd/DrD84zEPoUsuDn/slqFWQavjrI6E/rE7fCX1MP1JtIo9JPFEFddtuxYd5/bkUT+
MLf1SW+EXSQhUWdpfEwhvleZDJCrOuiqGGotO+mOBPnuUP2SfuiM8PUnJG11XZEbJszK/2t4sRG8
AL3Ekx6S6cA4+BKHG/R5B2k9ziBB8H9WppQNCOyAOLPJjus5/jggJmvL1gX5NRJYtba3kB8LFlGn
0TJgACMpKDOXoYd3oZzkg5noTIwUJnS2Td9tcJcJPe37eEMqUz3uTxLsmenl/DxImgguYJor9vMN
l01kjiIOGLbCoTsZv+ax/8oPxlxX2B6Ksi8txKcrdztRq89b1VfT4MhC46/bc0Kd2xYEA5a0prrC
ngjt5fSkC8tjBmPLakjKTnMf0qA+tm1X223s2R3mn4T4DJAU8k6DSV+++5mKjhR1Xu9/gI2gUgQ/
NMUjR7eXPEpoWpbWuaD/22qnMdU3bFcPCGcZEaoum+B/FJaht/VhxZwHd3/E+MU52pV+Iu974zF+
SB+H/t/EW/CGsOg/S6goG8jen/HhLGOXwheOc8+ttQwRiTuX67JvYuiiUShqYAak0ucUAkjhIwjz
8sShVb/E/n4dFVEWdZ8ZhC4hKQ7XM1B7tBEBtoNHfZN1mnVui1GmaQsvfZF26QDdCB9onp+bO65F
I49vyb0SXeUZX7KEY/yhVHCwpHppukUnSLU9wdiMHFYecr5IftxTAoJz+fe+56WNcwBXd9W7pObm
9ty2M/XlhRgkwV5sQTCf1D8QBZD1LHad5YvJSnlc38CtjhdZdGCC1/jjRr8iwO8Rlxwclx8FXTpH
cXtfQZWbbbv63BnlsoQ6BusMT7JVEEkhQfNWuLh8UPxypzf6sSWRzL6G8txKVgIAVFGuohXXqenD
uT28JKH8kaJ1SYz/GgkpD5AsLNqsk0dj+mWlx5XoRYvoEYlH+uW/TmY/Av1mLhCHeaF0f67Ju/xB
JtpX+mLVSVpe2MHcFZHlFDT9XMXYea+1+YGdtfJT981ZiarV6/D6GgwxyK9dR/QTAaO7tpcacl3O
B0uezjG4lhKFTaKK/WJ8fY+MSjAVtJ9ecZBonqfLUXrfc+y2aV8zXaIPo3C3oFclhIwUiuQ75jJS
ICEozf/6nRiEXOVMO4NqXBqfEzuqj3++yU2AxqXUAORGilQlrawRkDGzjJ45OJldKXbkCv5UM9YB
cDtl2N/YNdi2xfjbaY15SbNbhV+ZSCgrwyoUQZh2K0iEjVr04Ey13WJFtx+6oWtcqJ0lkrKe7UuQ
GOvklcf0LXhaXa2DsrPObJhC5qneqhSpmd62Rc7vlwYBMfQUHAg5E8bJ/1YElLtosFj/uWQUCiOV
+9Fw7zBsG3BsFrfjMex+WfjMD3CB+pG4k7X49KhCMRdmK85IkAHEBUEWIq0uZyfDLvq/e3OhqN65
jP8ooHxbndhrqDTOkm9TyNEsWf5zGPkVoIuwx92z+9wpykN9OOp1fGoJR4k17/+WGBmVkseUHjBP
SNkrueHIrDw/5Wy7oML51delgdwN1v7wX3/SWDu92ULftvhA2ALT6ERpfFx0ndpWaS8e9dnLLT8W
VJDpnPLzmwTgkolTi5fWeAXKkrq6ias2bkz/OHgvNiM6g4FFFKkP463aQxKPUJTZ3NpHVf+rYf9a
Ysjy4lJPHN2cqTfIjMnM/88/H9qOSLU0zqm+gSKvYwX4IdbKYwOEoyyZhulXTVkCdwcMSE2hyWVx
BTK+JcipXKD8DtlEpDkMKcgSguHaETHUi14GEogNQYDcFqFmDft+PFTU2inRCYveyHjvVmaJsij3
/0LcW3KABTrIa2yX7fApTAq9s+Efm3SxOBnjlH/QNdJWGqG1xHX0b5wdzmMdVoZwbt7NFC25ctnT
Biqkp9GtCwYGMVqOevtcR5PfjjTKhJFCx9+X25GUFoWYBbovAaqUJdra0JEXy5z/65HvtiU4R6Cv
8s756eCya5raj8etTUyilVoih20HKKk0Im/S2Vu1mOzlOkjLOLodBq2isWqzJ6BUUQ5D70yp3gUu
bdCTr8iffsFtLiisosZiprnaO6LFMXn6qBFGguF5PZdhIJ6Lq+Tfef4BeEKJs7dI3zOko45nNrTF
EbCHBWvsiXSAnVQKO9LdEvFpbiS5fnU5L99fdG/V6pH4mqERWD+rXfWRy1cG3y6X2xtp+fKbOzXo
hH7w34YmzND0OwMRG0fa66emJESdbg+ESDq4045r/H+S7e3n+STrnHWgWAqmUkN01hAaeoVZSoR6
HFUQhc5jw/uPaZOOeV4/mWD9u6dDOa2WTrMoYCkjJx7zpC6QJlFfTEVqjYqqkalaOIjK4nZMaH+u
JqdpBL60wUI3199uM4EkbJtuVh1EIoG+GAep58OsZSxGOJ2cxhKqqvbid8+MgC94Z9fgNFkGWqZW
xn1fTXN14NhbWKyUZp7/T7dSvqZl7sIUGL1lB+k4t1oxG6Itx/o22AUXop33ePqA1j1uCrgZfwSe
KbwzZzzz9nhX4fi8AAJQSuRLXKUw6DabJGUbymyoeRrtHFfeIieQQZeARfydcJn1nODCx//RTDry
TAOiklYrgQqR3YAhaw6UED9O2rWm/1PvOdIS75+Fm2bTdXjR4HKIO3F0gSuZXvdc9RZZu2+LgUFr
zUHmegag8BYN0mh1QNjQMJn3Il8rupFvDlas0fD+cGEhTgtP69tAKZcBnY36hBNB36H4jeXMl3pX
PDxQWUPBaNVkCE3br5OxxlgmKF8LaXY70qkoqVZ3XbYUWAWuJDAvlj9boaVovfTh8XQhgQFnatxU
3IMlTuva+w1lBc1OVfceeT0aODeD4f5p4WThDoZr+hSIzpU/ckCLeT6YrvlkYnkAypf2bXbLyk2m
jSy/sz75tBAxuYK6TOJzMNZPdsp9DAJnVo2V6+4GcXPlx5iiisIqS60PLxdIx9vsni2OQYDNAFj8
infN8KnPrkeTvImHoIXBc5Myfv4kkVRmQ7tXNAROKqtBKas+7mutPTMhfAscrTzEThJA/QviOlML
2v42O0OJ+ukJrv556UXS/lGTY1iRIO6B11hJKEvYU9gqF83LN/dCJ2oCY6+9EE1AM2PjC7Wwls4D
Jp64WdP6vt/XtKHsb3pIscFt95M1/NQqyCnUpsS5pIogvz878D93Kq+RXgrBjXzRA9/RySMo+59f
n3JrJL1ftxW8vAoUXD8/8da+Hp3TRb/ssw+EsbLcS2w0aMx9o3n+Eto1lHL/OkEd6HmqqMnNqLlp
8DBs5tQlRZaMIY1YmOKtyOZHuvG2KMFlcpE7DDbae00y6+Lm0Hev2SHSsth0D4ymVQtCkEAiEK2T
mwiyMbRFvZOtYCLJpX9ccwBx9WIVsoOj5SRDzal8MOTuUmhz1kzNPpf4DLD64NXmUcHXrNIIQdTe
nRf2vnIscsIP9tCsP+SDh6PW1jXgOG0kYLiJYzp6sbcIgIIuSvx58VDr/z1mwzBTcxJ31YO18YDU
ZWWSgIxcqSjFLiipOSa6mofNEv7UctLIFLk4fU9DkdixXKJ31Dh/W8LJIrpou880L1e1voCZFQRU
jCYNCek29iq7Mput5uSQOtgfuQ8xt7yQOpToNofg8wzbmH/7y+CPKFX0hq8ZwRImG581vnWd28GE
D+SeTzNpvhhRbH5v3KY+F/qik5i3slrPdmcwKPerwmgEgFG1CRXoJescl1PUkBKjGbLcVXjFvjRN
SVSqPpbeR9z5SLw2kwQH5USYaxHGWpNZsrV3vv18sPLtdulwgeQAxOslLHbqAhCtRbUdb0OCSFN2
gPs4TcrozK03wRScfW+yqpsrxiIH0MVYGkeoD8jy9v2iKHdOFB4KOwAlWagvZtUIyb3W209tHBE3
cKQvluPQmSVn98BmyqbbMzAfRMTwMiXsDCQGNn07MftgeZ0UAtsP/CAVs19Andy1kYqjx5wqIzhu
KdBcWAPV46H8CpE/T7hwlgQ++gJwLTwksz28q9nPDyImR76843K28uKbGe/UPgGbgU7GokyUmKdC
UziTmpeuyHAxMDUytzYaUCrRQi8h0vcqOijf1lulobLyGGt0Fsk4k22azMGixcNJMrGLo6441rPd
e2k/WrVesDRAU6jbzmBubLCpXUQwBQRvKtmLPfzUoWTuKJYA+HQXaUBZo9C9X0BtzG/ERNTHlQxk
aMkyfFTreQfFmuJJLREGH8aBrO25cW0iZF3uZ8CtrXdNFmeP3kWCGJ0OWAYIPQgfseu2Hp811cy8
9bHGtvsfaTH13MyJDsRPVmqUkLNhWKxNm5QucvKy/rnCCYcFny43wnpyJLaaxcUCMf3s8NyDVcl8
4vbUTgKHdo9Q+do6uRNCfrBVs9GOa1DwXV4c8je8x7J6BXWAMGCI2u7Hc1oPwv0MqyZtbawLOo1S
TcdJRXcqhzSI22RifRI3hWkiozpQMgrkC3qlt0jz8xfVBXukFgU2ON7oZKbRJxkuoDgnle+XmGjl
MFjZSQnkYl8Z5n6P/hDESf6Y+lxL7pwwawf3zkEhB9pQ1H62qqFpKfTUOgs5TivElITOpeP6t05J
A5hturfy/gVasXtkhVKsftnpqn9CtpvbwmtPnfHrxfmp2cGFl15WnhoGdrBOkVdjDR+5oW3ZAjWE
lzdauM2QP5tbEqwb+yEbV6NLO1Nk+nq/0BjxM+iB7BRnskjxsTZ8FH0PMXeAoX3cL2C7Gv+1IeJA
G7+9XWQ7Sy5rRprbPWcRCjhE4PALrCbmjbJI5rwh8yck8Ib32NN8DekZmF8Ret4X4uO/QDEIBuaV
oFMUcw8WuLRhMsmnlCrq6tiXRCWUDkeAGgQNsiHKK5qmbETXXDPtJ8tVJOTiq1ihIuUN2w5A0agA
g4ol6eXuakEJIkf3pPQYNZfFUMNHGM8ELY7wrwV9SXuA2bnFaVi8Dp+fh8iKkOQOawjPIaq3aobk
06zJTmTKQzZL5dTCOr00SrkqbRpKV/c7K3slQrFa9zhFz0DYz685xZyT7BlF8fphyv6pQgjML6Dv
H8dblBDyyFZQBf/N+Rz+fqdEbKPSVVUy+zwjtuMGRjuIf24jcYr1TwsbbKwIonPJMniZyt4T00XE
R0cMH1dY/RISEBGOP50hlhjh/fbFlvJDi34+LPH7RLlZCxeTrdTlEZO1xbTtLcCzgXOvr5DnL9Cq
2rx9iKGlG8YWilziSMG8IK+1u9yEuCbNzDCrOjiS/6Gb1sAR7sWfDo2yT1jyts9rDQfCEHEWFfxh
uW+wO+0CVZdoOixAAvLtxRHS9FR64wE7CSoRMK4QwcoC7pLSmpvrth5yCwm0VLhhbbqjFsWs4bKH
nXM8tGt7JLjENWp/fZa9Zwu5Sle4UF/pKwgmEbwd5niEIiGrKS72MskxIFZB3p3x8oHGtQwwe8J9
M3Q2bUBMbiy3zjdzTdjMh+QepRJv9zdAHVEWr2m4dusHviZWXZqhQ6hzHeBBykEX7Upid6Mwp8NN
aNIAdF7Gc67RU73iAP24ddy4VDlx/1hmqrhCsAYyWQvbtKEryEH3hymDohxu8E1CWOOjOJ2fRfJi
F9OiqwYsUYh4hManhi60fZ56eh9BV0OEQJ6TifezZIBQuwJehaG3rfzTr2dU77zIpfSe9xhZJCPt
SRyTvY4/XdcBwLr2ZhW8g01MIK03Z1555KwU+e10
`protect end_protected
