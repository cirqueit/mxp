XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[6O�4g�M��'� f~"H��A�f{$�0���|������@`�A�������2U"������lY�>��_���K�G���j&,k�6�;a6���!�y�X�jr���'6k��k�xyl����K����I:)k>tLHN��ϩ������^\����0
����v^��gpnj�����;�Ӎ�a�t�.g�Dw������{8�⳩�RK7�cQ#8*�ZZ���|�kv:v�QJ�ӈ��0���^Y��}�!�R�7e��o���4�оe"����PSHQ�nW�[}g<Ov�*�7�c���u����lW����b�؜ ��yu._�`"��D��X�&�^�,9�wENa�zaaTSæ���伣��l����8�16�<�K�����؟n ������g��t��A ��:�5b���?`��w�ƌ�K?��p�\�>Ǹo��=�ce�BbA���Μ=�s�P��䁻��Qaʼ���V�?�8�R�kOc��AAqI{�ρ��P��O�eMI�o�:�������=��DE�N�l�r��ӊq]L�Z��M~���`;�!��c��1��i�mV��碨��$����(6j-�;��p��j8=D!��(�i���fƬN���9E��8��
Q�1��+ OX�]*�wD��f�p�G)�ܚ�	�|��`ǒ7�(��50\+�v��ÿ,�"��~��,����J��֪�0=�&��t�+i;��˭�qk��e4�<�Ȇ������Us�^!Q1XlxVHYEB     400     1d0��_W����nV�X;��*,��9q�P�k�9�7�0h�F�_���Y|������zԜ�۲��ߣ�H���ص}����MR��ko�ų�#\��1�O�$������{FZy#�?��&�Kg�n��6�u�ܨ��7|%�\��$�/�ܿ�j�//����(�$�����R�j�q�6Y����i�Гz��y�*	�P���Q��A�����M+�wXO/ 5כ8��*]ܟ+p���V�T������UB/�p�"�!��X��D��#=է8!��22;��_K׺_�$tZ��%F�j�Uz�� �&8D��	���2)rdhD�����kυ�m���̝*|���4��>Ic1�d��:������K'�*p����a H�:��S�}�Ȑj[p|d�oz=G�ůxe3�:H\7`J9U�=��v�Z�	6F�>tǖ�	=�j0��XlxVHYEB     400     140�f�25>�ǁ	��:R����Ck��K �q$���~RQ����7��'����C���K����8f���2ͯщ
�D�7������1!՞	+�sdn�P~�rt����sE�\�_ĠEߥ@����׬hi�Hfx~qA���n�p�j� ��o	�����x����]�č�U�k/$�ovQ)�t����\��P�<��j���%��'�̸{��~���1��Z����_���I��� ��Z�.�/�!ޱ��ݠD  2��Z�{�����miE?�zn��l@Pc�:AT�Q�~�m�z�(�c�Z����XlxVHYEB     400     170���0e�U�� �C�L=�a4uS]��� ���<f���d�@>q<��;�6���	��J�����O/���o���
�45ZF��S��/˪�������
u�[�'��*M~3�yY��i<����K6aF&�ָ�T�>=�b=v
��\T���qh=F�Cs3�D5��d``��*zKT���a���_�#I3n�\�a�������\+��fl�O�R�ʟk2N7�n��1BŹ�@6u������d�'#�}Va"�c��J��n�g�Z�JFXT��1^_I�,�;�	8j���a�tZ��%`���U@5t-H�PX�^�lА�IjBK&{��U d�  9�L`�4WI�����
�XlxVHYEB     400     140���SJ	�O�f���<��CM�TZ�7��q��lC�*��:�I�J/u�(�ؗ�BPK��\�f�h�8�X_>�@��@JZ7�_�K�|��}�Z�Gu�?�\�&�N;{ _��K2�!���9Bc����вK���29�хf�d��<\/����f�P�4�������q���}�e�cp��U7�za�}7�T{���r>�����k���Fu	]h��xM�g=p%��nqG� �����c1���X�K�a��aë��?	����h��u���r�ڿ�'�ɂ�q���p_��J��]���/��*de�XlxVHYEB     400     110"@�:Д��m��]��D�b�B"�)���#��"��W���{xdz����zA�L����f@��.�G@�95��./���(�Vpq�b��1D���l�l�.�5<��_��:(:�]��o�y��"\������n/]���߾�i���,&��Y
3Xtn�n�@%a|�Z���1(�>�/$%Zx�8O�фe�)���-�q���FQ���t�r�F�D?Ģw���k��d1���H���B��B/~��Ԛ��!�@a��W9ΘrzXlxVHYEB     400     120�ř��tW��"� F��L ��u8P�q�&^�p�z�"cq�#W�-Afx�߇�T�������!�lU���S�}ʊ]�D~�PCa�V�6�;����쨳%��=4k�t�z��8K���sOw.�O1Q�o�!��>L��8���%�tni����@� �4@>K�˙�<FSƪ���]�Л� ]�*�v6J���C5�?w���ozC.oH�6'~��QE�w%6m���3P� ��
Q� �L�6��+�m��_��g�}_�<,R�|��d���4���:�+�1s��XlxVHYEB     400     140P�!�5�5��<�߃1ȃ>e��	�U�7c������w�q�� ��jN�.�%�����^�֎m�m�nj�xD�j[�H��c̑�����s��÷�*��)���U��@��>7{Θ��f��RMUY������Y��о}��n��;_B�Ö��(���R/׸�w�+]�<�j�Q�%������bzS���J�h� �/����:�#�h��禜��p:���~᪳��H}7�o���Yx1%�t�i�P%Xub���)c��g[�N�V0�d�Ĉ\?][|�L�C p�����$\Qq�!J~�@��T����SP����XlxVHYEB     400     150͠�:c��iu�V��:�Qb��d�V��X��@W����ں�K��E *Z����c�͊���@��'	�6Gpa	F%OR�tbo&ݫ׵ٱ����~:	v�9�(�N��R4]$SŅi(}�{+ϳ��T2A�5�!�h?����;�?��������i|/���P�	���{�l����Q���;�@�GѾ�}��I�M0Stj���4����������z4i���(��j�����
�4�|`��u��N�b�P�'��=7H�����BG���i��c���,���T5�����/1���ar���&����?���Īu4�������Sp�c�XlxVHYEB     400     140P�7��;|%Ӣ�d]�(�!B��а��fصt3�d��J�*-��+�n���Μey.�0kg��wW�;hF�%3aĎ�����SxEV��Ʃ���h0�q4��۲����qi�F��o٥,��P$�
��w��4a�����`[л�G�,G�=pl^���������Hwx�_�9�)�(M�d�^}'�#��ښ�X;f��N�<����-�A�c� �=d�@����v��ZP�R�fwr��`�;���V)�����]m�ғ��\Ԑ8�C~��$�I��sj�pOT0����ٻ��1���N� b��� �XlxVHYEB     400     100y�j��������`�,s�%���{�r�m����[�Pwe�O_�qT(Z��@X����_D��@k`G��/�1�� D���V�우Rhl�p��[��b��qA���x�]m�X�7*�jL��
� p�U/va��
J��K�|�
�B�����[�����^���������-���:��(�! k�m8q�A�����E0�����L�m�X�0l��Δx�2�)�Ip8� �L��)�M"�������!EXlxVHYEB     400      e0��0�t�h�KH&:�բ�-��N���4�������M���ȝW�ԁ�ϰ�p���慐�(��ڎ*�46�NS���Z�Y���cfh�
�볌fa��Uq�ƉȮ.#Sq��������O�0��/����b A��]M�G�+���zAĞ�kB�߮�Y�-E�|�_�����ѮO��fd�.�w�:&.����.X�x�0w���KL^v��j��XlxVHYEB     400      e0�Ѓ�K�/�FԂ�	�9F�&��5&�Tz�N��S�<���|���7Ζ��ea����=CY�!D���~4�����nQLPŒ�Α�S�	�g�� �������^o6�퐝�V��b�����T�������@���,19>���p�X�42���Ȟ�q��sz���}�o�����f�@�U�(=Qc�%�$��8�"w�i�6ty�j��� 3��a8XlxVHYEB     400      e0:���ˬ��b'I�"�]�+��\w�zX��[�o�eYX/�$�W��"hPe����g�a���?�����l�1TI|���e��;ј6�TK<v^�ff<8�+�c��C�Q����qW�}���P|�����Ȧ~��+c�ɱB�i��ꔕ�Z�3�F��{�OE�q��! ���ԧw��oIq�3�����R ��R\s��_p!b4~F�d>S5QXlxVHYEB     400      e0-5�xh�}��ɲҔKwt���˕c�ʖ��AX���w�eTp���{��,C��(�S� n�4YS�_���ֳ�_e�K@f��-��m6�w����(މ%�L�5�pV.�Ѐ�n�2��<[��V����KIt{1F��d\��aeŎ�Y�S����
���g�i�i7j�:����X�P��A�{9k�w����BH�1�@��y*.�(ۚM�XlxVHYEB     400      e0I�?k�e��yۺգ��4��|��l�խ���om{V�G�V�=�S���\[��%�YI��Uq O�&�Y�2@�)��}M�p�b������3a�wR��w]�2,��O�MZs�����r7E!nZ�˖{�g�c����BԀ��,���ྲྀ�d��@�~��+�tؐ,8L�O�� 6�V��k�q�F�e��ӣk��Sz��1;I븞�{������iO�0XlxVHYEB     400      e0)TPy�������W�P�L��˭�(��.?tθRs�;��[�e�3⤩��؈'�S�i��*�#���tQh����G�L��h��Rfn7�u��N#��a���i��
?���I����Q��yNQ�W�ȝ9���T���=٥l��»w=�ϴ��ۉ,j}Ϗ�wwL�O��I�����s������2 �g��
��acZ�r;��~<�}�XlxVHYEB     400     1c0,R&D�
��h=)���!E�>������&K������Oi�K3���� 쨞��*��W�͡�����g�tbrucnkؒ�f�������D��ؗ�����ClI�>��ϓk}�dKa��UVѝ4tr�t$���.��K����U�]G{�\���ǵ�5
yY<��:�Z��BҶ������:��^�N��uޓ!��h�EI^�%0XF����E�v����$J@���oYf�وE��Ǡ�hX�:���Aϴ������B��RM�#{Df�ϩ���=kcQ/�Tt̊�HC��ЛTd{xEF��.R�"�EB�}��|�� ��'*f�wx�s�|�� }�@�(��I7�+�mF0_�׍?x��YT��uu�T�L��$yX�*D�e	�r��܃�U��Ot����6l���0"߇WG�oS�?�C�ݺ@v>�XlxVHYEB     400     130>��]~��"cZ�ƅ��wL]k�<��)�*{M�Ѳ>����E�@��Ox�CLzV����܌�_�N���q5�s�p)?��z%��hmE��.R1fŁ3�qd/�:Ԏ� R88��ZXW�7�+w�[��ze3{ǝ췷�5�/:2W�
��y��Dߕ}욺H�!\�W�,Q�O����Ykp�C�1ۃa!c3Yh~��(�*c���@�KF��+Uu]C���kl8����k�ܸ��P#l���eS�;Վ������g�6���鋝�I���a��V#�$AR.��#�6^�XlxVHYEB     400     100O��q�T��E����[��Ȭ秛癁I�d��pY�@�`�Q��[��9�����uZ��&�e�B�p���R<�{;1�y����ư�r����׈�$i���6��Hb[�B �N~�%�|�g�z?��9^�8M�cix⦇ ��6��T	c]�xNK�~���΄�Q���򫳲3���Byg�X놻QK�qw�r�Q�mn�ɋ�T�m�\����<ק�6=�3�����C耮�pV���-1��5XlxVHYEB     400      f0۵�~:9a�Y��e��5q/H�ݫq?��F���.��=F� b~���K�zt��E��tiYq�q�%��Ln����N\�6�Ø8^RV�8o�(!�y�tg��A�N �:ͥ{OZr�<'S"��l�i�Y�y9��e���Ǵ��P�5�4�<���/�t�˃��3<��J�K4Lcՠ(�y����ԁ��E����Q��U�K��*]��U5�OZ��MK�)ZI�X�B^F�T�XlxVHYEB     400     140H��-g�|D�$�-G���xW�k z�&$��[o��Jf�_7�OË����@�`�ڮÎ�˧�t�];�͎Q�������@ �ں��/CL;���L0�ƟB/Ͼ��AJ�$��<�a{��ld��d��r�3��3�Q񪈁-,��rK����@W�>�G�W���F�!��s��3��(�3��ˑa0 Z���le�����J��z��ـ��en��h߯�L�O��I x�����5��>�\��W~��`NH��d��>��[MAB=�LQ*�T<��~j�!�N����O�9���Ȯ��K��(9�=��B5��XlxVHYEB     400     150�$�7�6��̒Y��ȋ�ߐ�{�x^jG).z��d�G���`#�e���=��ԠH͙g߻��7�
'?�*ٳw���8������Pj��/8r��eՏ����OԆ�l��@��6��}�q��������Zp�r���D�-��B{Z�����c<�1ù�"C�����#�-�Ώ�6��|�����cB�ӬL��A�m%��"�s[�j��L�����0$8���ۉ�^G�S��Z+��=�!�5ܬ��(����u_1��' d�R-j�q�u�5�Vr�J�t¸��r��I����V#q���Y��/)bW@ ����$X7�nW�� XlxVHYEB     400     170�^�3H<N�R����0�77�����qot��=lq�-6�3�6i	�����wB�f6�]Q���	d�a��O�@��!拾�<��хA+��Q(H��PF�3���rxq��^���!��(�p�ַ׈��1�y�\��LșfV��iɢ6/�!����,��?"�뾀RC)!s�.��yEq�k��U�}5��M���}�O|n?Q�G��A��-��ݟ�q�4�H:'�<x��?���F�%��(9��P�\���8���7V��|Zc�؞�?f����Nf��.�{�Vo,��3��w� ���#<����}��ܹ���`H3�o�ܛ���~���T�%��n���՗#�
�XlxVHYEB     400     160��,qOM`[7ȕ<���4�ep��@���B��	づ4�1����5��ݾ�Yt
���Ú8B\���#����ڬ�S,(f0ɵ���}�p;��Bm�w1]���co��ۍ��&��gS��H��>V�I�d�~;L��ޏR��#z���oQ���I"�:��3�{����7�I|���K�(�<���n�)�[9�S�e�5؀uh������h�j!�M3�@P�v�җ8�9(��C6�VX�C��,I�:TNGIa��c�,2�)��K�Ҩ��c	^����0q<��.rM�'�Vf�m�T՜��2"ׄSۋ�CeR㤙8$3;�V���'��na���ڸ��zzn��oXlxVHYEB     400     180����~����*1z�|t��4�w�H+�Ѿ���0�X��iȾ�\^I�DL,[������;�Sd�� 0A#��(��L��d�VQB=�>jhLF���Dy��K��_t���o�6���s��%������xu������Y��Ŵ�7��N�V_=,_����8�q��u�ȫ�NĒ�(��J�u��d�9'e��L��2 ����;Tu41�]t�X�/�CO������ы�ɜ�Ύ�Ɲ��>,ƛ5�s���v�H�NO6 �|��+Zo�旣�3�92��U��1h��Un�5��	�6yhπ�l�q�-da���}Y��S"���pMrR�m��OGl f����Q+g�HX�9!�������/Uz�����0P��XlxVHYEB     400     100ԅz�x �ր �
1� ��m-��]~G4�I{$w�R�gV�]�Џ�᳿��7l5v�l�SIg��I���3D�:����)���c
` r�����B�V���w��LzWG�k���ֽ��zA"� �&��H�d.)��;C�Ǖ�VcK�ɷ�_3WL��P�f��Q�0ս]�G!�/�o9=���+���![sIjF4ڊw�el�����*�O@�[/U��i�'�i��!��I�Aͬ����CV���f�/��XlxVHYEB     400     160�ف~g<��Eh��#�ٜ^R�N�vϬ�(s4k{!�^x���u��A��N����3�ԒC/W�̶���$�h6�+x��\2Ԡ���%*l~��}8�������)顎,���&��F�v�i�E�ES@P���\^|܂�CBR}��|,+.�(�O��M�+��~]�ى��H��f�A��_�L_c�Yg�D���Z����\4��@x�%e
͚�2����2�2d�Ə~���Nn�7L�CS�?/��3��,Q��K#h,ݑ Ń>&eLOi����H4.��5щph�A���ʕ���hj/"��^�{a`�°��g.u��f��������>rMN��29�fXlxVHYEB     400     160Ua=��{؎ERTY�̵�����G�&�-ԫ�)�^`b ��k����F���5Q��Q&0�زL7��x�m�`n�N��UM��v�U9B7%��9W�K.�Xٝ5���R~3TA��V9��l��ܾtw��������W�h�R��tD�5�m������e	�L ���������R�;�9J/�\^���I�E�G�%�$�R-��+�S_��6*��C�m��oe�̱i�\��va���rA�~�Ǐ8�2��Sk�1z����/���6�'UL�D]*�Ձ4�:�֘C�XHݧ�%~\��.Hc���c�$O��� ���e+�ސ4v�ݙA��2���h��yXlxVHYEB     400     140���7��YBm.��il#VxeS���R�|�x� BOa�t���̴�d�	EL埧Iȗ�P�(ޭ�K��j#��;����><��t��FKfE�|Tm��yx��Z�T��uA�;�[P�_�
ݎ�@�'�s��T��[ [I�:Ό����eц�|�-n҂ö��5	[�n���xM�R1��s��՞=��Do�K��%���7_�}iQ4���gc�]}�I�d�v�:T몡�Z���]�{��5�X�@��hg�)��H�X���Ǖ�WԢ8@d��H�b�2�r,�MK�9�F����\�g�XlxVHYEB     400     180w�)�S��l�d�M���g��~w��V�S�)�IJ����NW��m���um_��9�;�אi]J�2,az屧�������.�ک�4�5�8q����1o�1Tķ{���T�RG�Y�|LD'�^��y|�-��8M7��B��-n[����L������[��w|�v&		���96)\������`�k�ld��#^p��� a����Q'�#}O� ��ϲ|w�K�YXٍ�昇$__1���fZ�=S�)6�m���h�ᯐ���Щ=wЁ�8�/&���J�[)�m�A7�����m���AY9	��K(?�ʲ����$�%���h��W�g�Pv�-�����+�����Qm|�y�r�ݕ��ciIXlxVHYEB     400     140}���$�%_�=,րh�V��
���ǿ)B �v$0�K9QxU�l.��.���B�U#y�{��=Q\�D����yt��~��ܫd��J�2����V�!�\���z��CëD��]�t��{Ge�n����C5�*z���+�$��kP��2��v�"4P�A�Ұ��e�dϺ��C�0�R5B�N�����f��I�YC�]M�l&��cT����#ꍒ��0�3�T�}T=n�$�PU�I���R̙�	�c�3L7�,X�B.�m3plX=^�.��ô�߽>�b�4B�g�r�a��`��⒏�~��s�'��`���[�_XlxVHYEB     400     140r�ך<��6u�I��A/q7�$O�y��x驀L�q#�����pHx�/�|A;M���Zs����߶˛%3��+]�`�Ы��9�a'|t^N"�/�%���WdLK�]��G����dʹF�i!��J�s��M@m���Q��*�'�td�{~~/�|ȝj��$���l5wٍ��H�gǣb����h��?���L���&��1:*�Э�i�&z�qw��A̢��(�@�3������߮�*�@��,+� �n�Ѱ�x������Y[�u�!ZX?>��2Ʊ;���+ѭ�~h~���N��]�~zQ�}�'��_��n�XlxVHYEB     400     130�u���R������5?�h��]N�b���1W<����&����DsMUU�'-�e��P��x���T����$X��g����A�i��Tc�%vK�pc̖�l�a�Nx�߱0X��<��֎��VH��6��[��m֧>1��BT�6Λ2E�ԐF��Yם�:{dn?z���|�Q�`5������4��,�_a����3�C��X�����L7�]�"@��3�b5���D���
�j҅W`UD��*NyR�MX�u	�m�y�����j-O�7@��?���2��p|`���1��r��6XlxVHYEB     400     170Zz7}pۍ��Gp�3���@/�w�HH��/�wM:��O>% �eC�݉l��ӌ&%[�s�H��
Pd�nX�����c�����SW6����� �?��9�/�Y�c�� �*:0�!\�R�;ۚ�G��1$�,#�W�z6�s�`�v����`��5bg-4���mf�q��I��$������xXS��Ho�>��p��4F<�Tg��:�V ��C�G�G���L~<4+���"ќ.�����=Q]���H�d3��&鱼v�o?�
lB0�	߫h���/��qT��b���F`u���ў0���_ש��=�f=`�C�;�d	�<����2��
h���2��XlxVHYEB     400     170������Z�̅��Mi���H�i5�����T��M���]R��Ʀ.Ҧ�!�$��h^/A\+���q��%�pPNh��X���<�@ �eɀ�^�a�����ɀ�nڦ;���5�ͭ�~��m�����1"�#0�h�fMJ%�JA�J�e�e���)m홠���.M<sr�<��-�	�f�fK���fx ���m�̸1|A��=�>R5#T;�;���F5��ҙ�	\�D�]C��NW+����ۤm �h}��B�^��S�j Y�s�u4A�I���˺k��jB��ِoaᲙ�*�X?�)/q���p�/����A����r��da�C�B�S�ņ��cw,"!��Ι�14XlxVHYEB     400     190 �����!Y6ۦ��Vp��>H�u�I}��K�ڿ�pp��)��G�=>GM�z�R[@-ʐ>�H����t��`P���~0��ó8&�ߚ�>�v9i��[��q*����#����-�\ܧM0�8V���iC}���n ��o�Z�0���嵈C�x��]��T�e�VzߴfI��=�S �u��ŽZ	nʯ?����6K�?�f��*D7P3N���31�/6p��6֪\��0o%)����N� d�`��K�����WD��ݒO� ���˯��$�&�N/M���Х��'垎��T2޻sLgr5$�:yK���q=L���)$X�b4`@��f��֭M��$�E��8�"�22���}
����(����sNk�(�d����XlxVHYEB     400     150["��s��=($RU�]؟����?��m�m�g��dȽ]9<��ݗ��jo��s@C��"EQf��Fs�#�v{JN�w2H��0(ԑ�km0���{>E����l��"Kj�:,4V^��[Qv[�{rI���O�̷q?U�|�O��\s{F(���:"A����xDF�;\��9���(��+u& lա>�4)�Jd	�#�s�[!i�9��g��K�y^a��yf�t��pBF���Y�A5�C��-�=�v���!�Uܗ�K�a�Xܠ� g�I��.�ݩ>�h��6=���>`SV#�y�,D�.�Wb�`�W�"˟�0��� 6�qLXlxVHYEB     400     150�+�7(P�[d���WۘaZs��@o�ı��� �{ǆ�$���N����V����%�W�.O�r�� 5�g��=pT��7��Ч��9{�t��)cZ�mdL��A|�E�Ц|4LA8�
�(�`͡1�3�d��}c��-d�I�+���5�9��p&���朧�8��*�t)��T���[߄�rݿ_ւS���D�c;�ܞ�DbwÌ�%���%f�$�v-�H���WA5t�Yؘ-]�5�U@ڃ<�juϲ$�V�<�V'��v�W^
�U�1��ܸϲ�$��Wu*W7T�Lp�E/r���e���n��y�����?����XlxVHYEB     400     160sͣA�n�����Z�80kM����4�)�����0҅33h9+�D�ߍ�ЮU�;ܖb�� �UFa�`%���1��#F��]��H��,���N�/����z�5fa)���!H?g�{�W<�B�#�L�|��<���q�����VP(x���+��ސ�-����m@����ٞ�Vw�ZVI� ����װ���z�{S#+.	T��U�."|�%�#�ȡ�4����Y���
M_����9�*m����5��t,�λ��:D�4l�%Vw�w���)�d��f��(Z��g�\��6 ���%X��#�vv�?4Y�|9?en�Z��5rȪ��^m,�e_�S�6�:8�XlxVHYEB     400     140����.^�T��4p�FF�$�y�%n��@�N�H��/�xA��-p����;Q؏~������-)e�����n�Tva&��M���!��J�ď��r��[y	"�C�=m?#/����)L�ѭ��&���dN��8�[�w�����A���J�]�a�p��(: �S�D�W���4� �?��*01�S�0��H�����)��G��;��\��(澹B0��~$�&���If�L.����,h҅���Nk���!�}�����'.;��̏�ICI�;,����)n`�W vټ��&r
+�2�c��+ttj�#�QoXlxVHYEB     400     170	$lK��2O��f)҇����ayMr_�s��aQ��n��
Xm�J����+��r�E��~ݳ	��A�˹M�>��m��#��'$�]0�^�7ẋ/C�
�.�C��gH��eWo��G
���H'���^^j�q�$@�0�`��D���3mЬD����%��3"am��}FA�N��(Kow��k��$���j_���f�T��[ �)��!d�g�(�2S�gt_DpD�r�RD�8����g�7s�9�[�>0Q�yI
v!�pQ9�����g�Z*Z�`�|�J�hh���)��f1-�ߏ��͝-W\v�i��Y��9>}�
�4�5
����v�=���V���x�G>\M�m��uۿ-�ℾ�1owXlxVHYEB     400     150�ܣ�M�A�BĔx[tv�	v��i��>�u�1�V�!�8�u��{�#�̻2a��H�2E�*�~D���q��.�ϫ�������J15cz�8��*1є�+��ܾ�Pi�z7�pS���pe�������
Jex܇��>�b�� *թ'���p�"5���Cjl�a���4pC��8Y�������u��#ɀs�$���u�.FE�������I۫#��FP9�.��Ʌ��gzB����"��B�x��9����}�/�l2a�����b.�SgE:'�{�@�ښ��F?q���Q(�?s巊)�<�G|t���\�ﭘo�$Z���XlxVHYEB     400     110"�IN�(`΄�06V�1���~���C��׸O"���M������N&�rЦa�!Z�����i��f� È�(���pcb}�ގ2��_,9��pu��%��zS�����Ӏ m�W���Ѡ
�Lf=*x�[�� 2�¶ ����hW��ɢ�oK"�*�y�JHo�[=A����A����@Bk�� �%hF!��9�ϛc>U���z�3!�	��(,{:q/(�`���V/Ł����Ш�H^�P�9��|����_�HXlxVHYEB     400     150�C���ti����.��T��h����*�D$��*x+i@>�[�]���G��1�� �P��,�Q���VSZ5�;���U�oWU% I��}�m*&�g�3c���Ty�ܞ#v&w���iX��F��R���fw��r�D�z�b�^H Ōr�"��ʞڅK��sb����"^��w��\�7��<|SӼT=�jJ������9�}��oh��}���%�Ak��������q�=0������ib��F���2934EѾCqCCoa��Cm�Ix��� ����Z�],4��F�W{�K���
��3�i�̔׌��p�]I�XlxVHYEB     400     1a0�!���\M�WŏK�%xp����9�˄V+�Wm���$��o���ϝN�t��4�Fy���RMFz��nqb�� {����a��Nd���~��y�����g�F�A�����#��)!�g�4�DZ��t*�-a��+��B�ED���������9�>%���R��Rh�#^�o�O�������^ڮ�#�!�E��6�L�Pz-0n6�)��C�/��M!�qDsܡ0F�A�9�#���sf����'���4z�k�>X�;bBhD�7����S�R��c���Q4N�������8 $@��/e�ҭ잢Ы����	�XW\���	+�)�Y�G�%F)��p�f�Җ�^q	a��w�;�j���g��QXC���[/y�FՑ�pbؔ��#Y��ws�8���E.,�R�XlxVHYEB     400     130z�&�(��x�7sv�7:�$\���J�@�5��Ơ��H�b�r��̱��C�֛��ե��%�۞�Uw4w�H_���H
"9X{i߱�;�¹��� ��%u[* �t�G�Jyˎ�g5{�(l�ꄬ��/􂧑ѡm�c�ʛ�RVq/���7Xka����Z/���eMɂ�+��v@0>�s��d�:�|�t���4V�#b�������To��@��m�1\��*))q�"��ޢ�cj�V�C�O9�<tѨm�U�r�4L?��H��=����b�Q
���nx�Q~����x�HUXlxVHYEB     400     1209BK�(�@r�G}l��F���Eq$4����7?�9����
��ls���ؓ���	41��n�A�9�[��C}�SV8���[� ��/�����T���C�q�w9��r����/vsk�e�����ǔ���ϼ����c�s*�$N�w�B���7���أN��C�%���Ғ���N��Mz!��ɓ5�Y�F/��7+�3�E��?0�ʅLv��<��W�wmE(�b�����K,Ǖۉc���&.�&4���UO�n�+�Ux�zRٙ��i���ݨ��h�XlxVHYEB     400     170>�1���Yd����ŹW��(q#�Sdj�м�k���Z�;ZrA��A���4�2���֝�g��HŲC����e\Fes�V��$q��sqb�S�����o%��S9H�AQ�Dɐ�,��P��0���]�1��Yv\�AeX��L�}�ny�5|����r �/s9'�x����tWv��D�-�>ik�r�b\�;��M�� ,/I�e�&㥶�W�#,��#�=���4��8�F�#���h�E�����O���Kj�PP~����@����˵�o���2l}b��
���|�U�Jq�I����6���0��h�ǧ��#�^�Mz����5���*��A�J �n�.�U�5U�9��+����N�XlxVHYEB     400     160����~�.��iJʁ��n+(��6g��װ�ḛI5��Gչo�����BOk_.|��Gs�~��8G��eq�jv�/MX�^R���R���{�ͤoo:�&#�!�y���!��<�#������z�/\�/�|qL��an~����F "�Bc`�;\Tp���:�����rB�ˢ4v��/��}�PFM}t����_1�[,WB��֙x87~�4>���:��/��~X xa\��(p�
h2��?��%~��ȂA���I��/���j;C��9���'�'ï���hx��o��lVEl�
7���X����%�2�3Yr1�~XB�+�����к/s��	��XlxVHYEB     206      e0-��X������&��:�������O��`����g���
Oġ��=�3�X��
��x{���rS�A��>�ٯe��2��;-���u+�U[J�o�"���\�<2�τ��[��S���&��!k@�w�����uD.`�.��yk�/�"ͣ���:��`���`WB�>�ͪg�	�~�h���v��g�֥���>���HE�4}̥k}~OO�VC