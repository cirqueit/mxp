XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9h�!�yO�- ����F>(�5�#����Ɇk���R<6����֪ ��>��a�a��;c�4��l��aӿ������~����vY[l����;\�mL�d^��{Bo�+�K}u���h�(d��j�%F�y�OoD�uLo�QY0e���~�{���C%Z��|J�t��ڢ��{�K��,�".>�^� �����S�`�I�<��o����0d��������]ф�# m�N��CEysKHǉne�d]:�����f��l�n��Fs���6f>+�J:�$��v�f1v�득zb�<��P�R�8<�t�������&L�IAו��M�`��z&�ݿ	��S�[V(�
�9�������1��g��+��<�>^
��ܭ`���C�٫��}��.bD{nX�PBW>(r�ݕ�4I����|t��7�D&;������hR��.k4��Oҹ&X��R^B���,������/{=f��$f��j.P�bA��4��t�
)��0'HPfrdHkGǱ��o����;��M�I�K\4�d��v���{~V� ��K.ک���1��Eڪ��M��0�����$����u%LU%{"j��:�k<Kv����9�r-����z� ���V�Q�ۏ�9�C��M�rD������;Nr8^r<6⇥�s��Kn���ҭ�9 �/�!ض�_D��@���Y6���nޫ%�W��7*��p�"U�>�� �2��77������� ��g��W�x+�O��H�XlxVHYEB     400     1a0�w��5�}ZN��-�'�\w�"��Ŷ�Utu��7��0��P9Tm5�k	��+�E�w��ɒe�}n��`�x�j��ʶ�(x˻�(�=��#S}��H\�a���&s���"r����m6n������'H586}�:o�?J��<�g+~(���f����1���z/v�f
i~�K�5�/x��5�t��cQ���D%mS�[�4�H�O�D��W \rT�<B�oS��{�F��)�n&5������0w��G̨人JX�6+=uU��I�3��]v(����p_��}�C�JQ�a�ӟ0�%��}��Sy�ܫfͬ���i�������T&�l�����hѦ�z��0cb��<��Ԟ��"W%�~�Exvg����%�����$Kc�vX�CCs��⧈��XlxVHYEB     400      f0L�u��/���ǌA�Fuq��Bh�Ĉ��14��:�+o�8�8pɬG`K���:�Q��"�@g.��dέu뉿qi{�)DkIn�]��t���b�%MYbq�^7��O�Y��̗�sQYE��.�됀�1`��A`V섛�=+���i,B}"���E	p��gߎr�j����3�_���n5hm����໗��/��%r;3�m���D��\�"S�k\����t/9K����=�cXlxVHYEB     400     180��Ռ�(xY�!i�"���X$l��yz�.�1 ��B|�]�ː�2�`������Q���=ZY�����i��*�b��ЏPSc+�yJ�Zc����4���-].���oG�MB���>��,��:�g�(`�f��A2}*L��_k�j8�u�U� Q��pn|[��H9Y��%L���u|��I�F��62NW&PV��S������� Hr�6�DV�W��,މr��	��7|H[�V*܆�ot����t��;}�����D�vEj��9��I��-0����L� P~Μ,
�z�X�>�X��&���gV�ߺ�۟3A�L��sr��A5�z�9v"*-�.��*�h��P|���%ӊ���xO�_I�����Hj[w T�U�XlxVHYEB     400     230���)��/3P��E�t>���kq�⺑�6�x�m�sk:�h�ݥny2up.�\w:d�ƐH�d�|�]��*�.�nX�)VNşZ�^�P���Ó��Hm�3�|Z���i�]�~�[q��Gk��w�o1a7���:֣��E�`�|�W%��]�ֳ˰�uE�9�A�p�B�ω�*�s{�Hں���¨�MѪG�m�&��12h܈��3��@e�Ea*̽x�Q�XeBe|���G@\;(q'������@\Or��I�M怸Pf�&�
�%�RTJ~�M�y�V�<����Uo:��6Pt�cR�"����H
�U�I5
��k����`�\5fn��P%��D��K�r�����}{��\���"�¬��Q'v/��hM!'�vQƉ�=S�V�f\��5t�N��FX���T%�ڬ�����ݽ46�� �q?�Lz�-�p|�W��x����}�������U�ŝ;m�@/C���F�i�_7��� ��1�Y叙6A5q�>�l��o�~���#�#g�� O{��L@qXlxVHYEB     400     1c0ȶ���tZ�"�XTt�C�*��OeL�y���c�F��7s�W���?�p�a�V�+�ʩ�m��Tk�?7�\f�kZ�p��9��QL+�x��bJ"�-ł��������ʤY'���[!��F�k�n5M�"�[Ku��/�Sߵs)�����o���6kK\@�����GwX�צ&Z��M����U���`�1�9�/V�:���㛨����C��d�c[����p�����}1��i���ؘ�y���RY���vsH�>P�]}�T
g�<�<�>�kz��K��ه�]]c��T:�9č1��b�G7�[	�F$��T�&S�-'5P�ER�Q������N��M�,7N�<�*���>j���� u���@�'�x0�kG�7:o�>�w0���:w�X77WJ6o\TԮ+��_� ~�f��ۍA^>����XlxVHYEB     400     1a0צ�ei~�}����m+'�e��N�A֛싍��EX�lƸ����0���T�~��M���s�6Z�#�(|ӛ'}^g��}�L������M��*��4Il��?�8��"8@��Q�Bj�:2��5��\|N�J�ܹ����,�����5KH�\�b�47�<�d4D�̏���p�L?�'��NK��r$ve�L�p1\	�C��?�3@�b:\�����v�E�c������������6��,�Bj
������#�FJ�r�w��!N��?p���Dꡚͻ�%�㘹.�g��=�TswJ��W�\�t��ѹ�x�N��j�J9|�ƈ�1fw�P/=GV�H�}$4�˻eM��1��)��#�KF��ɷ�%A�7��P��〵�Z���|_�g|�7p��,�NXlxVHYEB     400     1a0.N���g�����oh|_������õ"u�~dJ��u�Kɀ�Z9��o�^�րW�փ24�|�S�K�0j
�K`.��ZE�u&�����Zvl�(P�)�}ӊ��	t}q`wlz6�Ҽ���q���7v뜠.>)�������>I��xi��٫m"�6��{���~ϼ�-:�1�B�Xo�W(A-�<���-��R�`iO�<�N��b���}��Qo����C,�n������y� sz$�'�	:7d�
�e0q&>6�޵\�n�%�®�l�*&��4T�1��)��$��� `ݤ���>�d 2<��Q�m��ph0qP������Woq�f��k._oJ*a}�s��fQu�B&���A��/v$����z��o��׉����*���E��א/d���XlxVHYEB     400     1b0������P 0Rɞ�X!'��x.ɟuQ耓X�T��cy'eB�r���5kOfnp���f�=��K��8��+Վ��4^��Kg��-˼^��:yNz�ml�6t�Y�f�LJ>�ٛ�:�h� �>:��-T�����"�H�a���Fu�6�h]��ܨ�}�|Ѿ�L����8E�Sn1�vu4dQ�[ ����,�K*#&;t{Bh��qx�dEk�8F�+]t�f�.��l}�m���4wA�;Z�W�*��g��ka��rsw�jό|y��'F���P�"�z8�1�����"@�oi�t�Pv����@G@a%)�!DP��-���j��4��9�Ⱥ����P��� M��t�I@��0�o��*Jp�0�Œc�����J�	P��,�dE�z���L�����2�J���A��T�XlxVHYEB     400     1e0����'WC���?�.G�LZ�!�Ō��8�8����`�Ә�5e�cX+n���k���j%(�mԸvɁ��UGiN�X�m���A�]	n#�Z�<	p���Q��s�>��z1T��������g��s��s#���� *�,,��e���w���W�FG�{cn��� W�YY�	=J]u�,ǈ5�>�~��)� fȅ@�>�6@	�/Z��̘v��3��u-�
ফ_�-��^S_��*3����	�`��qȔ�3�!�Ow^K_�� T�޷�]��*v���{�#����s� F��}4�Ku0��p�Y��>�ā�؉J.�ɉ����-x/R����P�W��r�߄���J�^����'}S0NÙ~�`�Q��]r]�1���3�A�ݷ���PX+F�P,�g�ߑ�cUrH.S:��q�1Х��R�O����Z?)��x�,M����:6�?�W<U��=���}�yoXlxVHYEB     400     170��:��_�_���\xי�Y���y���I�3���Ek��ʀ������{�����K��@�P���O����u�%���]�RnpfF �T �s"�W�u?��o}�S����a� ~��(]�M'�y�JoM����12�|{��~%h����djo`DG6JQ��6�A.�'��ذ_�A���~�뀉������{h�zJ�@:��vf�
���w�C�Q�(`�D	�p*� �^�r�UDFۮʨ��a 6��̵��d&|�:C��u����K�0����8��3�Q�	��牺h�
}�����.���/�Ѣ��h�k3�����h[-ԦV���0��J��({�X{�(-#���9������XlxVHYEB     400     140y!Ԟ�8�^��7Pݎn�QѨ���Q����l���:Fi�ͷi̿>����N� ���Ųj]zBo�fc����l�9�Z�y~����E�����X9G����?��&#�I�7_#�q"�e���Y��n�&|��It�b��qP�S�8�ݽ4�jB�BJ�A��Y�C����n�$��k@]��I��+!^w�@b� �׮

����j����A��4����2-�hpt�Wg�6w�A�"lj��v��u�贷����{� �*	:Y)��^�6�Ǵ;��b��~Q,ݻ�9
|^F�_,�z��#�E$
��FXlxVHYEB     400     140��.b�9�����7���g`���!Y�].�e�[H�Rk>�fڜ�6��_ 0��Oefōw���i�����e�����k�N�3{�'cOc�jzts&5;P?�@!����ڔ�cT��yj�D��d\��J�`�٩��1M�Ⱥ��U�z�s�mv9���8����OԧX,C������<Y�hj�����.��6CG�bw�b�l�o�e��/(C����Os���e�y]'=D�-Y, �� 
rާ ����N��0/�:�m�?-�� n�zj�Q�9�^������-jԭ̳��b5�=��3�vF��H��=XlxVHYEB     400     180B��p�,_Z�i��*%���Du����ztG=���Y$��F���v�x�V��癅�`���[N����lf���+f��r��!ؓ�a�>M��(o��r���yv�������3;�#4��f������WpO�|3���F 	(U�4c(��+���m�}ܼ��\sG����"�_GOXf@��JaaZ.���A܋v�+�Y"�����)�̮�7���������]��=�5�W�\~�mu��2�P��<��B��O� 2�g}�dLETG���K8���D�b�rM�.,�l-_���=�q�����������_���*�j��Ư5���h`_����A	�gR���*�~�8J%� �T�T �<�?</�T7XlxVHYEB     400     180�:�2���y�gr|1T�$��3�������+D>d�2�K1����6��h���߃��wi�#�{�,�%�4�ZÒobA�Ц�O�5��du�c�A�8�X���E�nW�	Ʉv>�҄�$ ǝ�~�Wx@��x���X6�>����o��P��L�h���/�j����pp+�X���03����rb�]��ҟZF}�7o��O5&,)�f��;�Pn5n�i#tf��3�1q71[ۢ��+�u7���ǡ`�7���̚�\�g^|�������RT���X\2�YBRn�������u���R������Q���k�͋A�Vٿ:R��pvD��i\4���Ąi��@�>�����Ã�e��)�q֌��+𮄃���<��XlxVHYEB     400     180|��Y��"5hx�u��\ͤ>.�Ŕ���ءd��&�~�!���V�8Q���o�?5�B�K���!W	 e�b��¾e����_w���[fW����4���Y��8�CV�䪣&A ��qpZv:�T��H�A-ڔ<�_o����58w$�4�n�LK��N�5 g�F'+w浆)��GFj�YUo��a2m�:������L��쌼�Dk*�ו��i�Btw�o)A!�ȳ�>O�y9����p|�(�Q(uHa� b%~ �	+^��քpU��BF~FP���a���9���X���f@���-&��=��ZON����*� ��ά�C����GBTtv!�R�)���9RK�����h픶��K�8I�	}�!I%ay�]��؂"��XlxVHYEB     400     1a0~�ՃsW��&�jB�8�=���E^q$���o�6����d��P��?"�����,�@EB��|�A9N<�lO�.T�6oƐH!���0$�(dD_ �D�r�@J0�J�\mơ�:=q�.�v+h|����*F�[��v����Z���2A��j���;!�����V3P�W��ֲ=��i���c
����w��j�$�����ք����{�����$ϝ(
,F<�NE>)ޥ��WVz�����7ߦ��pt������4�����_��i�)4�sQb!���X�ow.!����o��qH�ʝIN�lG��g������34�!�����n�I�ď�ږ�z��"Yw��߭�2(��7���Y�W$+oy�� �)��>�ϓ��瀷{�
l���)�1������XlxVHYEB     400     1a06og�'V�{8%t���|��U����!���i�#�.Q���< ����p~�	���b�$>�i&���f�e`3��N�uU1Ha�=����&qXR�
?�άȍ+������VM�![��nk/����]O���%�e&ks���.�Y�������]Y'1�}�򽓷m��Q��]�����y�Q��A�w���)���ĩ�?t2FK���w����Vj�~�N=\z����<t�bٞ��h�� �z�%v���
�7�<Z�;o�a¡y���=�������.Kf��ܸ�9#)�o8�k����R!X"7*���~5p����I�O� e�;z�,�^���V�੖	f� 0��!��p��a-������;�"�i�l3X�&)e���+�O�g?�&CdI�"Y��Y*�XlxVHYEB     22d     110Ű���g�p�+�r�i�z�A|2�M�����k��&a��t��R���%��^)0%eB����x��\�8[�M���������3�
�t�
y�psA��>/m֞��J���8P	�� ����4n���A^eb��ZmA�:�@�%5����\��tKc����"W~2{��z�m�мsħCH2�*��h�b��i�H)C�`��:r�����DIà�~��9̧�^?@��݄��-�0p�ƌVy�0�ɴb�>��E�д�w��@�