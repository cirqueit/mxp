`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
XxoB0UbvWFkLwUlk9sd0GTn08tvGpUPzyYGkTYbidRoXKaxK9UgsguI2slVmmIocDk3Ay5Q3Ylg4
RCj81jUjapLMdbRK26yORctd9NrNAIYxgTJOcmonGfYvccIhefMnnDWu4tlViZq/9tCDz1Pk1frV
bNzw0yovgXTGAPddg0iJ1mNpJSVOroPW6OB09Of4cAKW+0Ov0rq9GeBaFLr7C4bbaMZUGw7RVD92
u0GyxLPfMoJ91nCnyFT0DTunhAtUpb83Rw+pkWcCjA6wtSKyO6+m+XbDQ3owKPee46BlLd2c+GRw
+m/bdFBuukRc9UgKpv8vj4ojqREwdUgsTUQ4Vu83uf1bVFqh2t/WFz7XOy8rsGXu7iWit4Lvv8DA
ZLfeUmHDEVZCeTPYq7hLzLe7Dp/wrkNKPP5WtB9JzdOWFceB95k8UZHyqZrboz66y/J7+7qFsk7B
F6jNLiYu1ONuBUluJnNWAp6L8zofKoWu4OTZSUdicr79//LcgHm6Q9qkNKPyldub1tnAx8eh9YDF
ujBhA+7c2lsGUGrpJC2vXuGOhY30BKBeSUcUTsl5812R1tflBBBIbhNWOh36ZZejxy3ABf7edf4a
bclxgEfk8PQRMNm75OgE4zqf3vB3dpR4HPxhr71GHqI63pO4pw4/1kV+gr4+E/0MkenHUmr4Lj3i
FHYOySv/MR/c6Z+JAO7t1d+McskdT399tfJYPd3ZetPuCzJ2hDKcUGO4U0lSdhxtaAjwLo8fJLS7
E6hSx/dOAxZkKE6Piiwm7HFD6frgGyRe2QkLzZp760kqCT03IM4xod4uyWbHQok2EJA8ZC8jQQQo
YQ6FlPkqmM/Sl0/nl7rCQ5W+NpVq/b7fvMM4lWf+v7AASIxauqkps+0gROs9W75p9JYTK5JWrkQw
vq76JYsw+2jUzaWtBPBzdf2YO7pIZq/yJF2KNE9i8YFc0PBV9xIFNEXAJ7WXkRByqKy4al2DZ6sM
dLYsD38JaZC1VQByjq8FH3GcqLA8klg5+q9IRomWMr/ZGwHYk6oLwfSsqMMDSCavFKxfA6ZIXtN3
IlA0BEpuXJNdKcdkVlviqinKqijNgqBI2dEivI9nHmCkFbb4pcP8nyEdAwTPYS/jW34aKj3raurn
ZKzChBcU/BewicEUvZKUT7f+saCIcmsdwbn+8RGQQGsD08pTNsk7P9JB71fWiZUkSelQsffH2ekb
J0cCHEc6pYeqn168FMp80XxGq/+QAoQ+sdZT53MLMoxIZ4F1uEczBAng14DHarfn8I9TsePlfBdD
F2ZBDCNx4ARDYTHadvpVAYRNl7BpryWZg+lSCWdvBWr3AHxAQMJeXDMMHihm+vPBu+o28xThwRli
o6BMowmW+56Odp4KSzvNjXbIwOzTnWSaFeWxeNQkvsCbRRvyaWORK+at4lgu4sAoKGPiM3jEFrd1
PL6XqqldsKQFngBQRpundojc0iFBga4qTRmn3RmzY/r/uZrTYkai7vGkGicPcuL8npWQenDmaRLo
01rwLtIdzKK33z/qnJU64EzoSEnttpmY4N6KPtixm6kjenikwRu8EfKglQdbIWwgtKZ3lssJ0N5B
voWgyBlb8QcC60fdbMDTmOtdSbwpH9o8wCmvt8N/DepRDgI30GtH3vmNUs3EAkb1nZPqDj5OKOIM
fcwKU16QP7tlheeN+jp1sdhfU5mMY77UZEmNif/3o3sKPZkHFu8TEf8R0IH2haNpcmadPMRezaJR
zZCsBVYWW/9AjkT2PiCrcocsYSWA4AWZfbLm7/lnbx790N7ww3cNLAde3PCEZl5pqvkIA0VcAvGH
6BN+bF1FV/NDIAZTqTRaAYjmSot/Drs7p/l0Mi9YB55mEh/+HHy1jdY7FP2zLUC2Vowv6hCirA9M
C6pImoLI0eHGerzFtd50iREen/AWFccK9/SE4og5nCUhPZ/wC+9h2Zq0xmt1R3OJCzHP/ovsqcTA
7B/Cw8gPP5xfQsmTVEba1NPjH3VsmNRdrhkxKpqm/BDTviBuGA87b/dazRXw75gosXKWMG+lnXtu
lU2l5A+U9AdI/dKQ9fCFZwetHkts5DEKuIFhgDY9fMQveN98XeZlbSUzmfP97oUfZNRcA9NwxEd8
RjFjSnfQujAcd9Xi8tED/ZJ/s4Kl+BiKEuEAjag+XGuDptTR6Kjm5ytv1tf7Ij2JBRnkiICArX7X
q/Hr6BbQs7SM96F2CSc1Kz2QOwM8qBkoGbtNK8T6QrpXpFn43KvE9RKijEOpsKPYJeoURh/n2G6c
Jkw9EfltnqiJABjdRwQ7M6Xxemj0PiEGEpKya9dWfRZFwnDasY5MXu/rCp/Vd/EB3hl7OGDy5Yjh
zK1qLe6om5x1AYgMbnj/APP1qv6BfWVUbAkHbuDRMZi3+v8LuKJtxJatTgM0KKZckiYobubiabh3
Cy2NeNSpn2ymslqtlu4ohNnQ2Cc4CMxDNIgM25TvZwL3j68d9x0xXCGzEUT1Yebb+JcZlXCXxBZI
swmgzURfzhXsmnsWBb5hWwiaFUAZDYB5A5FyuTL/GrMEYFJjZ9HC2wMnFq7XacxoIWxfTbZ4coks
u5dzgkJITt21VuU591wwNqGcf9XIk0+D+47bLADqzu6F8yoKBk7s/EIBcKKvw96cUYus1HCEG/QQ
8Ud2hdSkP0Sbqq/MmpkZuTr6uYCupfaIwhDFUwsoJW2rp0on1l7KF/+Op86xzGXL/aFT4/I1HGzA
ptT0OFpFUHxMLXAKGEu5NHjWuYbkclh2KVvu4+RUjwun7ov13XuuX5dtecV684KtJt283vpoD4aI
Y+SCiLW2w1Eexg4fkXZmhg9H5StkZsbNxDx8RB1aPlyKmmAIhNlJYQUngl+AjRlsyD6KTk5Jwbhk
frOBLIVI6mXGXfD79eNslu4Wpq7iSfT2qnBntWo3IRGlQJIs8e9J9sLuTfnMs2g4DZeZ26ZJcrmQ
48LjrAgcU2cuJWwdcsUAHfG5ew8IgprufKLnHzvKZZbY+JEYubfA5YTS1GWHBcwOHbE9p1kaWtnb
qRa4Z15uuxRfBXsx/1Rc7fY9cRlyKP0NO9rq9NJWdXtZOns71B1mhjhnKG4Zye3RzV41bFm8QiS1
RU2b9e0ECzC8fVOK/AzP6i5YUXt5Rdk39K5KZ2QBApbnxA5bk5pqhQlKhZ/PiksDplmFyKw9kwxo
enVb8PlrBMAZ17eCMFSt479osNebrVIM22RAd3wcJxmSsqRWP7bQYl9CGkauJwBXzCXzJ0qM4DLb
sEXc7I3PvvKV8wzJ+Huj0QaBZpgnB1UwcQ2S+LDpU8UHegXDj1h7SNNacgq2XTBTpgJzYZPnkeei
gx/YrpiJ25L8FFc7kphG2G8+cNh8mOl7g2bcUoA4ZsMvpfHeBIgLFUbMxK3+x5LrHyS/uT2qpQME
7COT412/OPdOHZwjbs/15ugEjgiqO4v4upxq3ClZD0+rtY5oLAO4HG+vKy0QgW0iZAiGP4rAjSS1
hkLSiH9/1dzpoBgybUJP1agX2qXftZm99y9iaoJn+/ybm8i2DWlyVS+ip+iRDH4e531pSAFGFd57
yrR0WY1WTvaGI5JAJBoiJJdROSFpt8wdu+cIXe5V5Jbm7M3Gl4khqDo/zeYYiNCVtMx0YRTcuywL
Cg+nAQkU8y6ln8d5Vha0bIAePf1+r3+xmv+ppxpKX34eDCIKQOm6uHWmAbERlPgEKG2NbMNtnith
xYQzyZeJu4NSyJLOwJRhOWYrA//cKRkFJJpH96Bn9vR4d7+jx+ainSKmy7kKz1l8MoGDtrpvL7bb
jw58r+1rhjQhkteUXd4A+3AjOjy7ajNQeLeUA29yt62yI/Y3aRa39btBTTfnv5iM0LqML2CB8DDe
tPviL+gtgDHwNAbLmCy6g17P7/pEiYeY2FarpYdohYszkpO/MZUrGagCivQmy3bPs1U+w484H4kE
bvgmiooU6DCSH1XGYP1+WKwHq68z0n25udeIma+RHOEcGuc+hwzEpSBDjQpsifIzYXnciLLm5Dhl
YuzZBCX29NsSJ7xCx6MR8YXEo6xeK4lkgn1ynetRhgO3i20CHREL4EQNfmfur0rIjloKQSXCJAtv
clY2MHsUvYFOpTx8/LAz7onYBIiQnkwRxDOVuvh+FPXAfd15s/xIf9W/RsVp7JKQ6N8mgz3RMFNO
Mnjdgjm867HWkrTLTgbd1OIAqc/XWaCvKqMbApCNyW24
`protect end_protected
