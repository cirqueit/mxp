XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Zl<K�6*W�ޭD�s'qx����]p}!� ���O��1�w!݅ӓt~�WW��f��W�`Ky�C�po��vر����h$�y.�b�fþ�ȅ=tN��.d�t�ۨT�Il;��*�j?Ht7��~�-���(Y@Z|*k�� X��5�^[ZY���-ty��;�y{�>_O}&|����0fbL��<�͝cb[(�E�S���pE�F�[�$��$D���>�SNK��]��M��
*���͏F�y��ߠ�B�)"gz,�i��V��*`´��	������T��S��G�+��͹��������7�cJ"�:NѴ/v]w�1�*틙9�;Xֽ����MǮ� ͹,��?�&�;T����|� �U �	�:�PM�=�'�1��K	�ƆV���upS��0k�8 q��������h�����(��$o�֌�Gu	Q['�r��|<Ы��
ɋ���a�ki��p
�~ja���p�`�ˀ�%��p��N����F���z�۠{׋�oIuk����������l�~F��ET�[ꉅ%�0	3b��o!~Dz1�渄:�RM�����D�`���� ��'fI�R��s��Tg�h�a�G!;U¾�r�����0g̭�!�Ss� S��t�H��R���	5Ƹ���y��}M9
�^�
h��g�(SRِp6砅�U-ܚ0"�!�<����T6q_��r�w���b��]wC����� 3��A[�۠ކ��p��XlxVHYEB     400     1d0�g�a�AR>�oQ��h�#�=�X����,wV��;����i�������Y� -��R2uU��8k�%1d��$��]�tǵ�V;|򌌣��/��)ń]J|�e���p�+�l���D2��'i���� ]�v;j�ώ.fQv]vb������?��?BV�����>������0+�&��>��q�窨�h����אɊ�_A`@L�e�SoaTL�a-�\cX���8jI��L�-C�dIj�O��� 5IڤS���l.���û+j�榎�9��|�A��8z��n4�ꃛ�{��@��{�kI�mnIf'�i��L���M:O�؟̏Ѩ`�E����-g�S����ϔ�0�^f�.!^+Q@�6�1.��%�x���=�����`�W�V~Slq@r����rt8F�p��vh�^ '�!^ť��C� �#dB�9�(��;�=�7�N�`��_,�@�e�XlxVHYEB     400     170�[-�N�087(�_� |�i�/J�25�`�.������2��F\�G��n��͐#����#N�n�I�����i��vE:�����N�������i^6��e�k-.~R\�=[�@z���`����o�Z*	��`��gu�4Z�xq���l�>�qks��VN:�fD��Y�q�F|��i�Z�S�$b������K\���MiŢ���;Q���'(��N?��K1"BC��������yK����{�+��E��:�튳�O�Jm^�ו������S0%6�z$��YJ���	q����'cw��ԥk���9_�^���*W�e���ĩ�D�`�RM������n��'M����mC��8�L0̓�IrXlxVHYEB     400     120W����ҧS�n�)42.xw�1�پ!cwz��)˥����<��}���F{�RI�.wٌ��u��"T�V�J�<�+se�d�f�5sw��*�V޹��ոgX�Ad�8��E�'|�4����t��>\�5�&�f��Q�Y�*R<�=�i��:lb���>�iSB���6ѩku%0�ѫFmE�>e�I��t�Q���"W��r�@T�J�Ј�s=I���Ұ' R('<�k���;�Cf�z㦣�,]+�E�yp ��e����řj�һ�!@�]��E ��XlxVHYEB     400     170�"/4�uUBk슚��l��Q�1_�m(��DXh%�D@�y�+	K?@	��C?��ۜD�ײBض��g�	f���+�m�\� �������I�(c�mv�v����vrlgHk$H�#Gn��{�r�b�m>��f4&�v�!�
�-F��⭆�z�v_�"��4�V����_\��4����~}��t���g�� ��:L�q��-�"ǭ�3!sR텊n��C�6V��٬I�a'��_A�������V�-s��G��,��Z?�З^vIN��F��-����\�1!-��)��o_[WM(�oȽ��;�'/�y�����K�,fkQ���!��<�� O4R�Y)j�޿��±����}>XlxVHYEB     400     17005s�}||�����yW8��a$$��׊]���7LW,�VV�i�>\���[������y��I����D����Q�T����"a��(�����ͭ8��MF#��s�@��k}� 3�-<��_����a5��:�̃՜� $߮zc�w�6����"۲_�So䃃�#�Xyi�?$_�^��z�aT`U!���FL��s��@�u�j��[�>L8��ל�Gm5�a�f�7������a���#�ۀg``S�?&4��+:���-����Nk�U���u����ͷEkg�嚪��*X�g�f�PTN�	8a�L!?[dh@ӵ˦��N(����E��P�x,���M���7��eH3�u"#G#,���>���XlxVHYEB     400     140E�:��ha���Ӏ���N��7�3܁�^�CF����vNu�{EIS�2C���v�pD-[�^7B�s�um���������2��'�IwS�*�h�4}�.�CM&�l���!t}�Tu�&��F��Ҡ��bP3+B�'���g�1)O�.V)�q��O[!K��Zh���*\�t����h@�����tP>��T�95�t�U,+ѕ�]�H�eBm��v�w�Q�m9x��
�f.�%[v9��k�?����gۖOn�L&����vJ��{ ��.쾁[q��J��dF�x�ﳍtp{�a�m�C�S�#g{c�o����w�XlxVHYEB     400     100��_���uKdG�k�'jq됊��Q�(��-.�6A�8F���P��-
������fGtE�VV��#�z6�ȑ�c�D�"��M ;e�֟���xF�)=Hk\虔�	��Q0S�����7����$5�V�)Go�V�E��,؋�d�e�>2Htp�ľp�L�+���&�*�I����o>!�~B��)_��H�(�u8��x�ְ���$��"���ЖkA�μn[�2��T����> ���+���Θ4XlxVHYEB     400     170�6��Z���>*�^�[,�Z%��$N��N��yF��&;��Ə����lԟ��8�O�㞌��=I���h�������<���ỻ�s�"� �l���{�A3W�j��f
� ^QA�9w����q��2[�G����<Z���m(����/Ok�bZ�c�<��yהE��ѴUc6`W�$7�/�f �?�I��Ԍ[�8	Uw~��A�b3��@�\��Ĩzu�P0��.J�@�����`�Ô���/4IB`:���^��>��}$4h�M04{O��ĻZ�F�:�V<���
)ds��������Z�b��:~%�cqͤ�ぽ�*�����Ozՙ��b����]w
�VE7b"�XlxVHYEB     400     1b0�����:�3��� �н���ɜ?	}��Čl���,y��I4" �55�m꺎�'���e�k���ȁ��Հ7n�����x�UD�\�);���~��ιJ�(,��M�w�\��~�w�RL�����]����&�0�XO��7xCʾ	rn1O[ڀ��J/b��$}�h�y�����RX�6ɤ#Ckh�b��aPZ��[�Axz��{J�k6���#���|(�)�xs�G^�	��f��i�<�����CV��UHؠE����*��H{|�?I�j�P�D��zU �T��]p�>�S����.�l�#�DO��&���:E{$s�
DWG������j$�T0B4��>��O��#�΄B:�I��9�\���Q����x��d�0	��-~�sb�^�#@ް��Iǭ���E8�Tx.X�Ѧ�9�;�XlxVHYEB     400     160(� ᓐ0g�-�>�p��d���7k��9F]Dg*,TC��j��h��t�/<w�x�(��	0��ي�@Sϋ,DoC��̕�y��J�ׅ����}b�;+�I��eB13��f��<�čE2��b���ȃ�^��u�A"G��zf�;�ړEVj01�K�^#b����%V.)����֫�Ӂ9�%cQ���lU:��x#�Zf����_�KE�*�>��:g��G۽J7��n�0p�����C���3 ���U��W���!��sqy2�V�/�dl>S�=ds�,�q�i���O�%q�af����[j������l�t6�T�B'�XlxVHYEB     400     1d0芫gL�/&�_�%�r����i\�H�ZCR���V
��e��H�n3rg��T���٪4ͨ�]n�����_��=���i3E�"z�p��/Um���*;���A3���E�فj���Ȍϻ��D�2]|�d����R��>ʦ[i�X�h��{�p=Kdk&�بL
���m�sdq��&��1?M�V���ӽ��,�Q���rv\y���8�/:?�l�9^2x*�UQ�C@:ƞ�]lާ0y.���o��������ǽ{�WM�N�z�=�o�g0�,):�eу6rO�H}�ǟ �+��`ɯ%�:첤�N�	8�N������2;�cw]R�+��X������g����Ry蹁��X�� �ۼ)��2��fTs�1��"i���n,���Yy����UO�J��/����e1���:�y8��"�Pųk�n��)�c��׋�XlxVHYEB     400     170�"~)�T� 0-�v��W��v�.�i�S��?aU6�����Eϩ$̂���C��l�b�80V�������kv��=�+$��}>�֐�SO���»�3L0�;����y\̇��U���\���T	h0�䌒��ơ�����웇ǔm��6�V� ��꠹�ܼ!J0���cT��g��7��a4�2
����Q�:EZ��G޶������u[	�@�gl��Ǘ@�{�cD\<-Wp��j�=��
㓋F��g�Ɠy��m&��"7�q"�Z��Sx/����z�쭽l���H)=���7�wq�/���Cn���G�vI�ڭrh�MB�0�l���W�	�^Vl�2��o�=��bC��F�XlxVHYEB     400     160&
��W�0�]o�D��+�-$5��[�a�ۮ�ca�������ۀ3s�j*m^N�9~B���hO��7|(,I`%\��7�:��B���$�{Z��>�	�xp+����x��!C�~��dT��������O�����J�V���ĊzY^@Cڗ�ױ�r�1�����)����\��)��+�!Z�S1~9���>\ ӝ܎� �bJl��ee!4*1�ݞ�j�����W�^����I�Q�$@()0���A���Ϫr r��7��`�t<D�?��%g*�����o�w�N�e��V��+�J�P�Q���AÝX��N�nva`�ȕy�m�i�d�;+c�XlxVHYEB     400     180v�{����������S�&J�>�	�q�/39SRyɕc��@=Z_�9A&�o�{å?#dI$k�k���y+�9=�K��������s���	񣽜�?Xߣ�\�:W��8�.���ƍ�,���F���p����T�����B�I�����'������B�z��Ј6��]�x�E�k�J��*�2j�q�t���.m���D�l��^�Qۯ>�n��IL�"�5v���@Μp$�_V��IU�W� ��I���q�K�vϠ�A��	���E�fVF�6� D��О��\��V���L�k'�2�� Յ[��y�8m(O�r�vMh���פ}�T��/b�ߒp���k�yaAg�-���g�J���.�퐼XlxVHYEB     400     130]���臊��,�B}[���'�� ���Z�	����iM��l�k�����A��*3`!��
��>���v�XQe�T۳��+H��S_�2ߎ)�A"ol������W����$�`k�#y�]�vݘ,B�1�p��T+*W��QIz?�}C����{N��5N!�'�cȯ��;�T���� ���ML���b]��W�?~�q���� ��~:�&�qu���D](׾p�{H]��v���;�5�v�%7�K�,��x��!�C}�]a�֗��7BkL<��2�b�v��7]�XlxVHYEB     400     160�F��jْZq(�mb��&�H��5v���Q�U�sm�����F�E���̎��Pn�J�/�~>��&��:j^��M��/<Ü�*���̻iԏ��J�I9O���1?��"{�/�mo� ��F�d�q.�^HuF��n��JS��`�]�^�	��N���&4�5i��ޱ4���~X̙�Z�9��s;rc���X[��lѦ�`I8�ܥ����m����gy����������E�VcIA^^"��-��3�F�&$��]�Aؓ\9E7�o� j�����O���f�?6�ߛ�;qAO��?�Q	,��=�i��Iw�2�g�@K��+.�2d�XlxVHYEB     287     130�[W}�X��	��'�ۊ��8S���q-�[��2h+�����X�[��7�{��sL2����)s�B���X��{���`
���Z�ǧY�1�n��,�E�u;���{l=R�r|�`��t��q�"I�
�*�c�uhؗ�Bi��ɑL�,�?����r�F	l�,�����>wc�>��=L�D3
�82G=����>T����u�G�Ҏ�I�s�=��7~�R��W��c�s�	��6؆�n�
>�E�H�_��V��&�)'6�B޽	�8��I~��|���S}�