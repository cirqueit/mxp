��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���s��s���L��(�� J�0���M5�������R��S��Uȼ$뀗=��b�}x����2����PݜE����!�����pp���l���XL?8��O�ZJ�����gy��ͧ혷<6
���[3 <>���Y7�	8*G�d��teێS��q��E�a}.��L�"CȄ�(��]��PC��:8��I~D%�O�К㭘[yn��wŪJ��<.��z����L��
s~�Uһ��W�-����Jz���C���J����@��^�������D��9����g�ŶCa_
,	��y[����'�6Y�&ф� �%�PA��ꋟK�4\f�!�5��Ƭa߹�NR�k{�}B=�{8`��@V5X�F'��%\r�����n��M�@���t���,�s���d��pc�%�i�A���2hPis:�^��D�3�4�W�E�)�\�|d�L�mNF-���dx�G���͒4������e:y�\�o��\{��lEP��s��{Y�Y�s�ܢ�/���J�V\;v8w2������'jBD�ә_�1G�
�Rݡ&h��H�أ^NL��z>�\I�Z'f��O�dN�ԅ8��}�� J���r+q^@�Q���pN�l���֢��w��u�>�ԅ7\�Ěu�,G�@֡;�࢟���Z�w�W-�7�f(�������ĭ�>�smx����<�#���N#�K�F8���Ҫ�JY��-�Oc�۞�Bԑ/��U;yt����r�3�-��1MA�(�������9&)��/��BWH(�烉�0yFV� /�M��ke����Vvc�B+�%f����vCy�k\on"��s:|%���<xu	U�rq��L�f�f�̤]�l�L���;Ϫ`�A�#:>5`r�fX�b��	%�K87J|o����G��yߤc�Pf0�۝Z�`L���-��|�iE�ARn�h��j'd������^OGH�T]vfʗbȖ@�,���y�B���<uN�2x�A7Ss�����x�S�� �a
�@QαU�#OD�MAkH���v�̱Qb;�U5�{�b���m|�����.cެ^���"n��&9����&i�fw�|��4�L߼�^V|�k�d/�7bCf��)ojm�� ������g��▮�y� ����ݢ.v$����{4�'�m*�R����x�x3�8FÞ����� ~Z:������s�V)��.8�t�`8�"�����]ϥW9ߝ�?ס���P�L�o!k�s��W����PL�A%p_\k�g�
�ˢ} 
W&9��f���ҥ<|�sz��㵩�'��M;����� ?_�Vʺ-�Q��i��F���x'Pt:�+	�oeYK��$R�i�0�^~�+��ls�4�։���J�J���<�I��O�s@6�p��베@m�����|1޹\�q�'uz{��K��l�Ő�5������+�b��������P�Z6�8����7��b���=���������#�̢�'~)��*%4��T��5 ֫��}��C$7���b�e�^�|�G3�\�)(R���	5����J]r<}5L+��F�g�y�c%�c���EWo��!��}F�͕d}#?;8�Fz���dG�anc���8-Aq��[#������t���6w������(�93����8m�|�!U���0��t��q�ؐ�Fx�L7���L�ě�Ń:>�-\��d�<{&�b۹�|����lT��,��4A,c�A��y�/�G3�7M7�V�lX�͎����f���!8�O���5�`S�;�Z��el&�$��虍g}k�zGx� >�U�mH�6K?�ǃ]��2=���s��+�hL�*w��v��C����'�y���c�/��+=f�@�X��)"�.=��[u>PXtk�d��M���d(Mx�Fـ 2����
��Њ5��I��*E!2�13m�P-�Ln�̶������˗X�[�J�؁�kR~8�5���M�S��`v`)�T���~�Xa/�[ˋZ�(o�|��B�@��K���d-In����4�]/P��uB���%�u���sI���l��t�uNN���@�Q
S� ���aa7��Fb��32B���9|kn�n�dG��23&��(��l�yrD��k�f-��%����aS��Io5�r¹D��cɑĶ�[w:��G��f�(����um5Ֆ+!��*
��)�
�/>���XlJZ_�f^����{C$mr�|(���Vn_��|1��� K.��P�*��-��K���%o�,�w>�c���	eY��Gㆯf^W�\�3�y�p4�h�_,���U%c���@�y��i�ݍɩ4����?�ƾ:J����0�;�����,����'���ѝ���@oH�P$�k�~�36
&1G�a�+�%���䳈��ۙ���ݠ�r��ҐLf��o�e!0Yv���8R���{/�ٟ�8@Q���n��L"2K��a��'y{����gq,'���~J;�̅����b����6�����L펬	h�[������]�T�����x��S�l*��ת�e�`f������ic"��=-3NF�}k�No^�*EGy7_qi�+�̙��t�8�Wk�K���ۜ�I+5gWЪݱH�c8�4�<M�e���j]�g�5�x���R�\���^�V�RR>ai}EI�O��r;.��\�M�!z�bi��3�y;")I,Y�9=CzN#�Е��ͽRߒt.�-�9By����{G����X��KZ=�1׹�a&��I�:Eݵ�:Y��0~��N��ɟ=�zme~S?�\Mx�~�w�pQ+)��ft�*C�~��S��G�U���Ӆ;>��w�	�	]���� � �?�K۱�����&%�:04�aI�1&m������'��0TҘ�īǈ�+|E�cJ>� ���O_�<��i����C���;�`KA����S-���k��	Kz̀�FX��}ܽ�uV�+�tJ�,���i`A>]Z����?�R���#������{���EƱ���&���q�9�\���%�>^�p@��]���2�5j�H�<ɺ��S�_�,6c)޸}���W���s�ziZ$��H��8�#�|C�Gz]'G�*�Io��x�}��ږ@"�{�±X����(L� M���U�Ù`m��`1�[�}xVN��i,V����/c�F

�-�ۆ5F��B����-�ۦ��p��^��C���m�
x�g�gd�ȁ�-��2�7�=��/��!1�ň��%������p$e�>��:���ѓ��ĺ^�Eŋ�t�;8ŕ�(ں�2�&���J����m*�Gr9������ץ�M���~3� :�Zf)1*�9���8�1Jx�+�����J�`��t�V��@�).B�?���N��{�%��l{
�ԫ����^��~�ځ�yAa���&s���GǬ���e�|�G����ш�?ϲ����2zd4���
��b��vnn���ȿ4.�����*�Q� �.Ȣ��ӆ�ֵ��ybq`�gh#��-��r�#V�\H�r�'N=V��%�9�V�VO���	��(
*L�ׄEZ<E�P�\e�@�FL�����ҫ?IǄ�n-�!����!H����458�̢��z����=�KUF�k���
���,ٴ��\m'� �U��#��њK���.����EA��H�B[*f5YN9��Gv�Lp�� 	-�.IR��\�*�֭�~\�J�U~�É��0���+j�ھ0��i�'��/�Z�ֵ�Od6L=���_��2l�,0�9W������	\��g�>��wݳ��;��g6���j�� h+_��m�:{��U3�S�Sk���X�_=v�%fCw�h|�����3��t&Ͱ�I����
���+�+�>��~�.D@����e��K��뚮1>Fe���Kx�5��:l��a 	����}T��7I�h��������<�r6}|�	%�x�O��K͓K�og���U���VR�}Do�bv�w�>5<>�
���V����o��&E����=f)�0��e)p�Sn��k5�o$��H�k��kW�)lǥ-b��