`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
a2f4A3soPj+SsLUVjooF1PpOHlHZlPZ5owU5karFDvE0fqpybI5QvMJt/qTE1Gvmy/v+vI4aEasR
XH3dR0LftDiaaPtG/gzL81uVeABXgfoSO4QoerZ0yrk8B6Cp700VAvoIVSIBJLI0i2nD/07MIY0a
Z3STfdPtDB+N9E7aKgUNhTHWL+nk+/eU2bNn2B5cuRp2yIiAOcAAgaLPG1/AfGTxLFD116HH5IuS
Stxe7UsiJlKBOq60mRPGU5KA8tj4bUNXZ2nHMgZtKZQEECL/xLMyeJV/t3f53+llS3qCSg7Gsuy4
vTq2lwbay95tyNdrCe77l6bm4ufAaY68dmIM4f3grU8B1Ck0niaG416BKdlhmzKxA0nIlpC7tE9u
rbw5s2dd5yPbzMQjm3ZQto4oE/BVZH2Axaq38vspVYGR9jXZKqUu52rx2tBKacxbsFqQS1GbO9zT
CZNWa54CGGnYExOzT1aeBCb2hugg3KOfWmK8qjgR9gwEt8Ob2VB1K6Si7Gd5AMuy3t6fXybE1yVN
Ondh/upB/Q44lBm/0x9usBvvhy/A9KC/V/UEa2uqxf82DDfMmQULo14ZLleaman5QW80lYXh3HBo
Ffay3e3livcNECF1ztKivgJgCUf7ZoSbdCBQp0IGyDXyFcIWDEkA9yplghRN4WBBmLghp5DnQ+us
DpsgVs7AVsOlcyTQw8DR9WyNiBQNESZ+oq6lmCKP91cUNUz4lg3mWkdsVqRJ3yfKB1WNpSAj7hqt
qaE9XmpKL/oQMRqOw/KSMi2mqTmgSrDuy5my+sP5Rj65l4Rv5hgRQcRApmtEC28NIeEHS5SKh/nT
xJJz9wx6xszfhtPOgja8BRJm8kG2qOnExOiAvT06v7Yt0KAh0ASneUPlxA39xoqDTbPDSRvGTudO
C7Ghu61J6gYZnvguUvij4K7pzT2ZlvYr9BJEM20MGeGD5wjZkRhmBcHhuXSDYHgSEcFFKkP5M9Iv
WE4JZ9koXPKQ5v+tJ8MgVqIyBLvy3oPnRSb+x372WBsJIlNETh+u2iJgsqYTEa0IjQm6DASSHlsd
MFjAb7orfVFnJidO0TbDIaqvFUTgpGFJT851/IeXnq54Vb9h6FvYu0DysjxHkm8YZGCsiHNX+9vx
lG9cBz74a3+UJan+EVF6HMPC9GZVtNQhBp6siRrNz00vi0NmJh1teq+xBdXwoOHH+AhKB1ZZFkAt
4sl3rt00r+trgU/TrG2KEwf3EnCpp9jf2c8OVJpVvOTLoi/VMARVTMuxp3PoH2hgQ7UWnBJEO6Qx
ZCN7KTuQNxieSn5QCuhNyqR5O7OVWGCiECXtyL3XPRroHv3H7ITgB3NpUBGZwejD9rV7k5Uck0sL
ostbs33/V4txIfnHbkgfxxZMRpFAhmqmJm0hHdQ9TjUU9fFZ8RPE151+sObFo8Asi7kC4hMlYpnc
ctCM96Nbng6KhZs6YnXoIbb9SBKI8xjAASwKoNmUcXyezUwtP5DJaXvG4u8z/nWAaKzJwRvbdk6b
Vte34MTF9cP20dtf7ZM8+1YOqWKxtEro9PtijeLeQfPvC1BdeTLLqexYnB1uKamwigPu792YdmFJ
FZmuM2+RNTuC0P1YXgzjfdwZkpTG9ggpIdsX5hJoV1I0a10lViA1bwrBt2se/kyGgY933HhmUgq3
HcClher5i4aBl9b2ZS3mlrugB8JG2yjDvcXX/U/Hv3A8P9p48fwAASh5L/RO9m/+d7qk7MpDeXLW
TYVBd/o7kA1TtGllh45i4h7UuJqiX+TzMHHiZ+/AuRTnommiBBBVqIRY5rRkWSmcwWsFwrjaro0V
UrSKLrmgXH0RwhymSneGoJJ85knNc350cpS9YiCBM+QJdVqob9Ggduocx1ZsZoezESFP8OkpHIE9
bxpdgaP6ScUGqzRonU9tRUS4kSRa0baCd4yBdDByEQkQ1oUrxM4oG34A6PiHRrifdPxqxj6eKoyu
eu0hDDxYmJ+Ph41K9T5RRa8xquPjMin1+b9ERrx391qzZCGkBlu5we5W7N+Ngi2SWidB+6/uTp0G
T8eWbo5OLyuKQ/lxKFmGBfed3rlfP5JLFh9vBiY735HwM9X8swrpkKvW9gQteSlowzWw64tCyOlg
UwMc0WH2TG3wMpDYW2oWVAXvt9nRKaFM5pdnvCZTznGUGD38HnxVVDbRCQkLHq2teL9LUIo18XR9
IBNwdMNndpPdRonW8isAAMprVF1rjt/T77V/yL+VY18ZIW0Q+Q4Q44441LF8K45wb8RayPjapROp
ZB18KtONhNNh55yds71YcMmhDieMiZq6eRojEadZ3i7+gWVnUugFZhQmui5QUStKliUoUqpAgjkG
9hrXxBmJSIGqK94LWUFMZNS1SnsL6rr0i6kW1eG5v/GRpAEml/6u1nTsrGxvv8FPmCT9p18eE7A4
ZLtkXaV+HFKi+RVyLQsPOH09Hc9qn0rVw2fGrjrN6jUnfBUPV0wv/MRZ4Ab0MTVoLH+ayMYmRyPb
GOUzXeYo45mU9MzCKZ6N/hrlnl9DuBqOcHre4qBV5HG1D5//K6yTKdbsDI9fD0gQlVyFzYpPQhLn
+87re5agXCMZt/8+aXW0MBcfNP/qZGARpXfNx6xH7LktZsXSARKfRilPAWDYadKhAvIohFAV8sLv
hTXdpmIIyas5lop0hm6o7YTE00a0fD/J/oXtvADXvTZxiYu51w8xdAjK3MG99YEsorMnB+cO2tK5
+L322ae8qpN2Bdq5Bh78NncjbetGusK52+kSIftw4U+lrLv12fi+kQrKHsvKeSkRRp8J4NZw5yQT
GtuFG71citEtikZ0wLeuxJ5hWodkiQVR5cwCc3bEorz1qewxB4wrrOAcOiJXpfxDdjVu5DQN7yv/
HcZ2YBUNMwUSUfEzlvTJCWpT8P9ZsJ1W/x68GfqeTAATLzqiNY2DCuEAbMIeL41yYnGqgdR4LpZ0
iIqrlqrkXGmdDpq0j8BhLo136iwDMVw8SU9fQ5gya6XgpREzv6uLRdKkjLp1s/S+u2T9rGA7Htbj
kL1qUpY5kun9SjsANni0O2hb5MyK+dGfKbgrdm7IldicT15Hj5+TpB7BM2psfX8t4ZQTbACvb4fN
OWAxy8Ob75wY4SbjKWoC7WuFPWlHas7gelrO1qXS3QjH9FF0WyypSVRuRHKlAuzddDGlyVLzZD58
q+EAKhoo5kizWwlputi8lbIz6m3og/tjmlgFZs2pJ78A6nzqSOzHuJU2zPskQTNYI+MePukll2Ig
vFZBUkaoUpSVouZuLSgHm/KucfOkDv2hEHy2cVxyE7f4+vFFU9rdpnHMAwZWrBa7Aj0WR9jqRYOR
8+r4YnKTgLURfY5CAYoE+zAqmFUK/b6fw2jxkP6GyVQk99WaLupDFIXidPFlIGcdBtpFu+9gAQqy
AYkhcvVv1n/ZKXe8lCnzfV7IJZvDuTcANbg3f//2sdxJd+qw/yBGmsN2F4/NT76bmvzeJkh6eLd8
hreyZwHZyFvZeisiyoEWR+5wgZ94NLf/PtRJPz9DlXSLbii6L9x4ViQQi/NBTHumlaS1Omrs5PCi
8IWzTWcwxd9BZB7Kwe9jsiVfIUSo21FUOf2phgfJqZsouXJFwqvDdB+fKHVz4ZyKg+QxwuwpRO8Z
iyoHIguxbdmuWHs41yKk9I1JqKhrVVs6UMuhxGHlifxcW3UPsmhuyVQ1re511xCAaY6UTQDMwHZt
aXdyPcta0/+qprUexeYgmLQvJRE1txLDRFIcUAX5aB0ACHV/epCQS8wpRilnSbjDWy5N5FTMeHrn
V9YQAaXW6pPk56Cu2VxEtCRJO2TMrUsSVrt9h5NX+D0v9WPkeh++S33isOE1E+bf14VVGbFT30xD
JKVZj2XMaNHa9/7Rvg2ArRkJj1C6J5doUEvA9aC4dfZVGH0a816GT0fvhIiyExTZF/w+Z4M522/Q
+G50/DUPymJENnAbQoQuTLlurKOOYKaeLT721cNklQep5jRLx4DvlwVmHRGLZ2jxfZWm8l62ww18
eFIjGvs2kEkiJX9/JP4dR5Lpar/xF+UqbcCWsr5mNjvfI5l/Pq/PCw8GkbXk6+JBMJAFwxndbTXl
fcmb1AJFFkw6UFuslSgK4kN1G1QfvtmctdsQFfLu4IXSBupvkhPqxwz/UgQWJkXwX2W7DWpbmqlL
fXKLTbFusgKh9ZPda4JqHIfQvDEwqsdfUgKejy/OFUkfoiOeCwOQdfDYxinAcC5mzk4SL3rAhvAG
jk7QGHKqrleu5UNCRwIPNJfkv3T5aI2zzlxF23DnbgUKUJVXgwpbBaf7ywNY5OfECMRszf+E5HCL
wu+k2ZOtFr5wwrMjX2xrqvu2ElEvLmfV6Pt8sPKQq2RSHq0BZz/h4B4JFWGUdCkCg3j0jhG0e6rs
574cuQZXXde6yjUvW1lYTKPRTtT/pzAzwDtcKIafdbTeTRDclEbYFAfPFTQIW4zb/B5H6oBoIFPB
ymJh2QV4+4Si1KLXbEJFUgwdjTJ4Rn3xNmzCQqimdwGMFvTjHBtbQQ2vXl+b9MLJMqgMd/43SbFn
zSTJVfk/BCiPU3ZdzxH1jyG2w9V/3mpwEboEva4UK3JnDyeNfS9X3XJv612qlyAW4ja21F39C7J/
CO+XAmA4ueiNllsrd1X8CqP7Gx6LnQfv7yBATjeS+W04y/5/atqg8PCnh1MEziQ9gCU1UaSUcBRf
M6TwyoA4/D2M4niZ520EZnv6OrXjSzRLyzbA3lXSikUy7b1v320YrEbIDumvISD+Dw9WVLijptv5
sT8MQtVB6Ekla4d+DJO1cMD/dWRdgw+NfoSQeQBXVMN+AB/s2BBIxLQIulMup0G7yRmqzcGNNN0U
E+W9+PIuDG+UJL47I0vcgLMC8fQ6c0OInmp1is0E57NKLqE+Z6y+bTIX9dId/27eYDQYw0oaHJBv
sxd4DF0uFN16ZN4hvm1gUX3/O9N4yzfL+Y7xFIfp+jUf7j2aYuTBTZQJJ5Mf0ErqsbtccXw0b7Jn
9g/s5e8WdIkevmecrifwOrUGQM2EdK2VbM/9bxTfjmA2llOx3krXrcE67ygZafgQydNhRfcGIP2J
gxHvLWTYqZckxrCIIW/msdtkwVtRyQHeODLPnd6atNsYihCSq6fJVXGcgoWTnBpIHio/6sLsVBiu
dvBBPn7W9W3Ke62gXjFebU1nWAUv90YzI+VU+M82zdZVb7TH1Ew4M/hz7vTR1mqJBomFcBy81IFG
El5oh7BqBr47I5vxMB2GdUhpJMoDkzpfEsIgy8FiYtSFlrhX8UZljfUk53hUg30688bJTMr4dqQ2
1YxDCSh+WewFMwpVSlBijT5W3F54T+wxvFToxlE691d018r7G3H1H4Xz1bvK63jFkSvG8dAdkJ3i
MfF2OFfsWeAO9IScEc8RuBmWuLF3OzpmMDp/WDznrxLJJ3c1btH0Zk3y9QA/EsMERzaUDJSTNPOa
KkHBS6CTqEvH0oxxXL7nyywI9AEmsUTM3XVnhiEqOpO7FOUsfjPpaWk/X6rjKHpIfS1rO/gZDmRz
mg7n+P2Y8PdG11JK2IqO6K0IJhPuTZjiU1Rmk2VH6C9A9Nyl6FiTEd3ldj2JIB9tFJCiTSpIU0lJ
FNVSt+d/PYVmZNYI/Wxkn7Ouw9RC3dipMKatBw+GAI7KpRrNe632QsxS+1vhip2Kj6fXOOjVzz6h
Md3KEsiFJamH6pOue1acpOzSdNBeqke3lAl0EqI7CgS+dCu8ZujrWzbcV4am5cDsfo1+3rmRwUb0
/+uyTi2ldJLt/VAvgu4+6Of6sY9qGvLB/ZUeSfnmaIvPi3Fi49Zum6FRCBRNP55wlYlX085XkVbV
Qu8ZEP0CEkq43NuofcYokulLcxacKR7hq0DMeiUdwm8DnrKHmfikRyadz8qDntqLUDDOD0h7Rmjr
gDbB7e2DcUZhfE0/dTuu7lqwp1GS1ALHiyJNsxqxcBZRfpI582QZLVmy7d9dT+0gAdno7WJOnClQ
TdTOPFLl7UFnSsdeKMfz8Ha4Zsuf5tbQGBIExvgbhckL9M9C8mcOXAypdTpXeXo2yiwIQS3V9O2M
KAo/jHPMOQvZbQtpFZ13m+aJxUPC5IXychIxSE3KTsgupUd3OPDAekrQzed1hJwU2s6HJUGzthKT
+xSdExbNnAnJPXE53w3/fFjEHx9IM6sXqaIuw+MtGbHvnAC+kctTRNDVyQc+LixzfFUU/656EGiU
BnSSxjgDKJTSA8wF9pMhAxYlwCXAvtATVe8tRbnwcJUmTu0+y2PDMz8tobSKJD4w9tCJ0n+cKZQV
VZJRRUExL04jSQ1nswX5KaAiUvMOICLuhMc7BxRa+w4cyI/n2TfWQxPbcm7/D6HrNn0r2wprQd8D
SYw0iuuo1RximcAtSwwJXoZwRD6kCF882rrF7isAdH4Gjb4V1alukzs537zACcErhBFh1qjwxGnE
p0Dci49zw5XBBuZz1AwI8J8ogvCd74g/JvLd5h5onSYPp1pye0VDm3XcbV13jikCEXDlTp/LgqsV
9BBBVfY/Qpv/7ne6+OWCckyK1zg526C1+eFZJn7BrjoSW4iFDYbOP1C0PSnbMEbmkmlWvyIcxhDu
5uLpe9wtrELakkZr8zxCv4cEzVfUGRoN/niHz8k2OG6Ga6TvCY6flyC7hhddvOUgsOTHP1QRXguG
B4Finwfk4KPlxlVbOUrOJl9+QJkXwn1k44dAC81xFJv/B9N2igeUjFqF8ALkQLCh7hObKpGkXec+
ed3spV/J2BADjDWWd2OTmXhUa0w1UPQrocJubHhUYrfme+0S42aOaAAwMbjiBQ53rhn39ftuUwkY
rEtGqbfWBylKxu17vPZrxYLYKwvx8Vf99txRTTaBexUkkHHLrjMUub7DQQudQ+Ha9m7pHH/B8N9d
/LMmf6hgY2k3LDs/AdjLmVTOAmIVEkSQGaVJVA6yx2RwOiSGv81+jhCXi95+CHSPL5zgjRY2eiJi
gXTXKdBqAszZr/DvkreL7wqlr8VydDkMpbgwhJDt0eK/v1048nVP8b9d/g90yzdYvr3kcXbq0ybC
f0WfxQz3H197Bt80GNgjVbeWjdS+dpWgl/SqJsT6WHl3ceKNANG7LNdykzU2D6h16+HeGg3r+DKL
xO7UhLbdl+ypAlqRgvm2rfR/8qer4+gxjwDsN1mm3qKbc83OWDBgT1Z5/V6pOSJ0MNz2v+7qXEHD
yRPTUkEcTnHY5tk+BUsVcmvf9oXCqB0Mj3yVhavMaNMjk3GnbRoPfvQ//koEkWSh4V3HElKrPUvX
ovVrM3cp84ADQZS4L2txbMSa1cYqKygJ1WJp4+liLEuKU0oBzD/tofZptYDc2XAr0CHwApuzIcwR
6V0r1ovzVvAgvVWfAZxci4pcRYCd3SOzfAEGBoqzDRLTW4vBNe+xylHmxSi1EbVSZvNm7cv1dlC5
o7dynD0pXOzAfY/4SXR+6pxR0zW2fT7ZchBNMakegodMTK6MB+51ZCpDQTC8P162U4GzbwLHnGY1
QnCPZcHQjAGVTYARm/gur81P5Fcx3pawzxHGysmottfSDuqmridw+rshB9JMOuvlV8DbMU/Z6BVN
CYM/jX4Yy1BhNlyJ6Wlmr8gpi1tOSEBuKmJ0adPhMoWMa/PIpuJutsmtFRwL4MKW6MLbNLtWTOuK
5p2GP9wXRyiMvDFUz3HU/gQxHwGaqHTz0IGisxsgJW2oTReuHurP10ud9xoCwwTD3xyn/XE9DiUh
B1YiREC2y17ppKuZVQCbNANok0umusHT+YbX7JZjUl1T0bNIfLtoyd/ou7EraUq/U2tcxgW24mbi
RD5aw2KnIYijKVeGgMf8XSpj9eqQJY8B/xDZWXEAWksdkvGyOujwfE4NSvZVL1U60J1BHuCVM58Q
zGVauYKW/nU4PXwxOGDdqkak3IoWPYYoUqwcfhMB9XrgAIQJEM4WiRNUNgejDBJJnctlxbM3XpMC
LZqEV+/+xCgIw14xhmBDTVNV2L9ECwAJ70TEAZZurL/5f1BKWZvQF63Ld3J186JH0FdbOxx5CcLe
AtKCFrnFrLMc2s6ZG8+VxSjQHvhXbelRzh+VrjQc4yJnxeI4Lkxz2BhR/HeCdvV8s0TTqXWjICFs
lwQE6o+SxLD+YU/j993h3eALMWGaluHZMq56zxX+aiN4H+xyoCIkjhHgx967jKOQbZNAKjB9I4dF
f6zCGYi0vu46ZAEyOGF3gMfa1twMToY2OShCTRbzOqbccbQhjZhDQZcFtKCpOVF56X9SqIXXPgOe
HF9p0WQPVa8FrN7/hYexfoQzIPh49eDPDulaNjox2EGcQDxehRuOi35YF5LEe8/LNfjJFe10MZOT
+9QfUOkdRHCq7yDujS5Lk1V7HvYJ309RNDVJnWW9Fr4WbGiVfEPh7j3yTcwVRUEGavI2c+bwkwm7
6HjqXgfx9DF1ZQ5Pu+VVdXet8haBMdTiUUcM/wds/u63rXtX+FGEqBPhnF8zV6u1MZOxgVntpSEl
h57u9xTFEiA1xVZ9wWfO+Q==
`protect end_protected
