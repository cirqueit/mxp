XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
�ű���h��$G�|���Ta8�(��f��dVZ�<�[�����yz�"�='`�K�Vn�Y�7-����[[4�][4 |�Μ�V>�o/�������B�R�X{l\&�:����d[�d*Jm��΄y��j����hy!��Ȝ9���>mNH�YTzo��#�e�����������Hv-;e !q:��O�Ӡ��d�<o=�����/$"`�"�b�:��S�˫`��m�v��{[�&�
ꋒ+A���Ҟ�}�|jMh��֊mԨ05�@(���Q[伾���3�S�[Me���,]��Al�HӤ����r%j���~�:�
I�c=�����J��zZ�R(=��n��J�s(\�Խ_d'��>��X:3���������a�Oj���^01ɗ����C��G>�$Sn�1{����\u��#�>A���#ŵ�,��-4����#�e��{�������(B�ۗl;unlWc�"��
+��ӂ��>��R�"�k�L[�qMa�G>;��<"n���N7��x��ڽ���
N1�,��J�6�v�x�TK����� ��~�^��|���I1������w,���rp?VƯS9��! Ay4�
�kh�|>����R��d&�fHg��,[ް�G&dE6@t��X�Rs� [7�d�p���dܕ+�� �����Y�RC/��}9/������%��q�Qq�E�߾�n�kg�-�Im Mn�.�4x��y�&V[�JJ�pڣ�xXlxVHYEB     400     1a0��??
ǳi���c��2
�(L��͏��qU�x�(�!�/U蘷]H�JS�SLj�C/�J�V^�S·$A0P����_u� ��k�Tɣ�AUګN�gK����K�X���H0��'L�xu�����biE�ʛ���p���(h$ d���W���'��2����T��	�f
a򁝍5�����1RF��&�EO��tJ�&`�-��L�p�����8m�a��ڒ��IWϪ��x�S��f: ��?�%-��oP��J�Q$'#����������z�9i�ݞ��$�*�o ������h�&xEg� �q��]ڞ�̓�ͦD�?0y���S��R��V��z�d�=����m�'��h��a��:�:10��3_�,@s�h���U{���k�D7,���XlxVHYEB     400     1b0.��{�S�	{t�?�=�@J��H]1ڭ�.k��~LZJ��"����<�15��k6��f��z�Q��%�v���q8)���|+F�Ձ5�^�����֑޾����wr�<-y1!H@��V�&%)�2�9Vu�0�2�Pg�PG}��ņ�i�6K��퍞�Ѐq;���t|���#.
=��R���&ʅ���IJV��êω|sį�������Z��n�׼1$��fnzgn�)E0�V�;S�P&�e#~Q���!��e��	x/l�5j-�q��zX3t�a�j��^��He=��19��h!īi�����@q~��.��a��}V�����z���m|�� ���B����O�2��~�+�`�m7�X;~���js���"�$2��u�ʶ[�=2x +1�������ي_P9ҒI���CŚ߱>XlxVHYEB     3f5     130mݠ܎ث��?j�@���l܌֫�E�i�H���f��6[���!�����{6i���(\�6⟊us/;ش� d��ȅ~kDɪ싴OW�,��v�Թ��L[�:k� �:]�����Y��޼�?t�gTg\�,�|�5��K˸�������.���i�� ���+�Mr�━v��랞%"�g���M��[y� �r�i0$ Ϯ�o��b�HJw���Z&xx�w��k����P�H�Y:�}<���sm�=@yi#�s�G��m���,�.�{bpW�