XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����CF���h��(���rK���=����u�d�75�n���	�Pk&ؙ:��9��eRܷ����sŴ�S x����)��_�p�#�	�-:0R�Z#O|�&������tz��P�ȏ	�I�o)�x��ޯ�n?�f���#_CI�y��E{�R^�7A�D��?d��2VP!Rܣ������k&��Ig��&�m��u��\Ը�J��=h�~�a�h�*��3��7k���vp��B�د����,�q_v�X≻ja%��v]�ｴs�u�}�-��zBE�Hrn赱�p���Ov��H2���A�V��	���C��x*P��­Sh�Q�ږ*6Y�0�qb6��l��_���uR��\^RP�M�������� �v={���e*�������)�S�X�̜�6E~�@��@���z��t���!�0U�F*�1�E �YX-�Rs�}�A|-�ft�!�܊��&o����`�w�ڵ{����/��]W�.�+��`���M�S�91�a_U�m�Y`pIU���&�Qc���d��e�S�?Hog^7�ɑ��\Ò����O��N�t7PT|4]u��<�^T�[��m#yd��@�l��is�LL���
�h��f������O��F��4�]��)RR�*�)�������
�D"�>Z��Nv���(�(�-��9=�}��9`��8���uT����O�P��H�⨸�݉���&��$���R'�2d���l���!�1܅:u���w�����C��XlxVHYEB     400     1b0��8�-6�P�_-�ST�lㅱ�2��=��fn�(��]�����ӡ�J_}t�HYW�9PpY/=����.3ʤw/�l�JD>ʦ�|xjM�8$��!A�E6����a5f���VHi6�Ƶ��&�ᐄF���K������W��:L~'�_E�t�G���4^<N^q{� ��M�\CNb����5Qh�q�?�y��Ì)�sa�%o�.�jFީ��)`������#���=cG1H�QK��(��S;�R&&���<*E�1��+�j0�u['���BNY�0m�/Aܗ�6n�"��Qp�Y�Və9��OcB�LY�N��DK�O�u�m2!���+dn˲!�@�lWu�*4�Nxƒ���dH����ޜ�r��G�,~�73������(�U� N��?�g�>s�m�x=V�e�ϛo��i��
~�&XlxVHYEB     400     1b0U9$�w�.���
*��V�����Ed�{�����T-W�C����a/�����{ǂ5�_'����<�]NՅ��"f�)��%���# �<���h�=��܍��2��{�h��t���W�7
��������tgC��6M�L�^l7��U�ڄ��I��R�6/�]�O��5l��K���7�����|��`B@M���O=Ih_2{���D���$�l�{�0���v(�{n�Y�]k#��Q���P #�
�wp���f�݇��k=}�iz�R'A�w�R9�S�&��{�
��x�o���L~�+n���f[��|}c1��*j��]@��D�{y�����2!ll��<����|���Hc-V��H��1���*߬�(6�q�YZ�JZ��M�,�NK,�!��`��žώ$R�J�h�?�y�>�MXlxVHYEB     400     130.ѠX.�)r5 �b��@퇅ޔ��rUU%�����`)�?S 9��:Dm9���9��kǶ¿�:�橎X�x:B{���U@��҉�"B�~���9^���1��V��n���w�;8RY��$��+Ν�����,Ym����Ռg�+�	I(��`��i�Gh����. Y!��B�!����Zzߘ�hc���K�^�ߘݣh����)L��8d&�0Ȕ��p��N�⒒�#x��6������˧`���T�DG7����6d�]��!�*�sG>�G�a�=��BX���%}XlxVHYEB     400     190��^c�~U7P����^�<]�v������{�����]�b��;�����x\ά3�����}Z%�
�w�mV�m�̶���'�ӫo}�*(��f��Q���ѐ�Ys�ZJD��,��k*ԕuC�C��mE5�[�K��~B\��g}�FH���E6�~�S�W��q���m~/� �1���r��&�f�`�fĻ���MCg&�y!��Ǝɽx��M��3��� ��zrL�����$|���y�y3��J�؅�QvJTQ��������!F��$�x[]�`�V�F�?��:�z���eʵ���&,�52�Ri�h���5��Ϩ[�6e��vd�.g#=V,��C��|�s#�d�o!TGSq��ҹ\]+�Dz�H���d-��� ��gT�p����>$uJՖI�im2h�XlxVHYEB     400     160��Ͼ8Ap�]�y�ݗ�[��[�
KK�%��0���'#UG���a?Ё=�L��w�Ed�����vz"��z�yT���-
[k*��CmL���P�����"�=}8��T ���L#��:�k7J�؈H� �#���C�=�t�"���jf�a�5��x�������
�ͱ@]�����!̢`�d��1]Yw�{��+��m��W�1��rrv����i.�L+������T�u�{�p;]�>&��9G��xB7R�p6�dO���.�@��²�["�rD���@*�]��]�;迩w1��&=� ���P*Tv���`]˺\J|;H����`a-x�QXlxVHYEB     400     1b0U2�H}�6��s)~�2�h����<�5����\˨{@�W��szn K�,��0kߔW<wg�w5��.�TI��P�.i]Y4|%��d6(B	%�8۹�{{�J�?:.�n�w�6�R:.��dS�c���S��q�l�:��?�K��O������������B�`)"Jy
4E��:[��i�g0�k��������������<oi��/ێ��u6�$IX�´���e�7`%0��,*�"�O����y�E��7a�D ~�N�N;���m�uF�sUms��w�8�~	~<�+�]G�y٘M�V%������R�UK�.?�<l�/~�9��P}g��۱����״T���1+.����M5@;D֋�����r��?��uzSjFʊ���0h{P/@S����x?c�Ý�\lSB�U^x~Dl�XlxVHYEB     400     160(��Y��AxK ��f<�_�\�Ty����X��Ȍ3�i�,��S�Q�f�)<T�e�w��7Ӂ]���������0!�;,d�E��{,�;&�]�\���=�UQ������*o�����kxFE��!�r���h��J8�'���]l݌:��lsd�cө7��[d� ���V�O�R��6��m��[QL��s�n�����k�l
��>uzj���$z@�
'�N�P��?��㽲υ��˘?5�u`P�J���i���ûS0�N#���3;\����a头�y����	V����'�NS�J����rj� ���q�1�>���^���\�EJn��b�
56XlxVHYEB     400     120}����Q��\�:!��V> ��tN3�2�U�F��X�����>��O[�h�sF)��RE�jTÈ]�u�JI`�(|�ߊ���2K��Zn���<=>H�2
���W�`#ˎ���·�-L56�ʖ{����t�y�&mO��n1�rZ�}�ez��5�i��H�d��%��.�Ŝ�\��V�Ë�W�P�xw����?����<�Jw��V9��0�s��V������v��]���^���K��V��8X��]�i*�3 M��|}Y�L72~�\�:�#�(c��L=�XlxVHYEB     400     190z%:)�)��i{�*S�h�M���F�Ko6��i�RV�n�t1J���T
�*21\!̛�-�̉t��5dߋ�gQst�/e�4�-hH�^l ����ٲ��Qh��G��1a��P`G0K]+�:�Z�$�����/]��{���?��S¿���aߪh�m���z�Σ���<q��Z���L��\h�<��-Ǫ���t{�P�!�s1q�i�_��,�D��Q��Ӌn���AhS7�FptTtw#c�f���[΍�R#C+��8�
����N�u�x)I)jW�&W���)�q�OLΦbs��&��"L���$Ԟ.{���p�^�����a&=J��R��F�
��������BŊaE�,�bz�������HVKF��?�3
����1�IQ��XlxVHYEB     400     140�Q2/�Q��c�N�JFl��#%�i��¾ V��;3���=p\�v���pB���g��6-۴��)�b�9S��t��#Loj�Yڎ�ݟ��W9����N�Iu�Ÿ�]3(yTS �=�CY�!p���OɚaݰS#�P��r)�m�*�4����	�
2��tA6�PT��d�������\��x��@��ʍ���y�;�]���D!����䐓kZ����l��P �:�DEϡǅ;nvڏ����e�Xƕ�O�L��¥�m�]O��!8�F~?��n�h�X�ib!A�7�o;�ͣ�<�=���XlxVHYEB     400     160j�Z�����r-�L&q����Sg�@"n�/�+����^�.?���'���׃��s�2��*�@�^ՔdD���2�.��X* r�� 2p��!�SǠͿ�`�wd��}�e�Z�~|�+�#���L��dV��5S��
�0:O�~�h�}T^BJ!ϐ�֐�	V���"v�J�ω&�F�E���[��	T��&fٳ�n��֒c�ٟ:�-]��R5�6w�s�=~m���3Vc_�������� 	�YӖa��F��Ԡ3^W��p��0+�v�"._��w��t���>���Z0�]���Ȅ6^v����T����xu*���gѹ*��m>^l/����HGi���XlxVHYEB     21a     100�j��h^r&ܼ'�i����~�-r�%��5��V������\�n�}�`�b�X\�8g�a���W��\�����ґ��7�%=&����=ծ�G풏5&ht��b�?��Ch�%CkMJE��s�d�i�%Mr^�U�p|}(��`!���e�XǓ2���wt/C��([�~}p�+��<щQu�xuҼ]Af�v%|���8@\��A���<�i�|���n��w;���2O��ifo w�k�/6����