`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3088)
`protect data_block
iLcTaxmT0WpW1SZCvRXYofpYX3fj7r3qA2OhC2toSBAwXfawUgjC6psAqiyUGX4fRf8VdBBYmWRD
EzMlxnzPLWar44t90wbwQxMyBrvA1LDExnuZGYO2SC65UhVHvi5L1enC2bFwsoA6GL3/mg5be0bN
w/r9v7vVulPzYnVNdqPvRkz5O+xuBi6WElX7jCgSXFAgnOOKUifqYK6wLB3+1cXDZGHC4D74OMf0
iPxsoUgVpXNdI1n+ZjmNqiEpkYR60m5esCMIezRX2oI7qMZW72n14jb73h4q31tN4FLaugV9j/NT
0U75UtMQRNTwkS01yExcIUeycWBpXLzZaGxjWK57coDuyivnbbMEKcxM+tq/pS1q+/jtmguRrUdb
7McEw+YYx2sIN76NMtq8eE1SZ5+RHKeJCP9bpjbzA74+JdXMn7bDKymFxZu7D4LF55Jhmt5NNJy9
aRntyljGXc9EXqoEge+73vUtP28/7ZrZPX3QIGVqWrQNhTbdzNBYI6+VuWcbHYej1TRVyOd5Fnz6
pNib9jwQg7kipr2i4/vtuH9RySqLJWPbt9M41H5Lk0zY3ZuIGW3h1QADZW5zzdylZZ6f2PfKwTtN
yac8G9fr19H5lEtms5M0P55VDZdNlfwEwS9r5F4kPJTE291IfplydC15rMo2V7YSZgV12Q1NZ/RZ
MwAGxE5OSVW24q2JKmRmm1kiL2txUzzb+nEYwpG8rPRIbJw/vIrbpsD5/RqVnP2Kufp3M+3DAFeS
KwPQol4WosjRuC3qI3MWqCUCVSj7gmQtKUk22Ad0cp/XdeweS1mID52S1g6waV0QZRswxnWEZ76u
Zp34lJdK8JVK/xRx5zqv+g0i+BnzqL6yvy+c0aypQ1pltLXdk9eU/gNcobfIc4xhIhek/b084Izu
zuw+VwV2JjD4DMqEEed7bz8vFo1BDZ1S3LswKoXP1wBUN8G1LlqcDX7gzv71JJOEsM8PHvU25ujD
u8HhzPMAyJp/BtpRRIw6uruzo5Jpx8bsRxNFmNwsws6pG1fNB2ihOuEBWlNhaicBZE1ixeUJwXYX
xJJoEJBADRI7LPITLwhtKQjEBbxFmabctr4Ry99CeC5wA3PAbq/dZBir7SkW0cGO5ahuZNDDUn+P
Mvk4xKBQdPCo9qRxBC3mOliTp47alfIIm4iD5iEtRXu+KgN8RZszS68LIC6cOTJrEkIlbv22wRFT
zxan1e6DCrChcvhbJ+2tl0YOMLWLNNo9p8udIjjXovdUX9UAQ7B//XwzGBMjj71h0gO8qi1MVoYr
jWJIeo2uJejby5nv4fKcXtCTM/i8WtxdgSPIFJ7M17GVdSniLXu+3CmFBmlpVb2+PWmiKACIru/f
aNjVBSVgSqJk6Fxc2sipwMJTZFJMFj0zb1Yksf4CgLszDHJHMPlDalXEvVd1Bg2thWujKvKFHBAo
g9T99N1+JWKv15Vv4mNoYwuSA1Ea8BNaMDUUVGth2+yPc5qSyx4EFc+d5oZlRTckeO7PTe9/2QhY
bwF1lSTJElpdqa+dJ0xmRDtKSpCwhCgcf15sorDJk+XrCT4ccGmJXov3ujVOHGUbOUl0H/FVJrXn
Kx+PS283eDezUkeNC0QnaFUCZqiU+TxeohwPYiY1pwYHA6c0mslU3mKoba5muc4tT7Qy367b1Q/n
20rowfv9nOVbLDvKTQFpMrgs/PG+EMuhN8LcOM2ccjGzjutAQaxIqP/1RqmOwgh0GiamPBb6re8m
16zim3e/iunp9Zur5f5hSldv+OeOpt5xkmhTSc3w0DTkPeyEDolk7bmpe2FUNKDETv9k18H8R1Je
wRcw1CnnqLCWyCovv7EUS0GoILTpIk6xJw768PkFT4twD8YQFazPVdcQuKk2Eu8UM5GKK6KJhucv
Yc8c0CFzZmLlY/EpvmbO/jX0kyXmtS3u6zpFmKzNzqNSILrdRI3i/vNaag6Vnbv4xGYV7WD+iYvy
pAaTvgxfod8iBW/mzIyU9RtfoZ0IA12R11KkgJGQjFPNqNDF4VDKqbxcCEfhqG6zc90eDWsAcDhk
CIYBMXgad/f+5Mx3KgE7QBYfYqKjgTLwUf9U0xMjZWOJyP2qMIiRfxQv4cqN/s1YkTAUN66V5q+M
um8cZLH0ZxuZ1zyL/eXg9Wth5vjhu6K04lm9LJBOvt65ojP1acgRe9h5DUFMqQrM7EF9zH+Ml1Ow
0wI10yiL8DqH9/pVS8vUKYQcbYOONb/ytVtTBqZRVAnq0Zap0drJSmW/uj//N0vktG2tcnzZnsD3
T3GbZcxexMkmQJ2BFo8kHzgrCKfNuwyiPItFyuM13hWsGk4cNFV70KrI7S3lWDFhoJOl6DoaSfIk
i/NHuruMByCyx9hJgJHl6AyFMMUJzVIBX8ACPhJtxXzUSEsgOqkICNpdfdYyxe+a0EDs6/Xspglr
deKDfLOkvvS0OohJzJXDGVUZyMICbBMwoqazQi+lNOiT+TT4REkdLAvpl7fyo2xejhzwNvxeosUa
VSnD7BBaRHA+MBm54J/JQX/aVIFGKZu9+5AIHmH/VA28dZ1VChjfVPiqySmEzpuqCOnfJucGv3Rs
V2ce4qlMwv+hgqUrobTUxUphLF0dYrYe7U3WyzsR+vpjnCbrxOmtT7EvezaW2KmfYzS+Xp6QPADu
m0/g/v3sPp5yzASnqhXIT07y7b9LeC0impa6lykQ6dys5fBb7jy8rCOCd6KS4T7eRKDewOdZPptn
CMxsJrJfU5AGavYlU2KfiWTjhK99cSkDJHj8Jz79TTfTf60+bX2Omr+npkJWB/rzMo1XPpZWSQ4J
rcr5oYxg5JD4LVRx1aCXNKKQdFidwuymWbG+9qpRUboGYkkmO2sRCiAB5hy7cn4vd6Py5lNIwn4J
epVg4C1egQaisWHgwU20iv/ciq2t9WfZFhLW3LJ5Mxtk5Q1URhdPUikdWBsuZJ8CfeZJRJD8SQR/
5plekNDzt9KKBX3JjKU55VFfDxzb4I668tfQXHZmp3OB3S2BQ3oqkZFsaHQbJT+KIM23y/H/zrqV
Irn0F1BN0e6k8TLbYrRm2wNbjwUF0aLUZFLWQVBJCwLFg1LIUGeHn3In/r3V1dKyp9dkGdHelAzl
SITse3ormxWYj3bjae6+czs+I3zMpj/we0yJAFiyJj9QGi0ObvJZV4tPYHHcgP++R8zwRwpMQEx7
znCRRbnE5I1wD/0YDvic+eysErQ0SfDhYPaHgQ/vWCphRoqf+xNUguFvZqDCiw34lSdry0uRdieQ
NMnAp+5o59F8KS/ELZz8/eziuYTi5WrjK/NQPU9TQJd/nl4jLpwOJmIApxQUiOneJ1dZjxHWv5ev
HcuwDNmZjwl3ltcB0Pz01V6pCFeRfKA4MZla6gPtvg9HfvFewByCzjftb9plSf5tZDKnd4uNP06D
/yzz54Pdgj48KQqGQ9yw3PaNB0yxV3nJkE+BkND5kA4LzKw9JgbBRS3e6IwM9ZkKXz+66wJh86SE
ymCAcphoBW3lYuJXhELPo5TKASxOKhHIHfFRSawmOxvGx50UBUi3eevqP9lC7Ps4z2yQIq/0H1L7
zo7HOtvK5sZmbIeY3hNU+g83New8fpMdR1QrYLWuAKawggPVbWU8R57pbqhojG6PAenmLgy/3HrX
o0HmF9G12hY6sE6loIrwCywH1Pz9meIeqSMn4EOmtmvpKCmP4ubs5+gzYiNuoxiQimKZW8nOtuAV
M9WOU/JZt+Y3UMfDNP5e/XFYgn2bRkS904tENQG5UenUOcPQA/tcyVVKVT4dKQopOJwcuXGSrWkV
ttE5+5LknlRXSXNKrpVROe86VuZ0xakrWQSYFeTUaSjqPtsl1dAmANOQ/bciRi1tusi4b7b8M4Ej
KITXkxVzYEuyHKff8r59AhO9O7z2QzGm4oIw/wteyhH0Y839XV2S6fInUQ0AD9y3/flsm/D/Asfm
KkguOgvAbeGDK6Zvk9z+wd67l3t8xLoPymd904L5w1R9szj09Lu4pj4u2yAiPFmswqW2IZmoM7gi
XK76gaNt9MJzib5glsScn/RRuXJKMsM3We9flREmuVZzmxy2PcKVFdENoq/pYUalGdKcLKoGjNFK
XVWBNui4dI6KGw==
`protect end_protected
