XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���.��$Np����8��O��f3Y��Q�?0we�O\�|�����Ls����)@r&���
������\-$�*�d��}�aB�������G����v�}e��p�h�bt�� �M��HD�K̸��ʛ�����D�`���9��<?�d(��3�}��Q�洈8o��S.e��K,�Ff�����gҡ���^���;��B��G:�j�y�:}�sОc��¯����E��ޞ�Z��wx�����v���A)+	R��ƹU_�[���"�[�+��������J�M@�(lU��	rK�9aQ�
����I�ܰQ9EDI;�ҷb�e����1��H7��֨��G�'��ќ\��#�J�]"U0�Y�v6X(�x~���s ��5%�����+�]ZK{s��
&.[���y���A���k�^�6<�X����­r�;�P��</�c��w��jH���s�`��J��L���@�x!o��+U.0�k>�
 ,>�G7wEW#���U��j��7T��4-ঝv�%�ͨ角r��)�Fu�Lҽ}	��2�3��u�}��]Ĺ��	.�U "%Z|k?��>u���7dޙ �/�� �,���/��Lv�0r��i�z�`����
����u�1��(�?mϖE�+�U3:3m���ױt��)4��/d��U/�X�n�9Ԇ�1~w���=!�M�1Mk�J��C�O['JP�A����8�Z�R�M�"e<"��=�}��0#��	 ��OXlxVHYEB     400     1a0cQ�j�%"��w�r@�<������w��~��	�W��������i��Q��%��E�!��=�O�n��l_�Ǜ	�Z����($�[�����H�`�d��nl"=x]cH��I������������ǣ릂�rY�F�:��]N ��JP*w�� ���M�8����������vOW1G�����������tnPpͩ<��b�5�	�O!ȕGV\_���f�xڤ�i3N\p���u���~)/�#�AM�W��%<�b��3���[d$B�8WN��9zٕ^[F��� ���ә�.�`�unl����+-"��z�x�cJ0�֟��3�#� ?�빩XǼ�σ��یYץڜS���0GcV���O���ۭ�{^�dч��}����U�L�ՠ��C�i`$K�h�$L�< XlxVHYEB     400     150�fx���>3G������F�"8b��{e��]���Ŷ�{]? q�d������," �?4aX�E�Ň~�I?4\���T�[#P��D=-1I�o]'0t�~MF?���g�@�aK�=m=Wmi��X��c�q�;U�ùr҆Gp�j29�{G��I�ub���T�a��8y_q <a��)���E��笺�Q��Qή$�P�g�;+9�S�r��ڠ���)�p2�� !��&�1
k�Z�@���,�"�M�-E�rE�v�:b)���V�94���g�g�z�+�����I����_�g{T�h#e^��A�6�i�0f)e�Gz�jSJ;|pv��RLXlxVHYEB     400     190ޑ�	vhy
	w�\�8��A�nT��"Y/�,u�RВ�Z�Cz1�����>Zj9�7��Ne�zf#@���]w������C�����[+/.\��b{�D���M%�8�j�p�h�b��c�K�Y�3?~ƑK��!=�`J �����`�J�#�-�^a"H�B|l�������Y�2&F
������X����_I���$���4y�K��}?�B�z�Z@2�Ԫ��4H���F��W��,~šIh6x����D�[7��&�Rj�7�ͰR��=۷��֨��x�2rwl˂�_ZO�&꿽W
��;�v��~���E��\J�����+\�R��������}�m]�C�9��?C�JzX86��h� +�� ̛��L����>��I��l�6%Kfk�XlxVHYEB     400      f0Du�qw�x�j����M�/�����O
������E�늎�䖿Ժ�Y��%�H�q�??8|�)�E��������Ė��n	���Q��?�g\p�'�z(��怋 7_��"$ap�MEC���� �D��z������y�y��7)�]Z@��O�Euy�#�̰�b&��Rffԙ.�ls���Oq;k�/^B����������M�!�{w����׿h@�$1/����XlxVHYEB     400     120�S��O��V��_D|�d{5�4D�2��S�U*0�#�ߋ5O�����.u�\'w� `j�Îkgv<� u��$x�^O����TBn�^ݪ��uS^��,��"~�`�z^�ԙu�Ԟ��~YAt�}H�X�F
�tG����¼����_?vW����=QW��KH�#	Q����CW�;@rM��\�&h���w��~*�^��T��{%��P����/Q|Bi�Q�����,S�'�9S�=��Ϩ�3#�<��k�y���ً���yt�y�%p�u��XlxVHYEB     400     150�GG��/�آ$(;i��	5�j��G�����j��;Hv|+��{!��ӡ,���Z$���&��X�,y?�,6��1&^ ���߾��N+U-['��DA���6#v�����o a/�}pڞmo�mo���N�9o����3���š�+��'����� ���3޲�İE9�[RX㫴-�I��N�s`�/k �|�Q0���x@��3\W�=Bv�P��,v�ƻ�������_�<{1����.3�.��rGr+�����p%�N�*HN�"����Tn��$D�M��%�r�%ӗ�i�G�wbw��۲��E�'B���CY�j�Rm��r_¿�ǜ(��:rXlxVHYEB      ee      70�f8X
��T�P:��&�g���`�̏�Cہ��n��Ûr����r��D�WkD�8�w���y�X����qa�����9���8�3\Uҧ��3N|%��l6��X�