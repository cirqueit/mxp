XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����6�:Q,��w'�V���#���������8���--���)aϙ��w�Q�#�2aO�U��K`�k��X�"pೈ8�D*t��&�:��oM���OU+u[J��I�2װq�#D30g� nmc߿���H���Q�ͷ�ܢ?-w�v��e�/���A<��'��2r���mѠ�͆�2p;	ۡc�f��#\j���;����X��#�6߶�ĮOq���8�ڶڇ�����^�q& ��m(�R�4�h�"�U�|/|rzx�����/�����6����p��a�	���C�Y��L?�>N��+m[!�0�I_������/�3W���,�)�A��n��4Kq{���N I ��Y�Y�SW�	t��FDw�:�Gw�bM���k4�U���z�&��Q��9-�Ҽ�Ἂ����h��ٌ�Q��Рa9�:�EGE���99��|�BIa��NB	���)C� �@�`�x��14��-���h$�˯Z�@P�@�O���;�'?I�Z��d��b�˺�Eu����W}����#";�ı����/V
֯S8^���Ѭ�<Qڸ�xۄ��i�vAs�����X�yd��L*�%�#7�.囔gˁ��1���6ɹ����~d>��O�+;��zw� �3�mj��҄��np5LL��� ��5�!V'@��� �����|��Y«u��.-�S�=@�̝M'�7�Ƀ�C�Ely�~�[@��&�&�Y��� 群k$A�ݗxyV_8:XlxVHYEB     400     1d0�0i/8��a��<q�� �!*IB�>�������!�1�ӣL,$��"�pД���`H��8��3/	NL��*����%�g8h͖����C��^T3�W���2�xs��a�S���X�� owқ`����6,���'<��a,�YZT�}$@޻Z�����L3��F7˅\O�2ۮCM��Ma�Z��]o�YO��)���S?*�7�D96��Ԥ�� �e�`\���R�����/�3]��I����K�b�0͇VYRdB,έ�ʿ�KW�S��;(+�Y���i�b�VXpt�F?�7 �J-2LW�h�g�����kVG4mb:1�i���� �(��k�%W��<���k���d��r�n�G�މ�t@����M��-)��5���������5\x����Etx*@OZ˘	S�̧,��h��T�$(�� %
����K��	�XlxVHYEB     400     130�.q1�>#XkT����a�m����JK6�UO l�wt���X����{�����6sM5�d����#�揇��m�2-o��.z�H���ǖ�1N dp��G�Z�])qYnrj���}ϊe�b3���U��y�!$�(a����=Xp��Ϳ��8F��=� �zf7E��D�v����V˫xl�Y�{��Rhz��I_vM�"�U$�N&�P�E��K��`X�|���8�����=��wJ�1�08C� c�U��l�#}gfj�>>���Z�!+���X�IR�ڦ �ˤXd��QXlxVHYEB     121      90��JDEj��H�$P,Y�֊[�N�\�&?�#��d9� �/R� ��5��W�����Mucd�ߺ��ʣ�؃6�S�>��@�͛4��eN)o��ⓇiG�-�����xw�Xvfҋ#=ЕAջ\�h�3/�@#P�ӧ?�+v