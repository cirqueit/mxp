`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
9z42N6AweklEvzPy7Re8hzGBM0g+wepOKFYk5TxiVlHNyOv1fhR/v3TMvoaWs3OdGECVijdD8HVB
uBGX89HX3fez5tl5Wr2yQIaZr/CJL71LLb7SAcvpVsAd7wW8wQuJWec5tMXWbfmntzxMKO/a6oRs
s2pyLOiojuoPiQyZzYEQko9WEbyavDkCHyxaZ0m4/O5qIiZjyGvyfbHFkl6dXj8UZBWfFmAhdaPs
cDhGdLFc3YgFDmL7WDVQSpdD6QMk27WPZHX0rFKExnpQws7M/ecTmDVqTNFzYrP38WiZ2U4OVtri
WmIqC5czbz1ONIZGGbD1MUL74wTN39nc5lNm58Ubll0mtwsrk8gULgztttNjz2C3usi6WLPT8I8H
8bKwr4EbjXvnx1mqeG3dkbqMpFwXl6nrOkDhLT+UIIGxQ74rjz9E8n1ojZEFtVjE8h6q3MNiIVVA
8xRd0E7YICmkNB6S+ZICtcFAi91ryo3biU/FkdiOfma2kqQrdOIk3QAOutRysd9e0IN1/JzL3013
23oLGFctxImDxX7Qv6XFbv8/A6BpeKXoD3m8IZswhIVamkeNg/G5CYH1Don0sCPTYAYQiNIt/S+5
0d/ebWgw4zjUDR7qY4XWiwR8ZRG/QkLsksb6pu84ck0NVlOB9EeL8R2nhlf27EffAQnlkJfnu8kU
ktEEPLoS+pM4Kf2umtrzE8LNVbgP4MbSBiATBdY88c0XlLHfLPVm39vybhRSaSfKDmx2p4mdM3m7
wrG4xv7zNZ0TOUnafQRxzXqExF6JsWBbL08RT9SpPbgRXGXYsZmuqOHmHUmvNWfJBW/5Nk+WVOX2
YV2/j69MJWaT8MVPy2iD073mRE25vOPtc6/i/d7bRRISGcsT1XvcYkeeSm2HUU83/OhAm4Evm+UQ
MiKOl0QbsG5cPUGpzqutAFGx4WOOgruNGQm3lcRLnlMwY33+sB1mAh2wo9te+4hzgFcvUyyXvIuV
vjo3SF+K2OZNM0ZCRcg++hRp6XqhVt9FUPu0HuJLWHEEiHNhgsJXfH7nbkSwRjifDQQodOB4TNDO
VOpbkJ+D2dVCWYF33HA9CdgJOxaAlL4I5PjlvXJarjRLXTcZRRHIVby8qSXNaO76tfbkKEYVbk6N
QJGzAlpdtdF2kYpTxdgHiXf4+Wp0pt+2qBDhzmmkj9CO2MuDDUQIqS6+aiXt/ftWg1tG/lQN7Z/1
vhFIzez3zTTi3KJkSFT3ovRMUmV2mSv+yF5NtKZAFmnVCsvcTNmd75zo5r3xF/LNy+fzuC4E9Av4
++YwJgRgoLtGBEVfOcyoMFD+fyi/O6AXZPmW+Y068/gyKikmhi4pmAE4W8ujLyjVDUfdM0kPyOR6
6RrRLUCMy9gopKJLJz2D9QFXJf/8Ky7k4eItTtnPKBs0XEeDae4hQbLQQi5xnRPeauGa2RBTiw15
OKexvOco1ywJ4vrEHxbGqYyMXmwxt9qyL6IXZNueLntrVUic62xlIJVcxiO3Np/m8cmPtXxJAv9Z
D7xYdD4q+J9KMmDTIj/sTSIyQaQtlMg9iT0jBlmKVVzSDo+zGG7qJrzqcbso0e0jontPXagWCzws
g43OaT0Go1Y96rdhcqt2ZpAXL3eEODNOmLUKY2jnWIUA5F+WxH7z5u6ZINNlxfAHyOeZYLsKg4uR
+rXWh7qPMQG4Nzvt02crDlT2Ze0xC62KV2Jzkyip/muYcSm7eRH0pnERPg0vz+qgN0KHZsrKS9Kn
AbS9NQt3GBLaoSgNv/UUy6TNT+LWNargdJ+yIJe574365w+1bkai2A8Xq/Z45IIeKDOvSMCQZwqH
P5gEm2eH0kUBhBdeG7uOOmEWbB7X4COo2b6gRxIJr4TlsJfCji58Sz+vorCqjROnpy6JpAXpzg04
O4uZcq0wZCi+aH45V31xl0ciH2X15Adh6gyWtwFX8ZMLhDwioBgPhgb5NvqBksXyAup9Ydr2AMfB
BGCMRaMqANF0aGG7KZB+eZ7eokcqeKULndlp2k4BGpUI5Hbpr0zsQm7VFzxyl7u/3I+ekK+EoPNx
5hbmkP7zff4YsRbJRbwQN+fstvp25aEecInpiW7DTf78NZtECF7c/CszBHlI3GITQxULnyrBtbXn
j2wo1UZ2hPyqUvRHcQSlE1wJQwzdn+hbP2o1/W1moPLiOdtt8XURLQ5nL2NE5I9vWI6cn+hgqZam
+0IeQf8ynnOGPzSgESubfCB4lJz7UAihqhE7JoQzQFQzkpLO9qY+VQoVx2KQPOs+PXQof2cHeEsP
gOoxhFcgOfzgsgJPvD5H/59+3XQye/QWMgS25Pr1fN8X1MFGGSmcf2SA/dBK6Q0AIcMujAvoULa5
JLCYBDQLGhFE7coZZiMmTeEnAKlrjTgcuRepIrKwLipToMs0IjiMMbMqGz5+exXtFBRZ78f8HRyl
DMiDbYaQEjH7jZmZ3LI2qXYo9BXMRwyUl5AJxT4Uk+9rB1xL03F+7zWcbv56n819/3/LH9m6q4W9
t+/YCy6/TAUa/zslmqr95xXD9zGlXsiT5cVAWzFiEaz4ECtAxv5tLBZCWR3Z1ry40lD3depqO8Aw
bx93voqyJT4ypW3L7Wf6gAKO4LikKqvocdJiPTwhK4c9aCjFj3p2TjgK8qSkgANbn1em+Ge/qfvu
vR9bvexuZA9ezelDQf1zrxqacKfC8tzVtL53flYNo+9tax51cEEEE8d85l+BabCgEMcAVhHzWwtq
5LgtOlQId6MoSXf6K/o5WKApUH6IhmyzuRMksAlUZdjZadkz2UZtk1WygNw6URepwpRL+T7jrsrC
KqhaZiSzT3AQUzHPXYHlvpav5U9T9cWP621y4Wywjx4SjqVA0ddEKygsmEIVqhvNesH2BG8zrmFB
xsFHblqGpglmkMEPq/0grScZK5Oj5GbySn/gygd5a58265cOyFwhIcXiLSgq3XywWOUkeBa/pOhG
JmTab1DgxyTCdfldGErmSb5xXL0RF6vk3Gu3WnI8oiyL3ZdJty4DtCuT2mFSpbRJuoWpBLfU0iRj
+E9V5LVKnAH7nizCZ1TeROdB/GAtxW7I47z1s508Df4xm/mXwf8hUw5OgCm/YkftV0zhfWOxjS1c
ZAuecD6oY8MuLoa2/Ny99Gv/bfl3xr7WgJhcubc3p+hZhTHGTjmq8HUJiCXzcf+QKIiZvzJ6Zgnh
ASb7pcf9Ehz7Jch4NP/WRdQmQzwBHii21Gz5CASKR9B1cumDk4YkkNNULp0VZkj6SqTZsuaQZDDq
lnPIBQIapUklRWwyu1DT0fqH00FUSTAW3ZlER2NF/u7gds+D/mWIEyNK2xAfV4VOKjA9+l0x356s
VBg5/o8kSRBhHXIAIK99rRKsuQ+qKKxdyuYSOEgDZ0O19U/HrgX5a799oIuYiN0Ok/Aab+Gw++k9
BOMWVzasGtOMNaE/EP7MhuMu7fWbc5H7hs8vJF7xDwzygAE9zurPoh+gZGhmbIik4wJSRhxmutRg
wGdR6ssQWacNZV6YnpiJB+PS2EJ/PQZKDFqaxCRwnJLZlPGWeSxwK/GkPSOLuYbQXKIo9GuKbLlY
Wf9aQFoe8ehcQh2DkZfsHrCu0F3mYVaB9dVkhLohHkSOhbfYSka5775GMlII21o2WRlVK5wLVYAG
kKteNqT0GENw74Log1uXmW+3ldt6d9R4UPDICX/8njeiL65/7eWKAuESIZwWRxYYig+0ksnrT6Nk
4Q8bU7tKojlVrQ2bf/mc7Y6IhtLOPUaLPQ83k7cCbluD5P5HuhyJTZPyZpWCPLD6ApoLCLYAUust
tTZb6IEv3Iz+apnP20NkBVGymNskmuc7rYLCh5aVBn0qbZFn46qNZx+2/E2glHmSIKf29bsjGVxC
syqtNVPFZ6Y1nyzXGA61Ud+V1/OaIrDY1kfg0uYWfBKlrVoLy1ETHxhLPRd+6lchf+ks+2iOhXG9
Fm+azJSXamb1bXNkJuJSTWnwMWjDv+mqw/VCHl00EU6/b161OzuPjWP431GeJN0bYDmPVAjT9kH/
kwmEjlXUJvpYuOjBf5Fv85OkviEQTHzVGdDHndfCf1EW0uoogVY+cItZxVD07rdSW4QtqG5SEYXk
0/0YnepVXxp91MPnLfGoH7gtr65uLbWelmHdRpr30YqgpcmGG77KZEAfFjLzZgfdCyCggpeix3k1
dcIjz8zKS2xuJF9VN51J2r7celCAh/19U0Bqit5FPdO86syGW+mEH0jxPuY1YswSBXqmnk6T0KBq
AUrrf2yk9rduQEQqyPyJ3p8lCCOwxZ5fhmslPvlwRRVaSG7gLStAvz70SwuAiKnSt3qpkZIhHBO7
49nS/QndctoCHjTDnG+GSyOsc3GU6jVONHq8lFeDdhNvbN8N3elhDOM1vo4njgNLG1KbUYI4uV37
g/Q5PCEe6rNa6adn1UdKey+velRSippb/GPM21e+OiYmaRPOEU6sYWCMmXK1RWwWSVCzQZi/w8pp
ykqOHb+ZoYN1BNNx8sut3h5P+qDM0fvbi65zjJti92bnvtqMtKa3hWB8p2sMpKyziT4EO34IfeI/
ZzTDhZH8WN2Vyd2nQZ50L7QLIKdsTJUifRJ/dBP/hvR7Sb3Le8LPLBGnL/ojcTgfMGvcM3fwTtdn
syQlluMZ+TxJt+STV5xux0wiWnh0FReQydxETW+ntpJ0w569Jo37XIyDK+tVi7Wg1kwRU7aiWiZU
QTUS/pQpoZ1Mu8bWHQanJXgVUYbAO7t51/L1huLm66dHhm7UhOmob1dhtVzAyM0Il3p1qSKW30eS
q9KdETkMZqwwPjPcIHjCV2qAP9KoQ7sPxbsbZrADhEoMgK/Vr2+BxfQZP7qKKj81p0pJBlWZyQRU
gKUEWfWTgQ65OUno35srmorr/MX0IiF+NBhTWmI5hlUKytkJUYPlxTjHAWwuyMC1wdx/np3e1u0v
V6njkVrgTmG7sIqx/cng+f0j1pHuIQ0ZI1SB8h5A7QweIVUcQJqYG9i7EvkwqWwgjA7LOa6XA3Xr
VJgcGY1qWLiOKcontPxGbCZZeKSWl73k9LsRSV4a5KZe3il3bwIoxh8yqeSPz2NMTKcO7VwyXIGE
0N5zmg8pLX7A5Y++vO8+X1Mhcb0SIWRGj3u7fQk6A30Tw18lyqJx7q16StfyHrtgMJiUWFPmf3P/
ckyG8REqwe2wICOnuYmQlaq1B3KY6IyUebhJJi7vq1pkwjyMAdBYY6yP6Z+3nloKVX5+1aDKWCX4
WiTHYUJ4hrVAU5bOjzakQy0O8fSlp1rJ1cDVvLc3J65nJsJaFc0MpfoeSiXo8HRxMAHfr9b/L6tj
ExIS1YD/pijfle+TSzDzWdD5HJWuRB6uIRhH+Tkf6kwSgQpwwqbYzceycFkVXoyuuZaGmtqSAaRY
ETXg51NgfTKvHbykNrx6u3pSUWaYYcY6vVaffyKe5/lgFreduaxUrwdLBzaLIMJ43QGlG91xLG/C
Yj/Zk6As8fv3NhtR3QMqR7U9hP8h8TMxtMwH9ThqjYKHExuCwefgRaMPCBUKtuPcaw+RZEf1GmOT
dfcGuqVJTESdgxhKMFTRAjfl4Jlz3Si1U/UFJDdB98YRGhYLMS2RaO66pvdRx/v/PKu7Jd81Kji+
MLGYxBS6/F7iBYBx/rqQjhrDx90zPFZf2JPOeAxT9Y7GdXNAV1gZc3G2zbuX2M7lUHQ56/zeB3Qn
SWUHx9SV56TN1YdZeN4FbMZnxzSW6S8IRypxANGbFZcBoqCH70Cz02257gBZbyJqnjMpd7MAf+hu
WkFxEpTetc6lbBIL4fl9kR0d3qs7CL1GURLpkX4gQbX8OdQL9ANMABEi/pIxKaQ1zjaJArhcpnVu
T90rJyPBLjm4lMUOsfm7LIFbRKi7EZP8I1cYgjZCaW0MxZa/okXgH01gb03ibBLvTkTZdsA3oRFQ
CeHwgr8leNrU82m+yIToAyOMNGPRftvgDk2TxCtwTiRkJjgKSEuK6idf8+6DHyrCKFUnU+TPuU1/
+kTOyt+GSf/AlBLSYG5+61u3Gq0ikt2lPQu8PtMtpjkODgwuBKYPO4NqBJO2p9oXwKt64Qda1XDD
cKX1lqRFkc8c0+eUqFMT5iXRQV7FN4ClivCPYmiYyZ73zp+4htU8agZhRPJ85emK3eK36flAELGy
ICYG6wohKQNpKygO1G2Jk0DgUMJ/bm78QPEDyp+Ai0+iVytvwrSmVoyhTpWHWojKvLfMgi0iBQmX
eBYF3/6gPoVWqmNSP9upfSm0JcUEasvkqQCBj+LVGbMHSu8dPOyLOnU08dRVCMqVVtrvcNZLepC5
CaXX+yYDJe/tqQWPR5FM01FgXAVg1XPaeIkQeI2bZHn5rHZvt/b99kGWw8xNvtskBo/XmiXQymjO
Y3XHbvzB4gVwDjBt2uL9Z9oc8AP2Ke2/S2L5C/ibA+7ykMoHBBQZBzQYf93DIk6fqLbBruvPPBC/
9Um5KiwA+vmnuRue1ViO+toenzUGslI1PLakU4CmF5qcrOefgqsxPRXhFNC432BJiRoJd4XRsxGi
tfGyhUR3Cy+RVFAFRRyadZ/+PW5EQDFeXeuejoCYim3QjX0tn5CNX6UNyR8HFSZ7b5w2OM9pGuDa
uRB9ftQtBv2bL2ItNjyprwCJk1hajjSHMilr7eU26X284YMN//1wERsDvWnE9kd/tjxEqcn8SvFa
B6U89N7t7KSClYOI2LU4B1LyGBEySKDryHsXJGZWlfEt4L0X1cpLHZGZ5YV+dL+pEpDDJYEa2ak6
+ypW4e2z1BC6jYQWHnoiZzL5gQzVziqHuKeKBkuaBRp4Bg4L77JlsjVJ3VgrDi30pyQK5j1T7n0q
JTACI6KE6N7D1RjDv20OFBX5cChscTH+5FzR+/ym5dTkeDpj1ZmRheXcS0ubYYeXIGsi5IWqDANS
9zl7zmuMYzuj7xHl0pAm/7QJHqorKMUwoYbu90+HnQ3Y15Cov0AyY8ehdE8xrdLQxhLlpytAg8ut
Hglkpga92M/1VQHSL2rxRHo3wdiG63REfNQOw7etb3ZggTiJq0kkLwCN2g9FARV6ReRl0BQIEUnU
DfSxzTort5ZHrnR9kD+2WjzJhZzYHHn5X8Mtu5DW/KL8GrPr/aoL8HiW4YtJsHEibE+A6ks5QtwI
0wAFLpNJGZhA7Di75vIdFrTxId+/CI/Kzwxp/nJlo5cvXzv1u2SuNEZbIJc5wgXecpguAXt92OcF
Kvxdzl5SgKJvpxTmUaW3bctY8G361CtF4qwugfr/io7t+C6kK0MrgWbXBw+UmMO0+7B+R3vQ2GFE
4TkDMNFZQt18YRlBB19dpLJxhnPQgrBuz9cXHQx8Lr/ALBwJlguuaESnwd5ronz0YGY//zfnYLUg
MwyBmJifjQWKINjiYqF/ccaCUIriRDllBkEZcSPxg+mbA9NjIbmcOo5ZCD2m3V19/AIzez/0Z77e
QKn54HWkeLHojlxUBoinzugYpuJrPhD4t8ZNcwWR0B1YuGvS0T4/+GsKE7ysPZW5CPv0IgrpQJ9A
25sswH083u8rZjrEnDtSKXx3Ks211ZunwRLHDFJV1F2jqH5NY/zAZcN+lSoM0SbN21Gk47GskMcH
hOCJ8n4WcBxSEqDPjdDSmdBdapA9Zgbz0IATZvNUgNstJwe6n5hBcPUOE4oKyIM5ZuhVnEuI1SvG
Jket623lSeJfowZi7Uk5WnbqAYGd2sSpT0zdkNhWy1idbR0c1ksV+WNQpQWxqL9soXvCadwa75h/
Ohn8nBvvAOwmcslptil8y60+pNMTELkUFeptKK9pclZDg1D1eq76/c24BNU3BbDdEutS6TUbk2wH
S6YgVHMsKSuymJMQtWO8kbuGAFh+twLSdP/KEJ66YAsM/IMQOp3Q4oLI/Arntxpts2eDHNqtg6FV
n96rES/mpUum7Yf7weOU1Lrccg4soi4zMR8zBw83Xv19dbc5UenrgN4F6oIyZvGpECUSuJNC2e/1
u44dwjGEoCvyfsGyLT4X0+ncJ0cRwgK5p0eNbEJDt5h8bPhbvbgQ34C8FrxV5+oUvPire1c0RZf2
3Iv9pci7kpzXkMny0VYGoqBL18tYodrWFvM9GTtMKlgSg4nGQbHCzSCps2biTucNuavT9Z3qh8eh
OqwvxGt4Rjguac2NJg/c+6LO0s5IkKPAyRb0DhIt//z4ohIfCEVQZO17uCGXxaWcWAQJLbq/pu4y
cc3i3pl3a+3QntLi817s2jsBxi8bR/Ar9JXKizruIpHl38YHtIyZ2HRw8vDTxxUgEFGxALf7/21G
4tEtnmZbVnzQJLfBLWfZ6PKfWMUfSEeN9bpvPRcsV4BC9f4NUZJdMns4QoajzGs5inTF57QiIuu5
RwipJxQ8wFnpRU1rO3LBdy/DaVzhYlErFNC03hmVy+NmJIA8DcKJ4W0s66n3mjCObivJDzbyLSKs
ejxx8GPr49BDpmB9nOhzi4BdSkD0jEkDwX8MGWGXpyGohEidMh4Q838xtr2LNq4I6kRZD9cpLHGc
rHcujXgjci+WoWOT33i5Jw==
`protect end_protected
