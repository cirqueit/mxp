XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������d��*�$.��Ϻ�T��A~���%�<I7����;m��Ծ���'���w�M�Ë>$ d���8	ܦ����!�W�f*}Sc�0�0����&��6r^+-��5a���N�k5����෩�FgĜ63��Z��K���ǅKW�n9��x���Z]o���r�HK`�S+��?� U@�ֱ,����o���g���^!>��w�$Y!��|��H�;�,ݍ���%����l��f[P�vy0��\�!�VSV�N�����W��]��LY�
�蹑��	�rcQ7!��eF=��X�PqD�$�ӣK���n7Ű$�%]�J�n�"���'ܥ�fe�Cp' ;�w4w�#ɔk���Ďd�"��׫��ױ��̀����:J�{���!�K�l7��l@��͆��ˈų,D�����%�%NNJ�t�j�*]L޻���Tp�z�[P�˜�T�d�ٔ�
���u�S�����Ūi�w-^���'0���Ր,A,�Y�9B��w��=�bx���o�����+\�}&�4�Q�ӗ;��l)|l4}����[�쥭,Y���\!��/�&=1.�[�����,�<"w��uxK��m�K�<t�l,O�����<��[K�S�i���n�Dk,��G9��
��t��К@�������(��7���cb|.��A)�=@���|5iL���E�,�y�O���6O;*'��D�|�F}j `�����hanJy
 �0�f���-��XlxVHYEB     400     190��>U�y8�v<�����ϱ8M��p�{�������o��V���D���
����c�!)�̺+�9{M���D���iW���fJUj�I�Ȁ�%����Fg�R%@7�:h-�y�L*�D��.���d����Ԇ��L���}��ʌi`�����4�ܣks�ZE��Ȩ+/�Ɵ�w2Y3�nt���;;(L�`�iM��;cg4&b[��]��r����um��Fs{JG:g�W�YS���i;���G�g�"hq�����הZ�Y&2�B�羵_�If�0	��0_�s�2�����Ϛ�z�j�~L|����Ƥt��W��֔�*��oDMx��&��k�-q@K<���K�?���H|扌�����LTВ�­���{�7ϥeXlxVHYEB     400     140T�_Z��!�4.��%�#8FSfz���d�5e��AC��8��tIl��o+;`Vz1j�q��*�zƲ�hB���w��Çh���F��ٸ�K�y{��C���b���Q�@�↸�D>ez�ی!���)�3���c�	�w�h���X+�k&0\��:��2�f
H�Q����2���F�=���O�f��j��7���9���Y��ᘝ�/@,�:��B7yi7\
ڱA	[X4{'�fw+��k��6L�ǯ� �	�NH�V]���d��V�Ic��rP��C��:LB	�����XlxVHYEB     400     170V10���&�����`{4���Ǫ�>�'��|����g�θVx���D�>U�֌��qϣp�����G��y���y61z#)ijT����j�'����!�*�&�v%�)�T2� E�S#�
��KI�4�M��p���%*Mu)i�����'Q�!S��}��YXy�p�'�����uDA]�~��4�-|J�%����?�G'�P��Oy&@ +���̩ί���c��Y�FQ���lb��;��u���b�������:.����_w�!�b@�pTJ��+N�9����d1���T:&��.�cfPe�1Ԛ�\*��A@��0,�3�����orK�����c��x3Y���i=��� ��>?XlxVHYEB     400     1304�5�5�	2��*#�A��o�ի?�%�����nA��:c�8�o1Ì��v���B���}q�S��Q�:1�9YT4��dE]k��H"��\��C����.0c%N�m�����u0�s����8�d��G�mdRQ<�|���y��� ��t=�3��D�)����}Pj��?��eo*!��H9SzPfo��*�?c��>���x����@�C��_��XT���.���:廢�eSB ��JR\Jm��tYK�0Rʱ�!�Á���?��]߾��o��O3­����������'�@Ї�����XlxVHYEB     400      d0 ��e	A�&;�]��.���U���/]R�(r׺W��_l�!]%��Q��*�1���i�l6DP��/a]~�p�d&��F�b�c���;)�i��4!�/���"3�")$�	c�5+�XR�� �V�Ph�}���۹�eX]��xd��6O��z�*Fe��׼�9�e"I������)_�eA:�'�,7N�=/�=M�$���l��XlxVHYEB     400     130�v* j��M�|�[,I�~�W�hѩ��O�S\��կdљ���~`ʦ!�M��%��/����ܼ��f�4{�n^p6�U#��j������G�5��]#r������6���� S$�Z�~e۩�(��6��M���|2�
ɽ����=�+�V�g�U-�)��{��Md�N�'�G6�����ǖwkr̸��Vw�d?�0����q��;��?���H�C٩�S�����z��%��B�ŗ����9�ӭ��ܼ�!����'��r�s�3��:(�:�S�5�
:�a��&IM�K���XlxVHYEB     400      e0���Tx��(s1sb�����f�-ѫ���hQ.2���B����H���q� @�h-u�n���4�_�̩�M�)���J�]�~,8�l��䶾�l0F�M+��-7mQ����%=�=t{o��_��4������@���>Bx�^���;���:~]�P	@�]<>^�ׁ���b�Y�G�)�K��m�VKu�E�zx�*����[wfQXlxVHYEB     400     140�2Yb;B�y�o͖�`��>�w�N.��P�Ҧ���'8��nI�T:�ф���@(R�*���iG8_��b@��d�{W�&���H'��AB'��=��D��1�s�V(nM��x���#�j�pT'��r��9K-��+�4�SFZ����V³@�N�~���0[,i}�h��<�X�ɷn����Y�8d�`=8v�i˦�9����K�'�����5��GT�l��{&�Y<#;H,��:'�W�݅dI�z���D!t�k�����֣�U_�<�&E�@͆57?��e���8)n�UF�	�����x2��6=֔�XlxVHYEB     400     180u�����SU%M���9�,�?y`۔1H�9ϋc��s�\
�����Շ�}�~��ɰ{'���4 5�c�-P������â$��R$jg  �A-+��\��4�?(�ns�L<	*>�yߥR��ͣ�lV�еw��Crĳ1ݿ �}�Jl>�����#��M%���]��W��q;�����ؤBp,�͏ɧe��v�-꼪 �L��>�ʏ�Z�"��(��4yӡĳ���>10��?m��d�P�R�@�MF�$O������
j��c}����f�XC��mƄ�4��v�N8���9:���*�0��T��X$�!U����i�ҭ�4�`㶄o*J�ɴi�G���9D����k# �&��9�⁺C��=�_XlxVHYEB     400     150����K�6��d���b(#(m�E���AV9ʧ�~��A�G�Q����w���ݙP(y,�ۿ�5�y��K��-�e��n$�n��x���`4+^}Y�nI���
�H�uIr5l��iҎ
b�����Y̻�9}% ��/0Zt#u�
��#���%gp�,�J�3˺�ԑ4'�vW�$:B`H�Y��z�-Ď*�PcO�yȘLVε$��y"�B��wÏSftsb�:�J�]Yq2��̵=�ѧnz����;#W��9�!�26j��-- @0[�ƃm��̘�؋�3 1)�!�r\�^ZI�d%c�C�aڋFK8&��8"������\����)]�XlxVHYEB     400     160�R�	��4�"ح<>�f�f2	��:����3���˞v�W�(�g�8�����=t�q�����`�k�Ů�A�u}E�9^�g|뵟��);.�N�i�J��E�Tf�L��c�,�	Q}��7a����5����3"'�Z��
���ȃ��Nl"�)`���2�_|�	����=�Ġt2\ ��.�<(�)��سWw#�S���n`����������}�[m�t�&}�#��t�|dlS�O��{�~#a� �waM]��V\�zw�+wu�'U��5�y�/9��c��~�U	=�҃N���	��W�3s��υ�r΅(3�aΫFuh,e�|'d��(��\�r1�ah^XlxVHYEB     400     130���vI��I��j������	��SeX�G��"�,ye��\sS_�ƀ�&è!��w��qs E~��?�]��EA砵@�5���e�,�?Z�z�}�q$��zŉ�9���
���cIK���pd��v�d�_@�X
.�?�2����ga+�"�d/H���<V~�lK��*���Fux�\>>�.o�ő1e=O�<�e>��R���,��w�EۀZ@�"v��~�i��7"d��e�Ӳ
$V�HJ	`7x���|c�<a%����5t����E���u�l{����bױ�~�VC	��SXlxVHYEB     400     140��D�u�P��ǮF�ެ�;�=N��HD�q�id7�sA�. ׫	O������=�)��Eow�O�Ox�����]F�5K,��8��7��&]����[��#+��R�	e���V��uʟ����a|�<��2(��2r��ۙp��3kK�jL؝��L�ם��Š{�7	��8��tݡ��䕥����}��pHvO���y;ϊ �������E��S<b"���|���J	��u@Η=G86����AR[h�>8�`��G.猙��8�H.Z���rN�����3Wg-��b�$@��R�پ��ho���XlxVHYEB     400     1a0�"zf��<]�M���j��|FpPkî,���%r��P젞fB�n���d��73RSźF����ڮ���p�l	hM��9X�d���)�����
�smB ����EQq���ͮq}���x�痎ό�l/���&/���c�� ���q' 5cX��+�;Ej��AP�U��˯ioD^y�9t���s���6�q��'F���y�������4(?Gd�lpAhC�n���U$ʍ'�8?!֝��˕�,��/�Ox�T2�|0�H��7q��g��4����d!�R�̥�]Wn�5k��7p>���B?��Н�֚�I�P��S���<�k\ �Z��828�,t"zq#���=�}e�GiRb�N@W�][��n5�_v���>5_���iR�&J��]1y�mw�RYqB��Hw�j�木+XlxVHYEB     400     120r����Xq��rT��v�D�*ILj%;M$sε	�d/�6i鮕��J�$�o�J�)Қ!c��d��$��I<Pz*���N��3M��;b��asO��r
\Ȋ�^VBX�,�^4� �W�"b��	����b��A�.�|��L4��
�+�|A��b��z��ʌ��fn|�a�+>	^}v `,@����<�{���D�r�?��m J���Z!�Pv�R�����q�Y"^Ղ��5�c�!�dUY3x��*v������r���Ħ�U���_@�ؚ��nc�=�@�wXlxVHYEB     400     180�~�V��$��&�]��3�v��m+�T�b赦�56c�s���L2���^�F�Td����)��C��H��� g��>�.sM;����7S�5b�<f�� 悅��Ğ{���3��m�;9�>SC�J��y��.��	Y���&L:�rb��.YPx���u�/�����Q���ww���W?\�7�X�����0~��C�̎��]b�*���\@��tn��-AT��ul��W�-���O�Eң�]6�2���A���~��K�N�����i�YE�3A�;ݷh��+���M�A�6�,�x>�/�ݪ-3>|��w�Vg��!��D�}�O�ߏ�<��:ɚ2n$��MWU#8���f�����f��c����RSW��C���³D-;�f3sl�XlxVHYEB     400     160`�@���P\!�OfQ�K�w��Yq�2$M#ƨ-�����	�����Zڧsc�^�_+g�e"?���Z	���^�8#�����f�J��G�%�DF�
�?���zʉ;�ϝƟ����K�F�-T]��z�)_�%��'"���/�k�����IL#�>iw��%�������!e�+�i��咺f�5��1T���R���s�2��]1%�Q�ou�$�jF�߱8��ܸ[�;ÒZ[�{|��<mdRF1�$h�n��F��">D�K<V���RM�j@E�u��E �z#K¢�/��ߜ2�/A!M�����.�,_���G�cu<�@�B�'�VCc�O�Jk}p�ZN_XlxVHYEB     400     1b0��X�M�B�+^�R�%�i>�;��4��(�C�>#o�Ѵi�� �1�XU�*�z�z�z>��E�d�����Ӄ��+̓�Tلk��\���&�)��=<P�WgU�aJ����drc'xc���UbڢN���q�!�7^=��=�����7�B_��w��!��@�A�N��Pu?����=��KR�!��$b����5/c�v�*�By��Q|S��_��xQҥ�Rct�L��5JЄ��DC�8{g�6�V��?`{�߻��V�Y�+V�^��r��8]�\t�3�U�0@�7�%^wJ��7�d��T��O�������<��3`$.	e�Q��x�m��ш��YAg#�#>���FQc �3ґ��UD���*�Q�n4�g p���n!r	�t����/;]Q!#U���;-�xP��a�L�XlxVHYEB     400     160z��j-_>�L�J��	[琢Qs˷�	$a�%�{h�K�&�[�9�Qx��s5�݀��	��7x9k���ÿ��1����[Et�]s*TuS��,b}��#V��ҡPs��w��̨���^Ur�W2މS͙�3AD��N����xAݵ�y'���=J�������Z� �@�`�_��ˬ�6����(4^ecA�Q#���H���ǌt����e�/���D����O���/.�;��qB�W�;�AT�*�����(�q�@$8�x����o�e�r�L`"�~Ր���$�t�1��Ԗ��P�a�2� <i�-���1?��=��ə�T�k_QXlxVHYEB     400     130�����-�ԲO�U�wUm����B�<@���:�ڣ]1j�&��q�$�:C�{9����P�T5찊/��2��a'
+�w�v�U��i����t�z�|(�d����z���|�C�IH+��g�����D$�!\�0��.Dy-W��'��*����&y�ms��$���`��yrKS�����7-�0���ĕP�x��7ss�*�m������,���FO����*'b9EWE��%"fK�#"�y:ҴMHV��b�I�����ܚ�!�_ U�jF���%�D��iv�����)84��mXlxVHYEB     400     140]|�G���X�q����`>7x�8r��M�Z	�_��R��I��P����uP�1��o:�c��Q�`΍���0�pO�LPLڜ�c�݄����Eǈ�a*�b���x��^��s�;����>����ɪV�'���^�y��mdw�e�ϒ�b �R�s-�T0/������U� �u:�Ə��_��맩�<TeǥX�"k�cr4菋O���0�N�4�[@�YwzUp��y�}770Ϝ�Ϡ��D�ü<�{QE��9p_�g�,��1O�÷�}���)�&U�;9>�ê����h��4�D6���F��^�E�i�;�p�+XlxVHYEB     400     130�l��*̺
�WN�o�״[�����)��1&���/>���ؙ�QL�0��������:����1���ջMVS�"m��	V+k�3V_(�
mT�e�8�,d��We�bOX+L���w����Py����l�91�~�  ������e���%7C��k�ٵ��z&�
�� zP�qc���\OSqC%��U���n�h�8;�: ��
v�j��s|�77���]l~�#�&"���8ڣZ+�7i=P�h��PH\�h��P�ۇD�5f�>���uG޴;��f:p̼�{� AB�0�_4���XlxVHYEB     400     140vz<U��H��M_YȰ�8��1��"�x%N�� V��O!D��S���Đe�V�ޅ��f������� ��L8�Е��f#�H���dM#�k2����d��n CֆS+
�-�:��\�� �e����Y��ػ�e�C*V̕����(��-���`Ch�Ty�I2��}uA��R����G�\����&Ve��o	Zj [y!r��rV��۳�8�Q:�d��[mz5�l8+T��� �^;���!��Q%V��x@��x}�^���X`�?���lk��<k ���]�ʉ�'���u�����0c��Fk:I\ɲ�'��i6�XlxVHYEB     400      d0Q
�qJ�I��D�S��g�>�"����O�2[UL56`,�5�����u�����Y������^g�.7ch�Js�W=��6T��[�?�hA�4Z���n,�]���sV���j���l�]���s�����ꌘ�4\�J�k��9��6|�d�Z�nt�q�?�0yo��6��Ը����c���9륮γ((z��f��o��Zs�i��=K��XlxVHYEB     247      b0�r���@䎘�c\.�г� �e8�U,�v�^e�=3E:�-�Il�����J�.e�v�N,�`���x�3��X��=x�Q=�.�j1����#�qb�!�=�:3�GV_z�E�)a�;�
�L8&�`)���κn�8T.�U��.B�l��{��a+r<z��>p�zh�i��