`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
SCPuHB0FFsDrSzY48QmCu6iQWFq0p4vkh/4v8sumfmD+/0gB9nQjqvqx4G9IZ6oAVSFns8Z72MFp
/EC0xnazsHDWZq0WnFyw+MqL5cYVGJHYCD9HsWNI/KbgxW99fHnAm5r5MVb4bcOI8D54Zseiw71I
gwzZBMksYdZZy/NBemo3jMCzL4AWqubHmdLFFzA9iffF7Pr9Hle5tgS9ierd1x5pz9eyzClQk0rg
aL5XaV6fiKzeVU4B1+lgG7dvp3tJtC0LuAWZr8xMtf4kB71SV/eVAYpUfvFGC7SbaCtDVxGnbX3W
K6vK2w1MUdxW6mSwvF+IKQj2GII4Z4QtOyMDDYvZWCeTynacHBfANhytRKgljm68dZJkjVbWNLKP
64tyK8Wclk46iL7uxA+0fWbOD9Xz1GGFf06cJhlv05QEoa+lLcMxq8OCPDFjOluheb6zOUvzIM0t
X4zBnXvGugv722BzRLqfslZNC4W04QUWqmypJYVGgDHrlFE9S1+nzBDp77OGaPPixhymbGRVkAF3
z/4CQNFBmaSqChKjZqEFRiiXtEWQ16OfIjJ9kn2ApWAZ9Zf/RIg4bWtiE25q3tmpbxGlbULhwjrY
sU8R/xloEDMu4VnSZuOdAcTEfFas0rVhM4Lq/P3GVhtKYRDsDry4IB6Zdc7lHBJi+0QKDB9pbxef
uOeZB8OshBuof+aT+jpA8Lvat7eGXxSTdkJtNRy7A1m/WdnRjKDjkN+0r8Q0kS2D5usSGmVpmS+V
/Of4qQnMnJrUdceHpEwjCfslP3NjQ8Ye/8XltVghQ6KQj/FE7i/vBiwNc0wTTq/B3J2xc9NByOIq
z4ePKJV1akyJFWdPIIeBKxzC/CXvbLU/H8POyz1PICXN9GR559RSqr+6wlQPMcDbBWaxVnik3Zwq
s6d7BtD89eyxuQmFc1qCu0/Rh8wHRNSgx0r0dFUTHobS3fxu2bx7uyuwOL4prJJ2p2lanJvE9B47
mY6y5NA6urTWYq+uX0IxGOLYXrpU6xrtreqrsDh5RO/jKJVnVqys3+fqeiD111lftMfgdNPaeemZ
DNxOFlSM431mQQEf9iTCB2MSRjcUl/qS1cH/9zzvcn5dWnLLU7Zdc95J3WLmNgIteBQMTY+nOE4C
FiDj95/kAzyksNO3HZTu2v98OgjCFWnNBg86j0l+8Yya7tUFh56pX7hZXo8Iq+2Yzvt4m4j/ICEa
rlZ8enCIyvp6nzc5tOWuGMtqfBu6Gcsfz8d6g2+Ee1a+JSIEad4Y+R3PJ/ufArvGQbJqa/+tdIGF
ZYfXXA7DnJNXogn1hYBOrkig/Wx5qCFyqJjtLr+NdN87hKTlP2Fow4f6W7BuAgiI/1FsmezjFqk0
AcNmYXAxC3Ojy68iner178fe2nmBnA9n+6/BXtuz3I4297eFZgeJLDwQUDV1NV2L70RwSFBJGgR9
j4LevEnpDz2c3Z8pghtp5kXE8lhF1PXvXc4+6iynYwgRdLL5/BbfCQujOab822vbQPTdXrapQZ+r
7B4W9XPBm6NPxUx+yj5MuLHw1nZoGdikg9cEnYTAtDp8xES5uvt8rQ3lHaACsX79D+UY+lvGcCbG
ftI+V5POG0rrzO3JIy/H+FsjoWldq2GbfPGTIuXXDnTzcS7TP0+jTE6BzllfqKo+3OfxUJEXF72a
bcl73XIhMdCbdCdHEVmJ+ifZFoJDfHgRDVG42OPKsLftPlpppisWKJqxtRs5vJEvIiIqx1arbdeR
8/Uo8UPuSbR8WsJBFAYQKtRQ/NYxm/yLtdj6cr9sfiAykI6rUs2srC34dvWWOTMe5FbEIK/m7y5t
gaG273ZTDl+SiYuLn86Hm/QgFhP8ZsXTmK+uuPEMchmG3KkGLx9xwfayTddm6oExvRhJg5qSdQbd
2xU79DrX+UWPSXeSQLhbXS3+YHVRoRTuTWJomQCXIFmyLVD5uQdaOFOhSfPVKgpltGs1+B5dgk54
sDe/WY31TXrmwi2o35nuGUlcy7vZSjYObbEkoDOEonNjFMpVllxLojE0o6K3dd62/GiLEav9cJ3V
Q3hxkLsXNHUiFsI/6QbcQ0nAMKIETvtSW8Dii2uk7iu8IXRHLyof9zK3gtnTu/qyAMkQ8Q74M/Vr
0tYNveJSKE/uy4QuryznjFtBogwcOfDO3nbiLG2/KkCz+M2CzhOZH978oz6W4+AI/F7qlr8FFZ1G
d6QYbSUUnhkgpYZK6QRZmj+0Kj5U/ymq990FCUjcXsYRQWbUW6Gy6lkUqWHJMJcIvu3fk0ARY+gs
nU7jSpaOOZFPcsNbPRK8xOFaxhJW7OoNl6yMAlTIjWbYQmwtKwi9bu4sWz/wRArdusyDFQ8Pow9g
omPf5/LKfRC1Db/eqN0qiOIeeu7UmyW1UTnReV/fQB7qPa9tWDw2wZEZU/BpsVzBJLpGWYtbl5zV
IoNT7ITiApLGQzF6tI5euRRKPK+NFcKHEslhu5LRLi2LfJ/lFqZ6NL+5Z1MzWTcc24lnOhNleqRR
XFSW7ir4aiySrYrwzQYaDX2U+ZOYr/IdixE1DIaKLiuAT+LQ0gcT+o7D3vo5q9Fv9vJuGZdpvBY9
g9+aHseiro/0OzD9VCb6NCMEcZZ/rkjYDvF/fnzqx8qeUSJRU57C3seDDrdvxcX4/aZ02VbfQp+4
bFclwt2htM6sHkILzZrUmAyhA3VyD0qv8647dcL2xNX/9XRPvnypn7qlO1rc0N0vs8ZekyCH8Qgg
NE23NyFU3m5KLptBuAjfIAbNHVT81Ss8oGnmAj8qSPZO/XWl5XqbVaabqoPWx35Y/w05jCHEhh0+
RZIV/trG9iTI3WSZMklObpC91UzOj1/2//17Tq2234kIOB4gPhrpB+UKyW6o9XhmJZNgCIhS4rcz
gGajMqmQTXihYFwuLRSWSH0chTDLqx6oCiRv3VdKTzzW07JTCsk3lEocmV/g1h9sfmoJjdSsw3Yt
3ruWxcF2miZMBwfd7/498WMA6AtSpuMvNSWThTG4W4xH1CE6djrHC9pUHPv5khpRJHV1MacZ8Scx
Ty6s0uOtYDjl5dohwdraeDrsRDjHcRTcAyG7jE5WPIYRChEPyy8c3mGqZxvOoxgh/FiHC5vcBJEb
stlgI27QHaDLKN97jQ6Oyp6oOn703Z1leE3hI1fsRzfoTiyqleM0ALF1UYQCau4e0GQcz3dZePKz
HjE1yKnmQLsXgSyLzsy9uVd747wm1WQfLQGaRgvOqL/zvn50tzWLjKEk3p0JKkPUZLtXTJBm28bw
yHYIT5LaLPA4bk5jIoutJ54DeZSiqgNnfAAZuc3akerjJWbDEGsEWppT2H8yZrl5+vnDdGlIrqSI
H5t4nUoLPnosk8CNf3iiZUhf6WCm1uX0xhcTI6XGYNUOzME99lyWq0R3DhjJnd2M3JydmArF5qT0
nu2nN8OA48sTmLLf8/v94r2hFls6wDCLFPS3E/UgE6QlHdCI1p/0foUcRqkMZWJtzqz/d2RMmhTd
u28SYMgZUqoDuYfkofX77/gWI86bG3oS953WUs1h/SMHVdnbrDp6bVyKA2QpkXtjcZa+YOF11Pil
go3oRvL8HXnRQAMNbvxjfSz6ZCHmJ7h0l1dBDiCzz1VURQ3hpRvp5L3n023waNC/mPYKz7Bq2WdK
CdpR733oDHxRjSK85jhEkugS4HS1z9yaixhLY4wW/DVaP6KdB/HyHi5SKiG0uq+nM4VRrY6b6SZd
4BRQVWvpIEAS3+5Ys2dWi7v+Gr3YgeAt5wom3Se0T9Uj6Kbj6ISv2hZRasv86+ESTW1p5fy4LI0t
sDAiXC+cCnBVPFKICZm7u5oWrBmtlor8GKOo2WqtnTktxLvxuaYFJ473xR8j7uXcTJfy7mlszcnN
+slExShvTmUmxhw/ANOIB5yfWrtuftGrZ5I6tERA+6XtIeSqKGvAZmWN9QX0VvuZXuiIMK3wX0dV
1as7WXBppJ78Eqe9oNRkcSl5SpQzwGXhvVNZnqFNoVmiEKb6n+BdPeohDmtkb5SZbwbMkOoIV3S5
Dk6z/a5e3lLUh2DVgbKYd4fvvXw7hkXc8Fs9EwdRsI+tMrZKCdHVKE4KPrGo4auyKjMA9PkV7S1Y
pxbmewQ3NzWS/ZXXZEKtm23v2SPrI7DUTYxRFaydROPAz8yMaR0Hr/pHp2qZ5XHWAOKD5OHnLzfc
9SDlAg7FoYUPWhAcs3xFw68SNdH+VXLtY8qZXdt5vPW4deO8uXKCJMhxboER6EUQ7rMnKiytwy41
QRLOaR9GcNM14djYgu0bH+tG5eS4UnQtgV082k7Xw+lDSnXMXNO6vXueiQqPU9TYfmfM2foLiVko
Z12ojumfQVMOUXtk8G6GkJAeMdH86aVsxYbiF/ARqW1WW7JEC5B7gxqFzH83/N/siUBVu616zW70
IhJWUZIvBjKs0/VXSqYBjktTEG/slwSEoiEz1Co/DSZaFiP0PpjH8UljcLX7WdvDPIOYeYbcnZNQ
dvZJt5on0loAT+EyTjOrdxpFjsyG7la6bXbO+n0ZJqK0BXyByEUWcIWlKCpJ1f2O8h9RTBvYLWmc
DOKWAFv65JBzrvZs1AKh2NNKrnIuu2NfX3y+dlRsv2za4pmSO7bH0G9JhAV8+pd9TmpRJG4hlZIF
RY7TgpaEOR5gaTVT4hR9sSm6JsB++5ZLRSmp
`protect end_protected
