`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
P4Hs61ywXRtpd2JnuzyDpNG+GZc/aw1sf6FUAAbbgK9q3e9/JUOjzGNWCSxUeFWw0e3XxJwL8ONb
3w3F77tt6noTIlFGAKASUaLsGMNzEDuDbP/n6HWktXQfXh/x51jOPxazqvUzrV9M9lHJ9Kf+2bHS
q3l3ZJU1EUeydc/4HrmNM47ERlcb9ISpa7zns0CkGG+wpjfCFKWLQEk1sHbz13LQsEYacacB3aK1
03cdYeF/bThSOHSBFgl2H6I6p7VP4b7Vvkz5itxDCN/1JE2eWysJnTzZ7N3R0Qz+0FX845veaoXa
1aZN2vJG5k0HN+DBLQu88i1K6QyMrjnjMxzOLVgQ7SzGuKVwcBE18/R1JCF2X4vO1GWEEK1Ko0sr
Dx+EALMP1jy+vk4ZiVN1GeoJg7pc2rkNanUhAG0XPNrkRTKwiViTk9DjoeiyrS+yxU0KC+h4ajW3
2rsEIUdTW5xtg/Dy7GohD8KDrC4t7S5WHdTg7Tx/QrlXVpSQR5/NMiPdzEMNYzQh5b/gq/7dDRnl
XZjfkDPKTpapN1oPovacnOOUJFKI1QcxYz8UwhgbCJK+khzppLrS2Ec2mFp3unljZr1bsfay3/6d
7ifEe4r98JlsQcPLG6Um4vCIJVKKCHBGUg1LlIavinPP7FkQ9AahLPcJjL8iXH5iM31TGZDVwJEo
PBO10HtYLrsW4cW84QN95ViPt/xERkzNDZw2gzB4Wls/YToHFBENyOyt4jKQVvyNKree0J3UkrXh
Mt8h9xcemOnkfIelRXwNSVezcRAKXcas1ZI5bnYYGCCJ2GtbSoE5ers/v/Voz3YiMdyl8qd19q7Z
EAEQ9rF6TQGWwFoEOCAqQ1knR7UAJ9yq3ZZv7TQplwkiOHZVraMloS571gYJak56O3EJ85kwDrfc
OuKmDRxHGGygkicwIeT1VxdnpGa8GGWce5Xlc9dr6/LmDLaw3ZnBJIb1zcJGrV7WVHseqOK5EjXr
znkI6JVtDp0pfnDnkPrz68w59sidmG6dqRFlyNz9aew/sEP97LPRbw9EsWx3QyRcvnRCWRdq0SLB
VYfEttTIM09O7FvsNNj9NHNYboItNxbIxF5YuVkYydapp8s2e/RGw44DS34iaE7hfGMMfjkI8be+
IGgBwTUNhy4iHtKscC5R5zIaOWXf5wwGdSsj2oFnb2m0za/I6Omu8GKmEZdAph7g2WRaz5eAcMtz
QD4KMeUVhO33yciUnPq7/tFHTzwt0+r+OxfJbLl4VwIefM7zSyKB8IdR6QESyyeQWuG5qrhA6b0K
iVSVn228rfr1be4uUWhlyJ1z/x7b4i9J2rWIm7cHqOvsVv16nPIZ5HN2XWVY99eBvNPcUiwk4mhs
nb4UhQEzP1u/0MpKKrfTvo4WwGc2iGVNsRwwB5Sl3stTGbqx6t5Fem6qCVqCymhArL3Hj2CVvnnZ
G2mbv/aEeKWHzvTnpfRZRXVPLAlPJqu1NoeS7/DNw0HmmHb33VWECQZJXXsNQL5W/aivSAvdm7IP
/ZCVTYAyz+NztmiIshmIKTqkpvl3fTXJkvJd98g5EwKU7A8vy+X00am+RyzKYJtddzvLduMmLul1
5lNDMFw8c/CDX9SsgKB30UR/R+zVX3tVuGMXBbJSJrqIipjmZK7cdoPRtjWUNAXrf3Bu7UhJooRp
Ry1QbD0gcqsscCtpgGSrCv2lVp+LdnnGfkY2sG3GK0gJqi+rCTsnQbqifK2tVzMaURvZSg+tZYOQ
ugsb/6QVQR/xlczmBqzHp4iXrCN7Vvy0yzP+9/gHiAGM+BBTDRetEnzqeUE9Z+upJpHzyDMPJcHU
hb/KYHAx0MXKDZDqRVeyJuJ7L35DFHhVHjyGkwa7D9tsPc4DXSsNPTkTdXduwZBcp1mRIdZ9leFZ
szmhMfHrqr5D3iiU/isJMohhIacYLc2BJMFEh0Xu+RGctm+o9tsZQGivELUHJKKY0kcTHi0IWsrI
ZIW9vWf3xqMd+XsV9pUHLKO3LmJsBrSzatFbh7BmeG/2748B6ynQ+bNh5MYD+Yg5yMlhmAEcpCYk
/5nHzcuMlPYB6iLYOrRTzcavN5dP9Ey4t+kv1piHnlxk6kgm9fgsECPMtIW5jOnOpssERQyIsW2Q
sh8HfeB0zaTjJMPbgLhLzwQhiWsy7OgF9GzVnrEZK8Px+ehm4Pf3fIG58O2nAeaKKId5qxmltHLO
rcAuuM7MMciX5Oocyr+WMeidIUQb7d5c+mZVuvuogrDdK976T07YpkYxa/8kyPS+4/0NuVhvDyFQ
1p/bPKNK1s5UvIILa4wS2D17ZkFpQjZciEIaD51Ke9x8cbw+6JXyXnEpN0pLoFA3ZC/W0E6Ds9/P
XOd9faX20WqLf7xKBVa+fl/xsDvNIXY6jucHX6ARPRVbxrn3kHtttFi3C417aeqTbEYihEaaG/7Y
2bGzUBtGAfaC+UZjOJSMrGKRnWMmmJZ/xuWnzWfYOW4ryzRshIg0eFn6UIgFjqKiLNtnSmtAwL17
I3nrQFSv35ZKQD59PZ0QoOSyeXQyNUwIlNpv8nDHG6Oug3rcE7DMOiAGhqcr9dd+LrSCgmoJcuT4
t9XN0kxOr94KY+s4R6pBW0b0KD5xt9jvyNE6vLPq0QzQTJH4BZoURsktsPlhC+NZ5kWrqbxHdEII
aoafuG2FgZ48P/u27tZ+eaAFV0Gh9cLFsnRXfBgd4iL+UsC/Iv0YGxcZIjoKnv+GPpcMQ8wOx821
aqnwrusGRFaosCZC8QPVcWE9d/5dq7jssJwrK5QgHIRoLWAqSBC366RzC/u7C0ZYvZFUXtCvK/c2
b0R+BBYnrWQq9W/yYIzNLzoM48NAYl8eaPz3J61O/209mVcKdQr9nVOzJZ8SAif2Gxnry5iXBNyC
sN5bj3a8pzM42jXm6ld6pMnjNpIETflujz1/gljo3N4DlIDpzVMbFVgpbmwt6tA6NP8zWU917fW4
Iibzs1MNZFJ/014fd+LNQ5WAhV56jOF9wfgKxZ5qODf0X42pxvJ2UMxpVR2svLFngz8+g5e21el2
gl2rymEy/PxXo9RfAp5qLCJuKqyq3Uvv2oFB0JXxkOpO9E2POz9verS5SPVECTC4Qwq3Z+x6RUeS
YUBmI5GzrKtAJbbGjkbkC+30Wm1oRI/l0ilcKlABA6iW1gVTRYjRAindGF+eSfnP+jFx7NggV/Iv
Kue2oXc0Vpx/x3EaWlFlrN1G3YAPQvmiHPAjoBiSoW7On5ao3dbr5nFZCfNvkJmTvwPymLWeCneu
urG/Omyr41GBWVMMiw0CTmthrcWFfuQkFD4lW3D4FCtswDNcY1jmO3ui2eVoDgJzkHi22Ej9KP7j
nhnpuIvQ9K6f02V63nfoOF1bnLf4+BvPC3rxgTFysIxhRGtvFCZIDVofW2IxOYlNRX47hREMF2Jq
aj2L0/L+9bo53hlNfnvYc7V4e/LYiapimAsBHa2Rm502gI/iNfKmxvri36ULs4Rv5Bw0TkjgiF7H
zlW1pGbMnp3yqKoiR5QfOc7M6YZi5gZtZkuYk1zrZJqqAcP/D1c/qO0VxPyZ8h/2OvQqBk+4vzWO
WL2fyRb2zdMewl4dc+P8EBtjYvwTHMantimJ+3qzMjGLxsKVH7eOQaZSiyvMgm+eb8VoyiD7z3em
VGi1C3NZyAeQgR8pXbCVeUSIT2pMUYcNCc41IF1OCRhWqV2s2WyV6FVEcOneePoHqB/Pi9J6HWO6
yiSRJ7AXBMzznRbw9PIxbZzexouTIDZMM/qWPu66jctkeVI/bDQ0SLTqB2FEpKYJYMUki5yfmhtS
GdbUtZt5eNnNCN3nwJAlSoKS0HcOZRAufHlcfmsBV2h4CLBvw9ENBUsHoHry7hCsYtY5wxTOXFNN
iGR5611mWcBWQffmIk8gyDce9m/8aHXmZGJGpdPefo8R2Cv5lZ6hgH94zmnzSXUVpkdbbC4aawab
p6vYifpxKkN7qPB1qUPu0ldiIaSZXmXVkc5PzJg+WSeuLCKkmjsOQj9tqJ18pcBbLG9HMeKoDfvk
BHxbmDeA9wF8TWqKjEmJKVJ836SvH2DN8ZJ+hWrHh+4V+2YBlTbjzqNVm/ibH7yqq6wjHGL7cooK
FFomm3+Fnnudvpy8YLYP6i2uDzwaQ5Cp/3qqn733PYn8nyPeDKW8N8Ffkjfc+aU7zCnk+ORvE0Z5
tCOlp9w9m/mywJKgi6gz5rE27ElAxIhsvakyl4JeMtPcwh3bx5AIjK0TECmwfS16t+2UBrtEE8qK
ocq5RRf/mIywJWDgvroaY9nqxWxMX0O6xWBeTrrYtoniQ1Wmcuq6B3w83kqtbtA5b++XfNFu+nrM
8K2Hh1Fh0vnBAaHeTMOZeE7yEYLFrKh6jq2nAa3eG34s+yS7uLk8I/Q3RZk1oui0vq8cO2vt0pPh
cQHgEUIxu1+PwjUtNaIhsLF0qZM3oDPO5HWjIW16uqWLGKFzlTzez1X83bHe1SU6qPuM108Gyc6b
OYRPGHXmM0yzUH/VDwyUyTxtf6SlmIXRpgD6v4kZM1bV9n0B9Pbw4m7Y19RsDcXSU6StWwfezmCO
16GvyLctXUJ7YQqpCKYMUlbWBLWRt7QhwL/e88KmJMb/oJIR1D0DcD5V3huS6YAO418hBtharzSQ
hRmfX8oxHyd9Wr4N0OPaW0uWMzxTcFIA5OGGXI9kwoo6p04mN4p76ueLpCORkzFNhM+TbQrfL4kZ
SHeRrqXGOKIDEeA7F5J3mzQBUA6oK3c7jYwDp2rkyu6+bg3sQdaYFzL9MctTmGR93KvsYYI/XOMr
BXuHVqnBerzfS8IM9u30VoMG106h8pDEPmVYIttBR02xLS36RF8yNBFcHnj78ykc7o/VY+wE34SZ
LBWtqFnAc2vHhrzDCut/Fg==
`protect end_protected
