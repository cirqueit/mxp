��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l����C�=��31J����crŲW�0y���dalpp6�0�?�8��-���:��N���$w IbJB����Xf�QӻZ�p�����ؔ�T�]�0s.Q�8�sw]�5%��N�{��Qo�
f�TO����.�(ʗ:v���"]�#F�)�\]���6{�\�oV�Oh����C��À��pp�����~��7e�y�ף"<#���8p�Y���C����w��.1�Ȟ^��2�e���� �څt�2	8� ēF��M�`��}~�NS<j)ЉC����}p�R����դO�y�e�&�~�Λ{����$�Y�#C%G��>Z!�?ۇy�ӟ��3��5��\&K9�����e�t�%"t�����A����5�`�{FGU��7x�L������w=𲣇��^�����`�"�����ڏ�����)g�41a ��o
�ah�HkN��WXv�T}D9ke+-[�*,�9�X�v��F�X�Qݛ� ��Z!JN�àq�Z�Y%�I,����R��a�)t�Ŏ����iH���Җ�@��HL٭���˼���滵$_����ŅO�{#�*} ��e��@t��3r����1	ʠ��>�r������;r�����ʫ��b��e���\��Ӆ��[��Śڰ�f���3�;��Ǚ�a�B��G�#^a��#"�GXZ�C�%�B��l:?f,�:�[� ��a���[�S3x�5&<}�WJY;Q�G3��C�VR6�m������=K�r�^k��bWl���4S��ۜ�����P�)lr��
��F�1�ק�ud�ᑻ;����uM�=W�T�?���L	cb���p���J�^:�(
sȇ����B25��T}�hU[C��x����,x;�Ǳ�{S�7@-��=�@�s{�%�dQv����}L�	�[vpH�l�������G�/�νi6/� G���[]jq�� �:ֽA�����Йӟ�]rc#�� ����� �#���;@�S,|��.l{� TSV0�r����A��;�<1��`�sShT$P�d[�Ӑ#%T:l�l�����S�.CZϳ_�a5l�M9i�ڄi�n��K��C@7�i.1��3�IRm��O�NK~�E�T3'�� w��^��R���/C�(�n���C�����@��l��1�aA;,�1{�nI�,	V�<��z�۸Ѓ�JAWx�]�YU��i��m2�1�,���)�l���[
/�K&["YS���2�U�,��s�#����'JӠ\jM��d��$Q*?�ĄNz�7[�j�� �z��4����Ke$A��e�E/-�<�5p	\�c�Y=�iN6��3�~q<2�����2�8�8{0��!g����G���l��P|�ml��OM�o��-ч�~D%��j�pP�/�C���s����@�W���UX�.��ߍ|�
�6dM�;.�cw(�6C�4Kfc{��DU�W#�b���R��f���^x����8Y� ��M_���ubH���(t�����R��h]��"����o���P(��%k�Յ޾�,$�ֺr(O���U0�Z&�@`�&�m$���%��>8s��b��M��P����,-g�s
b��踍뛂6{E�͎ބM; XO�	�3���ʕjIa9q��b��;gY�ɐ�G���u�m�Ӂ�N���oD]��U8�,<���]�!�+{���>����1�+ʉ���<��L���D���#�a�[Aw&G��S��*e�������p��ۨ`4�_F�WK�Xx�����t=.\���V,�\��͢��L�GZ�:����\�{�8[�kv����@�Nq��\�f]��x�d,{����@u	 �S7	"��_g�shzp�_�:
�<I�7����X�m�l�Kb8j�''�q�<�x�'����u����<��U9|Tr�Ŕ�zC�ws�u��;�%Ƨ��i,z�i�Y�~1X+HHeø���"��yȭUH�6�6�[�=���Z�1�iJ�c)��q%�NFrF����uU��?����?���W}��E�ibS�S�o��eȳE�ܤ�_�l!+�[	4�$.��g����>d�d���
\�PK�~�b�)}��x~�z�0�Yh�&�o��l�X�Y^��O��e�S$��^��PcU֝�p��Uͯ�!�Ej�ն��^k��w>f��ظp�>������Q�sTVk�a詏΁�eCd��'��4�����C#*F��������#W��s�'����%��L�0( 1^����P�s�ܽ��<��O�*aC^��%A��mw�@�_��SDRr��e<�mty�K�{J��*�⛁
W��_@!BgoB�QUS7>��e�`?
u��}M�D�}���T&�xj�pZ:����$Y16��|���"�����+��)��n��\&t�Ǖ�k�>�� N���̫���{*3$�@�R�9�ʹVٻ�X'��_�PC���}(^�o2�+E��͐͊�2���)���RA_�YDOV��/��ِo	N'���<Lc �m�m<����xl�V)-O�sJ>	CL�:7 "�d`�`�
���yH*'��>�,U����S�D{i�@_�,�ܸ��(c\�i�8=8��|ZO4��;���׼��tsm��^�6"�+7����+9^l^�����0����N���QY'��j���v��DC�h�p�޼�`���~�w�c
"�{�9�j�A��d=B�ꠏa�a��%%@���E
�� it���Q�9�-�������N4&�!oW@k�쇣�����P�X������&#������� �Ɉ�D��-e ��(22�<M;�jy��n�k��/j�<Y��Շ^�~�x���F"M�AHa�09?P��I�LXZj� �N�m���D��PJ6艆T�P�u��Ԇ��[^�+1�{��R�o���ɳ13��%V�ұ�[�e��Vp��M����N� ��j���������w*�6���ί�|�`�~})6��a����ɄY>���\��sd�"h�-�oK����̶�3$���L!r���B&$��h�5.�S��T�6P��u�a�����;M(�jr��\͵%�®�H�t�_W�̦���x�L�krGJ��ᬌ���7�]���k���
h��s!%8��6��Y��Y�E��~X�� Z�WhND.�������<�Lv1��F���7\�*�_`�/�P_�:�ȑ��|%���N\�.���٣"X�)��f�����������{U꛸�����am��z{�t����6�,��W��Y\b^��
D�?��j&3���n����F�b��z���J�/e������k��/�U���� d��x~��վ_D@g\����xW��hJM��҇R��"��%r0m3����i��;wI F�62��̠�&QTR2@䌷�;4Z}�ȱnS�/sĠ�V����b�l�p�|��JTD�O��|T<� "'Z�D.NšE`+��6(.$]`�ξ��ؾ�T�υ����^zD����,Uq�A�lZ��$���猺��"���_t�XQo��ǛM�椈^�a�0�7����e{��4�]�� ���F�Z�@ָ��X�k�
�����?|�>
��L�MZ���B%v�k]<�G&_�Y�_���ÿc|]����?z���֬pA
M���@�`"Yp>�y��9a�ݪ�� z�w�c�7U�P3[��GS�G�Us$(��'��ʝ+��B�Q`���2)���VҠ�L(#�׍����N�iV��5��� �N�y����������g �"��p�+P�Q��:C}��{�����~�;Z�	��|�*s^�����?�!�F����d�,��/���S�2B6�6��(Ԥ{v��ґٴ�h9q3�W�\6�ϔ�`�Ah�;m4�Z�ډ��,����J�'D� <�|��*#_�r��U���h��:�	Z>D����1���' �|Rk-�IؤI}����y�`ALW���kH�hr'�/Z˜�@����"q�����'��W�ɠ�q��Mě����m��'�p�~@^���Fp�|n��=/���w���������]�뿫��P:[���՜�C,*��{�]�W����fE&:' ��䑭Px>���8������Q���TN�����^�ZF�یTī�2&���^r[:|5��^d��$rgS�S�bs�aЯ����5�p���g�w�ˈC@j~W,o<���>P�!�"� ѡ�TU5ʳ�*C��gS-�4d��n]"�y�gLbX(9>���]^b�@��ӵU��L��&/11FQvI��N�C�ڔ�*`����>ΞW���Y�ů`���F(�"�%�sA7�C��*�;}k�l%�N�\W���˱�D��p�K9�3��!��~ej!=Ť5�Ȋ��j͖�n��bH'^G�'���������Je���g�kt�z.�.��0rV��|2^����x��s����>�ݓX�]5Ll�ٍY; �Q����t5��-͡� b(�d����n��f3�j�Nď¯.Q$]E.���Dw���hӕ�������,�<����>[`6r��l�u���,�C2dq��	���d�e��s����e��1��x�si�៓�2�W]����g򞑱�����jS�{hS)�_���GHO���=��6c�7[�])
r(�GC��|���"Xр���@ʇBe�_?9�ykhۤZ<�"a]���h�tWO �!#�Lrm���mIÓ1�(R��0��r�}d��V/H�x�aՋu]r��.̟����D�&��v�4���Ƙ���Ȗy&���!>z��C#d]$acҲ?������p�V�bf4^@����[���L�.��u@-6����Y|1,;��^��#toV��T�h��w�d�"�*�N؜Fp�h0)�P�M�S�_�b,�w�'u��^��z���o�]���zñ���b?6n@�~ܳ @ޞ�(����=��"7�����4����bS�@>7�*�yTn)��2$��k��\�����	���b��6��v��ז:Y�M�z�g3˪6؇��RZf9����|��5�[��ՠ0O���_i(�mz�h�k+JX��j�m�{������8��B݊�t[�UKxWbi_vI��](��������x���N�� w�X��ԾHA�47Cͼ�6w�>�R��'e2Dz7j�d�6Z��o�������"��PO��������~�d~��A�y���E�S��N�X?�vDg�l��5���lY��w��qӜ����I�ޱ���*�ɞn6�p��T��D����+ru�{.Y[�QM�
��f,cuI���'�}g�3z�n�g�� �7��.������MP�J^`e�EDP0S!�v5Ԏ?�Sb/^<�s(ט��:����q"2"|$�y)BR֭5i|��8ǀƅ��ڤ���Y�r�Ҵ���9kT/h�77��r���f�!��Јpe/s�����0o��p��ETp�o�!&�����"��T����r�ڌ��$��&�J8i���S��gJ���4�%J�IIb�P�7d�[��� �fpt�Up�Y;��,�䬸Vh�~/!�ҕj����/�S�B9KK�ͽ́��:��F�F` rv�C~�a�	R��w���F�p��4��`H[��Ql��bƸ�:�5s]0���r �V��1k;�5��a��$�9qj9�9>j�_p����R�886{�,��n�_v\p��Gf��2�RqN�[�:H�I�݉�;��1�6CM�~�r�����j��(1ƨ�����A4pH�C;V]XW�%��h"M�Α�>������1�bcJy:r�)��W�B�J����Hs�k�'�w�ķ��<���y��A+�Zn�q��+d��_ڇ��Yտ�0?�"�XR������A�d6��95�����I)F*4�"�	�f�vNA�U�?���]�����P9�����H�1�Ѯ�������2@\�	aO��hዴ"���E�>,Ffpa<��F�7(o%Lby��r'��Ұ���K�b��@I�$n��4�Ww'��O\���L�wC��wV^�{�7ywHm�������������%�<m��6�q�O�O�߫��j^��&�$���f w�p5@���UO�Ri�L1f+�lw&o�% �av�N���r�f4h�#΃�c��M���i 9[I��KT���*�B�=��͈��uJH*��{[���X{���T㋐�6[��Qf�R��>�G�RK��� ��Y>e��{�m�T�x��|�j����z�MUd���&"�G�}��O��#�!�8����D��n�/��:�Zj��C
�4�@��dۑ
?	��봚�4�EBe�,b0Z'��!�AP'+ �����r@��E�D��ԿX���� ��Gc�OЋ��Z��F�E2-�[3PUȄf6���`�v���]�nAh��0;V�<&�	E��t�AM�`��s�k�. ��3;6dR�����Ȧ����'�;��Q���>����ӡ~@΁����HE�����<h6G:�E�p��5-t=�9T5ͦ�w��/�zM5|�� w?�٧2��8f�����72�k@�q�����UP�Ck�b�:�Q�=!!���TL~�_����k����u��s7UO��8�>\,S�#��kE�4C�`�FB�R�����l;x�E��'��l�=|e��o+^*Ҁ�N�S������_lŮ�⺂�3�M�0&Bь\��&O���(��ª��܌(�h���n���7��Gl--�@k`}�j�J*q ��8ɘʛ3_��`��=w7�N�1����r��^��3�+>�ͫ�=���M�w��Nϕ�4�z^(WDE��x���k��u�����`
p�w�U	��"d?/�ƕ�\P���@�-�?����ӌ�i\*��$�p�GʬK1i�f_���<��f;4���������`�S�.~2C�c>[�? [�b+r�u)ʸ?��2���|��VqO=k�:RGw>�HP�P΋�Ig.X����!Ņ9�Uc�����qM0���-�V'1�;��S8��Y(�n�y����UW��V�%S���n�;�P2� ���n
=�`��i����s�0#��Ov��b/ArЯ)�i�~u<�c�+�O����hl�C ��/ce}Յӫy���<��	�I�&��X0h�	��<s	�>�ڲS8wQ��z:��A����d��|�9ѿ����;y8�ާ�Y��ы��F���`��bʖ(��&��S��P�ME)û�C����`��0�"�a��g�j�@�d�h��|"��ٿ�Bv�\8U����Ӛ<����~�C����g)m�.I��KZ�%��#&���6ro�
ϟFi�i�Q��]�Pޭ[�g6+ku���^\&���"� ���V΂i��8�s�c����8˪�l5�Tgb���Q���ړ�g\kq�r����\�)Y�*�;K"\�%U����9�~A�p�?(��{,�.����:d���a���G0�9����M�A�CtI�K,��c�^�Y_��
o?Ѩ.��9�%G��.)���|Nꪪ6̕v�iС�Љ�g��	�m6i@l{�0A�p�w�?&�d��#��M$J�޹� ��۵Ǫ.咹�X�s�r�X8���E��Ӝ�t�Ί���]`�p}i�Y��ɟ���w�:2`Qƻ�
5��ox�p�^�%܂$���b�Gz!�"4�i��z��(\p�`��z����������<��Rr��[jh�Y�IK��b��lG�:�@�r�*��_�i�ȵoHV�����}1(?��[�!?g����}�r����C?��~=��o�0��tHq��qLOw0<5ֈ�4��������;�%�p*_-�3(-�A��īr��ǭ1�
I!�1���OӍip�귔����nL��bC�ӧ�?=����E=�Q9KT��~�U�v=
վoG�N�?`�^��a��g�,P���v[�4♖Rd����?�1V_U��ڥ�i�\�K?����(1�KL��'�K�v"���X���R}6��h xPCXC�'�q?�*@2y(fүx�&˙x�½�����+ȳ�hW�K�5��������]ތK"��,�`:o��u��o�96���(��V�2C#Bσ0�������L)ϊ�d
v�{9HXY6ߣ'�K�#g�1����Ej*뵩�(z�֦�}ot>b�?9S�&�~��盖{b�-㙍��X5)e�M�4��:��?�F�^G^NE1�>���WҖ�g3�̰��1�i��';���%ך�o�l	0t��ڎ��hX~����ƪ����sy���eR�*���u��� ���O��YP�e ��/�"_� �d���<!S���NZFQ�D�$��xl�U��~>-�G*20u���$/�� �je@�j�`X;�����?��7t��{�~+�~y@�ª��^��N�Yv9z
����YY�c}��h�Kt�J�՟R��?�&��>+<]�4w��o�ӵ��_�k�����<n+�.ຏ˙<�3��2|�M�H�p/ Y�(3
v��c֊{n�d�X�
!߅q�չ%��9�3>q2�$Db�@mtB+6��-�o��O9��T�4H��Z݁9��9C���z)��0;�n�DdB	L�}d0��/�3!F��$\W;?E��r�U�Lg"���A�DE#�@�3�";Zi�����.z�j#��u�����P#��"`����:p��(�
/ohv}���1`F�8k3>���R�X��Yb4�m;�BGϫ��g��*U�JuHө��o/�=eݙώ	��jg��������J[�X����Zm���Sn�'lL �'$zB��H c�|Nl�$2����ng�aO���!T�H\>�,˜q?��x���a�q��^��u��s��g��~�E�G���5�����U�� �a�T�oƂ����T�h֯�l �y�6��Bx\8̃�WN�hS/x��!H�VN�n��0���Z(��`�B�B�;�|�Y`3=��w4��M]ie��-����^�W,}����X]�m�m�+ 5�{;���,�=+��Tj��h���?e��	�d���H����ҡM��G�i V�,�����bX+��탮dq���$�SDf��!���:[q��弊��2&F��(G��d8�3�%���������NVcO�p:h/�*���x0�vT�_�;����[*(�����I-z�B��f��N�����M-Ծ[�2b��	�@H�4E��(a�p��6f6h��j�<�$�K��d���m�1��HE�u�����MW��b�Z�&W����1�?�굅 -�X[=BE��~����;����#�O(ǠNaƩH�Y����L+'_h)N��&�[,%��$�Х��̐RR������2��k�<p�"�%׋���j��Z}�6��>d��	�|lI/U	d" ?�$�UH��0nb.1+����>	/a�9�s,���@���gN~�9F^"d�T���	�͍�I2 ��Ж����{�8���Ս��0�D�xX�H��"l����Qz,���`�y��SG�ǣ��{I8 ��<�3$ʖ�~�$��\���?E)����:�S���c�[�5��r���R�f�Uu^���sj�;F��W�� @����������51�ظb�c���妳[�0 �v��24B�Me� sƶ�ieǼ|���ta��ۨ����8�h��uD�/x��g��:c"���@�ߨ�Ӿf�6@���K�yW����x�z�+��&�R`l�=@�	������"��c⮤t��|�~-eM
¥�C/�fCKwF��a��%�����;bڴԩH&���&?~Q��^�&�s5XĳFfݝx4��G�?�����3�5V!W��ADMA�\����1_�9����9D��]J� �����s�w6���3XG �a��c[*��6	Sc#�S!u1�M�t��3,�U�Zg
6Y�x[���mp�w���(��-I�U�L��5� 4������x���:�� Z�1"�u9���g��<!?]�m6/�]GtE�U92�m�q�}sKIVJ� :�I(�����e��������T��tK��@v�� �����vRꕄ��a���:�ל�؎og�.��M����N����6�R�Kw���Рs[���GW��kmn��D��L��mm�j[@-�0���"��MАLp]|r���dҤ2��~�.�;�;Շ����(D��'v�Jn�5���8'�_*� ?"nL�))��"é���FO<�h8PA0c�*z����������w�1>���0�Q.X[qֹa>�\\��.��
��9���	J�
�uLG� ���D��c�'�-���$;�C���]hn}c��>�# s[���]F4���mVH��B<G+F2�(%r�W>ٍT�k��Qv���z�-l}��M�+S~&P�Y�W6�����._���Ϳ��r�HS�spY8oV����>W]_E���U�H9q��H��Vo`0$��N�X|��?��?o^lcA���x��]B����`���n�r�������~�-� 8K�lAM�
�P��w%&J�ʖF��t�:�&�PbI������[ο�spw[�U�w#(��u�_��O�Jv�����4�u6q�O��.٢7�$��[eLPF�㈌:�orfK�E�`o��1�A�עk.FW��;�)�B/q������n���Q;Kw�Q�ɾr�q�����<4�a2�/�\ 	���	r �����0F�����4� ��1މ�{�p��cQ�G5S��X/6O|��l��=k�#���>����3F`%6<��q	�~���)�͙W�f�1�خN\��d6EKy2	憹��U��ό�j�h��k��GBߝh{ζ�mtG��~1Aa�x+����`��)��u* ��% �gu�lv��	��@���u !����5F{B�-\D=�c��C?^{��tI���پs�xj��_���]�/�|��n�k�c>a�������z�ƣ��藈��YǾ��13͝��c���T`��	���W����f\.�N[�\	(�Y�"pu\&Q�]�r"�ƴ	�X׬���uUX{�+������oXį9��P��k���W��0D��O��l%�G�A���<��(U�E:z�l� Et�`���Cv)��;_A�2��w�I��_|֙���Z�ޝr:CL�،.�`Vz�"z}1!�{C8G;��ni-���׫+���ì
*�)������:l5�7/k�"� ���H3�0��UL�J�,\K�jR~+�i���.|ɕ|�z�Ʉia������pGJ}��|���>��~�;t���?����s�2h��צ_̢D�_�$Dq��� �Y5��G�R�&g�z֞@-�K}ĂʪK��7r%�)�%�C�a�i�F���N�iK���<�RMk��[���s2 UFi�������g�N�ET�<������@d��%�����D��	�Hu�/��dT*��_1 IB���_9��nE�ӱ�<@?�uI�*��o6��%��8vݯg�m��o�=km�6ly @������'�B�����9
vR }�QU���[����o��BTو�"�)1�����4Loh1���y#o�:5�Ւ]d"c�'� � ���u%��I�W`�,� �E̕ogY���r������Ϫ|���=
xJ��+ok��F���q3�6�L��\��1?� MϦt�:��G��ͅ	�F�X�f%ɸ��y�R���	�
=��qê����10���A�b�8�Q�Rk�퀈��mg��q�|<EQZ�]6�M