`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 53104)
`protect data_block
buV3ALkE/VRYgj1uLxAcRzAw0VdSeNXAw6m6JEZHO5KgAIefsb2p72egSL4grN2SqzqL24ducqZJ
YM2xXnHss2FE9eKP80FbBOkLatR8d6kJBXbHrYAHCTls9x6A1z2GCfPDyhxZklw5GK+wG/ZGaHiZ
efPgvR4WaVtKaHF2r9rIoc67MQCmlmZwHVboa+2BQ2mABCoyKa3RHrvM2iZsYslXNbriTwgwBtb1
UvnwEZOmFl7gNQRGP3yT/iACZFfQ/AO9GP2ASiGVrp9P49wUAFQpk17pHYhhOHxU+BClLIfBG/7O
XQbbShhkSRSvi5/ZadvUkgUewcCb9j9S/wLCnugqOsa6boqidKZcCPFZzO7veZ4ZSx1UIMr5bDiI
hO6jE//XFg1AoW57n+365ohseRiXfHXhuZ0+ckcevgbbFJEQEBCf8mLoM6e/ohWfeErSdku1SzHr
hNJmqWp4B1SgTNhHd0zPRqg9mid6AZPK4bokBMXt3keEWQ9pe7HevSZCrUjQbRjQ/1ZgYRtD3EnS
3pXBxdS+YXmSNAvTBdXJUXVQIyFjE64vcG++DCuoIQWRf1oQcsapP+HePJgxrLZRhsmE/VYxhLdX
CTSsoJlucvzYXUNAh3XU2HCF4+eEKhLAB2W5owC+bQ+8VSbeneLcnsYUnvZyybhCPzswJorA6mjs
vqFJBxmTPVsLUD1GpbEb40jz06tZU7iUZ3tEu9bZtihXIh2sT27dDabJGf7J6/Sox6px/sfK7sge
DuHhU/Z0cDUpZeDI069o/lyAeCjZx62dTDcQTwxj1heUghgLxmCJu9H9b9JciIJcB+nDnWex10Cx
yxflMnYzbTjA/UeAeST0kUQ5A7yEnhh+QdR7NYdTIfKZtuJdwSYh5rWNNQfY2wur1W+VQg912fx7
rLJCdbqpLTCjLjBKm8zxDAdGIHZzDG60qMSxEzSWux6HRn3968kxDqYoINVPu23FeavObwSfXYES
yQcSPWnmnZdS7fxZYH+NYT1KAFJX57JqKQRcfUlMryY9Dhof5sGpkhrvriFSCJdaJ6fdW4iURewF
R41+PO0VbcTxv1tovcpN2stSyNiIULBBG4LVaVu/V7tLsyCSwPbI0LdNSg3aAXxaOTDtqZYdstHv
Aq7CahghVyYjWJ7Q5wWTu5IgoUlTg4lha//0LYYGv9GJD5/2LwcfHDeekXP/tOV1ZI8HPxGjDnLj
3pt+fF5j5Euc3kLG6Xv0U6Xj/2K/7AGruZyfR/Dpzz3okGiYLw5YyifHzrsl2l3GUFemy/yAvh5f
Vqqx+wwcg3XRsS+P5nYIoJ+4iSJvO7G3B5223YVjg8Rp6n0O1R5UqxEqTvns9Yb6l6QBpivJk1d9
PYSse55BnAMaCNOBqKF+3E+ZJnkbnOAzDvF7nRZZ4wwd4CPtJKRVARUOWxrWc+bdz45964Qjm3U3
XTNe7TfF9soCZhKXQIXq4to8vibGXUJOX6uhRIxbUjE66v7SciP53kt/MZkBNBReSoMaPyHoEDEG
6v+LeEmdK/lR9//v0BZxNuL7/r6dgbpqUUDX+zoD7RmLRqDy5Y9x9TKOcF9h3FOqqBJ7jGyN2mo2
UPAewG83tQeRJehVsPZdX/551eQdLsBV40Oi5xmjbsvMzD56WxqFR+I8nKyXAy0b83WWzxkXqFbP
cHAiZxFFK8OX3KyRPf/fYN+8kK3ZaRLD96t6PtUcxZgFdBZkSGAd5baRHkr+EVhfghugf688Ze5+
t9b5QwT2+l9G+kksS67M5f5oBzm7fKz34Xbug2HKUxt+/UAcC9I4Ce7JDP1v1gbc/0ElszvNALbw
ttKzg7bKD2lCAO1CC5aloKB6IKpuMX4/kk8RCYJKJQ7siilTH+Y57NWXYcju7aGD18FtmndcUW6g
OUx4mOP1BtGloHIEdIyro2AJGPJaQScBcqUIkmgxxyCM3Z3KWc6hkzibPIh71c0SINvVi1Xe3+BF
ePaEMMkAVeLI+dbvuIcSWf1RHkyaGIEesR/IJt95u8Rs5hvxFS+AV4Vkdpdss8YjYEI5ATKiWjsA
dxwBiVLJHztmO7+iYWiRL85QJOaxLaW4QGcmq2B2FEWdvHeuaLkQ0YlNBvw+If1O288MRQTIIoPU
/rPE5cJfYC2HVIYvUW6VuCUTK4gQbOUF6gW5swHUzXdiHCu5CdLoqMnRYk/jvrl41YDgQ48A483B
6OLCbEeLlf48EMFOts6bN7o6URMYE3JmhJPpkQeZ0mWfqe29iczuyWseBbgVWdb8VyfuU6I4PN+D
3BD1z0vkniQf+SAmDX1lfpfLDokLjlrZbL/XtmRavL/s7HCwgPAKUnhuGf0/iPgkQkcMlYAlZW1O
Mx7GL1JzQhVAgS4minJJegl1ujfNc/3nC6BcDhZF00VsAagf3dWg0neUvnkDrV4ifFTQpb7DR+o0
qHnGrKB3OJzDY9NZ1w+3EMeSBGnxAIlh29zUOCRd535PC1qA8S1JnQJtL1xycru/4euhQwCFHtsq
sVE5GQ08Ivjkx57VKXvAPsdYkdeQqypesnqMFM2bmJejombRgAbhWblCJfYploA6aERpHVbOMYNe
mS4KXCCsK414bGowX5hG4WklN9oHu/o6VU/czrW/DtXwBXNKDYUdJv1n/cFlgwtBRm/wDJzmtEab
vkJRnPmYTPbqYfqZDIldRfmXBJyMcCZfeagYUBW122sIgF60uU5ReZeoDgKJZarr4pnco/bfe47W
clGZ4hJhEQmnMR/CIhnRPZ0/Bv0/jUrrV6keuXLIyh8q1+QwA5t5OLzF793mOhVBkyDN5zddRhzQ
xghno1UEkw41TsOh9i+O/GG4EHh0qe+Yw+X+64Za24a7tYNi4QbsztRgFs+Nd30sSLwVP30e1jFa
FrAtDdA6EHpJ6EhI1IDDmw00TsPh1idL4h6qaXcdHJK8Rc2GSfrE9THOknefpDj3TwbbDdHzX46S
LqMMnLH+kr+RD8m2mW9sMcwQ8jRTVXPVxWVERmkao0gj1/5klxz0cUeNjtuJ0h3tF46yrnUdUokZ
6zuv+IBVtzAg9U+7FOo8nggxsgobNAWGysx/R7K7tOPPVczdOSnu0Fk3GO29UJRWspJEcvQtbQHf
y4fKtIC852FsfOIUWgT9iINT0RMUr99Dojfznn44fxad3n1vR0NMpQsZMqxOy3QbA3xxrcU3QkL+
ukRyTk9T7Erd7WXT+5SnuLv7tvxowJCBTTA0u9kk7SLvG2T6fmPg3Ob+87JAzzNbKhfcUT9pRiLA
BkndGNY3tbu84qjd8SF92+Q4iywTU7/Hy2/6WEBJrk5yTsPsWOsO+TuBsUpYP7PU0hCKk7HVC44t
F8L+g+RTEGQDaHKJUUNhsAQyaQZ97tIDjhQ4uIz+B0U8YjooOn2V7Rwcxzkmpt+DgJUJwgcAqSSa
/bXpprL1e20+VEOv7nkhI7NjvNV7BHHfwucIxGXfdQ846/eQaTXvgXoTSySKBjYdHtG3d1udJAla
uTAemVQq/JSKrwWHX3mgECs6YkxLOfaTN26xUdVuoWhDRoY0ZDCE180mYHGOFC5o/xdVUlrq+g8X
yuHtpJNaCW38SspSrRPoqEf0gGyUevp2cO0hlvI+E6pymdNg2kix+MHT6fsF8VmPfY0QEqd/83S8
IHtUxrvoqEq0yOO6dhXJBHDb1LkC2aZkB4sO+Edzwp9UrrYa86nBStE+UM+6Sb35OrKSCIH9SUXD
ybSZ2xNqoQO1FasHV95QXx8zlF9bPBhrD73/NQiuOQ44RDrK6mHGRsB7v9jfdgFAP9qgKaihQxvV
Quiq/3ofaXVO5GaV4/rE+gCjIPQlHNj/bjllek7+8sUA4gBdmUl727Lt7y2MCWrLQIsPVlLl+wgB
yuvQH9tjHMB/a44a84AcG4rI/EeyJTaDfzWlR99Gg1qRmx4Oi2OyWz9nSc+zuUEC0imLyaUnTSSG
+aG5fJ0OEFMnFbPO9xDw17BrpbVqFDYrRUZ2apQxPuNsSjMy10/OVprF8uEQq8OUnP3seMgSJYIt
HWsh1WnH10fQsGz11PGtbd3HEmZ5o25g6I7NNtF67A/H29QAS3E5mOwSe3q3aDeSi0+5eKqJYp22
6NytDmovLIWh+qW21dwm5lz4PKcc2ihbUBBnzh+YJr8LrG6Wz3CiWV5s+5V4W/DmWKZMLBTzhhSq
5M5+xfRPk5Oi+S2ryoxOsRdICDVk7V2TVZ8tAanQFATfwbV2V3jAVzDbDg8523Oa9gNhcnrFe6Be
Si7EUcpwXYBoXMBoIdktfs/BcHV8EEgLI5gxRilRT1oWQnfNF/TX3e4OeSbp27KPih0NkdPRacOj
hPc/0zOyjJf7UbPOavIW4M18GErE7aJ/7Lq8U9489AAdyTk6R7IZdrD+BBDr3br/HYnmhSvlcoxd
O+aAAiLkExGqdWx38Bnp1GkQp8hyyVEJZ8dTcO5qdTqEDTCaxstowyH3VMuOnzxS/a6TaNxD3Kqq
vANbJ0XU0WtJ5o48FTd0/ronZt83niFw9Mx5+rORQpfcXoJM3Eae/IjNqr/j67d5+yNNyEQ0Mvec
wAviIuEUn33eXj4fsFih1Kf7g4MXmnDF/OfxK5ZnDoJcAKFYym88M7Z2F9rFUhGQEOEFzzJuPwIg
qnFDI4iGPb4xxGyvf3Sk7s2FMB7Cyz/NQmYvmmwv80CKOQCAFEwrO/JaQSRYN9808qjwIqdmyOJa
kR7lIlSYaQzbYmCW88mwgn53Qb0Cp1o2++GxOUkOrfHyKl3RaHqIIu2jKb8969k2QfyFlkZIUEGM
7FH9nxXzy0T9ul4z+oBLooCgLO+i34SB4Q1KOJyUNpLOTTURhBSVqcjywLjc444d8q/bCls3tBDQ
2up2P7BDjBEAF4PabZb0RoJm9UEp0z3qA9LFSUtYWbTSsevdCBQQ8DgbB444VYpg1eQ3JPj4K2Gi
7gcpYW6HRJr3NavPPZpNDae4c89BIu7QB20v5NpHqjaFSeDrLW+cEinf7cGR8CMoY0IlzHa09Zb2
F9x4H7Q68ck9CFtjNgUsZyrrE5nIhSb+X4fAR1MdXvjOGLrRt+4IJY6QGBBudp7CUmOUcllENSzr
3AzAfWNmUg/9VbtGOkVzqRdsm3eYZTrFXd7C/2n4MMDbri0bloyneB7qkgme6J8Y2C6Pupe7t/9Z
FAOr4J/tm7l6HdjNvTqMsol4tZg6tU4W6xYiw4cm2FTww+eZrWvqZHn6l5Q9PJwrs5Raz8/Yyn6k
OlHiNuhaW3RBb/yoke5pAFiMQkK6oovqLCgKnb2kOeURNuwmPbX13u4pRPYn42ZzIdE242zDcKsH
nbAz+B64xaDfOYDhPheh96I1mAzM9wMTC35hkmZvZS2/c5EGUquIj2k2Qv5W4Ygb+RQf9KQh2GQN
yefubEel7C9oIXRjpNfH6ExmlC5HxTIPU2DhwfxyGLpIyWGgwiuxNsL5l6UJ3p3s7Yr37WqNuSIl
0sXN0PdQ74+Oz/O3nj8Dq+VGt4R7VBia03U3z2IaWiGTqfMi27Jw0fVhjkyStgfEPn1ytFXi5Nx+
c2aZINh0T4pEBSZ6mROGv334fIqMy7f9zCg5QxbiobWVMYk97DNfO3B9ibpsZS9da4X+Qu+i2Bdv
B4yRmZY0fVHqIpn+q+KKtCIs14jNR7PnW5ypkXXyWekdiS9VU+YlMi9WqZAaosR7bPMAhfdDgsmh
tzVOw43wWAwzOaF9B27eogOMtQVIxxbbISF+FXpPLnYLEaKEGovx7z1urL5xHKmITvv5iA1T/t/H
l2qD218geed0tPLD/qI/nlroBNSS2YmHm00Xqei2Nq9q2fYCOzvOldE4zT9dI6HP9K4SC3z5jSHF
V2TZ3PECXTRTznM4mEa/qgRVsNhIrHvUhldIESMlQ55YG9EUMtt+SqYoiOcS6K0wwy2pWT6GGB1S
hnPUhY+UWdjEqlhr3Tg013p1ir7Z6xsHPqVLw1uYTKcPjzi3TSWnCUdA1fri/jrzuJAECG8ZMMJb
HAXEmCz6rzCvzBrEDiUcea9hJfSkug8g6SVKPX7y7VCA9Uq+F/RqvsTYC6R/K8IIziSmgqJvvP9n
gFN3skMDqDpw5zgb6t7EIs0NVeUcavXo21HhKa1n4akzLCuDcLtgYQC9JWJPWdCr6w1UO/d/Y03r
XOYb4iNZDDtvEkl/Mo+kaqF9mtvp+qmt2PW6uG6k2xqXMWQVGkqxorRvkrQfl4nNsFjC2gjJ522u
9J+sm/xVhkjFx4XQ+MU9F8+XSGPXwuGNRZXuZl4FJjbpMWn2309e2pVI52qDwwoDJMTeVzLzvMtu
ro4QBwoK5uyG6o5v06UO4wR75KV0LKk6fPfnIx+4Zv+m6534Ftd1xQi5fkmkBY0iSA+xHaseYhLt
iV4ecCi1ze7FGmELag7XS09ei1gQvq4Bqt1qpHNIg+Sci9x9q2iYmQHHpYSZcibdjOqW2NnyRjQY
zOTUsYEPtQN5jvhbz+XionRA2puV5Ky90jfyuZiodSGbz/TUkH1pD49fyCX8d+lerCjGlbGLxLeq
DUm1J51GjK/3tfIR2lKBN896/c1dw7bhub1NnsDA4M8JJgw4VdBVUG4ZxJIXEk054Ox5I9AqbQWy
NKHDuHeyDFzATk0RmXebgyrO83HFWvH+W1LhF0swVeFbK4chfXYzbpDExmQJWPtt41V8IDqsh8Md
cCfpzyTxKlcJkWzNTrNHru5byKM1YkhORy/PWHcPU3vJA9nBAOicXRo+s1BsePQ0UURZ3DUEqNo7
25J1+FJ6SHi6wiR6c1zCnrJlTLSP4xiKoDznaOrtv+kTiXeOaSAymGvaGSD7usbuBeHwc+psM87/
DTdKkQsK93ywUDrbhSMmDu1zmaG5CTUX5GzUGLrY5FQ6ZFtn8IDQ3o6Fz+8+gyqASHljenhIvsoo
HFp6j+s/FueH0eqWTWEYkSPbZUrsa0BPY8LWdI4hxsGGSktH1bslN6l+byjYkDdQAqe7ceSNIJdP
q1C7nXou8v1tECdwbA7HwMKaw4nSrVJIdY+7lyg4rhiojabgo08Ohvt1nv72J2ZpGOBJJ5vFGa1a
AWH8DmhAnnL1x1caZzP0lg+duL5Y1Ze1uIgTyssPZ38Y7LCF6Soc6Op59SMyI7vgohLQ3wH+JWgy
q1BxNzWPhe6GsKpUJr5QaNbFtPBrWYmeJ3S958fdrxI1h+hF3ItlVSvgMflOh2Msb3AAluNd9DHR
VkSsUvwLrm8FG7B1L/JhezrSbj2iz2S/9N++muKSciNbhYnMNEsLjDWdjXvYfuLrlmPVADBi9b8Y
Wbtk8N9/5QUAskH1A2A+pRTN9fw4Q/f3uwBR440B/Zqe6ojzwzrJRaWOZu33wjFGjGHc8lq3BdgX
72TfIuf1FH8xf/AukBJsrKHbw+SNSVovDCExCdDcRGoJMg66NrDxuzgQ0xt387EJXkM1quJH3HRM
vn+tbPOsLqIa/aDf44WC43p8Sf9sLy9ulC7JuvTM1TfDV2MQnKW53/CK9GPPabo2FqICtPRa0R8A
d1dJcIfzMAPiPJnYp54n9cyeuRBt9DBJ0lMbKXujbzw0IVhLBiUOmsfJaxtOvqIxaowmItp4l4I5
h2an0C4pjXsFuVyPaxHDbstCF9n70+94C5kNCDhF/F8OVYvPFFpVhnN6aN9rh/sIXCrI+D9+aDjA
uu+2OMD7w+bDQiOEqi4j5/JdItx6OVPTmgAV68ILR5NIMvfP3Vxbvk6wEqhB6TODmHoyK8df1Pf5
xV+i0ON/lgCa9nXTQq+dTFprRyWAEu0WKs4XD60a3Vey5W5/kGcn/ctv8xWawDzuSw/QtKA45T3t
Grk3fQa5dctyVEj02punJD7EhBvZPtnljkncQcGbX6Mv3ISx030gWXU/2qiiJH0tnJNnE7raHY5H
eCl2JbGbSoKcvrPDAqF5671/TNfOnGfpTXCE3mAh+SRKtmYkSaOjkNHJy3kER78dphS5sDS5xduy
iDScIrq8hC+dAZxE0ZHNPsU4iE+AfF3RTjjXskaxv3c7tzI/yNa7OcyCl4ZMZ3DFc0vGfiF1lZsN
t+8vBSu87sAywhfqW1omODFHCeDwkQk1XDy5ywoz1ctHybWKNIcs9hAoz9JBpaze8Gi8w0oKHFqy
B7FM7SpjQxacukTqQvuHtIZ0m5qWJq2NtZ5jx7yw/JY6uMrcbm7kMgCspLIwoLYwyCK2pFmxEgmw
D18GoDeDqbzwweor69f5hlLu9PBHBHs3z4BiQLO21YsLuk+aDPDvZem5lnTbIjEbOWwSMuiO26VT
18LKYaPBZDxwUFPsL107FyRfXM/f3GULBbmlI41fHDHqFx4AqLJixKULdNnWZyGPalLlxytza4vv
xMtby8chXExosAYOp5V1S24etfApy4+wLA4L3YN9uBUDRSZ73Tq65MUAJEPizm/jEKTiFhu/pR+q
7Fxz51/1dNNXagEsP346P4I+FufcU8dRSb0g2e4+Gzq9aEZcyaxWd/MzvpGd/eEwvh3TyI2kYSnD
afxJhCfomMQKYFxt3LH/nwmSaEn8s3cU9rIae0E6L/RTHYOinfuRi8PIBj8wk9cMYMjfbm2R/XOJ
Nq/3qt/cePcMiwt6jGZXWdv19fUYuRx1wkVOpGLXcLMFJwQzEcoS+qIgA1icyyRNbB6kJNAOfznS
DAxsc+mDSxAs8N0cqzei+aUDaXWRwe4tgJtZ+ytlOi82zmkMBBuCrmEa9bstg1hXTi5z1CmcvFlQ
VDUdG6BB2IKoE/REkHSYMuxjtHjsLIVgf3/TOWZZvjXMDeQpOyub12B0qCey0OI6muv3gHx0QUp5
GSTc0aWF/vs6A/2n4KCl0CgfEOguqejY4nFMCy60zYtIV8pwmysEBvP+Iz+k7o01oyKkvBduh2bZ
9M1+ZIeEJxzf8SFGidq25RACIMj4If3Dk0P4V9CqOMjEgdCFZ3UxIG2w5iLxRzcdwkVaguVPm+0U
NVetGTLZKvS4AamXvYs7JDdKhLNvCU3AHLvfzi4LV1ZZLtF9J6njOeTnhYBOjuWgMgUMfnisS9Ff
ESrXElQhSqAp3YyNFut+zUmu6c93IsV0FIWOeyjKfKi6zszQ3WgCG2fac+97GzeUqeBr+Qzk6WjA
c5vnkzvLYlTwhZh5q0sO0+mk4TqzHPE4Sxd4BESon8kE6Cv0fIWFtLt76As/1eOAn2tOjQtMZfZv
pWJ9EuNhz5YPn/fkU7wDs38Qhiq/B1l5EClF9XkkBIKr/mLsbw2tkYU8mM4YA/ZGCikv4UXeKYhA
r0XsvzSIqgWTqMwOMexy0dHSrouqQUSmn5yHGHl4Nj5aVXqHplI/OPBXThuDcROW8qSAfmDgkrYJ
dVF7Fjt82wTF05wkKIRG0YLUl1CpWZEHXv898lstuOVKRWuw2YcvAmy7DEhy02g2KGi7YsIKfcPD
8VgesQmXfXQ4SN7QYXjSNQQ6jrmzbhfoy8+cM+cjVnMge4Qx5V2WiOopc+u50BR/EbnC+0VTiZ2D
lGdfTtViUmEdJvKly+PxTLmA7BzJl1SU4lbWM2uDXEEK6NNjouyQHmaT4aOox+7ecYrGZ1kW2uzn
tfwIOG0ESwUHiYbaelMoWIrblocZKS+PLbt6cUxzkpiFBUYZKnOw2l8IXISsBQ5mn1VeUzRBXxBs
HI7nEggN23Af3KUvB8mn0mskY/4ih1F2IFMiSznMJ1xz4JJFCexsYtXAzv8BQHTxHkESB7/QvHV5
ld1WKcvRxsZvi9WNHBuBhAY/h7xaTtaexC/Fni2O9nzFmRz7XgVqdOL1+KmXqrdaYAwV4bXaZVVk
otlj5pLr93og8o+WxowzrKY6WGYoPSHVuHX4GwAfI9RJn9vEbiIt+D48GEZtVjHqFwbNp+8bRZ9h
VFc1EVVIPLr+yUFX67kZfw+UYMheHu0sxHIMd2xCWeeV5VV524SmGTtO3P7OG/N91tdADEEQlEAp
9IkrxJQ3AlgXVoaJvYR5KRHmtY4B7YtVqb2Qi4AmKe9TWXB/n2QFN50V4vH0tdFk9K3iO6JeIGrm
8reyQJ3hsNYevmFYa2CV2MyieP9b0RZMT/GF0gE7Q0OxGqabVi+APIQOtB+H5sKiDeW9hwFrql9Z
2jvoHI6P7n3+2h4miExmED6mN0p4ZyBBpM37gDCMwxkaMHT0Ffr0Qtbe8f3kxO8gCab4rKG2N6Rm
/lultjI0PczvdcyKjW1hXhgOGkHCQTAA0M7h8aKdQdqjm/ty9HmvgY/LOm9tOEYTmdo367eM9yU4
vMqKIEC0u9D62OXF9c6AiSS2rAjnGJWMvp3AZA1tOcNNZDQp5CqqFS9qyGgHPthEn4D/8f+syHit
+2QnApah7fGs+vESudFz4xueFbPZtq/vBCtE2oftgt8I/r9tl8UPkFXjQuwu9cQ8HQdby/jNAiTO
Dqb4/UAlW8XPftJ9km6Ee0IeIrHI1/u6vO4KC41iNKaAumP8Vh0NGIfNl4P+5/0F64v59cZSy7ik
Pi8R8TqCNukkfBpO2KsjIJLHyJHb7v/bIeVyCjPFe3QbXaq+yYpLWzfRsbLBzm9R60o4EA7yWY78
Ai5sCXvNmBrCHX9lcU6bqY2thHT0IjmFbp4j6L/ajmirtCvjdYT+DW8wtzSr02xKz1YCFJkItdFF
XU7hu1UrAETmYsZ5o8TVIj1F8oIuXjUi9/Shda131IfgBGcWQaUIaqjEgcTtWYyxbfsi0NEpFFut
QmWz68fqZ3JfrWuf/RdrQwR0DLzFBftfEueElXUGUE1rsP5ZHDqk/iC7yonGGgRnNLl1ED0YSRHb
JwlwvtwFIeo6NvMn86N6msl0rvdMKhzuWDqeyCJf72EoSLuUZv26/ZTqZr7MSAAT2XE77u4xQlfD
/GSjigcq+uTZsTy/BOg4uLLCEcCY4nV1Lv0SjQJbEZQZcy+q9EtNdowiag4m1z9fkItjK7BmTqRp
JtWccXmHBqbBFl72rM/FsuzOUEtS3owxxVm2VmzxbF98w1je0+jcZZ8tRH+useyHR4SO+sCWpGOg
HAuZ0ItFGscHC4b+4lXUWxUeL67qYLGO5PBdf0HyhJ/VQIzWohwfD5tBd8zB8ynIXhWW2jDRFSYU
d+SlZ7B+sg5pXkm0WlCCP8T2lxYNzP3BwjTsvXPJ9Dk5+Q0n2omQx9+WlhjiwXqamHubZ4TdSbkS
JPUJmInGcEZULewnWhMW6P371HOuaR/TfsgQhWEWcx2PyZUrG8H4O/4z63mvSVsl0DmWBrZzf983
Ivq2cAbumF/S0JwB5tgaF9OWzxN5m7Tl1dpcU+FkJgDLCs07cv7dIrlxlSVO8ozydyJ1QjpAeOiC
D0+ZdTo/ydxI0UZRxNTj3cerXHOceetJtVwsrdR1cZPcF8UhfQUhJXwSFFrbgp8/xEpI4EAcYXUw
kCX1dbPQ1GLCa9BbYVI/B+1Yfb1g99MbKwtRBFGx8dpb5i5n1qMdeR07lhMVLuyIYvyyqCZzwqBU
U1Uexh8JUhdj2D+oVTcSudeZ/nLZD47ovBMje0WB3KdfeTcRW/atEqcp67dgl6WZZonw1xuFeuVB
7jtoXTOAi503/+a9XYNLi72BqTNRbhQoh7hj7pYH48VIVd/DKjZy/xZlNfO1S5L7nbMaN96RVzQH
yoDhAqUJa6zCC9K5zo7DyEzZ0QI7Qwb9L6/gQm+yGBiLxgoK0QLohdOcnqZ7z+1dhWGH9yimHmF0
qOClT9xZtlm7K0dJaP3AYQYwiRAh7J1DAiieIoLY6fAfbNHq541erMsSDHfaasnRlHYsANjHE4yC
Re8gxUbjmuQhVwK7FDegqaIWEtB0mj5BPeVa1zIj2pWOzb5DeFXLD6pl+uXtVQ0qkwo5tvXOyLFg
l8z0ACEKA0VYPpbuoK41EiawA4D5pmr5XZpEAgL5yE56SJK9mvUEa1T9xBP1rbkDOwmfKXFaiAHK
CU3HVOheiiP0fz0wdKeAupVRJ7dd5iZ3ieSG/KelqkjReLPkJjBpQKSXDWeFgmzzwohXfj/exim5
hq6/ddk8ThDP5v6E+q2ixKDSq6xZMBf9zPE9aPzJpfMYNX31LENvsP3CKQ+HPWhlT7wzaLvBDek/
D4rl0V6ARgxCtuL8GwoWijNumyhGgPKLRJ7Ktj5i7pSE5D4ildppcEPjAjukuNbW69QBbaSWJIJ3
WEYyvnNv5IXj70whRKJiBJfRj3qPdx5mWS//srm4QwKHMkb1uNnTWyXwqjqv/sO/zF/0P8XGWkkt
qW8hoyVJzEjLV9qJFPytZW7xKmzInwlhumRMoVt6Top3r5DGxhcmck/5Enk2XxnBdjvQUHBgeUKd
//kto1jCCuXPyyQxqf3Aou50lsdyJA4DgmmiMjjyn3R+Z1Ylu1MyN4ynrILQ94z/3mqi9xCLw+0N
1varluLxgIn9TiDVPYXl9RIVVwt/JbGKxhIOE74ryRLuGhQovgg5GQJpjN4GNF6OgIZiChb9F4/e
2RqkjBQvUUoOLr8mNCzJA4Bi47BxZjNDQsRHumeDiCH6g6hRtnFuEW5UTfY84jEZypdssdHrI/F3
X+BkrZQh90a+LFZLi4kiRzu/oks5zrvzGZaXpsuIXA9/iPYwFOftPQgzHATydC7xjqUbViIiw+uF
NfrpleJvjKSKBdCm9Fvsgcc1FsLkN4xYLxFmO6vN5Tl0wBDZpBYEQJ+yFyoZTMGvBT0xlyAeQ21s
Da6vzdrt2z9H7uUI5vxaH8xFInoKVpEllrDjX4I+PsCPLX5ch2fvijOpByIpkSkNJ7/b55mFSGDG
9x465m/w5f+wVAiKztlaC4qK27Anwnri7uOKm8AOGRynjiS2b3b4dyJ3zeJ0BT+a4HCMSArmyX7h
Qc5kcTpF9iTE3p6jRJqAIivgSqmVAv37sreMISnAyOKXeEoR24fHoQVRWoDkV3YHmoGyr4wv7pwi
IU8RbYU3HlL6NPBagwfJsH67yGlb9z60ZPzx8wp87m8w3dzzOWssDmqwmvCR6sTNAeXdaTgWTDh/
x3KlqNTMD2CgMrchN/jxJshWw44dkQFdxXXMLIlhc+7ialrk3++RbvBsD7ZszuspMxCzJLyfISSx
nul5oGDLIa4TDytfj7vmfJb3GV5Fz4BXHagWscNmiHj8iZVfFZJeMPX66JGNGMcXRT0uRqlF36q+
2seMC8T3l9fObWPlL80J5T5xI0Q0AiAL6iOcVz2gF/7np11psLFbe0CB2H30a+gnx6B93JSFJ7uU
PVTQ6o1tnHF2S++gEL2roAgHiysPbpPjWvVbp7yQhZ/uY+iV/IpaAqipc/jW7nNEODzfuX1T3Wb9
GGVHFEspgBbu8vTCAkNLBVyyHUlMszBjGB5qc7yCSFv5gXfF8OqTnUNCHXb3ooNN4UE0FIZ3sboy
rZ9epdDWz3kNwsCjt91KUb/AcpudxSkf6HG10fsb77qa+U32o+oen2T5FsZ0fc2ouOyxpA9F88bB
bUX8Mpmykd2jktLXhXTz2n6DFT/9gF2N8ZyuhOz89S2BNeOZBokRbSY3e5MCMHO/GkU5sAdydiCE
SguOOEW6pTOXMh+ayFT6a0Q8ai+mAbWLfU/YAAIRC1svfg64/c5GLJYF7jdgNfwtOoVvKxNUdSGQ
J/rAvd9n1jm8C3KlHPpXflxgvJivQegShrWx7TXHGfmIeopBbXhp94MtaWk1LC6GKl0tDtg7uSTw
vhmgQ1zJYMPG4ECTZyLXnWjEDWNa2wkvWUDhs36nBwC54mOG+EeNx0GYAdB6k/t+ZxKYkPblFBAh
ZlUBXhn8/A+35V/7v1HMk3mAnsMBMhdiXyq88EzNLUx+aq7wYZVlEiaqzdXDi46a82GMEZktiDDL
pwF3eUdBokNKED9SJRGwWp94RYGItllTlrDkE7UdDBt5JEKlhANlMPNOWOEL2K6dHWaInmF80oUe
EKKSKl2/H/RrIH9EiD7bVo/dvu8k3N8XNdUrXyIds9zQHyMA1069r0c9cCNkYDfDpfLMEzr5+fCK
aQLDT4Chi5R6vMf8YsbSFiR/Q9h1MIWfbFgXxsIf35+VFVbuJl23lVh6QirCDKVSyQFjN8ueD8GO
U1xRWdIru9wPOjzizJv1vS3LYrO9E08Hjt3pq3AalB6S7Vsbqopug/Iun2oe79vKmIGHRiJU/BCW
7LE1m/0xr0eEWibqpQ9GeTOU54lNrBQSTrXbNfET+cqaZPVzADh/N0jMz/AbLFB53xLEf5tNoUg7
X5Qt+1s6ToqYIcmuDqyi6Ym0uqAN6rARDSgUTwBnKDxnpBCl1Qe5BvluTwEM0b0z1uU67B7R/21f
seIBO9CISaS+/lGx63rQkpfwExvuot/g3Fz8eWR5fSBJx16lw5+s7WMtZAmu/GknjLSdE5ay+5vs
pkdMQbA9T6HGSJGq/J0QRsZZW5qy7tWun3wg3HBi6l+XqjPKzLCyfb7pdwfGqzIlj+YtOQad5PIE
mh8NuFScoMXP6ZWn6yIMNh+7aokQi6s1t6r1fVT45KkT7NbpaZQkVEuSDApLTsgQMYWiSntMOUYU
w9knVFA787RirdDQziRGdG04fBQp2MYFZ1OpHTnHlI09KZJWyvVTdkKZgip5WViK95fx8J5TSCMj
KkL+PjY6XJ7aOwf5yY0NaFzWG94YunRoWLVjnlpAdgX8sLBjCeZbpqPNUhNEb5gUtfIT/yKeTik3
RQ1eiJIhSoAiTNRRkOAfixcYSn6g9z1JxyvxwWPBDdJn1xBkqPtJ5iTqJdVai4/7lUxrIQjSYhvU
TqXDce+WtyqlqvNfhou6HNWJXJ1rGrsGWk7S16OH9iBbFxoHUHT734jJ7V2O3iXfd64G4phGbnxV
E8ShqclMK4It9+4RvZtSrx18Kxle/RPlZZr8NarfTJI9YF6R9iSlNP2ogV91mWEDjQb+TGHCPRJi
2/Vwr5pltZqVqO94xsr2MWbJIL87IXky6yUKmHWaalpamSAWM5A2ouIEI1k814Py2hbfv0OxbdpM
H2bCkOPmZnpDTFeMuZvKSy3q/tpVsHNX4Qqr2yC8KcEgtEBjKgddUQghToDMddJtyyGEftVaBUt/
yOwsutcrzUYeXiF0w2CLYvJGHpQFinT7FLdY7ImUL0pOYIOzqAtoVybYeCpHHV9m2u08zGhjk5gz
56t7uLQa4kjIfJYoFCfV+oy6SgT5MmoZ5d6p7Dh4Z4RGcOIBBtwwCidDYWRv730hPpqIermCua7J
qnif/AyRYL6B5JqGH+uSwBdAoo6goskToi/92DsHJB1ibYmyPL9Drq78M3WBbnaUPVItdcTsJeNo
9csgPkhLsPmJM1C1JGS2uwNmTKEvn3n4i3/1oOmsf2AIZyd+TThZh32bbkIAnDLJgfjaIlzdi7cF
3R8XUsk0q9CQ8d4nuSWEUBTHIopEWFHbHdQpfqp4c+u1QRtTqSxHwU2/4P91h5Lmkds4iVVAbVwU
fr3b+pehKQpDkmWqhGk6/R7oRRTm1YOLpDx5YEWsXdhknuoCUdC3s82kQZRLg76GzB4CPDl5VLZB
KhlscCIs4ZU8/ZLtZPEKYRm6XG4bxPovhssDg7huHhnZ7iaOV2jxR3ftIkCzkKGtskjcPL2kiJze
RyEOYpLext3dryyTKwGrr6SrLYkeTQJG7MJPGs+Z0uMJScrXgbNXlLgDjylIYdTBRS2o9R+xk6Cn
X6kS44DK2+1IH/RvXptGEO0SuxvlRjJX0JiDPpX4s6metuwdoqYmjDzbeRK9+fgVwKxPKj/Jgzal
Oc+gRXhf3ENEmMIZC4w0mgG257br8rmlUgQ48O2NPNUQAoeBeWrrRuF5FUCVc8LmTFElS31zD0Ny
zGt8dOUZ7Y/PhYmTmmvdL0Y0jPG+4/XEZwrFo0+fg9O1/uTtSkAgC15filE2sUF+jt9Ins71mj+r
2RWCRbsb2rihwd4paQVrd2Hro7HxrHe2/kJYb0rZcBhIW/xy+uRDTHf0zTue4h2aVQ2T7Wfo2oeF
0Gt7p3QpMTRr5SMgMb/y2qQp9Q7uu6p4fuZtb3eEx0nuxwNXZihdAlcQjx4GhjMenIdS2FbRhMDX
SqYfISf8ClbJIADgWkeP+Erf99M5hy8NzKwwisMboEDzRhrJVZ5S4VZa1lr7J6eIb7fCGpKiqyLl
EcM6dH478qhHO4p8mGut0D5cd3CZgngNjNEJ9lbK+DD2OYW96w/92+e8sLrrLBNLLoyBM3qDLwRe
nqOPANRZyLWPoMaXH8eYG+HZUGZ+6uihFDpG2Ms53TV1ewyqoVy9iQhkN7Fl3rxvsGLTfs3P7nOe
h2zaMu3Zp0Df3mJJ/5l9An+PrNZ3M5qXXxiviLY9CrpMpY6do/RbXVM4qinKI4BGUarQmXXbjHqZ
loMi8nOyclIHezAnexPpiJXqdepSPc80yYsCQgXA8GfnvETtVV/Yzyi8KpGdMOs5f7W8ELMVd6zo
8ZR0xw/42J9TkmvpT1VNw0lBGyLnw+ROJ4sqSRKsRMrOtD3V3wUaQA6LOzX0AgKfLY3aQR/fnyqv
qSYvOgtMe7YMZiKj+BH3SYZKYF5ju5tTTBrQkzo6IIsnsz3f+3kJpvQRKO7PGV181KEu86QMzZKf
+leLLiQIFEjNtgvMUCyfN2QGCcOu1xPepe8NB/eAweUkNr+t/SwG7MwGvN+Nks6LLbwCE7IIorJr
Br+XpaSy6l4miywBbdIR/t7eZub/1S5pgIZAQd4EJy+JaX8Sd54r1tmI+wieBa2EtpE6HWJXF6ky
IJISdQ0y7G+kxTgRtqeGgu4MUTx//U5t77O1bu4Zi0znqWQBFiDWgdmArteD8v9c2l+nq3s08aTT
YBznH+QMtkDdRG99dfI6X57UNSaGoQMs3CmBEI3TZeACIeBwzMwU0vCqlYMwkmUaYNJTvkjQOKW2
Rqbc8PmqXTFeXbLRkc/SmExq5wB+kWaY2AW8++TdyD1ZRIuqOXbqPT4QuTRNlg4HlgjmjVsr7+9T
Ho57xNNnAIv0DldEiDz7brDDmuiS3l9+rOSkP66ubRf7NnuCG30NXuhc5KCW0ysqY/ezm93tvQvB
8DyeBQ2DIZk82hOQGJkE/osFG8GkVCqTzMrc2Y1xu+HWJwSIrAam7PSLrq9m6LXmy6fCELgarioR
pLUNNmyK/2JgMjHxOPzYXHlYPLUf2vVeNK6zWNofcgCGufajKoKnD/VudAle62bEY9W7x5NjIckL
tm5XVJtKGj5J5HaSAcadH80huVIZr7QvgI0SKYhY8pQ2QOhNib+Ow1gbh+w0CjV86GcyXCdDkBTJ
koaqYU2TC9nLhq0m6buRbI/SrgaGFzL2W9E9ORwTNZgy5kxOeNQqgMRUJYnxlsCFIeocauldgVSQ
hpm5IbSBz5kNE03SCNluwvTSkpNohr2EhgpudRJNdNWA9jAkRCezvZIyQ8CQZd0VckBMsXcIRypi
s0orDF7D8Gh9C/st0yGXU+tQQelmzDTZTZtCZJFPec3ADJwvVJWBc+nrINxBz800jHYfizWu4XhI
DrwC5i3rkU2WKcS/QjxkWW5/2INvfhR1t9WsPrunAfk6jdxeIST8pQirN0I9MVIHL3U5GcxTbCSi
fs7yJxBEJ/dqHR74/8vJQGo84M2etpfJ0h/0JCXvETg6oF14f94yrU8DP/xSpukm5TOh8WeWh1Pf
BM/dfwdg6xNhOtarwpM5qFp+ljdKg5zOP9NEtp+3KHGBUu+sfDm/Nd7C+IvfZl4wI7mPOyfTohy1
H0NFuyrYupVdx2RKTrEZQC1ttf1um2+L1VZyIGFDsQNNF6PJh3J6Eyd33D1V0PODFbsK8AHFR1Vq
TEjiWfWSe0Y+wibrG0OmHC5KyyrfOTZyu71wsu0DLITrEbBWNoLVXC8F8SaT06Naeq2r0InVfDAW
3VmUKANeMywx6g356jBglv8OnC5tSeu6CBBaWgIWFfu9obTkjMckoRC0JdlK3IK0mwW72h8oOZRm
PMP+Ku/gjjoXnwGyVoPLLw8n5fYdoLuEkeYpYQge0rdEpO7aWZxk0zuOpKUzVGW/CLLCDPo7rcdM
3mWDtYDiUfNK27s33h/qJVNw6hIUTHXYHFo1kc7TUF61J4mMzOstxsBiQbnPhxHXmDuJ/VQDolzs
TPZ8vNK4BLvWcyapUmlK/x689UsahS8CsJhvt4ExeyAW8SttMUa4N56DwCUlOxwyl6d9nnMP0FUA
8x874Uoch0P4acgmMk6nS4N+/UlUkAA/8GYKr1zyeAStCQxvpONj5SacVk3s85Ojk0bRQ7oY93il
dwZwPbZmhYGhAAfIuLdfDrzba07O+I255YtpZo54k9I65YzB13kfVqTUg8rePBGvDiRBfWzx/H+6
TPy+Zt7wo4y0ws01I3s0qCiNq3p82/t/xjjzVt8lPDxpEI8JNYef/n/sKTFR/Ec50ld9LOEJ89bJ
jOQHEqYdSQ63sr3/7NZWkQt/FB1sYmDieQSX561harAND3dTUq0GEwHoyP8q0IImw2lyLkbgcRMd
hhX5pjoqF9LFTTBfbqdXs4p8qnLpGWSIaNFfoWrARrsHvi29Yz54rHZ2gVNpfVp3SS2mGHqGnkvO
itjfDLVUQt3iCwSHaKstO14nyguxD+pbSQE5Y5FTQrWjMbcLU6FTPcH2DjarLYxbg6j5+VGU4IKs
z8EWOSNtmoevW7Ns59h1y2RHjvmfucEF0FtS5Q8peB/v3YZkBe0QfzXH1byjdf3/ebpb7GdSVg7f
NA/0aOwLBOFdvlRXK4s3VtR/sEN5rFleUJneGxXTMhS8Tw2tsrREdMppF+Sr4UFqgukIRV4xTjX2
H0W87SIHzRvuf5WGc9XNJitQGb8Tnlz33SXCyRwrXiruzYvnm0wy8DVR+ghwEBUdwRJFR/TJkM+X
ISpqIiG7nAMO2/e6HqcJ9zlMYgclYO0o3EPN+swQ6wq6xzsGpa11e7KIZJ3jwH2lFg2poWZ7wd9P
bCQXcGcgbIs0CBbox4FSio8wOpDuUllaB1tAuVb06Be3FYg9trd6dmKHEL6Etqz3a5TOnYcqmah3
CrIbE3XnMQUhz+bLqqJeKKkl+4DDWmPW02GZ1g10b/Z6/JxaL6Ho56gdVe6zgbL8wlh+5ZOSLGP7
aou8YeE6Qz6DCKBSmgOI3i2rIMPXeBzSUyGwYP7LlZgFqEIM0vtBgnW0taAU8eEEPEW1i3+xUqSs
06+PE183Q1qr/FfqKB2VxATd5Jya99pQMzmeAVoB34F7SZ428qfJq8B7P+1zF4dydWHQFgtqfptj
s8KJc+TSWmRiHv+qa/kV0ao1YJFGzBiFuNBlGwdigOr4f7tt0Z2R0K5ekUenQHQ/6sRF5adDHL4j
927NUxhw+YRRTzvfEvHFFMMhRdSq76q11AHd2kja9JWZbmAWb0zkrweV03gYzOEbOIg1WmCBRtg0
xuaLZnrF3PGAFK8cz6EujNoK6aj13TdpB32GHzHDydlAh0he8Ss5/JSpNHa0y53RGTuwmkoBNZEn
gpcyPTviyY/0QVe5IBIH0omur6VP/NDBxHlCOCsejxfa1cXmUJcgFG5VmwvVS3LFYFu4MANrof0W
eIM3sjoGi4Fi4o8soWlRmfC2W0XdKvLO7IasYEQ9qNeOQFFlS+t3i1P1EKER0vnBG/7hj2ynVaMS
DXOQlOz0Gr53FmBQ8wF5MovlL8DREoBM/TD8AGOZe1tf38vkOe4VmGlM8oSBr8peaikhk4WavAgw
A05vZmpTJ+/MPOFueOMfhQ+5IZ25IzNwz4a6tX+fZpyZCG9vBwtMFgrQp0qvZOWIELQ96G0pdfEv
BKsHjqD6Jd86UqIf8eqc+LU/a3VwBKbmWdvevJiEVo+b2HPOs7uKRYnvE/btlvDIGMbSg3lqvTWA
FRWQPCR/8SAK/hDxdtUUi/6g3NHToQ4ESwRgxsuxScSxqwI1PMp5YnkOhnw4EDklflbh2XA0mO2w
qB8uR6SCwdXCLSD2WPbpErlkBtS25xrTgb6YNSuD6VmK0YtujHRbSwTPzTR4M/R+frGGcIMuTUUF
NP61JhXPgzp87MsDZcH/TNq8F3VQ5y478uYFc83ka+2/4sW8SPuEZ171nGkpaVfm0kYwzFVaTA8j
pjRrKxxGd1aF2Oi37zxjAqRALUoTNc8WgKBm6ioz6jsM+dSvJowEPnqsTUeLgpHx9RpY56ATQOa+
3ykQ+YJr7iTEkafz34CMr9TbSU2FxcosQCuScbtiBGSssPgX28CLwceanHWXKbTHzkUraV6InpA8
QRyp6lul9A/1AAEo4kUsFSNd3RBqqI2+xMS69CmE3H7l1emLqDZ+QydKplfK4jY6ekHsr2M89mMa
HdjZgbIHdpVHKGsZkQMsoeX7QIo9u6DGhcfj4/OR4fVFulwa2Q6nksllyJFlNTromAbLJyYCZqT4
0NGsBUbYHqMmHM8aBCvpXo2UFeR7N3DLB3TElkqyq1DRZvmFngwTzuZVl7bGpR60SPwxICX6hFGm
UckUwie56DTGsAoYD/tS+IqtkYSOpQNOb2PXyH9h4wEzHjUiWRqKc682QKzF7R/V5eujjLxT5h+W
IHS/1UIJM8BZH26eAswGioFFjVNoN7IUevcDepTYtFAwwsJtH+1xhT0BgSr4uRIAmNqvF5dP7wp0
2aA069CNMYFtU/B4LZshLrwxSW9qNOaAw84YyCpe2eJGxPwn52riDUhB46ra+6/0mGu7JDWW28/+
4264cfv2NL+6LQbP4k5nx9UIvP5Lld7JzxT8wHVvPPfsHrFwLaYxUvmuvwZNuKZf4qG5voNUkXb9
4o/tpiDkSyfJgLSHKkm2qPToKuVKR0mP2TlM+v7nqa5volsStMDXztLRqW+n/WLeqilsiLjtqIXK
Qe2xLO/M2MYGCwsFfbo6MObU+JkVn+Hn6QXJ3PqGdMxXH9gQQRBiHgkHISrFTyw+rT9a/axYfhV2
grFWz0XgdNNnF9tj/CihIBRjeW7RtARh7ZDPx9vGLKQLKyNj8mnRE32IRjGGkENnGRYS7GLHC7Lq
MCUtTOGzn9p26omKn/b7xfT6tc25lQrmfytH720Gsi2k1FkJJxOIzDGa40h+xog1ugc62BAwQADE
yJ3VPjyyfUpPCg68iKsrxQuuaYjoV3PZf4EPX7hx0oPAHOLep+7tKF8NLfbNvOCTKCLV1NwLG7Aq
wn97cAEgBZ4kRmozD1EibdMso0N5cJoUMXeSmnOOWkKoRFIuo0QZGJL0zOxTgrvqXzFxp470yNNv
BHtBUBsscmYarf+OAB2RCXSOlw01APItscdAG5+phN+JYoRIVbGpyEb+Q00tbhKTqo4Ak8KCbg4s
X6y3PoxN6oFSBBrUWCLrVjn/7dj2MVaj+kMFejZcg62SGFxOHFvHR4ZxXVPuXIhwHtdGIsNByw3W
9EfplRGOgVjChsjJ2YhXXpoQtdh3Unu9JkJotMPCy6AgaEb7XKYYGzeyTDUhzOwSGxPPfUaaVmFj
7/8oABGiwVevAvWeph7LE+GJ7W2Kr+h+hSmXLePQHFPUJ2mFhBZlM9E0JGh64L2l2ZzE305i4FDc
b9GTceY3Cf9YwJ0p1nHXnkpVWes+NOAPZAqZ75xg6mZJG+lCiwu3wv8x/03v+fqiHmruE0DMykb5
kHeq1/rVqdZK0aKi22CqVbEcWFVeniCncW3Wvdjwmt4Ehpwf7Q5GMowlIfzD5S9KeT/tSrdYCLOc
E50YQ2D0SNp0gUMgJu6uPMgipbRAb43T18n8m3BzWxIk0B5PgQ9zuK8mKdF3M8CYSj2uMkW/BXR+
fFsOdFHSX6FvgWAtEYeCMXbhTy3FZUvpFBJCZ4687b+vkfdXQAEd9LkruZgDwV+NXVv60akXS0MF
/4AAPG72Yq3dlKVFRKvJP0Froq2VyqPRzNqkcyZQtf9FKaQE1es1mBcEXvR/vKaNKpipyucwdz/y
SXIzLfivC/ClKUufxcASYl6qOFUmshVE2KiA+yg6KqwwJHUIu0//M1fChbIDmQATwzqjjhB5DyAL
xu2JAJX3RZhS2Nl2VmJvKAbG34AXsreNJktfVMUtvPxVWPL72XyNORdDCZMuE5stlAglcZFGbl2r
RrpKtSxWsDW/A2Nmrx/9Xs/bK4XwlPWIXwl8LD8y5DugKQ9htsCYa0cHFRtoBELq33t2+64chQgv
NollbgtVUs/tgWqpBtaM2FBPx2i6ANcbE9cTN5hx1RS478IulwJB65g9uCVTEDJhnlbdMDT4Mh2Y
SxxBxM8rkP+KVSeJqIVyKDRWZ3vXveFVhPJbQdYy45DpLYNub/zm8DaVY4mPouDRfqRga8FhLF91
Pxzw5IPGeGUOeCaqNwi680pKxWMyNhI5G6U5phd0SoOhK7eZYJy3fP7MfRp8FH7n5fn6or9eN/zY
bLX7LwZoThwB8AX94s8+uUyxN1lzqQJdwyRZtfxKJ09MChr5oci2KENVPihpcEq+pI6JyVjfEfmi
JsJzwsBbcYxFIxrrytYZ6flvzwFq6z6mTcUwPqz9TZ/0fVXM1zu2HT16NRuMuQe5iWfLXV8lMzOv
+Ud5EIuwErXKLLd6J0Oe69kgM3MPtz3yM3NU+C5MJ5/VfF2MiCsRIvl6mAtpC2Tkv2z+RCtx48Hb
Hwb86a+RSHAkUxJwMO2svUdt8FBG3srltll+Q9n7pTrz6vShUG09jXa9bup5mXrgmvqfX7Vl/+Ia
GMtlKy8vlXYcEYimqndiZku8xQfVxky3zl7dX/NmjlrwmQwtqBgxaU6Cbk4g7ZgQOUxM4p4zrd0l
dYuAO/io0FhZdHxhWmUM5s4H7algt3ToGcqRvEHO9cOPZPg7rB6HP/dpciawm5RWHMSa7S2OuktD
g2QIfmdV99nEMfnGuvd6zbrXi7Z5FPnm0VIne9RG4/PwfloI7SB/x71bz0kmtQC0GC3kxFV/LzVA
4DrXJdixRhe70/WhqOaECWlQwXI/O7yorjQnFGWcWtn9EzkTOukqn2NAGmvKAIn4QESlLOKNxaoY
1rjbdyrsxTRQtVsc9LliwQxFSmo93tpj5QIO2AjtSelvhzmsfe2b8tZhpUaZDd6kcFyi9se1MGpe
Lqe4zyGRqiFr/8YZ20DEQVa1tjNSDiqQRtC7Fw4mjFFyMzY6kfb0fMNzJ+2MMyZwaBYHcdHPzIZ4
IJxxjb5eA7qJ3Gt5dMYCksryk1VFKp/g5s0Q7lgDK8Iddoa5tUHzi0x5G2GWhiNZ7dtWiN1zj85O
ZZLL6rPY+reHlIbjCdOBWZ11n5IU26Fx9s3xS6Nsy9/sdHlKP+MceZceU0EIbPfsP4GQJ5tjT3KW
hsyC15Su1TuRoIRf4Mj0janAB9RTw9GLgsUQVATcY2X7nqeYCViIalTElgSVXtj1t/Zah1YFKG8+
kAktE9FHCG++QNvuEz2R8v1Pegk6Ex0Xxwq2BA6pb2qiwtadn7JuelsPH8VFq2eh7tmTshElw31O
CjMTBVpjGiwecd3WwBhMebcNz55cMTF5FOULat8jnnEubbPf8IdWJ25SqYIuuQ1or9IV/CSu3xMt
j1s9fFbqUWDA4SiD1i9rJNOSDVfCe7XfoKbzT68LQW2/q+hb5hRBRr0Utr4bZb3KvhjmggYvSPym
szrflmf3mtmxydRWh5T5SfgJkg8M+DI9SSf6ZpvgElRWlR9FmCB0gaktucQg14tAKKS4PvIrMsp1
zob2qXKB4U+xturqAPj8RbqHlK/xYGw9JADOo/N3qFGZZw+O/o/2bkkOyOZq5A2Be+Uk6llLoUSN
vAa/RCL08U3gwIVm88oRz7DIZqXKzQFTIh5/eFUlMRzPijqJe3u4bRGLbbX+uISy2q1+BGMwVsAL
9qiz0UxxDtTJhS1jUe9xuvZ6ublMVsQE9P3vMIsD0jn+H5fLz7XEAVsgy8a5Sk+2vPrpOUeDKzoE
Mi+zBxUlKuapJnHC2vafiLwrKVYhSBSqwVTjQzGe4eoPYz+6VkuAssIWSd6hs0NqgohFtmTbXa1o
0tmbOxR5ryqQWGVqxA7do8aEDn9Zpp/3vb7dnmiaerB54OK7KU384wuUmmgLOJGvfhNy6EZTQXeC
P4mEFJCPlWAlcCmk8KaZRj25bmY+Q+gii2Fa5jcotBj75X75T4VnctP2D+vN1CibclgBs3FaKxOy
2B3wlhO8x7tM/iWp7oBtFamlEwIFcBwULbXbVLeiNGjDtFezNMItg+DIGYpTmOevdBomSM65vGKY
hFO4mJMt53j1XAA2e6MKzzzk7FbM/TLJnFJSpBS6hCC3BE8cAztloU3EOtwYO5Rolq9h7Od3NAQm
cEKT70R+f2+tM6pJ56kl5tSnRHlCL6Hhbw08/CJuEFjscpbqtpFHreAad69ZH5tMESWReJRGo11C
4TMWalVenS1aTjKzbxh7v5OyqyP/8EwbkExnprdR7pnTlU4uPrSPPNGBBHLW7wIRbr3mGoxWlaIW
u8WharOKnenB6FaqLbXtfsUJxU0Y+dKwM7a30VDceBh2Fu97zZl5/oiBn7F5ntnYtorlvGP5dhC4
crbpXr79gTJXvJw5Mc6cp4/dHDoDHaxReVGG0XATLGZSv+Tn4ELLCUwM5bi/ebDmb4nMJF7JY3Z6
E+6qqOedLpBEyQ9iRD+OAa01i9ErJzfqAQTUoAjJ6Zf2hIH9msy5wwTi+bWAzsd4LD7ikpwfcdRs
bsX2xJ6FZSY6d1jagYGfFxLXbAiyHkJ35sjr8P1ZTtwq/wpqA7qLndBT14J7ipkajAEwU/r/U/2P
o5EuoU//4+sWyofGDFA3M5zyqdhjl2zOrFI9Alsx8nEBkOXDxkBWk2VOLuV5XISYoXfmdxZn0WpJ
wIyaomuyTgJ+SkXPRG17M8wie/hE2r0ngDRJ4+LYDDETwvbdF4bi4onS3R50GZeHPwek3POHyiTj
80ZAELYSHZe1uP/bkFnwcPLGE+dPAM+g1hRCMw06bu4e9fo6dc6tOcQ0XvHT/MaJlNenpx/OJ3UL
BHJRDr12JGcbt6N3sS51REb0Fk8SEl91zI8HwcR9lcmLW4j5khbYRjzNr2oEjTslOTocxWpEK5Tz
7kMCOE4bgaTdrj8xaWCKOcWgJzSbDKhsp/Pjp7tdOxGwuf+R6ux4eiuK9Ex/IG6hzLRa36EuN/ac
lQ5K70Yc+XKkAzh8J/1Rdj1yy0O5suhUrN5SwC/YPchTZmyXuNPHxCJlvb89XpZbUK9zD9su6t6V
vOP91iYbqQ/bvc55bHiIkyMlaylKuNtj6KfM2KZy5fYO6xQaNWj7JblkbIXMJM1tzpy755Ezi4nY
sJq/gfG2PxIs6KuCOOFo8URSQUIyuYtWoSqu3B/q9EhURlv8icqs1UCynZBKLVMp/qMTU/54r/vL
CS86g8d04uICwNw+sYhccVT12p1TtEwUyylAMfpEzITbXrhhcWQlB08ZfMe0RltePqTn0sk7DEDv
+yNDW3MDb998m5sFlITrRylr6jVBMbr4kvf74mEoX6u3jh//es0t4vERs9AKbdk6vyVSJ7GNW30B
bMreT46DjehWiYUFSeAh6oYXFtGnMsak31GttkkgN59ubzgL/t3STW02pRR4y02KuTHEeZFxVLRS
RCBNuUc76RtUTl5Rm7FgelUg85EldAh4rwnpTYbs7pgVJIGlvO0nirAtrymjxHqM2vCGA5PT68/P
Bl4jeZ02xX12uT+GZY0QF61L7lcxU37MIsGBZyI9u0+8GiERKrCtEXUSJO00Ls8w5IwpzaqmpnlD
ctq2ckqS3J6SfRgK6jjBGHwAo1NbF40tHhq157yXWK5KYG1TLQ1O/R7iSLxlMhjlwLSAZeL1aQLJ
75z+WjRQVqOaPxu81X9qx9af8eMvdzenTxeMfOCCJPLmtDqpXPS4vevMEizzLOcVTmi1pq0fPQA0
4hGWAaSpHkThFxPOUSf8o3AOxVxd0uke4cGGiRPeJaFe6p7pNxYE93ssxv4THJn9uJ7DTuceEqWX
emNO5ramAqE+6Ys/ZCEVSLH/Ui0VrSp3JsJhEHJ5GcM0hxQlMXeaWA+J96Sws+bbm+X9h9JIS2IO
cDN32+P+rSShImRvJHqRMSI8s1Wf5YSMuyl9gnwqKlioptWxLK4xJ26fnMTmtEUefIVQlt6ytFMH
WXFx3UmTijEylicJFyCX4C3IBWuOxgE8fcm/LLvTt87bZ6KP6KwfdOeS8KysfJIF/qN4cJv5+Czl
HitukKj2uljJr89tQ50/PNi8D+lfNM7Z2FAwf7FbkuShXjKwQ2XbfONijmwN1TbRPgGGMrNUHd2Z
qK5hgBvfyD32k6v+ZMULsPY44sbmVn4tpr/In4UsHxz7jaSFIUYJDh2WMkchZwcFNiD7fgiqgqOF
LhhD9A3IXCaYHWSCe0ICQBBZz3hctBaCYUM5b6kGJsBqsQZUVB+rF3/cgA4KksfMrpSRkndn9AYh
J/rLdJzbWIZHZRz4u2VS0RsbHDD0qH8rcNRQbzojOohGYrNxbzGt6X3auramIq4PSD5iqqB8baIn
91Nj708MFiv+QSzmf3cCgsYot/WJvBBRwlsa7JXw5icTrjqv2QsXwS/7DB2LKDYIJ/BvUz/1lZxE
9PR23TmzfRRJcKxWZwlNP7qvYhGcaGf3ZOou5ckX5PVedoA4KETdQWu/qd34UL3czDk2mdbhyCMR
3zQpEXofi8f75Kj66BHdB3FGP7X7ffOrbf0YFK8ModPNYY2f3um3Q9g1mPu5R62xgJgkjePgsJ4y
8S9lT5P2Ke58WwGkMDJS37ZugUEZ+FZQw8kcERZGj1egWCYdf1KK651VzTX5IuG5hZI+EPSowX5u
eTfSJ0pvQ4GnMUTo8cls9iKClp5QOZsX4df/DVYzZYGasKRAug9MMuF9iIZiov5vmdPvSFaZ6Qj6
q6QV2l+xf990rf8fvAgHfIGnl6Z2lxInaMj4SJQzPz2eqOlOI10QiEZDQVIw8CYnf+TuDAp+75kC
otigjlXOiIBBJhVZN0gnjjklCO9E7G7QPixB5VR9A29OdMnqzPeIVHgplBNC3FtLvoyl7EsEvF+Y
jh4HDs0JzV2TRlKcq3v3qYaRDb7qfbk2/9v8lqCUf/vIbvnedtNFy+8xjDk+11rcI3SCr3Y5fzAT
92G127zcopTDSi7M3iiqHksDZyeH1i0y0J/IRjkl48QZrI89pFADDyqYw6qgYLjXdxFOIj277UD0
drZcFx4YRgQH+PfUdg4+bgdcdug9gj9Eo73KRw2IMfHaBoI1+xlCt/0/kFHH2CJYe/NW/ulrAp7U
GVtp1L6dCp5jFyFQEXojq55n+dMv5OSPHYi6oYUbn6Ib+mClcCWqTxKeMiD2/CO4vcwHdSQmFfqS
EftQUZd6cyz1Bm1GBpfyvnLfg9SDz2j2qnjuHXpU68IWdMfnjMZY1cdpBmkaCeP/gmFEmDGS1H8H
AHOqusE0ppzzM98NwRHUwkU7vc8h+dL5VBCP5Bqd+izQwZdk/+Q+VhZYC360pf4z0TLq7rDqrX/Z
2H4nJSHhTCMQZ9fHIG0mlMxaZt+sClHnuTEvj3Fz9QiFnsI7myqp7FSUjcFPh7PtTa0iATtctA7V
2+H5HRgIPVe4Dc8GO+jgn8vg7gdHKIC845joFQChTWQhp19N8/vA/qNbepTDX4TYiY72LTqTHnW3
hPNke22ywQ301JKyLX5ga8vj+OesUhpXcywexVJJUHD61WUm00fIa3nuB1aVNihVDM5/afoYj9Km
MaJKZ2AsNQuhLnStZRRSIg3uU1cc9RU4C2079hN58MEDXAxc3PGS4m/zujKYTdHDxUY5sQqiJM/x
UgubPAeVWZcoomdJzYzDK4O7/y56eGk++r1RQs93wiza50lIOOWydBYfXwlRXm53v1kZSqFFL7WP
Oi+JHJJr7KlRTFs32DDJuTWUOGsghJ2HhDJwP3gCmYQ9tFe/WQ23fKT1gq3ulOZk11Owzs+SpYuq
iJK2jQSaHMcb5IXlhGYI//Ge8NvMatXapm+m17W2GeEXqourZkEPrKjykCpPsd5q1GU03ddqlAOG
JMCZAC8NZxVFunD7KB5AZVSdLIMI1Ron9KujCqXWxnWMJoGFRSaIguNQufISn4b9uE/bona3VZ6c
kULpkMCbsRYqogJDRqKBdWHXjdP34GnzZrMxuHJokfgFffKWJTJH3f6m0fDu2s1Ufpgwj5m2BK0R
KhkzUQkyA0nJFcDGs3jgYfcOuVheWXcvHPG+qeqVvJsuDd7oRReip2/pnRQqh12/OBcJOqXMjDGl
vlRJEk0Wie3b6ibK4z2BOukn8zwabNOawLG1Y7kKbS0ZCzL8C8tyGf5zEO/o2H+znj3GRexuiNJJ
YWwcQACl9h3VshEN4SpzCrBvu/1VGcDAzMsmeQTL/0jOeb0f54+OigYCyLifVEHxGbrHQLEfrfue
eVSGYl+quOrmbCYe82jC1lvrKJBtEcYKKLkT+zTyooCrr8zWehNauz5mXfIQ2zAf0XbUAKEs62D2
ozPWxZ3KOJCZyn7ILHnWQrxpVcMvfi6fh86M/BnVsKVj2p4veB7y8YfnF7FYdzV5XRD3iU2I2/EV
ljiC1j6Gay36HOXF5EYUMsQWX5NERwpZ9lwIMC4jzF+z+9t1m4JztvNv//FZFgAs4aHDUiIIX2CM
L/0OLYhT7uu8QMTJ+kkLWanhvX8eHzHea2+DqdQa8rUOraHmTJQxbCrh7ndkjPZeQT5KNXwiY7Nq
FWsl7H1preATF3ODwTlkSLkWwHC05VpQ8gKcwtQG7Y0VtBX2VGJXA/sXPKUGFD7aFEHH5Lz5rm3v
iJ4UcPSp7dJMf9ULbLuoFKtQLiGilHsKwKV+zj2fWWTlCEdAf8k+bZAXiTkZ849IfLBjQPyMvG3U
XgVZKTAoLkcURhNFG98js0HvTj4KxIYn8iuJtO+C54nguedx6szvXQLPMavS/77Ltjx8gHlExfKr
JtB7HPdgff0uL01gCHQacMgf9tC7OlvgPMT07sfHCn1BMz7klGUFKq9RNWG3r718d3NjERoaEQMI
NPFhvH0Yg99gq4ecD8yOs+91PG+oNbeApKz2fFCjhOyeDa07OXQfsLtsUNHZYc+7TBsnSdlB6sQg
iEEoqbvyIHMFQRx6axHGH9KfXWcF+x5j89Cp94XYtd5RsaE4DjrDReqU9iwWRpb1Djae5BOzTc/6
9ldbtidAWh5HoRytQolN+jl/fEDL48UUZboqExt3tSbBpIcnUKyy2ph3XxjK/dK+QhYbN6xE8nV8
iu+MhLDUtOFKkpsplheQCamiiF7xWgdeZcPbcGL3U4r19zwVnZjziARayOYPIe8p/9M77I25Iqiz
r4zRQF+oeNGuY1AlfT2il3vXIVGY66ft0Ihaa5zg7oFjkYxMgT7BounJa6XJItDFzzhqNCNsfxxe
6GfQuBpSlwh6oJVMDhXZ7J6jft/iPz+oGMzHcAOfqQXM0t1ZGuIrioS8CuxYTjtUV5WijRIkP+J1
E88Izx6qgwI0YDRypJTpi71CchGNysuCK+F+e+f6x2VForo1YkHHVXwnO31SgUx+75eGYapEj+h7
yeajvRUigqrr0/L28KUrxkQxq90cS3dlvoumDN0yDDoIl6uRgbbzfa6YV5Zi3qsocyXESKcuFotb
6hv1VK5hDDNqjlpg7d0Esj+oSDkuv/2nk4hW7U3BDA76iprx7jpwsAht8ve/IFvnDrulu1glpAY7
6+kyV6KOXn+WtshVTOmME1b0CcHRCY75uBrjWK3rqDty3SAXrEbmQ8JVjR5buystnHf3KzFUQlOr
vNZ9Umcg6QB7p/SLOYyn5BEXGizop6bCcRfBcJNEuwN+8bkca5zXynRcylSHv+aqm0M4+RYhsf8n
IBDbf7iniMD6UbzMSsg0XID9SrBYJLa8kVFHNpSFDUmcfVTpifDi7EpcWs74Th1e5KGBFCqCPOPX
cioiaGmk/AD8jTHPqGGB8MBx2VjOh8HpLnaqkNhWt6FHoB5gHvNo1wPYLJhZjf3/FZkB+2XG11bE
okqEjydvdWTR6qYFHTndk+QZzc1h/UGBL6CdQTGhiPPSg7yhFS5Eubk5gdTedydiNCXxxTAuCtlQ
vSzeBYIbtEd1Z8QhR1UslcrNYnWGNeIPaXJzEE+WV+ojUtbiXWCSXNe81zmN5ijAsN/9HvdFBDQF
mEMz/yYm4h3MSy3S59iZt00ZM9H6aVAQl0tcELDC3Eoz+4KQQbraC09V3r9F3yMsnthVW+eqae8v
EJhp2CH+2vmPbfPkSoOnol/Wkj0mZJsVQu73jgH9nCTlx+wzaFI+Do8zLbX39Ok95x/hqDJbUiuh
/OhDpnUlEuezAyuaLWZKPD2RxSwJQBfD9ibA8+4ftAKDJ2Uj0nzKOsRXHrYPk0bDvn1g59paoPqa
K4OXcGGgQjb26q2FoF/jKMqWHKU49QFTggJ0nhjW9esMJiCI5aQvK7ZcK86rB4NgzFILxTINy66N
JFk6PoTrHP/vnzPfS2GVHDToBSzPpNk06nl6IO668uTF9F0RlWXp+eNYj6bYkoFB7mvjlbRqyfT0
mDZyjVLKGaWj4B6j9b1g9F+q3hxtXQAA1vBSSW02YEIeR3lx6lHLO4hQNMWVlZp7GZ4Bwvypocs0
XfD4UHKMF6dNFtqWsWPqx25JhHhJ3+ghQ0K5lj7Z4VVwFO0yKKALIwvjlZRGl8HA3nREhNIkwpbm
zm2a/Bz3nrpMMA4K0shu4qe6OwGLdSKJq3YDn5xqoyYr5akcx8fKA1JIeQUQ4QocbO9O5bxQjz03
rxFznqZSdH0HzfuKOy3z+b0ey4zNxKoy4UXTwAsWt/ovCEK25FJ/Q4hUDqDTdOiPoQX2ZhPKbnkc
D2McJRgIqMXnX7MNv80WcJkElRHC3fbfV0SnZGIg8zJDWerX2fDDpKQKCioXiIVNvWVw31xPM0Q8
AirrblJ4+5Xh3lsjsWimmh4H0lfZivoissHkYbOqB+LkFhlxMScIw77nWbyOz8fwnmvs2+3xrlNJ
Rb6HRqSOyb+CChjjLN7B53+h9mx9sRlZpkVAb8dUwceuLQ8lZPfK7bqDqj5w8cSpOlaCrJ6J6gq4
4cs4MzoCpovCIhP4/8MZSBDU4uWfgzZXPfxuq5SzJkrPKMttAdJCWxnsY/LxpTHyUM2DW3CQKLH7
Cws6GzCZ3mfgDwoqEGhFMPYaZrW6Ncdac/wT2phUDOIbDINhFShZwyW7sgtG4on/sFEQ8Rli/m2B
BaWag+9jdnC+OtXanQI6NDVDSToIqBbQnNdmKfePqhP+sbj5NDUTpTD9a7Hz1CwPd8ltzh9RKH/D
4IbCap7iNUyIxY5dRKfqzHvVM4ffhE7WQIzaxLEgu65NJruxCMh99q3a57zfKoSiG/i4pUZmpYQN
v0E3Ezl/EsKhcGomJO+w5YTKZeGqAY3cGe7bEiFU9Fk7hCOcrYEnJvNsnGmwoHY3YZ5ZVawZ1EPc
dT9UXZNpMkyUP3cGSdjwTT0nLbPF7waUHJMNkK0ps7DBDFCi2xCuNa2s6wSZ2uHUwKYwjpCo6l1A
5sfE2BkYwvqPMuXDyTktR1fAztZJypO/1XTlENgMYGMgAoWy/2M+Mhm2TA/Lnz5dJw3XT5/QrtG7
mG+gb1LS7WjgTtUeSn4UQo2B9PbQ+Di8j32+m33+HeT16NWdcOoWNjiFlAJzrCt3xxJO4YOn5tGS
BVKKPZH7k10NMfF5WtcuqiyRT96djYEYAeLuYmEtU5A9Y+aoZtv/61dx2uwpd4d5+g9vlkEf68GQ
km2fiZFns+4TxbK+XEF4XFPRpNIy7sLD8AWlp6p84zMym39YTQS4GCPk+gjOhsP6TuJpNOw71LuM
hkvVpSKRXpIaCRnbPPWkQUaVyq+/sb5z5iePGe1WGCD36TJLx1naO0QWh46+hnebrIbjmTsjSVMD
4ZI1HQd730BzjV+qnz0uSGXRuMaykjzRgBr07IpTZ2aaSMxchmsf6oEKAHMWryYY7JCnl14LdDDD
OZMzs7B3ec8luKKKONv38XH77IQd13EQepHNwpr1xdtQJoRIKka7B42gKooxEom4q0vXmAgQSDOq
dLOpkQs6nArO3xXNwHGQtmgBwNy9tWPe+BUVadhwzbbn2WymS+4/ELAj/FveMstRQloCPXtiwHM3
yJ2H+M7vJfYKDsIzt3OHy2AwM7RkBbHl2vd3L//4d8xEugoL+UnfacEosAnmMxc53d4Zq/4uSPiH
Ka2XHbnFKY63Lhaokqq+8V2ytqrPAH8q0WPLAMlxk26KoEFTVj+sVBHSG0Pf3wTZtGd0hSW0RJyk
zXvBdMNXKf5SIcEWuV/sWd8wERA8CLuPmwMLK769tXy0UmCkM9hFAUu8MHE1wTRQQJAEXVVnHfg6
7SPqIRUUArAU24Xm6JSUvCf6jCVbrAufOaftFvVmOVcCphNX2hsbk10+Gr6SOBPnfv5CSon33Poj
anF7Qdw7zL0/7l3rgF0DmJAXVN380X/Nifiy8KFF9H5ZCrleKgLFRZIDYX8+LH1H+bAYcM12OWGQ
VHR7GUFwyhxdyk70SZl4rAXcXUqLT6i7Ksx+Idnu09BitcAssvyWT50r5rcp9fGVIXtJ+Y4iD6Aw
jn/LkcrN2GSjdj1NZispxDyh9Ozrf6OGrPnzrr90PJk/+zByWN9aRg2g39RI2FpqAqW9RrCSKpdy
vy41Q7v5oUt2NpOXba4enlpH3NtJ2jc59uOeMSqAoq8GxkG6vCHWZ840dwU2+UOtMNqyAs4gMbSo
9skRTGXzaKtjwoYCYTxgZMCPqik2qwoZBAP9V6mujFRpphbcCIhKbseRjMhqC0hioMkdiWtlDiyY
5zJctfuGIHmjDCbjhlFWcRo2NEZZhA7i87XPOVoK4NzC8AvnDv5oGABAA6hEm2cxdW5kSn0CeVh7
lu2uWZX6b36NNfJcXS40nXNesBirejGTQBAM4MsaClu9CsB7riaiGARLrAnOwpqbM/Qcdj3XbeFh
1WBCXwtl5Of6sriWc3Voz2m7y4o5gOcnN0F1FsUrnbHricUVQeTZJ5LkZD/Q5d2vcq/6ZkHNB5ks
UPFJMGnxPfIPW+7/ZdcXyf2TzzpngM2BUrRKlM5ILm+ABVoqhu9lHpWS4NQeQKtf8RIgBdQ94AuS
xg6MT9CoA7B5M1R6/pFffZBhC36rRark8jVcMgSZGsaIiqEfuDNcHHheyupS6hldtfB2d8VYtRz2
eBbRbRv8AFRfJrfalJMIWldEQIpdKO701j0wXo3Y5/To2ePrXLlkp/xUCi7rAtWOEExw4IwwzCAg
ObICIcz30v4Xg8pqTVPZknXF+WyHHnajP1ae00U8jLU03v0sX5xARritfyIAYboDyTEwhzbFY0nU
X1jLOdI7Zyp2A5+RldlHvWmt+advkR2LMsyJ+TiYEd2FFtjHBWD0ZwBX99WKeEdi1fw4LrNsjEOK
cFL9rxSW2AO6vGkWyVnhaj8BF9cH3FSvc2XRZAsvuP6lpe8ZfTVJlYARcT/H4JqcbjyrQIPIqzOa
baCUU3UbZTuvnlr+CqllpOAZlqo/FDdzdHL2qR6dceyyOkhePbnylsp9Teo80QP4u2twCRSNrTUx
kvf/LKP6qwL60XkmK+gkPil1tk9yRbacWRlB15H41XSnQIb4cF/aee22LYo/p8LG2Rat2Y/Jbp+q
IFUFL+zhPIaYgXP2IXpiP+Sf+bdTbjs1P0MX3J9UXZhnzcmLhDFTGX1e8BRnpjiZNzmSrUyosgb7
qt3Q3Q84BnM3NVUv7o2dzjLVTvuPUGOx+lV2EKSOi3a5zX/gaJO87Gg6gzVsApQpmYkg6yu1nrnG
txi/ZIWT66AxgE5foa63oOmW2JTmKpqA2zkAngJ4KT5XgV6oDaXBwz2tPb30MSIy1SCQBlLA6uK3
MQihLx6KEIEMGKGIuXtOcq3Y9yXQMTsr4y6bL3ubDW0B8jsWj75VnnMPwzhgWEEGxuPnucMsfOnK
pWoRRMzOy9Ce0WyJ2C+p8U9Nxj+rAa5nwwAHCbPTz7g+qYaHTP/8apN9Ux2m01spzwFKAhF+OI2v
+h7G5bQt8CkoRyKEvR25I1zCYLG8L1edAWnTkHihwYnSWNgtYgk8FaDw6+eEUEtuKBaAedMMXPyX
KlACkZVXvBWr0PbFIJkTFbRTDPtylAUZshW3kRV8/Qc2wc2judtCMgzMtPOOquXYFj5FyPBSq0I2
6/8Y4kN/vVZFdaDCyz9qVydhJhxV6Y14dezKpaMjndYMVEUsTo6MSye3+Huy8LxYusmZJL+QblrK
djQ1FI5HT4FMCBw4ObcJbQlq+NENbq/gtQqUBWJ7xrVVAp7SqwtC1rHBXGKQ9uiFaMJ6JTY4zTwJ
RiKoCnDpRtaWdwCUqhCIgN533nKBhxfHimCMzMPsWS/YjoWl0mkDhqZFjKnE0NrJD3IL2j34mpEO
O/WW7o2P29hYOewE13EwR7jaMZoPnwJXo3ZXu9pBVWEqK+dq1NL5KswaGcrIX6jKF7PffhrBb7cX
MFCmf9Gf6iGQoApK8d+T4npKPHliGWLh/lj3/1hBO3btS5SzpfqLy4MP6DRaPTABngc180HY9GQa
7M3ZC8tOASxLzgVyj/8am+4SDIcDy4y4qGPKYGVgZp1KDSEamF2ZOsCFhj2aswm53GQk/grphYro
uKVH1KwmYmy5aCaDnJKBrinXBlyzWuN6HISa8tzX/OHRQsudXvttH1Xtwp6TerGDLJXcZeWXdIKA
E9eZOW02VQNRfbUNnrlZVw5at1LayIVUZ+GYKIUy0YMu3lFPLZS8ZFG+crQP8pMBhAM25EzwUKod
H90WHtTxnZemioi1KvbGykXdt/KptJ7oLTL9rDxXpGndY3ZHlXDUyLY6a7x8X8P+yjtegiq6vImw
69ufdMHuBfLXWWYtyZFurwM57HdHq6tq86tvXKWhjFGelWzOJN0C3ogrWjq0R+bXunUYQSzNqt5d
TKiZUXveOSwdcrvLrg6smtGye3QjCKEOAmrwEOwgiL/75QpG/ucORJLIFIk7qVutdV3fT+rVnMSr
zaLwFcTBUd1qKJkaHg/tHp/9AtBhZvL97UBv42i5M4xNpyHK3X1xc6EdM3IE8oqZMYobh94y/F2q
IY5LPMk9Y+WKLhc2O33wbUkSE6W3l8nxMUPN7piV8QVr+D1Uw0CDzkFClcsFtxXdFA3006V+QLIM
AGesqsT3Nbfs01Yo0soicv9VCyURaiG3GpkByoQn8uGONPni69HucEyl6xSNtkuf34kLUzQfomHk
UwP4iyM1407Mdk1ZuXM0t71X4D1C+b9MirGT4Qzbf7sBxJyigz1Qw2NqsBXGl+6lFmKH21WQfzK0
MKcfddrgV6mfQG8/jpYgukYBcHAjEH5KP7RDFyunaXVkbyyK6E7Jf4mStcxgtrPZqvVdr5pEN3Qj
Yosly32IwmoTdjABgqT5uke40+yPuLGuepNyf/mYH6PmLBHNQBLok1/99Wh29GH+dIKXuNXDevXg
U128gcr1U+Uhpd36SyK2IHgBtBgKan7FWLg9Ea0yyiMMzsOTwHpoDeF3VkbV/lSCm6vj023aKE3y
COEB8eQp5yhsYtXDkHc2TDzm0uLvVZgQGbD4vAywNMXoAH1XXrDm2Zaw7+oP4dr9BaUFg9CCAtFQ
3EFzjQpvcaLCmtLTcJoq2mgyBSv2yvycvJLYg8girLYyPA3TGI8LdBLUT7jOAcp0ouPZ8mgLH1Se
QI1KjsQ8atPXUu6qmM3kQqUI5LMRN81h0y9xf2wYb90YWWE2mrFaENYTgOmGa+JeSy+FmbwWHA+T
x/1v3IkJd5sG1XtAiowFnXMWM4ypEz6ZWZ8o2e/xCdnF8NZqqS7xt/hRh2TCPAuY+GAtq00yOFUf
NA5GfwZ9y975H+Buf3VQp5lqqgiJmlxjeENPk8dfL8O8xjGKMLV29L6NE/XRwTAld3c7kv9QspZL
x52EDE+mXXxKPG0RfUWGyNv5aGg1Zh/rKCpv8UhfeWowtvMN8j8WjKbBAiy4/WL0lld1ZqL6daVX
Pd94xXpvcIzt2kKamtA/XY53OIe60X4ta33KJyA7nWfIvvnVYYZLO3sX6DVM38TgjYu58JI5BPgC
cggsN8nK0JBOAu09oU28JNEk6Zvx4SNqV7/X+a4LvfuE3beZQdyGRCtWcW0y27DEm9x7WbArSsrN
ksuPPVNHtNWAtUy1jg95xAZkEd3qKAhKKTrE4PN9XBpxazxpfOTaa89nrsMO++CfAO/Vcs3PnzZH
Z6l4UIrVGnqrFShAHdN2rFe+fadLb/6XpYVbtZfVHB2KnLDuxOiI0Kdojm0I6GFxeNO/M9dICfAF
iIh1br6K3Q1+w7JWGdde3e+bB9WNrlaaVQY4oS6iNuQe2mElSO0gncCRxX8ACBO2CBuwy8ACXP8R
382LCCYrhN/dv2uk7ronkPlISWwHJPN9q71uRxuKqAGkShHeRoj/cYlcAz4EBNPq48/FI4U2F8o2
iP5QQIUlJCjWWmZ/svoAn/lqBwmYbSNzmTbAPsi7sU2r6nzdGckbdyzjqbazaKKfg1T72Idh1KJw
sSRl9QOqPF/VoLpNz+EBB4hOhzradp8gw+ZyJhYvVV3vhAEDgxtfpKd7zdeBT0NdGSLZvIa4DLpV
1xW4bd8h0fDa0by9dlYoi90jKD4TUlVISCseRVPUQ2Zd7JS+MXaG3CLol2lYgPai8LQbVutyYrYo
JS6MoytpFGbj2Fwp3a9ATKR/ZkvHC/qx5SY3XaMmABLZ84cQ+4eluckAgMnb0Eekmk6v0qyQxFI4
MeKokELRCykDLt7EN6DxmsVX4Q7bvV1QU8gjdHIx4TvYi8Z4sOLc3+QqlAGQthw+hZQaxMl5lweG
eEl03126CKMTztgcnRfQD7khGGSDrB3KBVgwVF5sX4fqJcEDyrIQPo1aMYsvB87dZhnsdP7zs/tt
fdfvAFgCJnjEVIQscjzuo2EOsKJu1waN/xEHZn7EitJ4WIztbGydM1yfjgTOSgS43QZ+Dz66GIVk
nQvaVXtF5WR7/fAI4zAdyCNzCvJlxyvEvCw/fTDKvXoHCpJtHrNP3gS537OrRjd1Gr0uVXXYouAH
Ak4674+X8qEtdq0XJDEfoMu9wuH32tx3jsugn/03wsHQ1x3Ow8MoY3vbeLov9DMWn7k5aVN+WpAq
+IJzOKYAdM3Og/erk357YgHHkEsgACvvzF5FT/fadvhjyutkhUPfCch4I6YW0setBnEStMaGFF/K
duLni8ldHBCnw4r85fmape0WmgaxUk4jZjjPYz13o6dA746QxKJ+VP2EhF31SZeaJHrG4IQ+dgFQ
Oz8nzc4n4+kWKteDZNIPZ3QXTIi0FD+q9B5JwjpxUMnKhk+uyf+myaRsEXEhfRx19BCPgc+jBKfn
Ctt/E6jCZ9zFR/G6/AkjCY+ctZlrzPIq+iO8fYPQ187kQbPHjrc1+tK/BsqO1UllbnG40MiEhcM7
LVLOOFQbKdfMEjJ0HgQiyNyg3CNbOK0KL2WbPobne0LorRpJKnLJr5ZXDEsTfjMWRozy3mHSjvhK
L5sO16hanIlafpqFCWjXFtl9RlZL8X0AdnzIbkI/ktP5KVftgXE06KS3TIBHGAp1ZZHmPvvEWGfn
WFDXSzGhqJtBNQVTwF51NBhlFU1TcIUnWm3eFwiQnmZqtZsx56TdCs3Lf3VoPLZOkHFNGqsqIy+J
cp7ijgCsA9wYhE46WWB3DskfcRfn6dn4A+QM5NVK84nsId/5a4MgYYqSClJq3JIyEk+1oG6z/eZT
ZJQN3oJvQC3NNWGcA+gHHqNTF1iev3tHYjA5kupwYqm9JhoByDbGEHx5pjPll1BTRRIuF33tw4oJ
Rn4JS8p9Xij3WowUOgXHwcoa+XTVqa543HhtybHSt/beCvE49t/obfHvEmTsqsaoTuiNAcvQrXWV
bYIPSuuTxvG38IE+cS4hZMFX4LNjYqVeuRsjphtzHg46gHKKbwGk0ctrg3ADepANoop6yOZ88VaZ
AmAIoAE9RGoXlWxIgUT6JV5Oi+Br1zqfQX+0XHmXpdNoPXtBLmGf5Ud70xwVPBKH9247y4azClYF
5+LYLtmBkIbGSxo5o/yiD8NdtGDKkhilHaGxbK0i9hrzyZcG7l0iuMbKZDG+gs9+Ctkv94ye+Kkd
zarbTGLlocdlYrSCZ+zlP1y0KICrbe9raPfu3mKAAd/d0GpBm/PGZE2CeGaAXf4hYocSY6r31PJe
spoDUrSE9VGKvkT7SjFZTC4WWuGd2lOMHuTNrmp4kJbETPpDvtasH6opP5I2YLNc4QE10jIcI9f9
Ylolaelus18Y1VMbqlRmOXqJ3o21buaUW3dFgc9am14QYycjt2wWZm7sCBd9PXAIWDxU80Tz6DMa
kj5WZZF6dCfgEmQ31qerf+qcnbZnc1GL2oDqCCVvEqzmwcAY2JsIIKnb44agYqQ+jhRImtL+zURy
BlXwRyoVHMGSwb7tf3pxSy8t5gOD8HmGA975QOM0gz4GHPSZ54E/6+WfJ5oGoPwoQxLbvFCNRPFk
1I0+GAhOdpkX1oexqVhig24xzu3SUY9nhkG1Oem0+RZ8KPgsJyuixqca5qjhXdDHi4zBVFeshqLD
C73M/ARVFwDIuYyPhFnub00Vyz0VPYE2u5FKUjuSq7pZ+/BcyaYjlagaIC6RuAJBOp8cl7eefSMc
NdAyiteCzpWp+HqrD4hOSoShCGpeeT6lNaRR+jrM+4FK1KcfmjZ3DwYMWdjDueZwxmM9lwnGsatB
WMSz+3ECR3FmWYEa/kZ7CP+bPQiii1bvumjg5+B5dllS76uVCAtdRbGRRqhuHSx94jhE18Qf7bJk
eg89jUUFDVdqVNahizPEjavGBzaZD9QKzRBml6RrhwO+jM8nKourt5j+PJVxHlmwWJWxCWIsHcqr
U6lWjLLWg2kxh6ZV2Eo8wzqkCamTGd8xBQoFTaVEC2JajrD1Zo16EPKvO8bECJTZEqsIewdrJhDF
BuK0s+w57iZbWgh/yzORoJHSVsDVFWGJwcoggH4XVOT2Ha5rkdiqNxfG2slUAJBkVWyo0XBey94O
irCYSKkkUJgQg2w+0TMx6l6lZrUHCxS1oXXoxW6tklOBAJkHqcAXZgJRdi8ZR91oARR9iwIJA5Sc
I5UfjiDwitVoJ6yDgEkwci6iUj1lyeeCYPvuStZzFGrsBfd7fvjZ61PdUXAQ+55pG/EPQyOyfSw/
R06NTi/PpalbqwLxZxlaSIL0USiNaoBsfWxOnW4SkcVvqQ1ScSye5Be/xwYNLzMrNE4dkd/vMIzr
++0ROkT3WFjVpI16UNttKEW0qEGcx8D0l+gJYr5QvNysMAdnbmvdLZCjQgUMY8yTkjI9Z9xzPGQC
/62mkGDW1dkTYNpSDehRPHdgufLvexX/X/NbDrrMdH0yMTg/RkYWw8Yqfsg7IGWgJWJMLwp2a9Sb
aTHSQ485yyssiVaDVvxzheXssDtMR9bkEQ+vBSC0eI5fARc5bt84aNxtOvAWuz0eB4fSPYGrSpeO
+Q0yGx4ySFtzLitlvPfFvqNE1b6tiHLKzdbSub70z/GxPslBSpPKXqW/wgQfmO7u110TsEwKazkN
KTli1Y1n+ZLoCtqrDtQuSW+og7TeR4tY4pVvBoqadWv7CIhYvcrnJWQCtX/HZ3O0SZJy9Dp/Mm0+
5OoIQHbu4oZllIx01cVzEdTfemBJdXNZaF6cdklbVpNyi0lqHk7BIal3sgnpecXkF2d1zFKuyWk5
Wnc6Nc8DZ9rwHzFb/Dn5Bs1xuDg8kNuCldPLeQyGln915jaYUan+WM6mee8lj1b8t/I8dF1btu5I
w8l9H1WU/q9dqGb6LdWzOyghVzMC0ihyXqeP/KL0G9+Aiao7IdRdA0jg+T076023LuyAVtcuCokt
Xc1wyzqnPUtdRJ3oxc/8l8J5snvLncCkVs07Xhzzhnwdli53VCLGYV25MMchu40YziYUqKEu0PR7
jwau43t+yp857q8uxFSCL04jP9WmW0zQWizW3gp9PdJ20qywCAQuMjw+ja9ypqFg/4QqKBsiPulJ
8tsZ+vp1E64a9Hbne9dTPFI1BHS334pQEG0qZKb7u44jfQh/XmrZUSVSSxTNUuW8nXRYJyid0CZD
nStuaGNfV+78gmfRhVYjORlnte33hqduqhn9SpZsD7hKr5IFQpyOHCQ2hUQf/7u8wokMObgpsEvc
XCa89Xo+sj20NcoTA8peJq49PV8MeOU4RtEhDhLbB90qJHRPuFF5zW/lg5oEK236lNmNHRpb5MX5
h7a9JnRq7cGCktUvmNEupYYrso1wt05ob8WKsbTDUEOqH5xPW+29X7MelvWD0Ogh8K85Y9lOdt0X
HuTaypKgWhkQDBS1HJH9sfNGNsANwZCT5prZvjPhQ3eaVDh3AjDBS7oIBYh6mot5lIIWAy7UQTg4
UedZIe//KxdD3aKZoBniJgKybpQ+ytlOHIzCqrOtLEr+rOSCCLMNasTR0xpihP6UYWwX9Q5zu6Py
Ju3gjof+NxZ/d2F1oyoBE754tJwZ6Wdcs+R36lrx0ceCyrd2muciFja6KntUIUDhMzKo3qZe7rRu
UjcxSWqBUyEIkzCv72gtpjt1vURUC2GK/Q7s9fzn97epZ4uS55Kyp+8nLOsJeOWJYzDFd86Q9+ty
QFQDf53etANWdkvbyJCwOlxRzDLX8j5LwfvwCerDGgcgApdgew6JkWEcyzPQbp0qGaJnVljHiNKS
IELkLq3UG13L0dDNvX/sapZX3rNYpw+6H26mmfLQwtqWWgv5HqAtunYPvMQfCdn7ST7CLiG1q0TW
D/yVEJ2NtINR4jEdr+ye6m3DltCIcO2C54gHCB3HSW9FIZ+2jON2u0pSSCJc05lHhh6QuQ6iUEer
j95b+uBAu752/siPLvUtxOBggrYKnas2r6eWsPm/ppLCk2WfN4Ene6jX0bnZiw2iXgU/+s1mKNA8
j4GUSjWD9KhuncZV+EZBDsmOKUSEnIsNUy5y0bZnxutSnYDfpArx5HY8k9sOjsA+ohqkcgeUaA5M
gFfhNEZOFrOQIwAoNUn9r6bYEj6ab5z54xrFg0N2CkqyItPbkB232IoUBerW9PHr+FHPx8qiLSmo
VEreXsncEjwcoS8sHW9qQ2Uaf5s0m9GE9fvKFAndbNuBCxWGNJSKxduBKI273EbktmSPX85j2QxB
WsyptVkIg7xyL1hpBZjqXCchzOzHGzllHixnkf1AnFcjGjSBdUfSotGawq0MOIni4KyROwst/pU3
VRF5Lve5Z/UgPF22CisOO85Ify2ThXdV9+uHX5UTRKilBEEKC4fifeoU+fxToqVw0NuR0Qb7F6nf
48K/9jKt+cAL+RE1dzUFU4goq9LinQsDbfELo9Qr6jVzVaFPfSxItnKbLmaT1MUFg6etnrUvuqnM
1lUYngv9HCGFRsepcNIVR7C/pzGlDNsJ7e6i8ZzVGmIGTNwkocIsMtuXFgEV0iFuGGVhz21vA3sc
KQK63KZh72+ElfrfKs9YN1ddPqpb/3VN5spLYwIgBA/gyev7ZDcIdfaIgj6U+8G767uFFBdsSOan
+lZTKEWzDfU3iiPSAghv2xSoEopeQptGr6xlPOl8ijftp0cVbeXWOHHrrjS7bpcpfV0GzC4yJfI7
fiJmMzmJjS/ZdDHXsZMC5CHEjNQCjnjcrjmeiUx7eUiicixGPrJccozmfPllQoq4J60GjOIFAiXk
MzAPLmhRay9eOIHPJlqeIR0pGH6JhX6HhJtM0DbBZo3ef7aucUcKuCLts4VbDjqajb/Ohmyebd1q
TL7K+aimn/4l7f41iRGK1PLwTEyJWAZEkrqt3qHARZ4kvaBkQgUH0+nVcbeDceVopAiqcUR5w49N
IejJmEpJhgmw8mSmQycZP1Vg5lQFstQYkUhBClHnuwPTP9kkwy2PcH4q8CBo+rfQefrEcGBqn/BV
Cp1f/QXtb3mtsA2xEOI48mOgdvMSIi1o/lJnlYixN9SzSCs9xr7bZOZUW2bjL2tsziLbwJMYilwN
FBIEWjypEEsKqG7bVdn8fdlVfwsFbcVv/eEOnLmR/8deFE7Mq1za5z84/GfFLowYTGQu6AG7gkEc
NlNuryQfUwoDCEoQTdDbe+yz1OjvmpX+Gguq+A01JBqL1pFAricFIJ8CRrMtgj9SwjFaBZ887x9b
JLPc16SRQjHXOG0uLYlik4p9VEJEwVDTJb9i7FQwWQy2cDtPLBYtysfWJqcsyCGU3+Fol4OAtHeo
I+4Grz2R8i0doe79wCbr6ZOHaRoM66UzBwn9l5qu5bTlEWY92Bx03Au8p1teXLvKQBG+71HC3ifb
uaD2lCx/JDNGx+kd95txIltxgegTaUpyGVL7UJTm6wGFUVfPhJVGs2aifSddzYX0T3hWIn2nAK4D
CM2d2+dF9SDEbLLw9+pCmDvlBJKTO/HrenUBWcOF7lpzi2+YbQ+MPaMSHSTbOQJBwpp2RjECCzbu
8oY5NUA0F9/nhrzrMDPSc+X+hd68XIBRSLqNHVbkSZ9OvkF53A1oZvA9gH42pXF4YVB3IPKU0Fc3
HL3tNKhKZSedgRTZfp/ugndCtuo80eAfMS/pB7/dAsavC+2o/QQI7GiDuV1Q9btJjYOXvP5KEwrs
iRC4FMMoFJKArcDXd3IXMvnUPAKtlLB+LltbyvoDVBheluJOOb0Rjb0PN2XIYzO5YB/zBGZ5Rr/M
5eudoRgnwmPIEj9WocWqa7nID8nsYcJeVUk4wKiWKRoo39Pk2H+L1jZFAV9Go7Fdq19E6Ji91VAl
4JgD0GS3/gBwiysAJ6Kcc0q+6mQERLHuuM5UKqSljBhThrQy2Bhv7Ke7gGQJrVBUDvcBq9gzMci2
pXxeN1AiREYVAaOae08cCx0kdPEh/oByV/ykC1s4eEqcV3xTzZXSDDPVLTKifku5+FWEYAWjnE0e
lu6qGuHOdtrTRwtLrGzWe1HI5WBLXrOne43U4Pj6VRfqySh1MdWWBQtNlyau/005+laTzq4VF20h
SpmjuOPepr258IqWvoYh/wdpXIT4vDsl43t5hTiBIDGYqOeF8CNWSbbu8pkYkDOPnVcIYK8ddG+C
pAMRBB1ldSo6nRtp/wxowU0Dk6cr4D3qGGVDtm07NIrm3E5fTesEinK5PmayyRgO6AzLRdGJP2Wb
Ga0yMtuSJjdTwXX9CXAI+xwOTq6U/bQCvwsimX45xHGqf6x5f5ER2sgPUG4TriqI9u/aAZyPTEIo
Q2V2d8m3CxNQ17VJpYslNNovm7xpK98ZGMYEXXw2o2uu73zSf9VTWxOdkKIkKNXQhiDAdMFJhrO3
NgtI3HUgbyTqFUcekun9Y1D2GuLnXLN+JyC3aGW3ED/XlmBuC00uDI63ObDFQ5NYwkHQwI6LiawN
yxBtJjBV9clvx4nze8mNEiOcZshDWBqgh1oOtH49+LrRxWSXVwT3mygEc8PjqM2+CtnvhV9QWT98
jEaON6UoxRzTrvaK5DXUhY+yapxDyPOq3u46g9+wLl15ZVWmIT1IUTQ8ScM7sg+Ua7LIHubM5nJs
wOMHeTZIaaM2OB5f241Ca672yMyfMaG9uQ7I7XgodphgiKRCXKMMM/K9Jh91HsRaUY3Gi3bxcYsB
EzsVBUJo0UQYFzrAqgSKXuzS/lOhAM2Utoz3Doldsb1LYb5WpNDP+5vXnaZuzxBHeTkXRiSQaxj5
8kqzFnkPbtT3hSncrIoddoZqL7aeUjqCs80sJWEkL0b35VGfpUCwaJEP5GJ1pkSKj/1QhQB8TkbT
tBTGgvY1AgW0ZvBSNIqAqVC2UZOK1o6y2B1j258xa1Dp1gWMgYqN1s5f7MkHxe2I1bBlIT+YS7+N
nQvusxaEwVGo7GDYH/+bYBbXJ0lr1GnbM41/JzbtilH9oysDrk3/LkTl+WxA2APCBjZ9OFfTxs+p
cpkEjKPAqCyASW/04Lq7dsmx39KvLZqB+P2qsRTX4PpJX0IPOeoYOD83qRGsZ4ClhHduyyGrZohN
6pSf6MbQYtkvl6I+5j6bNPs5pY3Bc90NxBZX7Cxtbx6KaWl6bsdBZlWhQJpBpZpayYBMlqq9IvUy
m6Li2XA1614DgFCxxW2iy2vQ8OQk35PgNi+XrOdmCQy4vlBy3zitqY4jlog15W9uicJPyqyTJLAs
XmsylFBBM7XE5Bz9fiYD8fbNjZ67VMUpBQM47LkKqkX2ugocyfkIIxnY5fZfqabA/zaM/aFuoZXK
ShjizbwTzWXcHxEeidVHR4vHWsCNuX02WKwdcn93rc0RgV11hdWaKahs/oOcmlFnkrkbr+xEaKlg
20vmICcMzdauDane0uknpP9fF9sQ+AmYDK41a/bzKGYRuaxuAuOWqUiJ6SFDpLcX36WtOA875ALk
FCYCdoqOnhAP63fQ1+47yb11LaGpIIkirZPW8WxSiOsFU8ds32UIeD6iDSJeXi8OUqoSvjgcUf30
ZaFblxB7KkOXEqZRi07TTtPTTKvZ7GN34vM58/NAH6vRaqlqoEo7e6YJGOu8toOKNDRuRHi0+qHv
BfuMPwIfBPjQjBnOqdQRRF+P61g9w/nRO8DD96vXeiQQz2opLFsh5F4f45XvW1Z4+zAV5L97wgsl
r0O6FT3WjgtVr8ANKWlHIW8/VAvX37A5pFl1H9KTbtomlhSr9VAzEHy9sgbm3rSSx5ZMWU9FJ1A/
h6O/jr5qCfKaAfUboZfSDrhR2Epk+Jg5gu/znY8Uxh3jGBYD6/vN8mLao6+f4LE4Gkp2FESK+PhU
6D5FVcMiOmyR0GVt00AWtx7vQuOYcOLRahiAQ3zXPOKe4MqdXKrSFjoIKFrLT8ki+FAGmpmS5J3Z
5BYvkri8IYbjDZC8BBK8hHdtdd02wbb666n45mVwGGGDo7rguC9uEPH7xhQc3AcihT5ppf344z81
pSMQJ0dK/oA0gEZ9mPG8Sc44/sq3R229xDhGdo45uK02tBUWYjSpYz9L4qF20tA8yqiPXLxCrJfZ
NRdHC/5I3IEQWcVnGIcr7PyDbZRI6bDFEKfTy3z4i3RnHITymHa7AE7Gbj79J/MYzJaGaHlgq/E5
p6HUPX2GwmrPYRqe/Tm8KCAwrR9MYTHPs1bgOyR10IfUL05M15mp0ELjpD55ZzaQ9d2HBmjGFzCy
epkdHnYozLX4toqrOJ/MyXz7H1mFOHmTcn58dV1fBFbRXd4Jl7V01WWDx1UfSO28ecwLgeKXSasA
OgyAK8oVKauqTvpbspZbqcu75C5comoGJuE3m07NmuCEtShmKoWMUZVdHBQCqgHGCTfywO6ivisa
J76p79wDwu/mOB7rrn37UVj7STvhHn09eoHHkN6VW7xurSs2Le6Xu+18WynNBWzXhwLdm2/bgA6N
jqfeDhP4Pd2lQVEopVoX8N8OeVP0m56CKhpyahjf1jbWYRi8JFvLmGQCZzLyWCpAANxW3UdpziLB
qMfqdgM6qKkMEhTI5QecNggC3amPkiKtH4M1b3+z5P7GbtVkpn0MZ8FJcHpSKZ4mhRu1qDH2lFol
JL0uPHqgk3Mzav3IWAAj2cF0kv0+Q8DnAMf/I2fG3QHmIbNxJdM4ERbfU+k76nKtFeMTI83XdGxJ
OVT0v56OXh8zNSeLhyrXb/5SeH2Hf0V4QxuqXIzV445MKyWO0QSFDS77LVi55qT5V2jAtjGSiR87
/XS2Td/T2Efs4Q0ZD2ot4d/t9GrSr0SDmgVWE6NXpN4yZWtCteqA7IztE9l9pUWvV7I2x2A7wSs+
4cvtMgYS1DMz/t90sbKwiVe+zYq+nFqsh6clbOtvZBVo9a++lBQKJhSB5ax4L6APXZ33WJJJqtIq
5D81PbKP12SsJ2+7IbvzUprQhZb6ou1u34f5VicWOWD7pEBRCrNZVvtYILgu4L+tK6y4g8rDPlZE
zoZlSwuQy0jzjrhhBXeAZx6hSwWV1eeeFUrx8rV0DvCUdEqOCbU2+RipYge/woiYUUt1KZqQxl4R
TFBX6UNg3v30MwshwHkX0BWqnEWBwrFxnfrTVhaYFTbjq2MFc9lOY2iLXRd951AirYT2SMQvkaYt
leWqnNLg/I0XCEID/VCAy0NP1YmFVgHsSoQikYBVpkyE7coDmRBSEEFsonzXOMgX8qWCpVQUL0aQ
JqbgO3FrGMGHowUtfQVJqfjmrVLEklXLdRlKk840bz1ghnqTU5L0ODGqA6/Y0sgyAcHZvguh+5An
DbcHiqQ4xSCxNityRtqu5mLyakx3raCwjrW8cEf5Fz4Sfg0ETM1KyawPeYSm9+IdSPeZukkMrgYE
39L9IXJBiUuUvgTZci4wgfPsf0wDkHGIRAAWI0cYmjnkMwO/ty6Cqxje33dLGIMTxv9jhm4e7bIZ
0HGanmBTuRQx9v/h3azKzcZvxmsoNr4zUUOtKpUsONeP5ySQzlV4jqPU/3xnLBm0aMrtbxDG0rHk
ugED6FondaEwbKOgK2N45jOvvrT9THKNaALacReiDjloYzd2F/B0HEHNc6C9Ok4DQ3xKdmJv5jSR
udq3n3fs+oxAwr7fLckTCydsHrrugQ/932Wlx/De2mM9wbMUuXBjxAQst9FCnL2DlOdDF52KGH25
AA+KMnrHW/0DuEcRKq0AxG38/QO3SG7hozWcNc0xwpIQo8YXPTiYdKDpApOb8zetY/rzJncjGmH8
LonoTv5Xxnr93dWi7UpMmNSEsa/su24del/DCs9LWKMuM4ZMeOz0qnrqkJoe1LH2xEnjZBIYFz+q
th4Ap04LYaAtAhGDANvcmZbkITgOJ/Ac1mjZ0tniA8IM+dDflnencTa2COiNbLvqzLuEcSjk4ULk
Jllq1OWFy83ZOgYEcqmiAo5uhCKe40YB5sovIdkw3yR8SSRu9Gym6DIqburWOJpPMmhTEgnLrOar
7EPVwhlojm/6JfcybzTgz+8f2jIM2w0ECY3t/571JHxyJ+iiaVTnO8a/zo2u2ILFqQeLmSGGPK0a
4zTvEV2u9xs88/raEQDJPPYvBQ2BJNKMtaPD745POFRcDYwCWeWYJCIPQpdyOlAADixPbOFzlKY1
T4AleyAJuZSEKu534HbiG5l3iVoIF1nHpV5e9T9QjmEet8Wq8JnnhhSXsmD1p8JvNKzM5MjaHaIX
aM+uodPxMRCLQ7kCJcdtcEYXOsfY3A+yXLdDf4tMq6qe5WmBv1thxPnCOyCAh5OG30N08VMKLmYt
bebKj8K2hEFlHzzGYJh2sUkRzsve4+kOPdI1YfGkOgBf4MwEI8xYJp49x5qo11BoAALWZ6MorCYj
pYLgE4Z4cDphDHGa1qp1v3k6IvpxuQ8yIPzd+RP4lKr+qT4x+DIPsqurOl9i67K+MBKH0wrlaiIy
E4pvPvaKWOlvq7jeQNL+o6dS6PyAbxurtVRo+HvxpmsJhMtYA1wiKo6PAXuHCRxl1O69H6T/RXSA
R1+2twGemIM5dnqys8+CEzXFFqJQbB7PcG/i0WB/ye1bRrkhS3sQPO/odzdiRPsTCrGy/AKw93AQ
j5HHKWPce9QW8k+tshc4UBKstFiv+tMRMnyjyRPo1Z2zhFDuCV5gVvQUhIWQEIhWlWOC0hFmt+MT
3vsB4Ud+VhmdymLlSMc4iO1EXPQ8QC29P6R52AeTTz0LmxvHAyk72RhrGmDrzXyf/Y3prcdbuseH
ZZW8RzHhziZn039thOeuDncuyWmu4kbdnTn1RuKwzG5MeMoc4oTkc1k62L+JaXB0NklfBvyzpw6J
NRYEi8sQ6f+a+ZLg42EOjLTJ6R9iSifCu1YnV9U51/ExNZOX8TtsnPQDzRHWjGSOaWPrPH3FtYOQ
F8cmrlj3t1R/DCvw8jmY2XEnBwnUpEzG1Ssp4C/YRaJLlcsAbpHSH88u4TimPZHVpGjJsvvNRLAy
VD/AWppYMQZ8cpoTMg+92IEvgFGiHIknA+6hNcXI4CgNbusbiEmoVollTCjxcehFhZGqIb4PC1GO
zE33lDRAKXM86Pb590SFXZmxFVhXFrJnROzjwDz2eiFckHw4r6Zl7Y9tdGAKmZ05GwLRpVor85Bt
cgqXX+pSiFtdhcNGef41tJ3A4JkWosU66wh1co/SbhAaxgo7RMZSwhR/ajUk8b9i1QcDrCoh8XUm
ikUJ18nObvl2aCBYWHGNWkFMqPGubNdIT2Vb2sTHUYpX7jSYn2tuYDjgy7+IhCgHtLw6H0CWcS5x
MKkKNGsPqqEpXK4Hz93XpeWByB4ijGYlS0jPBB1dz70eXixqTljugLnSh12yThJXzsZeYvFJzlru
ovY9p7H3QMO0fDYS7imd8jHW8vco2Z03zajvOB1Cw2YtuK0U/OdoA5CEfpZYOIiUwMBOwHYkujm0
FCPPgRv9AYKBj8qawloSdhsLw0csX/dy04Xe326DSNkRzvgAUQbGUm1LzUf5MF9USytatMPYFy5p
XNp8HrGmh0C2wOW+I8OTxILQKgFOg1YMzJzcSm+oYw7wXLTIesbWc61ipIOzS/U+u9ak1c6qGTEN
hF8NiHflHS6gCa3nQ+Fx9J9RY4n9rtFfrs5k59lcMHofuG5TRQkDEY+9P/cIRbhAkKTwNz7OlRpV
c/4hkdxL0/PNXijR9bmVa5URVDwDVWEVEnCIxlI9mR94Uibs/053h9kWFYfVDNge62ERKMtgGoss
7o592gCpCFfQWKPtbpEvmc+yFbA2zHvZp5APSWL8TBbSDs338UvvTo+JkG5PRYO4i1F7Um+kOAQQ
XYoJzqgmaEQymDCtJpQ/KVHHeutohaWeE7IRICeHoI3JMAoyH0pdNgYjcwLkoEL8huQ+vNuE12cs
HqGLHDBVRLi0uYUIs58hN5b4trSH73NtdC5jcZcChg9jXYOualShqFH0jNYuNm3Zm853UFaWHFXj
VD9/MyAjKy3jNegg76j0Sb3Kotq2dX7m5qSAkdYhh9JdZIiyqiGk/+vxjx1dosZbjxJfVLCzwML7
NsCuzYfnyiNFFbf0vpndd/zy2x0MmZVpYBSyANzuIyeouxTw5LTBnFdUfbxU9yuci1InkK3qfyMg
qXqKVoBZwH5APpQThyH+KDmCiNNRumREqwELa6eLDhTxzmV5vcaxBBviDIiw72JYl0B9kLEkdGFY
9n1gIJcL1d9NFQOSHztukIHhWNiWGdgIZ/QD1T6uUYl5EI4hoRrLraPQXfw8fcKwv399y3ioz/Qg
y43dIJn8vVKOnkWPooKe1RPdpxe2Z3jYWxArZLJlQrRJnR85PvxNWlEl7yjHwLg1JpQAyiGjRqOI
Mi3x+492M+C05sQypKVK/GXaPcbGFlSTIGBsDjO39KKIGMIRXzqdc4Sb2HRaPTHi6fHH2IYj7Vaz
xroMpi56HRIZ7AA5cQ629wc0nkzjq5pBXBJNzROxyo51tc6sfDn3J9qIeH8PPA+ZyU57sNmtYk1n
5Mtz+7D6Jew35U0h//hnnN4qPk7isvnuX9ji2865XKDvlrFDBvRD/lj8VsBJ8Oo10O+GzZZIG5Op
ZqlDzS7QrZComYFbG3Z0NOGKTFVVTGcDU8VOPkjpoKqnE123ZppgUvtnVWkDXghQC7K2+GsB5kmM
qBP4clIc+2xowGnSqKqFdxK+Sl7youdQr/YuJtq+0PDVDLx98ANypJE0F4YxEdNboCJrdfmkHDxo
y1e4qMHQ0g2DdNXTkygfdIBLtU5Q1AwdFN+upIGbxq4vkq3b2d4zYkPXclpcMjytW51gThb4Nv1g
WB45c9xNL+PKl2JUK/skF0U0IqpS9fFpHaO7qjY9/efsn7S+vFkhQRQZv9hoStBbPjgFtnmXWLg7
S6obL1DsuOWAj0PTZrA1I71DcXDALn1Wd0FcGJdjmsyGw6JePtMCVX6lOeYTtczYj2Ziad3xWyUO
aySQSwXdhNWF8vTHambcqdME6k0AzQbKGX4n15ltj4lQQap9GUpDJC9vVy3QnCzTYy02TGV1HETh
tvArXULIEy1A4xZ9Ymmq3pG0BLBluWXyKUBDs5BwH9ACPC9eKrrGSh6huaKOYzPKK9/JC4ML1dDW
Bfn2zwBiGoZadAfA0XRpr6cAmU+/N0puESJAIgsYYhncEpsvcn0OvsWaYtpzm4anTpF+kP/tobwc
JEpaNXMuaGI1L9+Fa+Lwwe3nkUpphSQM4LojT1hGmcoTA+EVGwGADkP4bcFS7s9xg2BH501QyPo0
y/e4D0uSClg7OpRcvX6SvSwomw1pNyqaa4ioxujxsJYHpYsV3+DPlQZNVed2zZnNp6WbHNdBVvkD
OL20hDM/uTfNMSkvfZyfBsJsTFmGLWX0bSnbPjRMKALh2I9cBekHYFAc0BKpoKLbIMZ5roJjAvo8
uAnnCNsj0fNgJqHdl8kk/I6G5Z3B4Y5P4+xOktK8d1dGYpVfczk9ImsgpueC458dnBHe05slLMG8
VsszS6YfF5lmmCNjrrYF4igyRyM23TFShMj0mZh6cdvlF+x0uJdxFskbZJO7FU9vhUgjHnMdqmSk
0EyZ2KZXgQzohoYJX0VV8810GHgBlk9429aku4uSXeRn3VEl/6Q8DuFmJS5PJ8PTCPxZcGW7ccC1
eXFXApZEj8VyAz++eK57Myz13aMplGgEzB0E77ntTl8cCND5Nj1umpok8x41ubFaN8dYu3F4jTTv
1nfGxwITvynqA6dwgQ7Wp/xmQ/DYcj/zQTbgDLzpzXg0M4NMWmrSBVudestySL1ICTa6XtEw/fD3
m7Mk8mkwQ1lhgMrxZgoXbtYDNF9B1RcDSbhaMY5SIeI9LcRL0W7LCqAXh1OKHImX5kwSZWTy5Amh
C6zgk8USi+NHySpC1aC8jqR4v5182mz+/e5B/m4rIl8WgRuINYDiZVDlv3MZoQof/rfQ0GKjfmrK
8hAr9iquIYVKXMkE/s7FPVwLiE3qJWX3320VcpRY9sV3CCg/E+lEsJHVw9Pr3XX95cWY65rpCtEx
K8W3TIJD04+ZQiDYxbC5pER4/SnoeCgP74A/KkZEc/7UgArMuAEHXyhfXygZMrrK9roVkY/pxTEU
UOIjDjyRkzc46b10FCeZ6Cb+l4sN7hU0byWMe84AjRuWEs5JuP5ZbcHmzkjVeYOS6f+G5rVt/K5e
GEwB0V7sn0Lr8TXdZYD5uK13n9R5fjfVrDFrDUHf1rYpIKdiTkQSSoZX9085qrHASmAd0ATofyoo
O3B3iaCAXQzlSr/QeuHHr5NpIC9baiU/Fqs862UZeVlGTPwW2+bewOOwOB5wZ1SJ47zoydEDT7to
Yg0kfv94hTM2EDqnPaiXsHkVAV/4mHwcTcXS/2eN0VPVel5SFuBJLAyLSAUlSto41KX80GspaqPD
Y8JwGFaYu5tDF4lt0oSQ0C4cFvlplvleOUUSzExXCTFB32tV2mJ2NgV8mJLLELmgfIWOKfP79EYe
aN1WIe+tNZVizrSmL6D8OYtTx2ZOfUCqkN14xNLjdayq1DyqLO2cR+3FpJNXSfTMCj7NUZsvV1kF
9E5H8ge2566J++yxi0iG5FSN1BkXPZBKC62Gm4gpnKYwHhWY8wMYTkW4ZHJ4GNnMFTozbXf1T/ZZ
mX7Zbblmrh2nMa4VvKtWfroVXfUvAmeT12PYP7Jye4hVAH2pLoUicrWOoXVoS7+rnogaOkqXBVS7
n3L/pl7vdZASX9b8Dm0lQkA/5G6lGJiIy7v/rbwUrB4vQNk7V/DgRCKaLUxA27IlII6740k44rW6
e1gv+GcUkXLdNGVcgp9+klcko6Xca2MNYeHGnE6p81KNsGvAIv7tJo38I4JIhME/jgIY6Sousywy
GkmPIoAAHUWeEeTHEda+Sa529jZSkkkKq1iMdu8r/HoIppsXGFjocEpyLZDE+0VqgAXVhZr/GutZ
2ZrhYJLqLX4QsixfhqCxENC9ecFik+PYooRhr1CoDOyVvhK9fcdbssl8YnO2vlSZHJOgfxA9vckt
dKB60k+BLGXB9vQciXkngmaoD0IHJLtOdnF1REHzP4grjfvbRI7GNInukI9aqVDhOtvEJVB3IS59
xvkkk0V15Nt1z2WjCGR/o93R63g3aXxT9c+2aWv495+c0iFZJhVYREeqNCXNjtXI9CcSCTB1rOCt
XULsEQcBE6kmb9+74Y7eIcob5ZumlfC3tLmmC1ZpBDKExhif7o9clW6Fto9bgDWAs5RgFtPGcslD
uAui5/mHYEH1g+QcE94ppQY1Dmx52IWer6B9CpYV5Atu+YKXdaacYTrBNot+7/8kJizOmomleu+Y
6DIkJxN90lXDCtUjAxdtSQ+8hhlCAnClpvgMd37ES00v/B3ENDaMiAlfMtkIbj7e/U/qYWiadDUR
/0lmzqikqXrphZPrfq3n8GeiDpyROkXRs6Q7rbPVrfAF3tOPKqAImoPRCMpmXkecI2w++rvGkgUG
5w9ZHZEdnZsZcccpODkybdXiTuiNKEx3LTw8FMYF/qZqdHC4mK0xD2nVNNaQFRebRtrW9VEw1Zzk
eZ4jY97XGWF3J99v4ybu4tkmQWQor5iMyhlHea3z+zLLr5QWLysE5oSEkVfqptsQkf/gQBe3lNUo
J7qeGuI5g2DEtHFycHgPJW3GlANP5teZKnvRk8CC7ZjS0kP69u9925mB8OiJ/TT420lVAv5NtGzt
w8XFmzDyClh/Xrp44oWFAxtuexdiI53C7RbBYAhE2sZUrcAmm7AFrV+YDZxifIoNAOlF6puFMY1t
N9GNV54KjRuICsPoaKZXze9ihrYf21mWxQjkZSxqMIrKjKbynccjJQMTxwV3yjiP9meDSY4BINDq
3XbrRvVXNAzkYsjB11bXTWiDyosJvhLJ8WnaReDj5hggy+VjGZPswR9GtyWhlYNU54nRknw666Fo
WRjqL3oJggzM4gvMHIKP0FBZzO/0bZ1oTQps+sig8K+qMan7NaK5OSRuODILjNee7BkjOK9D+yL/
XdVyim2GqhSRsB1/m4XV3EHS+k0tZIi2NrL/i0kjerux6DTNTAFiwK7/oQCfbK6PgAkmSk9mnnvY
IRsN33VrBQldO3TApddG5IH1RA10uGhMUa3Y8+3vV4fT5PQkpWVeI2gK4OLtnm6eVjdmvllI2HfP
SiB98KpAA/Ybh2elzo/Gzd+Q5iQqVpxiaDeDgCPATw5HCPJvCz/ieDTk9bXyCggKAlKS/FYxpv6l
asET12gK3GQPRv1xdWXyTAV6iOho2l/b/kQxtCrNXTqgwqjXERQ5BxjXX0g4S4bzVY/nxKpAIN1X
hUg+ybzB7dnjCUp25LXxHJdOAac/PwZSP8cdRoUkYZddpHcH2UcpORofEbHCbhP30yMqUhwTxf6X
pJGPDNAJ5dFbmyvYE42Dpqw53cUuMZ8sB8mFW57ZjwlE2b5Os+8SsJsvAx4JqK8/XNrfb4kYkqOW
3w96CNerOHhWPCjUfsoXKBiqDHZySwedRAUQkcQB3StALE/TAqPLxNgUj8GujJPfQ1eat97CFOXZ
01i2wcPCeMpDPvdYLamx3f8lZ1LKEA3Q+5iHbcmqPjDQ3ccuntOwQer+d17Ae8qaTP5YP6xQvNrM
jTCQGR3Tkvjd5E6ibQ2dqhN4zPGCvtXsuglYNQutPZh9p8LvgB7EENeoxbyxRuEIwrMlkCIUGzyb
DEjgIXhxHP6tu8bvM6PJPk5MquoX3/07/w+E+AEYH76pEBndx2zUil895rXTwnABBgAOoUtu0Atd
E0QSUDYYIrmZgpXr5j30JbhfypRDu+LItNx94tXGvIaeNme1a2NesTuClb4MLqmpobEO+VreycdS
gTYGyaH8tqvAg42KOjE36rqvvPGRlkZ6ltw88wZPNSCdkFFPVA3K6CFS6aIFSsHvdqYbShgfeewv
VtSGz86GjvXBNZRk2RRuswYWcYa6rKcUaELKeWL28HqiiFEjE/WOm4mwaiodaVefVBovHP7d2ied
epabOXsqsBYCW0qE5NEXUeahbBFf4aBm3pFNn64N3ylheSHe/xw5si2ORbltgIqFqRzTfmYXwUl/
LVaCawRLvxVD04pYWF2+mivOpEIoOJhB6xwE4LKU2YRB5MHOYp9PwCbUuPBS2jmOUfe71k0ETW7y
lZY2cKarDDiKptbAN5fTBujy0mlgEfINTiHclTs84Dev8ZAjxBi16FZ8CRgn13eEBglmFRHRKnJV
fuxEOQq6WreqKQGcqTDWNivwItm2YHU9nTvTAzy40B0TBtnoGfj5PmkOvQ0BcvCybuXyqAwYgAVH
ZsCeuFtrOnVZy2EzThO4PZEdYT8Jl/JjjhvBfq6l2kzcYjEUbDZFFJPwqSaw5SEAlkI04d1iA1ff
DMFf9TyTyC5sHzOTF45ud/SxN5NFDF149MULqhFbZ+ArTq7mg3dozQbJKutY1LZGdMIPjuuvD+qN
TsFP2q2cETmqTGWm7083l2Ee28m736z4VZTsMmc5ztvZZqexhUT0x/uuycJFK1tHKY7CJu0ZIIff
8wjD03e+AiYSc43nm9v5F2ZnLCgXKL436qSbX+fUdd4yLQ31GuqFM7wvFvoPZu8FSg8Bz9X6LVx7
0bhapZJh6OZONeeMcHdOr+LMST3jHq80n8pOdkzChNeXV0VVVXI5OROZUgo4W/dS5ymvzvaHW2ea
o8fbRcKy/M6p2F33UbhqL4rNJ+HVB5ZmSdilbRD3nEjSzNHSv88Ahqt7nBygz7HT5Vj+CdUhNUtK
8Iv4u8blsa/4GgsstciQ3gC4EE/+0njIWNsQYAFdO2nFbTnT8P7saVVJnkbHR+OjNtIS/Y/N7cMx
m859BfPAFzPvykAOdgA3zV2jFxP5qUfU1KMqr3OOsZkp6phb8+ic+zpnWxcFwcjybykKfRpT7Zoy
s/QyBjBkWSWf+Z8iIp00WRFllwx4nVFq0OujRj9X4Oa/RQor7nBrf1K04soTxZErao8ViBBPtjZ5
Ajrxy7r/d9PKGzvHmbLb588jqvHWk7JQch4bHfECW9F3L4Owk02J74U9RKSFVR32SthIqX5Rlu3X
8dyifBSkEeElpZIeIjfbmmqcUVbb9nyemye/P19AMl/DegAtioponcW5yY8QyfEZogo28/8qy+KL
HVraWQ92hov68Bei/abhi0rIde4t+Qhewhqbp14Pw5ijRGESwXgLZxvhZ91ARphuysefwHItWD5I
9m1QddK7SddPeEX5jdfDUQUH5aO3T4kzR45292HsDON6/bi5UBJFGqLsgwmnJYbe0Jvxn2GR3c4Q
Fwuq2VKfbbek2SJBM+3A9rztUi1FiBHYbDrc4v+B/+jiDYEAU/Id5kua7k3S5GWqNXq4dD/Mbwhd
z/YzY1eUT+R88AuRtN5Pzn1H2kU3jLT5FRAB3HOlQEvV2xlArRNe1bN4NKxDqECYij5fLzk3aQLt
VRhasKXj0WWkWxzHOUPxUP1EyQOFZfKLEDolrp7lTVP39sdQoJFQ9wxzUem5N6j2QFzBOBm2pOyC
8Awm9bbWROpgAHo7xZ/s22d5wYWqXAOcCut83y1f6kL6Ic86wbsWjdBMUR84zgI0/Z41F/1GMz1R
snpgwcbINaj4JOdMcqthzB/k4b20Vfx+jVMnoAC345ArX4zEdNAt0IOmq5i0ud1xzPnwpuYaKXEf
b1X62+dm7cBwQIc54jXS0aj7W5a09N0+mw2VnuPCSZqr741vBdsmxSoUO0w/WNmHDIweP8biUjBT
lWkLy7blkuteQ/ULQN5+QtQDgq/6drZKkJ4SZSVepvoBNFrottDoz4QEY9mDda5+HguU8kX732eg
0lvq/dNm2MUdHgNMvQGJf7CBSiRmtF8P58hTkEIGlDBBPw7JmwfRVzdDix4e5f4j5/5bsmDLB5lN
bxEDGwXD0cd5anOQSfpyu3RYYQDm8IyNb6dgdh+dvpKK0BSxWm5HhAdzedxk7SDbHpkA9byXa16e
U2W6pnKJP9FSEgFdaDJ+Tf7VQP8Jxg1m6xtak9/qO6xjRzsQPk4+TZsXb1JpMEt/c6Cqtxcrshx7
XJuETdiAc6++gd9J9h+3LlPyNjWsg2mCctiMi9KfF/TepVMxzLA8o3ZHRsT64CgMs/pnbc0bX0D0
l1oDD2DkWX2YErSnMzWuIwj74bwnQJYG10NhDsjiplaheXkXLKxvd3ZA9A7DCV2XwIMeUY7tihX/
qS0JQGOECBjKYItuaJ1hb6UNRP1OekVFC/rv0ms9kjbVepH/s4kmFhp5bSy8QnQlp7nUkpAChHUL
68v/XeQKKjS7gUO/iX6DnVMal0tTdbZRJw8DPfoCbXTv2CGN+XhJl7mdfKUYUfx1Wve5K3dOmwVP
QQ392o5A5wmLa8xkGdUx0zlVmYsFgHVqKpLYIxHFyS4HhBgvmuzE14/sZeyNVFqjPcqTaC+DOj0Y
TrNSI2lVH3TGN5BmEsTSzzPtubw2wdfIbI22G9NcZtagNtp7yEoFW9yV6qv/znCzxaDOGeTO46Yo
bIoBPgqCr0Ja55m/ljx4esNnnEi/g4B9OT3E0rJYGjOdKC+gNkvvG1g/A271lk5wSau9aiwan7h7
vVuuNzyWhZKoLusC7REaiPqMGR+/Liun79JQT9pu16ac1UC1H/aiLm5xqAFZ7j8Pg1N6TTxM9iUK
8o0pGuG2blREcUyyIjCl9bKeCO3sxf+BMSNbd0saPMwI72HZXy5dGKs4XCldNb3vAoJQWSKNN9l/
k9NThjyah/78A6hvKCDlOsMH3h1FEmlhPvCkBnaN12V/ERnSOiye2757ntjuEyUBQL+ILXTLRuq+
yPHyG/d3mP6mderU0kemQVGXugMUNi+J8e2+nLmTsGyS3H8z1YRzSOKiJq0kYGgphiwpj1wp4Jb4
aDb9Gil2mJiorOJ/8kKgZyWJkgvmjI9ObmwcG1MaNLgZo5IWBPIrVU/PrOv2eSe4UNKKzi1LYlUR
TlS2qmclTR4rEmeUOyPBl7mvvRSS94l9P1T0v1PJljXyt8gNMSnrHlFHLTduNdpStIQ77JNgd5eZ
gft4VlGSIStMMe+UtDQc2SceiihtinS6Bnefx2xRGBWHvKRoyf/ay7TXyDl+ma8l1mgv9YTVoUYT
KNyb6/q6HqUn4djuMGuFN0T8Ozjh7i5zaG0U5EiMMOklizEDCx3OcT29bvWxNTckU+BFNM7pCdwH
CC1kbZteGC3uQ5qFT9O9ZxiflT/jdOhvgrSCexCndSNRRY/5aUblE15q+fSjJnoyx3g8okSqBKeM
enqOamUyzTPAkoxgi9m0o9MLfLEsnuSvzh+li5oR2nDi6BvIYybFMEDLzXU+K3/4AF1I0cGqEBr9
2RU8WhXRCmS7Fq7IIYw0hiCP6lZwlBxa5IMTKVTxbgJySwpQLDpSphYljZTgaWr7aiNg3Afja+Bj
WA6XgByl0SStsl13rpayyDsWN/saUA7/AP75n+3SajIfWpIisLWz9L98NnCFwlBb/U6gx9xjEJBh
+rV/xBXDD+Kc9UfwozZArKe07S9QKFQXTprrLwr7PNp07nB04PctwzciwyxvKqmJ4khfbq1L0C0v
rulahFBFDBhpyWuONeoRj+QEdwEt7mUJQdZsby6XtmQinB2pPP8PW+TbdwGEwZUX1IA0dBO84/fl
JJu+VyskP0Mo9Y9tqe48hvWe4dkvlJTmIckkJOKPJaZV+BzJbmpr3pucZk51tAZq1NSn8XKuW9il
77oWFWj/grBxAR7S/T89a/eRwhSstgf9ReYIjPkHfJt4cRBiNcfMQXEtjT85BOmPKoklZUKJnA8B
M59oncHtRNeZ+Qp5bw7A3n2vb/tirTSAGPZYbqbrtwv3ae9fPm8WdoRTkXKcnKgb0dZQ5CZS5m+N
EN5qf5/jx1JCi27USZwrvYKWBaRWmh1j8HTq+F3UBVwhb+s5n5ZYWGOi6J/AQ+uWHJ0HSPt/HA9I
HXHJP7RhaSa9r7qpzoRfw4SLxR+ZS932JtQL1ZA2Qxnqgi0gzirJYD4gGRPLrAZfG9gRTiucbpkY
9NHLCBT/n8FcwPi5XhSy7HwfPNRog2KIa8nz3Rk6HnKsufsrHFibyzFnyeNXj9ddq4MpPxrKlxOW
Kk5FKi6aLF/8UdaOdbzeGd/E9ZrIq4A2xSmWXCSnnzxTRTYS6Acp3SsCXJqP9Q7ky7ZZI3r8ASiD
9aEUnIMTIiFmt3AS2rIh+0U108qlqf9ijNCDkb+8++Wvo3Y/RXTIawarAXU1tl7kI4NAiPZtzMN9
KecMkItC5dwF2etw/j3JLVT+ZX2HFd5pr7MemCEo3ANM2xVX25baJFv5aLRR3yZiEp8Wyr3KZ03h
VEaDQ4uKHauF5ggnoEB2LUADu359w/eXokYlnSrPdKEkripm317sfa1klnE7lvx0NUhaTitBeaf7
b00D5gfmk2DAFL72zMaV2B9pNAAlf35f2Pdicn8L6bVrjW2gltAGtwTR8BAVHmlCoVMTGg1eUKEX
jQvYmFQUHs+fdAXPjByQOyFqk4+LDgVL2uRYwMFrqhO0JSnA1t6/mzkd43ckg/Y0jqfGn0HRbMJM
HzeD603K0ttPBgqipTfNw4NpAmghNseiMHHAGJhwO6lfR7P3Ko7YT7vp2KxErGpVXYSlmvl1tHb6
m23ZPvTn5+RigJNVAfg7LhIzkGg95JU0pQ3x2wnX3cQshBCWD8sZtDEao0z9As1cZnt/80e33G7J
ulCH1agqyy6OaHwon+ejx3Z8X0HFY04ss6pnT1oBVGhsjUDEwHxJpI+M8yaV9OOr+KLU7TTD3Ukr
y9j8qGtM4I9uVpMRubfv0fOEqI0HBq+VZqWCwZ/YflE7Cyvkl/UZTAF3bOWSKGUHLM3YDlxiP23t
4Kp9xKbo6DV8zXYSQsyLwEXCoMceP+wRcXQnFJ+VMJTu8pGS/ZEjACaUZABcNKZH2cwiKcVXux5a
u7KoTXamw82ZXLDzGTwsXJGknPPBcOE3iObGmnftpBvBVCY8uY4titVu8WSI+eiVJE5wO/cHRlZL
LfwZ2v47lSjTHHB8/FC17YMQNQedpz6w7x//9GzIsGPYcMuQe3LZuW9VBhBN/q6LTjoot5gP49iK
H3T8k9fmqYhJNMCdAjfPH3W/MA+yCssDCvafOfKE26J1kgcMDPaOGXORApNe6swUs5YEpFw/UCDf
FADG9Secl2zYGEkvKumhqLQel4w0aZwKEtujYXxr98/jov6WRZmpporepycjehIi/yyiyN8zDahi
gJjiFU+uPZeBhZi8IcpkfTmfXOU3VwCYWxNZN2M9zt58e1+eBvcs39ZcG7sKu/jqVDFeqBmWdlGF
hNKUYpQ0AYM5FYiPc/9blg42Y54/bqNblWrJbZ0ybNYY1ls+U+fo6Z17UXljkqeyoCny/IT1Eoan
i7Ky5TQuOtBfRSNc6nN7LHagB5X7CZu1Gjj5TYb6UrL/ZP0m4DLz8r7wYOduimS+9yKcocULguPb
XeWqD+BeDn0ykpUTrpVkpYP4RWmX/gWKRLEzb3mbzTTnj/yf9aISNY8evLgZo+FvW+QXC1x4rQI7
OK4ldmG2eOeeF8/3dHVpEkSArjo90it9Ro5xZtjgZ05vS5T/9x2az8TxbIIo8QHXhWxvDB7llSF7
ZgKHe8JXBhgbKNtvrt80v560ACvjUHKD+4EZTAKw8r6ee8A5aAHhjRQYygDfQL0O+SRO0jwpe960
c3Jb6FpkI4aIJqYNl4E3kITQ6onos4UfCuErr9C+uFcFHfG5RaiBXXiOzjZKlUjn8JE2mTFjeLbO
f74mAw0Grtwi+VsZVhIe77MoMgH6GxQm9Qp9rBOgESl+hr2PdroN+uBct5A9kB1iFoJZdbzBr66y
izN7TTcL5aEzI1ChYfmB4Oq0fzghwl6aHMEfTTyLGgoijVo8BzgKaReMTbjbyY72bdU88PyXZOcy
Uc/Dh9nzL4yun0CraggXH0JL6nYnx1sSIOG3HkCEnRpEKp4K1tmK+1gDLyO/YHNRsYmlbs1jyxCt
mjRazsN9FLc+JG3nby+JbDxrnyvysVDjOBERZeLf0XC63QQAOOFE55Pjt7VmVBH2VR0yz9Ql6cvn
Gohj5vjDjjJWZhNE9ARvNLbOrMQVvlwqkGwHO+3EonYIjBYHF8X/ktkgZSYyIhb8YpFE0UQSzvrJ
yHtyP3tvTjkkOvTkjXMOeMjKoZb9V5zkAXixThNCyGHefJh6NDm8pErJ+RJVeVP+9/yR21UsxgVu
qtDOSpldOR4Am+91LC0h7ZOsrtbUH7Ao5gyoPZ8Jw/Hj24gHQxFkrDnqY46v7OWSm7c4f1Feq1pr
BMA+Qbuhn3zw/Y/Jejr2TSgdnpAyRd83q4VCvbRT07lCuOV7pI4h8lLXyDtYBQHMPgGUh2lsiuxb
K33VUwJqTOtmoPkChOS6B8Ya6CW1ieTTLCsGiOZBMV+MiLm2SCfL6iTyshKwRckDMqv3PlHr1KPI
NNcgOboe13hQQ3gNVMfBdNdaQt++8IqLjKHUwx4bOBsJ1wtUUlIP0dxdaIa4eUmD6DSpOG3rWqvu
Q6T56fsWV9llaz2Z/5FEOiB0Axf8LL+M0FemnYLJ5nhqWlp4nDI3R8Sskx114430Xcyk3ta0e8Dt
LSreUp45k1x4Xem3NRlFyT+qGR/ZhTnyBA2KTKau3KucXcxuIP+STHA83tpRImz/yLXZROKcTuih
I7P8NKqcoYDvXhrcKhGKtShm9YnfIBJZcRnAHg8gPcJbc2kPNcycNF1miinA/aY+UkeMBoEl2xzR
+YTdUMV/kelJKBRUG3vs4VrHE3Kt4nmvHRU7QlP2/NcFBMyetSH2hQ+UaRRD3U3GVTOgpXR1vx5M
AsCEcA+mO7lIllwRM57ZYoDY3158sObmF4cRdrc0jYit2T884gXwcCe1df1EGLAzs3VQO8Bq0iQR
AMkjkt/3upG+c0PDE73qlBhoHtRD+sMVshuwPT7TeqvjQpBkiILNVd2RNmwu2PeaXT8emQPmMrHI
WjXO11w5svMO90hJvekPKz9hS4sXzTkJtZeD+ErmEG6Ogb4s7w5AgY4k+c1LrnxwC1fK20i7nLiU
W8Bj1S7/ZJedH2f7RGYsme5tTFN1OOgOdKM/DFhCvsZHMjR+vJaGM3xCftm2wmr6foFnGQexBOYe
tfrc0HZ8m3tQvmWnzSqkWI0EsHcDskBgYuvM334YPOKOEndNyJH5UbKDYN23OwtUnnq2yIH9NEv+
h7lhKQJ+PkzXHGxmyAS+fh8c+eb9alN6GCqzclqOrwfvwqv9+1jmX4tQChfiS5nv12cBtF8H751f
xGTXH+tcCHXKU8KxxUgR+sH35sRXuWzcn9GShDpMZqCK7YoM1zxG4lkSlFPcL+SdK5zwtcSckbKW
kU1h4gCQMZ4dkRdd/50RK6p5Na/E30aEuYFaqUnQNBFXdrXoIPVcsiYtVx+7p9JuIhf0f+cH6TOq
dLbqbZWTuJoDKDDZaB1+gxG0r1T9zZNHSIn8O4z/8zK5o6Wq54YqH0sRyRE4whwZp3wUjYWSS134
+OALpDjKyIq/T3bzpTeRAoJVdYey169TISKh35CtJbMK0pIGMb3+CJcBRqUIFyDYFvMJeQzb6+eJ
9N572/R13cEQphN7mqXED5DR7Z0EETVoB1hVc1+/31ZVNBz/G+UGV6Nk4n58JvkKaR82aJ0iyXfL
OQ0hvYih+VEw/jFaweEmMZfWQ6n24MeOz/Wlirn4XYc42CzQRBH+1993feTymO09YqSaSvqHJwhC
kUwoOQYJ3Tkp0s6aCLwmjaz6Ge4WovBOvznBmrEvtN7sFoIu6N6pO1Rz2q7tuKNOex0rfgVi3Swp
0PXyimEPh/esxr2H2mQEqtZbVrBagAYXQ+MDKzhRFU0sDxxCNBzlF/VRaKYNxrmI4K4ab5u2ka6I
nof66e3mOQH/EYyu8hY+q37J6iETAEinVCTSzky2zf6D66DFdKS+AH4TNa2ivF+rYdakWnn5CbDe
SEjsMMRaEi5QK7pzuLEl8ACd2UtnHDVEJTwnnnH/6QHtf2KGg7p2dFeeaIbIBxI/hru6Nz2q+KS1
ll1yb8pb0nd6U9doclHJ+a42xvf91gjh3HeVCP1xMwdOMAz1MgjZUYK8aIaCU8/LFMtrwc0jip6Q
cuOuK10qn7C7zOTHInsYC3hIYVSoPVcb9DRS59tOH475cWEbxCOnHLvIP1Qsu1PsYkyH5jBniBcO
ODM49+f6chUZuGma3mMmF+/9PHEEnS+0jgIs5XKa2c4jJaCjctmCnqgyKN1WZawGSauB6feLh2Wn
UKdBu13hVRZSvcLSf7QY5y4V08SXAGl9xlsoxMu/Gl0NLcuD9+j24fxZJXEbzK4jbSTptYPtZwEG
PWkkENOOeRMyHJX6fY1aaK2Idnj3Q8Okij2D9LEqyP9VAw5KZURYwbUpf2vK7xXZnSE6EQQ+b8JH
rVhs1uJ+d+mhMlARXa6ra8dlmNTSvwyvyyjToRkq13+OZJVaFn62xOIgR585XsWqNmnIgmoxTQpQ
HcrVNOE7AWra9l+t8EIsBCy6I8L5cqnuhVggd37t15zn986Vok209fc01XQp8CcGSUR8zT+Wp1ID
rfNWEbpMT+SC+0KqyJmWhaoJH5VY0S//SI3BZRB/cTzKa1Qy8gHAgT7MFKg/Iuf+nz6vDkhD2uI5
pjw2Akaughysc9YSxIT0+NPlZUm9E9y1+hxjhVOytEhC+rfORVhoHWJNSc/ajNgdWyWxMgDVqdkb
QzZJg0kxWl9NNHLsYuukt6u/ElwXRlfsmaIIFB8URoPlqUQp4evmMamtcPw2w5aHI6f5Uef74vYO
fwQs4nDMQeHYYD+ZNVwjp7whvE0e5k5R2hlEGovPBhE7DCg6NGR8Y+iaJoL5srlxjzo7vMy9zYo6
gvO5jac07pi1P9WRFzxmWUbpDnqRH6pWCWSHl1MSYMxjn8xs7V0xZQq6JKOiHrg689U44wJML2sS
ahiOPqYgUwPg5cMlOImIhJ/ex+Jlpc3c4d8vF15cRHK7LFYJVImJJomldwf7/SI5qQNEfqElmCbS
OfI7XGUHaGs1EItTmFeuXckEeR9+ytil7z6JjPInRKjMcOa4Hox0NvjkBjdhgKKwx6VtTSDf2MAg
6XWH6fC49mwzWTk0rejQxHN2HYFRiVM9j/uanD+V+yeiZ4lmCD+mPlzPtR0NYTOsaCq5+ADzEVuh
ULNBLKh971jwHAQH0MOk6zVfke756lXuZ+uKQ0DJiRE7JQ7FCaC9/IdEwFhV3r+eA6STgJOcD9gu
pipHDbPqpmeP+pX8z7xBtWiL9R8s1kclYYPPcoyb8U8fDO1i861ObiugxU26UfJ6K36Tsh6UPbB2
dWydxdW/678UBFnp6Utl1tqdu7ffJvU0tp/1Z/onQnXJUpzdfYfQ33gVhFm1lM4nZrYMDrq7TMz/
S2wB6iah11yBNrjzv9FRH5XE6rL51sSSpbRHsQHkj8klmifihGEX4dUpcblQ4MvjnNzpBc4QzI+s
EtL3VuWK+biM9lrz9gUgsOYD6YlIRuqqJ2/+B5OZGIJLGq5Nq1nCIFR/WRP19Z57qspuMBm+WMUE
ZU9QlzedWAQl3iHR944R5O4XZxxUZBG3qKr9yTd5hM5johVpfSJJjF9jv1fCS3C2C7tLBx8qxpcx
H4IOBMWPYULkDIsC2Q63natn9Ddqb9VNEGBECHj5jSgvAkd6Qq+qrk4URUMX9uK2yr354Wvtv3HL
19rDzZP93jqgvRZC7Fkvad74fQsvJ2cztYrEW8OxX6t/7Yaz/zJfH/DJqEzj7Qce3t6i9WiR8u09
9bvpTLPUdCvOdx3m/XKtq/3gnfsk6om+L7CB20QnZ8d1ydeRtkJr0k8aKF6RFjZZdXI2zNSGjFAv
OIX1lACTcEkCqs8mnftcctiJXKN4jgwP9D05BwEJC0TYa4t448zC0Oc6AiRepOYhuD/Vc2PpTQzB
r+b/Z6LsbntqhbDGIWrVCydLGe4tliSEkVcVz8SsS3vkLeZAu7cuOKJXjPMolSFhThhN0mtWwqgN
90tf0NmL4LcMrQpI729zZbPfg/5Mzresviy+LEIghjgvTn9J7fP9KJYg8rT+sw991prajfyE7Hqz
00fHa8Od2r0BoZ+ZHfeV8dKgvZw0vYDwND9pg11kK6U9hfn+wTJCedKtmOIwIvoICksmiqC0MLuO
G90C+PmdsGzhRT+F+5uqONaiHnK7FMF71xincYejXS5mlgT4kfDlRmIshet04rHlqeqLencBxovt
bHuDGypfF0K7Yzl4G3TjA3gFb2sGWi0gYPHGY8lbX+oYiif6luAPU5LyLN1XdWZLDs6q9tFqkaty
5Jb52pINuSt8QqIGoxn+FTVdmQYX87r0oQbxxcIa/MVFBEraJMhzKtfkKUjYmUVKze6JF26Gujb9
OEWi2bQ0Q06Kv1+XnzM/dauiVoCB2kIAjJd2IfuDztKWSZQqEp8wUsVXJ/hcDIkNeCHasxqiQF2f
/8F8wqFj/4mFdkXAp+daONkSV0a+qF7g83PTgc6fhL/SeJXJOKXpjQDzjaOt7ujOLqHx6+DzYY/d
V2GL7vCzymWZCCZd2hP0hNX5SZPbyQ/lHVB9jKx2f8s32XTfsVv3DcQwq3lC653mbh7AJUZTWD5m
yTopJmgJ8d5mbNqDuDA5ZBiL5imt+UONl1w/SfVOj1IqPQvD3utC513AkCAFigjHho2dgLsnj9M4
BOrXemJGRWastiPsqU/x70rfp6N0sKxRzlH1D9syQCKbU+65FNlxEqic0emXPGBeKHtPcE7t9EY+
srevO8zUZ8vQQ/BFANuweDzrQGqxGMTfGn4cSc1/YjVwN4CLLsBY2LBJY93mRRsgGuqsmjJNvUTQ
tnSIkvyC7E1WRaiInWzUQEfTAgu4KgMGutlIVl3Nr5Bld+/ZHeMfJQEvn1aYNVC52JXqhTyVGkXe
lOcU6ccQYrRzf0N2NcdB1Rk6unxvKJm23OlwV5xuB1sbqQ/0lUzBqp4ZqSuww7z//m/IunZWXDIW
QjFecscas+OZtgmzUtT5cMp81iQU600kr2QMZKJA7kwAOFajFBYdXmVOtMM7uYwv7DsjOr/qbnuU
A+afPGed9B2EOqwCS2MeZ+zm/7KN0oo/mXNKPrWcI/JRSGiBG5SecoCW7oEscGcSUFe7C04mfym7
KTNcYb4Tm817kzGhN3/jTKzORj4OdAI12M5KgCMNrLery+EWXxwcyfHJJbzy/b0Mwhc5gmCvV2tf
8ojN6GFtTZkBA30jFvZrZQ0pdjkuhG93tZL3bJqKMMzeuHRpokM/AXBvrEUg1BfWSL2F96FABELt
PPQgxuN2mQSrL3aVvi7/KdY3whkJmT0UoMP1zcgCj1FEhe+IfeWikz2AHCrDLQ0qpbcpLCL3MDe4
xlHvvCvjAQsJRfGAc8JYBCnV6sPKyC0kQkXjGAEC7Iqbu1oGC0LaouS485qibxhFQpI7hFIRdJG2
CtogEk+1gYrUnGDaBcreQIU/8/CPGYTjybKmNTiQFDkEBOUDc01pr72LUedjdsyVblM3+LF8A1WH
J/o15fctGg0LqhH1lpMZhNlQd3r95wPvPvtn4z0TUra25gOfvyHP6TH2JX0O1CCENx47/guW+a74
s+dwF8VhrCLTNLioYxK3H/GNKle2y8NqStpRGgfZ0Y6pR26aEf0ly3GFOwt9AS23QDam/RihxVcb
gS5hYFtGwv9yWcrb+682fk5odt1dA49BKtB/s81h8h369pYVJxaUBv+DLn+DOb2jV1dkt5It4Lj1
6U7ZE1cqXJCbZBW9b+3U+uAgEpU4ERFxWuQRc138CJnsS/AfS36yYutrXh7X7Gp1yt9K1vMIBDM0
GgScGsnJEWgEEeDVjuKWRGUpwB8wUtJflnEtYwcpEvDd2dj1xS42haCCL6AOUYk61MPGp/0BkZCH
suETAiAwNHTajzpnanz6AomrExImRu6eHbQbvRzdnnmZEVpxBEIdvljEHcB7KzzAH8TzRCAsvl4k
Ug8clFrTxYsKJuN0rxEn9M+MDJCaj9M2HpVZFQPT4MRtHfa4myBIzkWbNtvwaU+X5sbMnjYGPn3s
cxfdhuTbKwcX2dWQgeBBOgw/rrNSDH4FqPLXyUflZxGf8W4M9r/8XoDMIf9jsFColmPNYoPOmjfO
MyTdJ0nMEd4Aq9U+0CTJOjWLW53LrlzV9OvEqbiXxhsvS3CNP9p1ncsk4hPOSWHKq4E+Ss76zETO
6/Ql0QhofQUIyHOhAxKdNvrynPqM/nIRxN0A9AsHCHjJ+ti//1hAVIDN1TWMedM4rzZxIW7U1O42
egoNh/OlijNdma/XfirCcoynHtrSZLI5faW4UL8YNTdrEaMc0gJSYmx05ACyqWJlzGt2N6UkUlq+
x2jrIQvCOjWi5IuffLm2TBEvK0UFvMTXaAGPZtJUhoMVt3aQl5fY158XiQ4TRmpMtnBSs/ucVVTo
9ssvlRz5KxtG02BFHEet/3KASQ1qTMEQVkBbU7opyTRgPU7G4IPkG6B5ZOSaIVW0KzF23jyAki9s
SKXtB5Esmfwi4PaOOiDXKSbPx9mEzQktWEYTi3rj2h1aXN80ZedV3VI7z++ms0JNuJYf2rQUv/HQ
Xquj4fkGd20rF27RHGvtzHnMQTsUTUD8pI+tRjJYhj3yxTQV5IK5maFR7EOUqcbgINJ1XWEbNwkY
pFr/xzSn9KGo0r9pf2ATuEpRboNg67CJFU5t2FBK4sqn7Us9tMvyGbjmJkmyIYPyGd2n5xVNKx8X
t4T2D1LyDp6u8BXDOJ0gcvhX/+IU7f2MEETKu19+wblmhncCR/nZqsg/67AHZLncl7fTQwXDRD6T
+R55gT5C7f5NtyThIUKX5SkHvnr81nqACvWzMhuk2Y+RzuOd+8Sggpaii37EEPLvgVst/n+01Y1z
UwBOQOdi48qC5sjhXgRtjraozSxzD+HgPFbVniro53ovnyE9iWo9MpjhLIVFnUdMKcTBre59oUez
hvQfGt9iTl0ECvF5pfjQojz8amBLODos5eewVSr9u2RLih8fcWJaCuEerbp9N0uUqo6Xpi46vnOv
TASMrKbJNVvD9IzkkOocNNJhZpSJxS4cCli0tv1EG2USM48aYf6kiy3yGjhd5134el84ddASIAYe
sDOZ+4lszNmTmEtLNMvPro29q/9OazZf+3BOuGKis9hOneIw2pe3dE/w8YolrDLsvGmcBcJ/wIRf
3E+jzVNS9l5JJmvc88fn+eJiRt9LdwI7SEd/CIMj3tz2D3rELahIiIzyCXHTga9/UJmxhgaNFc7s
OSjUt6CUZpc1bvM5P9WDkuZIaz8lCBVxWnQADsWYyO7iN0xOVzn919wLPhKOTRXMD10yrRdGbKp1
a70KTo7ee1AViTllGqV3WmxdiGAUtYY/E+9C3HW2au3u3hwxwVhFxCS4oC8Gg4y9W4gwbVUVUyHk
b8Sye/hSUJSFgfcYueteRoVecq8T5Wv+91FjrvRdmOYYlXxWutCX5+jx6GzdTCPeJ0FrJOY8Mew0
bPWHDrlMPh602PTQ50B72V0/9aKSbb8nQQX41JDcNCffPltNFy8zMeqEX9GG1S7qTygPXdQ5XwVf
2tSXK9g4lMQx5ISLtboNyRIb0lXUYUVDvllGoiEztFfdu2DQthSYC+3iNn7XUJbMlCrcZVwfkY89
CDuQEj9DHu9Sq1JC0hlnWoN6ygDqOxf+YhqE065XfBd3pF/UDsPsxsz2a5hG5d8NAf31iWEZ9+F2
EGfkBEAqDR8byP2oyxJTnXqRgpChKXbLbsLhyzUwTbwoXKq3NTFZhkQDGTcq2P3HxQevNbaFwZLY
TV3GU4jDezBd7BkwQwCserj/WjwcZRtvyowrQZk27MorRRF6GIhaEhxnBAtkLxkp/isKEq50mva/
U7L51d+FF7uZUO2F1GkkCF3pwvnq3UOeiWe3L25K1D/97d07MrAiscoO9Jt9G26bC9U9bwnGnnNf
Z2P1cDX3hzd2hHYiXO1e0GamJUeDrpkPQ5bp5gEUDIBCtgD819Y5uqlJu2DA3CrW+J8w9BFlMqsm
ZTC5jWa/Uk4mqrXo+KkSedDh7NYr7ExCig2KTdmrpyhkXJXB3YD44DhCnE9INseZ87WCcmA4QuVu
YszggQBD5inGuR175Urk7oei2cOAr4Z7+gROTlNRt6hPKauY3lqEs3eWWFWzRQAQatPw4wjaT2nG
PmObTiqyLmLuLkQR6D7UcK9CFmDjQ4RlaqYTprwco6YVfb/scg1xvYf2ay+yblm1WWAPGzfHAcSX
fMuAD9aXSF8hFwBKGvlfO6/EkM8QF0eOoEwXZgK4g7Gxs43KaL5OF5yJPspoExtlb5TZ4+TxuK1a
FaBAvIBspsHfZYG5Wz1HEfxDNU33v9sLjJDZS+XvjHO+de6S/j49LRUcR/7zaADbDwZDA0fUCwIx
74+Bq1ej92IL/QZkcEP/JxGksMyi0Q7z8GFvWuLzvlqa9dIZMdghnhzjTzeo1ohW43iYcR0eM8xJ
UoNnifTY10nVtFW/rFEOYdA338IUrM9KDPvw3/+Nw7W1t60oX0KVUNaKz0Y2li37oG8xAZi1fwJl
vl1IDq8wTFWwbo4AndZZhGF2RigTApR8/g6auQAXq95EayG3/vZYI/i2VNEwMRQRJng04VUfCK6S
NYAQ1AgSHLMGF6GRiu5sIGP2vwy/HFuv/nTHW0XNstq1UIM1a5LkzSc7elNl/dHl1evtHBkRfVdk
vn1pJNVovHw6MGG/1uad/i4ekeb5p1465lWUfFMb4l88VaBbjzz0XeGD8FHGHbn097qE+cumamse
BwJPoC9lpxOOzw0cNLHAkcw1rIz4pjr7gZvuZ+lFrchmKlmvTDpuYdnb2c5Bt89XBLoNgXT7ro4p
Me8tm35P7tQQxtUW96vmMYnV0eNHsmcsqA01gkOa48p4I1IUxxhRozKtguBIQuJMu7M2iMAqQued
AEpkjvTRF5o881CUx8jNyyCxL7TAScjKr1Shzj8feckbc6SwLvBzDMMd1qtwGUagzCO3ym0EGKeH
xMiQ2NSQQlZ6uS/kfIrP17WQ/r3U3VoBUiwYzfg+xMd/vkLu8SayqjVECn4SfoaHctxBR50+IlhA
XCLoNgRcn7Wa+SDryaP+TaEsHxPwc6jWLaX9SBW87bMU7CabSsQ3nYrJsEbtAjXFoq9G1jPINkJf
prdUJf2uovI2DCiRfziEXiR5rBrPeK0tzIPTt1Nesi59Ms/I7nS48cRGFl7CqQdQsUggveql5PyJ
BtC7Ag8E3eI4luGD8JJxY6f7g65Sm9Z5kM9Xy/pxF17JyIZO09VL67F3jmi4VUh1fd0O09EnNcp9
WD00SlnxU7Wcb56Wj7moZXGDja4V4u7WWbwYsR+R120/PTk3nxUeXIpOJkeCQyu4b2oI5xV1E9HW
azcHt7zwVnVuCaSVtLpzJ2hg84wEDIqeM46TcdmFZdMbzwyhNc5D2Ey2IZowyF0meSlvB4kekpOI
s4yENgKkqkZpfCzfNVUU4rCL4Jru6ezoij4is44TCrnaZSp+C/epwXQUPPJLVSLeQDEmFebNqlr9
7uqF7fc2tghLLU59FER1NxRGm/QhacdOkx5bu+akBTxt1otM/6sfK8u+lzdDRvKVasp0LyW/hjQC
AUHE+3i4TIO8yFUPUwIEwQlhuhaKu95cm7qxGoWSJjBKyrcHrf9eJ4wK42gK/hTovT3S0cGMJL51
0A//0ModDKq/xT2tNQjrvylCfZg9LkY3jjFmVmWlNbQds+5ZvGTGL7lCwuGjjCEoUMRbnqpmWK55
xipWjTwfQGsvOcXX+WvYzJ2ke4ABxND+MlHQizkkrKS417N9AX9avgHncVLUAxZZdvYxG4CxYHl4
aON0zaHkaH+HhLysRCNlJw2Dv/19aSW/21OiuJeOWurMvp2l8bEJIaH/7fbmK1YwvdYwVPJIECFh
A1ZaMBalxMBGSlnFwY66yA0QWM3tO5wHrr0w3fSeNjKRtbobwTrgq/9dUvLhb/QEwIXcXd0wb3wj
1f1JGC24MET0g+qoeG0sannRDXQUVR9dmzFpZxYmuypNMtK6nic9qZkNd7d1x/Br5w8KlrPVZ4IY
TDwvvUPxFrzbykVpRMQD8mU9V77jAG+ZrZ8p8rWSYsfgSSQTBk/bWIjPE3LT+HkK1/S/JDw8o+qz
u72o/D+C/Xd7uj4MBQiJKy8cWyofabhXDVZVcK+TyCV/MI8URONkb4TpXjUFPxuZMh8+7KzKa0nE
mWynTEs7+yZxDN++OusAEqPJKnkBICe8mAT6zxydtEdNonUG74a2gob4P2z452gs5jvCRR+HHWqd
vi16kEGnaQmNvJsNhaGdwbekufHVlXl9leeaDMBqEhXS99RQ1CjT+elUWZNQQ2FFYp4Em+kSi8z1
XDc/RcoeRhGf48a1ETenZpOlaVE6CK/YiRxHYhkgWFficmEo6W0QQgAKRuwjBNh6+ktADOarm9uR
nFJ/MyfBAEO35ObpCzmX+3e8gKbb767313pMJolwJPR05XTW+iJ2h6ExaGzUQOeteZ35U17D/w14
gaaD74c8tcNZl0V72J9pLMcOC8qJc28mDB+mMvzlJsTU9NbIVSffqR5kpDBktiFHYqSvk3WipFV9
EAcVUMlTfXjpocssRSLPW6mFQdYLc0hGCOBAqkyqjGskYizbmcBMVQ3f4F8N2Sat2/xhVdhobZN9
MJXPc5x7k+dR8yDQAlJg91a0WrgBnqFd+pk/k6muFwtARCT8GV/wxocg55RwAnQkCT2BdNofI75l
f8vQkmoQ/BQgfM5vdegGWYbmLV1+LKUrDmt7dKV38aeqPkZsl8K/E+x9t8Pkd+v4d6abLDMM6eyr
R0Ihw3A6I4+NcxO9tEtlatEBeLOjTOr6d27OQo2ntraykmLsQjpG5HsBwWFmxzzQRNs6UwsBvq4k
sdIXUXoF5SuUyQfjY1iN8c54kif3o7H3Xb0ETM1RBHbmKVn9dg==
`protect end_protected
