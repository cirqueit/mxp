XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;�����EG(d�d�8��,��1Bv3X O,E�G.���&4�Ҋi��B���խ
�F��$�?;��_���b���t�%���j{̜˰� �RmX��q�J��~��&�E�Ƙ�5�L�-X�K�Z���6��x:x�^�-*���x�"B"�.��]�}z*�\<��,���� �+>���mp��Đ���bH7�A{�C����Ta6�)�!x�3��g�����$/��'��m�Wɠ�1bT��r���r�	K�'����	ޅl��H�O�KB��f�����!����ӆl��;�|oa���ڲ]y��Ǽ'�l��	�������N+9)��ox6ضn�1,
SBMI������3{o.o�����+��\qB	������&���vܢ�P���#�������iϪUv �{}�4oB�Q{C�N��Ϣ��/�cR�V\�Y�����~��^�{��>�U�W�g&Y�4�f�@GG�ȁ��㫃H���ٮ���&�F�n��Ě�S�=U�B�&p��E���+�S��7�ц��W������6/>bv��(
����N�U���dY�c��9������"�'/MkL�A#!�"?PWDw<�|5�4�䇘*
L� y�'��1��嵪�vQ�X��YlyI��d�r�YN)����MuL4�F|��x!+Ԟչ0�!�� y�IX��U{��H͡j���Q_���Z��6���FH!���E�m�֮�*z�hXlxVHYEB     400     190<�j�\�����V�K�:fA��b���֧8S������Т~	#d=� "za�e��<�>�8{�W��ȴ�L�F�j]\Ћ����9vVA�����.'��H�F�1(������Sr����D��z���/y|��3�.:ԭ��}\O��7LH&��̊T���[�F���)���K��ꈋ���5ǗK���0v�R�7��7�r��5���?�#�2�Н61w5�d��K��lŦ]F�M�����Yǃ� �;�ۮDAWD��q-Ӹ�5V?���V�ύ�kj���^�q����Tq��BS�%|�{蹎$��������VY]P�nVj�����6nU��}n��OF ���R{M�L��c��)�<jFh��w.������=HRg��VCߐ3�$Va]�XlxVHYEB     400     1a0
G���gu��_�M 2����93���wܴ�$���ӵ��WV
����_�`C�s�FmI�vO�qL_�9|?O�:�+�g�`�m��J��}Fg ��{K(�a)�<6qa�5��0�>]�?�-�ڼa�)K�3l]:����V��IO"�ubo��o�&�<p4�9�8Z�e��44?��B�%�|��4�c|i8Bx3;��,	&�#�
9������M�s��*)��Z�"$ ��S\w�����z#;��q�]�M(��*�Z��}q�HK�\�,�w�3)�?���dz�hS!.lq�jz]��p�LWaqM�6�M(xBk�Vg���K�	�㓑���w(}>�!��<��1¶�	D���/�Y��r�/^Yy����x[�%���认߬j��|ĤXlxVHYEB     400     130,26~H���a?���5	�I��I�/?9#Z0���q�}#o�/���I�<z`�U���S_y��{��jW>��.��x��R�=Lyo��ۜe���˅���=�Ȼ.JZm��4��C6W?�'(�Y��US��nk=t� |������I�k*d�>�ʚ����d�gᓃ�܉�c��1�.s����=��#���(
*	�{� �-�Z; ?����SU��֌��Hpm1��	`��U��2C]#`0���������i5ϼ�n���E��ɔLNђ�'*�>��]]�`�J`����XlxVHYEB     400     160��h�l4�xR��)�jp/���P��f��uP�RUJ-�,���~���}B{��rn׼5b�� >zG2AR0 ��a�������o�]*����،��c2�/�|^p�Ƚ�֫�\���]]ܤy�	�m^Pԡ�9�9��/�5g�����h΀`W��?��K��l\^]��MC����I��̢�Adˡ�+��n��0��z�2=X��8"������Y���U�9��&)�3�{M�F�k��Nr��^��R��0��-�~ 5�\ڷ��wk�Y��nS_�������]��|w>�(]Q֊'CLs]��N���O���<W9ZyE$)�h�и��]�k'���w�|�7���XlxVHYEB      3a      40(!��4�kz/#4�Im��0��%�L��f�FQ�8}���"W���N(l��=6����ݮ_t6��