XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��kQs�߳����F����B�5k�U��v]�tii*�+v��I&̅E����P��/��&�P�ؑ,� ���������m��ڡ
��H֖j�.�%�)O�.���?4=�v�m�7�*���1�5i!�+^�2hkN04�R7����n�;�'�lX�!����pvbD��Q8S���h0 m�xZ�������:4�o<�H�31��q���#����w[�]�@/ay@g0F��Iv��gFQG�6���ДxkJ��V��|�(ʇ��%�h@AI<����y��I�r>婤^���lY�p�􅶒
b��c�
�V`	�]k9ӑ!I�ڔ�;ւ����̂N�ɧ���L��N�Ĝ�Yh�Wu���,�^v;�����:u�Ԁ&�0@���Js2N�[.�)�nPt� x혓�Q��
���m�N6��)W߻.ݧ>� �1$SL9OS������a��R�,�Ƨ��as߅v���.H,-��;3z{3}*�61z��}��-�M��>s����|���{�i<ʶ	���~8{S�WӲ�2����{2׭!�0�T��w9�
Bۙ^0�r�@�A@#yِC6��/Y3ݜ��|���yÝ�{}��W�&D��*�u�l�x����1ӦY��V�`#?���GZA���:�jَA��ǁ�x!��[1����8O��<��<�����o-T&��4��8��yP7��l����I��ޡ�����pl泰E⢕�U~������nJ�!�PXlxVHYEB     400     1e0s��o~w
�zP	�< 7����A)��-�b��;*">��P�h[����ʍ�@�%�ѳq-��<>�%yp����a���
G�b��Z�ۄۜ��pڧ��n���C响'$�Mq��xW��(� ����i��ƥ�٥k9���(+Cu��1��BU7���!�`pem��r�P;��K�l�`ʇ�������C��ӕޢ ���r���0��"zXA����D1���-k�!䈸mʄ�c��Џ:?��_mW������#&'c������"�0w���j����*/<d�-p�E���4[�o<=��nκv$8@�#�o��%�h����"w�z���������KK�+���S3�4��f:�m����+��H�M<K�2�u��78��Ai>���H\���NAe}�?���	�<(/t�p�h5�A�i��)M�)H+�h�P�����A<*�a��XlxVHYEB     400     140���gS�h�@���Ӄ���h�Ӭ�Q�),��y�h�Xk�����B�53,���Pn�BbDM1'`1#	�"U����ٌ�wtQ��RY�`,�P��뿗)9Qtp�U�=n�fe���F�o��G��A�JC/_+IA}�k���Z��R�R��F�Ֆ+HF(��[�������U6��wӷ��_�i��o����k"]�:bݮ@K~H��1�߻��	A�W���.9�UȑQq^h`H}f���͍�#z������_�ɴ�#)J���?�X��NJ�9ɖ�>IW����t�)�K��%����*��;Ϭ�|ƒ/XlxVHYEB     400     140<Ҋݘ�&�
�i
�z��:-�e�׻p[É�����}7ѯ�L>���M.��{��ȉIs��q�C�
Y�zw����FQ�Î%m8i�� �~-����j����lp7҃%(����-�2���gr�����S)6��R22�S')ax��E�qcV�x�S��\�����uK�2����������)3ޝ�>|��r�e�>Zԭ����� �H���%/-�l��_�lظ5m�K?u�=�Rf3�H�%�9���B���t#�P\�{�x�cT8��p�}%�F5�Z�l�*�oiO�r�Y�#jY�?��E�F^}M�mXlxVHYEB     400     1a0���?J�����z��h9�YC���(!�b�#T�Lu�S浠5��Z�7D@%(P5���A�.��k+��@w�P4�Ҩ�¾<���d���~�{+#W���b-A�P��4��^�c ��bܢ1U�,8(av��5E��G@���,:b�'�_�,����9#�Q�I(���l���ۘ�(��ry�J�f�����s��g��CZyrK�L+͉��K4?��|�+�r:�tw�Aܠ�;��g�b�����;�:��J���ԁbnP@��Q�������F��t����w����\�x����Πҁ؂��v?D�Ώ!��%���(�����(�-�.�S���	�IԼ��	²�`n�}� A�j�����ZTc�������|¨��#�˖	�-�	9�i�R�m�XlxVHYEB     400     130�~%"�/T���ĩ���^��1��z"X�4��A6���|yz��zD��<�6�
��N����i��ւ�r�|�0�ͭ��{_,�0#�F�}�)���_Ҏf�3�T��������S�w���B���p`�5)��{�ȼ��7,[Nkr�ΰt�)ݞ��A4���;���n�A��34��7A/�E�o�ʤ�4޶?���/*n��>Rb뙿�eB�r�3 �#�J���S�����2�o�N3Ge
y}k�k<�.6שu��9��f�Ո�U�~�8>j$�����gӬ�=��� q1�XlxVHYEB     400     190� ���g�u�Ko�I�1㬶��8-���1����di+J�rW���A���9�cg[c�����9ɕ����q����XT��`�M���MQ�	EV{�$��XV����P"���k�d(-p�]�����5F/��_�Ї����	��i<J�^�Ԍ���.��; �5f5_h��2�����V
�]1}p�gΩ�9Q����y*����w��h4�r��疭�⊯g@���h]�#����r4'�e���WB�b ,)�tůʝ$Q&2G��+c`"����3��B�;,�ݶw��al�(z$u�R.�7�o73+k�_�����]݉w�Q�Z�{ִ6k"�
��[�$A�B$�D����|�[�,$E�p�9{9�#.��q���,Z���XlxVHYEB     400     160
�lH��M#HT�*'�N�t�'l��BO�nD�K2<��\}����ZaU�5v���W�kF�~A�D)7w���~�^�Ά��=�o�n�>~i$8@�Z8m�wjp�yt���A\wX� �p��ٹ� �qT��m�Gk��w�Ã�N=��4��y? �6���m�Rw��k^�Y�,Zޤ)�g;JK	��R�?�@��������m���F��
��2���v����>�a?M��I�'�_k��a�e=��K�>��4�կ�B�.��Vn��A�%�&ћ�*�n��~�^D���0>�vg��̛��Dup)����t�j1�6�ݧg��W��XlxVHYEB     400     150r�a�)"_S�:�zq��Ц�,`ᄝ,�_�O[�<yk�*�{@�b�����g9I�b�PCP2k�Bg��9�=f@QX`�P-k܀��c�,�O�OFe/�򤥞���W��-�<W�~b�wz���v�O`'�,vȰ����+��������4��!�H���}�ަ�@��B�<�fr;;Q�C�/$[Nj��W�}�Y�)�`Ț��H�3f/H�l99F��Uq������b~�SNGD���H���*��j�"�g��Y���3Ȝa�	���U��������3%1���Xh����[0��?m��8%��H@�I��E�;?XlxVHYEB     400     1b0u�}e��=��혚dGO�eMt���]��,�)����G�V��J"�C-3�(��V_�/-/�s/j59#���o��/%@��� C �k�Bږq��wy�תP]l_�f�gw�Hvg��BkW(g��m�lnh�!cI���!co�3��9&�L�[�1|�t#�W�YQ��[6���CV��FQ�|����ojS�Xa*Ÿ�yy+<�l'���AoArS���w���.J��qS=�_
�J�f�������C�@�;�23�:nvU�P>P�g���n�b/�_ �+e�s�*5n{)�5�������Hؚ���#64_�*�֝��}� G��n��(3��:VD����Q�/E��KW�L�?Հ%��� �&h�әb�<���
q$��)����k�V2�S'�*��6��s����wXlxVHYEB     400     1d0��#g9R�5F��b*�f�h��v|Z�W������L��y޳ޜ�=P<�ل��[A�_E�ʄ���!�Ln@��g_�}���͙���5��� 
6Rx��&���I�
�̂����9F���+>E���c�^�l;'Q,7��i�o�����������F�bR�̎PhR��U{J)�@gqV�t��p������u<6XZ�:3�J6�L�`�>����fs��r�M�*aQ�%2/�ͻ1~^��1m�SEGy���<�Pw��(X���)���y��IJ�::.	o�x��rb5foB&L�oɥ�O��NF�sj�<5�L:M���h��IO�!=eu\�:��<!Ŗɋ'm�LC��D����IgQL� �](�Q�ם��0��ԧ�%��|�='ڑݜsKG�� ��h�ϙ�Ho��40$�P�;�_B���P
K ~f`�u�"�A73�Bn��XlxVHYEB     400     160��d���̏>Rs��C��aj�5�i�n�ܐ��I���'�κ٣��UnI
W;���B��?$�	BH�o����[ﳛp��K� �� AUO�z}�#M�֎hn��>��/e���i-�{Ǯ�e�AK}
��:�\��}օKim>���fC�o�Z�JB�J�(�o`�a&�!k�Ě=K�o�-�K^���N��{�&���?���\3�K�
jeRQ�� @"wU���ܧ��ڤ�_�cv �w����� ֳ�i�k5Gq�~gi��G����Л�n���+��h�Lk� ������e�p"?�69��[�����]�����C��	p�>A��%���XlxVHYEB     400     130�e��[Ƶ��hS���_ �jJ�|�e��؄���;#(-<Ȝ>v���i�G3Y%�g�{%���}E�Ϧ�u�i���Vt��(^Գ_�7��G 2?/���-�Z�ن�(1�E]���<�Q�'b��7� �Ǖ�d��ϣչ;%f7W7w^Qw^U���1n_&*A�w��Mn�M:H3ȴ��So�p���EJ�z���Gr�i�O�h��CvVd�h#c��&��WtN�j�����I-�NW�Iwϳ��i�/�[C�^�g,{��6�	q���|� 2�G�����Y�XlxVHYEB     400     180	\�*�,#mL�8\駱k�DR��y�C�o
<��V)9�:>��7F������"��"q�:��z�Be}��Zg"��.�󧁬	{���t��| �|Q�t�4�1H�.S�8Q���N�aՆ��ɤ���?�G�P_�	�b*�X��-���lq��@3�SND�u������ཌྷH���=1��I#OD_��6K)ޑȓ��A�����̛�F%Iq�WZ%�ԃjk��)r��r's��rU�27�8͋�?zf&��;��vN�5�5�a>�W{a�ՉH(RN�w���#��5�Ta�y	WџɁ��V�s)a���qp0q<ۂ:���;g�c|��_(E������1���Gnxf.�?Aƹ��?0eF���Z��Q�9`������XlxVHYEB     400     150D�}7a\�`��W����ť�<����[U�M�ܥ�)#��~�4�sɻ|�gV;���$s��;�cC�\�j�4J���k���je�Q6-��3$9�o	Mu~����׊tH��}x.����������L�	M��ॕR
�VLx&����]"�]S"2����y=���9� �=C��� E	+��|ٝ�r�Q�ez��L?����%��؇d�1���~��,��F>ZWB�@H"H��R�"���	ͮ��S�PV+~`��jg�"���ڜ�D>�����i����c)���UҔ���R��^L_!X�j1�E�Y4�@f,�ǟ�l'��YXlxVHYEB     400     120d�3��Ԑ:��z�h���z������=B���D#���D�x5����P�a�S�xV��}�[+���%��ep������ݯ�_�����(i1�z���^����M/;����ƻX?�z�M�%�_�� ,��r*�Fs������(9��඼(DYs?O*
��p-֋��J$�(4�P�K�N����;"W�<r������O����#�䓇c+�:Ʋ�hί-��R"�k��ϲy�ѕڽ,j�O�� �� �&��Lz��WV�1}\y��}��bUXlxVHYEB     400     100�֘�϶�K[��Mp]S&��e��N'k}G#����u�������+����/�ε�L�������)pC
<���q����WQp[!�X*��U��i�$[��.�T�M6j�R2}be؜{H��d��h�<����ɚ�+���u�zU�K����
P��v�����W]'N�"�5Q0I�	&�%N����K߰5�M��;�o��7�K�-�}w��yc�ڝ1D��?!��ar�Su� r��}�EF`"�;�ciXlxVHYEB     400     1a0�Y�rL��2�l�~S:�<5MC�n�0j��5���7��0ivy���h��*�l����C���N�
�>�H��`�]9 `o�z$��4�!�b���0���%��ہC%����W5�ʛ�uz�t�F�.��x	�݄A���sxCY�.��]�$-)���爷��z��F�5�S�MN]'b�����,^�BM�_�Lp��'q��F�y�B��ђ��������=�����Z16�GLZ�P����`�����a�#;r��1�g^��;��񫱗Va� ���fJ��Ʋ*��D"o�ٳ�;��CI�J��o�7U�f<{���%D�w �]`��d{^����v��u�1U�rQ��v���d�F�I�eBx�"����J,a���J�S��[�6��ml�Dx�+���C��C�XlxVHYEB      27      30��v妆�M��G~�WS#>	,��=�3>d��"�V�*�	�{x�