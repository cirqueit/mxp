`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3168)
`protect data_block
kmd4+h5RRwfivDnQLcH+90tgKOp+4MvVwmGoggd8NWbwo+m+CrF4+6CedhxuCbZHm5llSWqXsMMV
titeZUc5YZYc92CL5qsBX4pyG9a0nigRaXWFBWjGli1z2/P3/CO8Q0izvm0EPx2Td4KVLuUnFHhu
ucQ65DElF086ZhW3IiwweWD1q22LajMGHH4UuR8QPfi95BXI2gPKKT0lj4txWevAbcCMDHcXLzkh
BYXVpNshXq1U6TX7bcnbtlKgUBlRfkdxV4Z3aWWu5GKeE6+TnYsjGkQC7DmTv9KpvZ3dA0ehPNls
cZyZoI4Dk/P/m6HPTbRJi6rp/KS4WeaR5Mpb15WR8EbMrdGvsCKCKB5WGaWsCVB755sy/7LuQ/ed
fJ4zCmqrB8OlCmofjJcTAS3IY1vWNWvP4kcoCVGWJbqJPg9ZPrN2viLgDo0rqUcg/0DlHEkrxLbM
d9dRKL9ivJvlsDwqr7+DxMlC3jXI3d1/+SX01JXJmeb8fmGBV769Rbbu4MjDEpi+zTullHSzBfy2
PD4Ig8j7T5lGCS30jz8GmrOgSJI9PyOeX/CmXXtHj5m+KKJm3RnHlXC12Jmid8/pZn5c2NSuonz5
v0bmFHTrJzxE0u5iJpmUGX9/rqdM9QaCc/G8gOjH47HIQ4JcYxUx82CLq6sijYxba81QB9uj6fkW
l78F9phqmVvrB3l3tUveBibRbysFiR7b4GgMUGkhqbsTYVDXnT0I9URwZ8nkraKRPbrhpE/PXBRK
AhbtueLCUncVdF14wpY12mWC/x8tQNjl8o6UWu0zWqn/McSqy82ZK6K0r0XISYgbs8aEipILTHyy
XIbkHLws3ITIoEGNsKsI74XuRjuSIGC0Jkw8ffri3uaSo10liCwdCYDQO2C7kPprJ9kLHOzuepIJ
p4ArM9wzbnvjW0sAbVxmEPuXyM667XM6VwJRzRNc529HugPQZQfLa1uQIZBHLUPM/5e8mmoKORb9
G3J1nZaNzsplHIr0rtQqZ8OzfWSAS2CpOF5BY/0XCHYuS0bUdzYRHMUu/bSCFSi9NEw3M/bh8qrG
qPp+MXZqgjE35anGa5+wFToCAyeyBsrv1n5aWOX+QPg9LqF85hG3EU8JCsgK3vnAsiX4H8JztcwP
I+3M6LzDyMTzDtBnXMJy+sYeMMaSpzPqb8nxFocPo1teoFBe8fJGUqQumVwtOK/W2Z+2iIckn3rM
jW+lo9Xr4sGBRt9K3uDxcMwEfqaXIki6uddjg2/51aGolCQaKVd+kpRjLTV1JTZvLVpi3ar4trfH
9aDBjZuMXAjxzMAgnHjuUANgJv2ZzGoUXBR8Xq8/0PrORp6qzTtVJngXtFE0dktksl14XU1Dfff7
Q98FeuSk49owZHOItWZ8u/wh+Q+j4PyouTXxuq+lytqyCmY8qs3sVR0Y+GgqeGxvCQbMo652lfRI
4+7dKBTYR8ZztmHkViG37S3Ri0Cif/lHZwcegUhlVJGfcgMi48J2W/n47G9DGFVcsknsPx9vho4l
5ruyWsI1nEzerfIZFQ0xIP2CkNtyKBoDHl3r7InnJwb+Zg67a9s55uvSWMBrdxDwu+IQDXXpxTHt
qGH0Ow8xuJ0i9EIE0V/oZ5akcrfwMZREJCSUxwtuc5wSIaJ4a9wGxgVmYB8mNy3RuOHSbTEkYIsp
tp4JuzQWSV29dLAjNBx5iBPC+gDSrk0IRXkPCp+vLn5I/4nqxua7duCyu7qbmf3KUQAgs8c6C0PL
qsXASNC95CeX8qTT3JlRffBDP6KFD3GS6eP9p7Uv8YhhbB3l0BAnGajLVnmVXqaMp7Rlal4GmMaK
QRJmZE9UYRcRya59HelThqXdoF1rc4DXia4Jr6f/l5dPtAglY8NsIBXCRNG9etmpIu2zYbmy+iNT
6b2S3HQIa7AeDa/Q3TmzcdWvOcg3es0pKIVapBkqVIxwYTXme6czREjAXeMmvslnxyrBd0RVr64H
M9R65OKLf+ofngHE6ldRWSLhWySgJ2f/H0eCvBxMJayVcISw1Wo3c3x7fXO2W2mv+9rGePidiQRq
YD8r1CMQSFVo6U3FTPbrfzQiqzWMve82vwKHmW2eSWPRSq9IjSmJJEZ5mi+FOZlitCALsZxU+P8O
Pr5UR8kfrNqoqOoJpLd1GC1auR6/MicSmvIoG53S85QDEfr+HwxQ0MJyId663vTeMgPfw83SfgaY
tU+LVQ470PFGDpI7esyVVCLe9gDHYN37vIJR1GhDcQVHKU72B+x8NkmJLiao5AdzfvMold68UWDp
z846Q96paa466idf148aOxuWxd8xI94b7E30D7c/cJ6NDw2WpLzHfHVT/zZ7HHb1gO46K6HJvGDP
0OcUSRiIG7a7UYMZ5zSo9D9sZCVUdQS9e6DjgxldJ8SBuYnMkkFylYCfzHUFWmAbyCHRpcFw0dBL
lERAWJypAhuYdJ/qd6K7Cyybu6kH4YE7qRxyYenSFwosbk97C25xW7ZUSxCU1C0/O5n3iSPHaZHf
Kc4S6AZDaUU6qv6Vmz/fyMix+2b8tdp3Ji9SwZLW5Cpa99nwXDjXLSUnsWGG6CzBakNdR87f1Af4
dyOQXR/CNUst5b0AoZ19CMf5QBRmqpkcun2+YgXcQ96icH7j97AxY1jRaFTNkWKhUShe4XtvkGBr
JtGR5/Ov0W5D7RJifYMvNe30Z2SwKacxxIVaIkDNd9/VdJ8cGkonLlwnmb+xa3r1DDft+yXblV6M
qP8POVfxXFVY4Lspc+BVkBG7ZqX+hAnHW6WN7sUpSE0QaDIKr0FX1LMCAj8z7DDebcxuO8khLjyU
mzfRspZcXQEQ2dSO0w3eAemB+lUgmqWDsrBbQIGsqidfDEjoWMgDg9rcP39mlEq1/OLqAdZXFcUJ
RMhhSZzDTGGEVrGWBSlK2FeZu4gMRV7XYGOhng34OxTRmgBOsbe2iU+RzrFdNAvHRBNmU73/zaK3
pA19rk8peJgnnI6VLVV52VAgGuLUl2ajhOMskq6TkXUgFTAK56A0Lqw2EKhy5GwL1N5MCsJLCKWF
9iE6EifTLjSNM8W5RYgGycPl/SjPA/GwBnNs4Wj+WlRaWBt3zpxDY3JaYUWJ4EJfE9X0kzQOQWrM
57AJuMwitQwPhelSEph/J48Ww3hytSJpKwxE3aAygJDl1t6BBzEly208nBNxflcgmQmZUtX513kO
ZYaGB0NqWe6nsaD4VJx0EU0u2939qgvt7ceIBk/NRPu7nfC/PZYopvzmqfJ9upNo9LLK0wN4Qp76
qXi3kUWADPYFJsnqqO2BGfzjnqprBnNYpuq3XNynl9RQ5LfVaOTiSu67znYrbGss8jCXF5/mrP8u
lf31OcY26jGoaL6rmqO5NhwbvujLbdpXfuJ37QBpgJ2gJFIc2HKmD0pE+U7Sa4nfCLLdNwWz6Qe5
jGZmunIaXlTd33QCm50GCJsfp45CaGMrKeuvG1ElnKMSdZaz3bhlphbM6kVxi7HA8w64avflsdeB
Eh5kr+zRFqd4u5Zfwj/LgEGgdYIIG+3Af7Ueu9ZsfRT+IyY46baB1q5QdRAr7ow69LLrbopIl6rs
NI4LSAk+i+L58JWsxiUfx64T9HZn8MQnfHpOL0F6ze1nH9R/oxauayQDISAp0XkLDyzFVqkbc8iZ
Hin/56z1+XGk6/rFZluy9IJNJnS6k2hpuhNS2K3De/wNnuKlp51CSd8znzWvmRL+auv0MalzNVZq
2QrYCvMf/EjqpBU18YTPEDrMTKh2adDw7aWsGKwAXjHEm/e39v8JIh9LwiyIlq6GG38z8ZHjlHt6
eJMgAy5wgmT77nBfIPqFDQTDvoKKRTgB0P/VRWopkaNGQmPOjnRtO83KG357HOrDXwB7ljmvoX8h
OduGSi4qpBqEB3TMGm41W/cvMU9DItoIqfaIvHbYND7vNoQ/dXfYkp/BU9T6jZ3nbWIS4/AP2/Ap
W0LDmak9YneglutV696bVWN73hL2XyBFDFKOQuMgdwk5Zpm7uz3kmZ6m8W6bLPIDC+M/hshbIkKa
ZMpnaVOtYeXiznr5c0CuphnIS7oKwL3TkRVJ7dcrflFfmiQJ9lK6SsVI/IqzgQ8khba9yR/khxoL
7Z2zHGX+/3Iqd4PRdtKnLDGPTFEh16RvAtz3cct13tmkB8tFvu8DNhA5d95UnnJWKkGFKs1pWIHu
WIV06H9Hj/s+uGmzPqxzoSLmUjiro8RG70A9SyF9Wgb7
`protect end_protected
