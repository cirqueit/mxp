`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12176)
`protect data_block
GWzOsV7xEzilf43jUSGXR0ad5LjIQrnBRrRmEI2dXZ0ToDjWdVcpK2ejY9L/+609uRPibVeoktvn
xugqUU44O4nW1lyXQvCEp5fUwtIfePZK6uIxYah2Tc70KtJPPgjziOwTcfsGnleENoVSbRjG9phP
fbcJUBto2EqTlmCFw25p5KNpQzHXXSJ6YT+qcq0hXCbwSPXdsEJYpGbsWrHU5oZGdchdiyVde8LL
HULFfZIcLbN4hezv8puae57hxtuCcRtn6aoeJQDav1obhW2Q3MU/XzF6VGOtS8pClNivKOn37XrX
b+vyvfUuTcz37wjKaGDnFrBDcx4fXQAqPi7plxxExzBmne8SDySsxgU62fF3S+a124cmd65TVY3M
8+e1cWu23ieXbxQK7vRGEZ0a5elaWZ05vszQQHqJKO7CrJqxZn1gVUYNmqBflF3UjbNW1u79MZap
1yXiRxN3sjYVU2lSj7suutU6MqB/8nVXpq24uORsWayPzuRQTIvEp+eSPtSOPUHEjR+YjNFlGUK9
Og6KEJm2xKZ2XC8I3TNdXB0ABG2WZWRuqfZ1jPHIOj9+o0inW6sfhqvwHWQ5eiAL+cVgsNu9yDnK
2Of6kQDkVYyoJSh6QluwA+5YdtX3HajDMsyb3kXEKWPP5cxnAvLmtWfBj08wbzOQp1SmW230ytRV
9Sw+PnEXYwHIr3tka2PR9bYRM7SrYyoW2TTUmHr2cjomTmCKelqE2vQEfGMxVpfXqapiIYL7hu6B
zFcDri/C2CkfkmTXVNUYxQQEsZ/SuxwVfI2n87Fwo3uEXyjh7GwS1VPalZGmiZ/r6m5P4EJnUu0n
fK98LtkOpv3YtIJpADAn+9/XdA/vP9cDGUFbINis9X9zJa/SQIxsqzv5gSz8/aFFd3yIAyDfKjeK
FBr5WqIqDZVucRsEn3PqNxpKzihmjPUDvPdRuBRv4GSZT/4SiuFItIBbdhlt4uck7vMz0tOyfjby
Cu7ywq9GwL6ngJvWGCn8lM7X/tuFaeVX0QcfBR2IMGBaPJ6JrAkWbtCVnWrlQWr1JFP8NOc+srjC
BwDGPZ9sbzXoSYYAGa9JzCNtt/NZgyghHYOWHjpUv6bdmfpBo300L4wcsF5hCKDreA5y4spsRGof
wiXXBM0U7qR9RQrOayH4NVOxLXj77dy6OHXpbSxcnOZyV9w6jC0YfnUzswr7BqOll938QisByz/d
FywXHZxwuWxgK77xCuFkKQa3ylUXEdsSbQl+nLZ7wra4lZzBAvBBGUMkYMWYGaU/ii2ZqTRR6gd1
IBKu9WoTV7svo6vSVXs6KinZw/5X+U+uZ7ZSvJQSEfwvVStv5D2LV5+48mX4w4+ArFY4bVrFw5XA
rue8I1QfIi+Ii6J8AXwbRN47SX5oOv//bTaLfy4KkJKPCJQhf0gdEZ9ogxxacEwsBdXhF/7PheVv
d0mkGQXK+i03wHKWROJF2OiI7+R4lDDD8YrhqJ0b/MC9eR5MEcZPrhKtVexhK31ChlWofebReW08
OASa3Shc6myiu4HPx9yjCjR4vTdVwFiqQskzhbFdjq6Q38B/mPTqC+W7KO+FNpLGEZbieOeMZPpT
RMTO2sEFJzio5MXhHOW9ebiAr4HuzEaYGVtysfwwIBN2kEUXCwxvR/9MalfxtqzxbnSRztqQNXKD
jsNDrQV/i1ckVQLLA5tnL650/TOqQ/NAyJWBeTlYYxfVW5l9VcGZmsES3xYci9OZpvjEqp5dp4w9
61uUkOHI0AwNkEbCaMJlvDm2j27fbM5FvBuW/2jRmcv7EkTnPdYHW7jFaL//hmixWI4sLWAG4ChF
WxZuH4vmqJdE1J6G4Avozns+G1izQtY5NUcxCa48a8d11wPjE+1Np3rZzyHHLUv43SpoWignF2h3
BTXg7yj17tk5jT1RXN6YD4hPB9XCn9ruJRubhFt+P0TQEL+vIuLcKVdWgJAoPNDK/NRLCcUYJTbu
mytSBNxRQRVh3ix/ijUbd/uNNdHiK+6m1zhFGVef38tCwyva83Ca7loBg3ojg+Hy7z5ojHUDz6ei
l7a7OtYHubhzBZ2M03OdgnIyVk+DedF0KDdi1CZSU40h1G4+EcQ7DVipddMMGu0Ph/vljPCljcCz
+LGV4kedA6hSx8Cx3qgiXd9ewY/+GO0IMQikRo9KtOPmGCPGnCv16ggMaK8YsuaUJuxC11WUUA+a
KYU1p5BPSZ5BpU/MLVjXFckoFeGsvwq1XDGxr9Dyk8rj4kWWDRMYXnf5SZOqhZz/7fWv7JlOCy40
vaYF3OL2g+2rYU7TASc4yroG0cwFntaDe9ODy6R/LAJZk1m/ohVfZRezYD2kckG0cQq8D6JCHcSj
UCMroxWsLvU6IFVCoDVpVImS0nmHk42BepauSoCCAvsDo4O7oZYenL4IBaQncTo9GFcHv3JFcieW
SVFouftYmpRxFRf/6eZMu2qHxfqdO2PuvV3iyge+YgHxmpmnlaBNSB/W7tEiETsrxxCQlm5d7WIB
hHaZrcTWWgw5lMB3MDZOYHWRP80KIfQbSIzvh0gS/0n5dyB6jEXr+j9lf34Q3BJPkn5XfbmJelO5
X89gQFRym4HOP4DeUJMR6jBa63Mu3MxcnZH2JnicZI2Lrek2iVEfEzCpTvFMiFK6xgDZHsW2I3Ak
cg/gTv4Dg+QOiiLoSP/VTFSpOTKF8BQpuga74clmzvumICgF9qDMbxHUYX6lBwjHCKC/vTQrndWK
vjjplJVm3ak8mVADhc+Rx9zlLoIPYOrYAzK8ySu7kHoqHmWKoWqgZrDHS8CGwxihJW+TLt9dPh0V
WEILMHStblDLBzJrfiIK2H+AjXq9OKvB642sJXlaQNTDm4Tcy7VeT4FGGAWrVIfPlzbyCEQfrkoY
CoaXpEp+/9uMxk8DHT1G+SuAc4hO26UHG2tH0kFcwH/ShZmyhi3RwkytLZNMBpzYqCejRx9Ij/5G
AZPG8kb5u+0bvJnJv/tp8l1KDlekjfZdKst7qjCsctSLo81Sk+sho/faP8Lg4bZ9ZN3vyNQySZYw
GENoPOD5OQPcqSlltoJSUFBGSZO/Kn0DHi24sau0Ih9jE4F4bcSDhSMBARHZytZ9Jnn2vqczwWkM
SpltgfoFzEDN0pQ4mYpGXyGCVyRqIHBJMawUMXgilpVENoVmr6WWb6d8sOS2RqcJUnbGP/Ptatv0
CRnhrimiBkfA3bXx17FqaiaIhQrJ9NTPm3j72bdWZr7oCPifc69Dazfvr3eorD9DYWnv9M5x4+Gx
U8f4R67qdt2nO37TFtDDry1TyLkUj2o+A0hNcMr4Hu+Jr8K6VDHwd2R7A7CHlFavdEOiqGkPvkHg
u1sw7cXTM47wq7M0dAIxmhEUIJYDvLLk/u/Vt+MCEB1ZqTuLdE8yvxXesyD743DB22jjyHq34p8v
b23ZRgI0Z4BPyZl8TeJyabcfd5OhRGOJ/+vgthEs733KLuYan7HwUSfq9HRqHifqS0ZpTR9aRJof
88N8iGiDkOcbmKak9P764wFcnrM5427yGNww3uxMoaw0owrAfnt3j7AR82UuEPS4tZJhR2YLuQjO
5GJOFHAl0R+vM6g9PL2j/h5DuA4rsAx4t4iS3U1pKlilgP/tyTp2aTX4/Y6PVLMnzXjXEaklOngr
q635Wvdi8kLVYwmTxEyg3sGVsPSvUx3+ztjc3Fj85vt99GwonN7nkxyVeWEzruw9vgxBOc1rl/Es
bXLW/lborkQPbxzdnUDIDfmMEBhNGyvv4Wx8ucGiCAgER8Whw3g0jOwZkGnK/MECcMgWuABY/Qze
IrjGvR/DTKV8bg+h0vPg3UmhHK7ZCw1ZSjkTXaVZemI1QMP1O1Zd7j6mrq8SvKN5WaR4wmxY6sqV
l45o/iNzls7h/sgkh75UUA5R/ElAqUh/w0nQf4pUrwCbkah6yLX0/XZlr0R+t0Sf0tt2iq9ON+86
kUbLTK9+ubeUiXp8jN3wTAjv1W8qbvD41pfBRya+0OANUXQksasnEIFMYrVXUbtnbBP7cm0Ngof1
2BTVxxHGA52tsfreHHdUVRygsxoULKMVHXH0pFGzpzFdrelPpjYPCV7jYKJY5EQ1jjJebYvO9BCT
d8AeFlXva4ct6zIHW2ilDmJtb1qIu0RzAn1VlZquen1qPA80Hua6cfD9RHV5l4AOJL2E8+bsKZYf
pynq9fBmXMjijQByyJpr6gOi2zRa7hPkqLXrlEFtsyzlZ+oiPivoARlTlqIqLWFwGVpuQ5HQTcph
VLYXYSGCXA5J+TtaYdEBnj0lViE5aHZOB6zVcuHrvEaSsYuVt9DpBt/3kUuQtJIYtSbvtdCR2pit
pyd8wJGEnN2Gnx75gNeySPSJowjoZoaeuZObXP2bw3uUANHk/JGdrHghZrrKoJcR6/3Ukd/ION9x
YIufh3h0UabEUZf8SXQmUp3LW91VfXaaiMBboztRayFtnPw/uTpNF5SaOxM3TIMHjE5heDOh3iYU
62tcXqTbFbR+lMCXmUv/SmuS7XazP6IpoFZNpWYQuu6yBG0WCWQzvuilXG+agOGNZwBk+rCWGMW+
uTURf7t+BCOXWp7zbGOi2iyoDAn4wXMtrLOnHLZTIC1ij73UuXoW5yPUbTDlcIl/52L7ThffXJ/o
+0cv+6I/ET+JJgsB45xax2eey1j8u1ytneajQ5fVxIZ6BHhQEGt6LvBEGJtFXabqP+5qa4YIk+ku
Hj/WJjUdGmunVWo0G4iGsLqArSYb6n08bdsyUL/ADGYG125oC7Qq/rJWDiAtzqsjR+P6PkWEwVeV
pBEuTO2KIWnF5Zwhkts0rU3PYoJmVy71LuNXhN3qkTuTpbpxr7YRMxmORAD9FX6wk5av/s9JgVad
KSZbPCFoxqzNrULvFaBs//CQlYhLSgoNWbk8l91OH7/6TEPG7n2cskJXEizGTLKYqG8KpxE127gg
twZsy1snQ29DAauLmqzDvfWdLFRo329dVgi/lTmqKfCVFEOy0OB0MNEu7Anh+CPTIlIrZRe/Mm0c
aYcocJcq6ZWOK+zv2Ad/NKMYMiITRngiWeqYXfMXTC2Luawv9QMMfPgWhpBl6hV3zdt5FPHI+wgr
hMsXwA1wrwGcaZU6aokt+c59IqZA892hom04EIKuwBIPKLb0EUffv5hUfEdXzB2wL80eah4Ed8YV
jlvVO5SWAgzkvpqfEZztCQcKkPysstK+A42ybWPvAx08fljSMFsa7r+LajKXx+RKq+Un+PwhK2BV
rxUYpuqIpptVdF2rt8HSv04maoUqDgw+Sxztn6nSphv7kBBrHHQ/aODhD/VN9IBsUZ5Nc/3JxcWo
R2jQsTDW0EV698pygpmi5qfflma/VTGUi+Opnwrkq7ho4lZEaMKn9gotXBNfM5GsBGccc9GzA7GG
PoiiTOaoy/qLbCXgsq9AsQP0Z33rYtj3SO0ppPub8G7ua9fOH5z7qwPADWV94ZRdy0WhGQgQNFWj
mcg6uXfSM3rDHFmJPZa7gXmObXKM9DQWob32/v+7BEYvXAOxxUUWv3s1YhKk16cr0H3onBvfusPH
Hk4yFcbZXzIqImKQZQNuJjSkpWgJEb2BnYSZvoHdf+4SNtxrwM2v9PnPMLkKcIqZOGDGKzw6LUze
p1IltPUV24gfxLKkdQVW487F2+Wsp/0+L0aJvfqlTFhw1FOt8Nnmg1JqJsuUI0J5g4IWA2r009zd
jCoH2U0rYi1+CkxVA/9iu8jc+cRmS2wa1a99V4TQgPbMO/9ndWCTaigdaRdvxPAhH1LGbkKKeAAb
VWYKufWfTapNQICa6CmPBMM9UOsp/7tjSeWVZFejaYPgkNhAdjWmcIQ/05BZ3Xyf1CdOHUgR2zy1
scyWI7AnrExGyE2Ewe4PuJ8wBe7vBJsnnuLTXvikp4H4LEI6YiNFc01LZFx0XPDvjqPXm5tisSs6
9AOBctx0twnXvMqid6ZVdUVThazkfFh/DNozksZMxrEHxePB8pRBkWPR0JP9u2t9JQx4ORV7ajGN
g+UXnvcidBQGOmTB2tHGaranvKTTyh27gYhJO7f3m+OheU9ojuS+RwDIXK5+n3UjbzC1oQV7XTK5
TO1AmlotZpQQe6fHPjwIAXRZPDnIYRU45Lw/ticLnr5nSMazuW3aPMQP9ZleRBQf1HurfCkjP+5S
U0dkC4fHQJit8RJ7M+Yczac3kQIizCLgWoN8MMbZndWaPtqh6erGClaLCrGobtC1XwY5/+VGgC7V
C8jgtJ5P99pgMd8fHgvEiVhSfse1GHmZ7Kp7Ptw4e3bHdEDinGHc0AalHnEcZ4DvlQho7yTcknKi
kixOH7zAnTW2kE4j7BZavROxSj2wXN45mAvbLISlNBW6dACraLIkwiWib1M1xgwtknBlx3f+aa4i
g+YsN/Kf2n9YHH6TmMxaKdVJT2xtZaK/4B5LLw3S/mLgE4z8kjvMABx/uAAKdQsx+nVg3V5ObIIE
8Qe/DersWfnwhFBK3mv3h6nUWJhVTEJSUTy/x8QRRMT7Qq8kj7naKHULZQw7mBt/zr5zcmCQcmV4
Y5fsvbgP1NtnjDbCAR2qmhC8ZVck5O65CALXY3vO3OoqE/hxdKL6gQ/NDmHF1fWnTYAO4+xLSmB1
XdYn0rvkJjp+KKiON7j4RrOGRthtGEBgPSbBOCkNbWcqNZEqZ6iABwTUiLFSylNTGW/qCdFnAf73
3+Zpa5mpTHK5o1q4GsfbgWXCsvyhm00a6RGtaqsOjcwKauctygKgOTdTZssPiMyS465G4copozgN
QjrpX8ekNtuTx9tV0n0KVyOkZBozZ8J15cVZAuq2b+xYUS7vWgfKA5feeLdvWbuVd7+V/dgbzdCE
HiuAnv5WgJ9Ug9nRkwuGS8Rlyj7+5bHyzdFGrz/0FLk4+q9yponEpLSMg3DY0D9pYz/gtmiCLZpp
QT66V0ltgwlGFviU/uO7GaawOM0ljgldykYIhX1t6eB08Rd/axtFJIMBzjXAgXvzbjPKls8N2awh
QrKoPhwlfmZ1UMmdsflZwfpPAvDnTPkaeSnb/M+f4LIJ15zrLEKLN2707QYOUZUUwONMhla8u3Bm
9QLalN8nAVzFc1rMDsmeg4aEqHniCt5v/GYFZUb/RfbgiF+M9LQttsLHid9eXUoOAzGbrllfuWEg
KkBTlsOaCDC091QUrEzSJgFZ4xy88nqTijoJeJ6MO2/jZFm/0uHQ+Yaap4nDVKQSWFK9l9x8en4z
W+MuWGrPRppa+cJZRRX18Sn/CWu8W2TutM1/zR0M7Z0U/sAQh5XtjlQ6enAw7R0FUMKGtaXy8qUm
+eVHutvjrLvkYqiRO1DK1l50uYfTmBJeMWQuqFeiasrppswrP9l9Al7bCHo2W0Zv84vJfyYpEbQR
3bqnf1jUwGOInSJHL/BPD9RJhsBs+L0yjrEx1Nqv076FuwtEQoZ54JimYHYcVbYFPynJq1B68o/M
Sos2w9BgHpzNktwRjqzsuwBis06aGDXaD25NbGRZfEZdLOcNV69FhSID+p2p6hbIFubrXlcS2a4F
R5SvXhBmWM8noA/MzfJXYurXnfUptXbX6ABGPR7e5MbsADboMfFV8jzObs+ywlXdQSYbX5s7ARzF
iK+DREJMEOcD3pIOqhvD3REjbwCRH0LbkU21/HVdK1QwnLfbR+urQbITXF/CybgmhaiC4XLUe6xA
JTsMVVVOj8f4pLqEsG+HzjtQ9Lbx4WL5Y4GN02W5qv/08koOff9m437eXyaUfadvJgWsqm/xpipi
3KuRrC+KRzgPXDqBBQdFjQ3SQnpzHFnK1QEHwcK393UVQ2r/pOCGuI3RWJX7IcFoyXIsq2t2/gM9
MgPybR+lHzzwhJDn0kq6uU5B7yKBnLitKY8ZSeB4ruXw9xrekRNPv67BOA2jkqYlpxwEY5d7LWxR
AHTOehCLY2puXWGWfXDH7xapAB6uADsAJx8PFZkffrPJCAWiE1hpvwNRg69Za7T4cQ+ma8JVujED
PwyFCSCoH1wQAGYlEVd5n5sBZfPEjIoz1gLKYUNXgkQDscIcRMdUheYIf9wK+168vlL8TrYTx5iu
RNhSe+IbdcgniSrWD6qnm3HB7q+hqZN8cbdbYIJ5rbiGYr6typAD6EXEumoDtkCaGAR1Dz8BzVZu
lnFPzWGoAabxNix9M3i2s57UoUMsvBYjJLNxNoGaQea3cF9/k67SKt2OvTSbPd9Z0EQmj5quYzDe
8hmoiqvmdbU+49yuUXY125/+PI6f4MzY3RyGrR52iWd8F97+sLdCNc6zfRG2F4JD9qXjFdkxIKqi
1/P771PYC5C0EkoHZUoPs8yGZ9Vm2WwU59I2tF/JUIbPV/Fpl5L8XYBtp3sXNtc3ncs5snuz65VW
5S+1td985Zv/OFPa+6NLVTQZl/x+JfizaMhUJCYJDOw09HD3DyrdP77jM76P9DC4u/eFhMnJImkE
kskJWrm4x3ueakypykyZbdVYfMy21RSlmTYCaJQJ+fRkf6aDa4iATWyL1PXrAEw4vpbqsEoFR4fa
pLp6qvzcATZhukvEr5IyONt4O5omH/SZJ1UPY1Smjp08uYG9rzqCjz0U+O7Zk+NsPr5LgwLPbTMj
2bsRmt4WgAJ8O0dY99CbDW5MYG0cMAe35rVBcocyz/Xp9LBnxEdauzx5+F8GqTbEXtT7sFDyhIq1
et0dnjni1jnxK3vT1muuE/8o5oG1hrTGwESMm8CQrygeF5YPw4PxwikTVucKq2mrprKknkMrVMwx
/9y7Z2mvN7CcP3a76s4vMUXNWmsWH+AycETPatZ1j+lUWr/n+981ocSQntGd8mHiWdcfsX0sU1FY
u6ClFGkG0M1xTC/fHYiSnKrySZFodFjL88mlTzT4FZ9mXaLxfXvU7y6SGKRQFeu7Z7m6RIEHZ+YR
fq94I+/xnhy/TNhSSz9BCDsUk/ooHcfHhPb3bFuBmp0ub6bzb14ncnvNAyaXRpRhhONYr8VUuNgt
Wmu9+SDRgYxgqQ4lKNmuSHy3Tbhxpwnyg9trX1O+VzmwopGo7qDxrga3mIC+A05VSW7HuoRHgsTA
WkHDy9c4U9OqymM+tuLRUaqs76lWLpzo4eVECtb/qeQihaDKfrjGNtKgGi/RlQfeTpeLz2IZNVSw
JSc/jjtSrJyYiRVYcHGgFVoIlzW5V+aKewHoRgV2GcSE0dzQ0deWG3kuTC4z3Aq+y/o/eFUBnDbF
dyJ3tIvs1mwwKLN2ezYDFcJQePP2sdASCztPFFhH44Ia0yy6rNOzPew8b/XPkIVmNQ4wB5SLHu71
PiXO5X1yaAXsQjasfQFwOEaqesNZOoLzUWPPxM23lkGjPaF+ZRrp3jXs7zvnuehBv5NorDvPcTcH
+cd/m/fF7Y1rxC0l/I9TPCNYJmLLAJr94LgKXSev6QI0R21njhW1t5NI/b2SJ/xGWxeklrc6Gmfc
h/VlokCIy5OrAze8GXuoK75YabzbAQ+5Kpr1XM7xwx5/VYThSzXbJVKX88PKGqdmyLJYJw0wkOoh
GeXS4KqOsaknlSWuX4JBU8G6xJrHzmXvCd4a8BJUY+kFXBFjVVOjPsa6uwaCqWyGpQsExb6M70t8
GrZT/Wqwi1apIFPDoiGiSQFyf8A2wnIQzX2LpsIc85o5hIsgHA7s7u3dXn+byuy7NAZF6nkAaKpF
qLnuFYqm4O8NMPQlyeWcpsWjF6lJA04MmM03osqHDBPGIByITytkB0sR6pDa7syBTLGj040CbecP
hP+qjgCWQoQsRbc30RtGk7aAklHo3y/MyEiM/wHzyBdiszugg1MU3UMc57xwVMM+mXl2HuuteNGH
bR3AXdW6nUU3OGQBmAlc6YlMC+KLqE8GEi+ea1mgLhuGprpm2Lf02OJUEOeVnJFKvGdZPGaxnn9Q
42HWQvNIzj5RC7y0Rn7mxxW7MaCD5op61Mqz08poKbLg+EEnnHSSpD0pt3jUE3kZCLDw95XoT/TJ
yukITnIVZf3H7WrCVBMXm+MqXYPSBfiv2LPp3Th09fPEPb/vUfJL9ET2hafFPzvcFGo5Y92bl1qD
SpeH3Jd0SWzc2MSl4dw0dsd913u+/oU4XnWzg3IVtdRCSi67SMn6JhmQnbslLomfniSK5ggt5XSe
f57EWi/b27I3x+bX94YAUc7FAPn/4l/tmF9EA5YYlkgZONGNYpOhwDmrASkVLd0Rp32j/Uhlt2a7
bBCdn5Ng06qNdOFPNSEWYk39KeFkEljVCCAQ9k5oinaTg4s4eC1pGZauTDFo+9VlgG0e2dxNXb4k
JdsjbHBoB8SMg+xKfESKnsRL5OR08MYjHGvf6voHrIdHwo8lJKffPRuhE1aIN4IEF5GXZ8wQtyib
xDBJaWOJM0+cS8eb2uh95wMrkR+hvEJ2ohxaZ0tHmQibbIh3t3uy1aeW5OvdeQb6L4Fi3EfKlKNL
CODE2clY+CD4GX6kLub/Z+GNTQg8OpFPCyHbOtUELrbn88qp98dlXCcW1HOqjvZut2+ovs1KR7oO
mwSKZMOv9WH1PiPrx7Olm+BUSB6Y3oY66nLI8VVAhNp0tntBo1oDNmRRizJSCtQ+7hi/ZbXMRyQK
CQcqvbUHjqBC00ppTKjiqFP888MmvH8125SJBXFdYozsCrKex2IUT/8cZTV1y87cJPArw2PmjOrj
e+uo09tcGtNVa/PW/vja6Esj25u6xkyk40xnmYEmw4OsqXrGn5HHEh3aO/8ZG16MyD4E6WXeT/16
+egJNoZYRkY+okmq0cF8WkRFk5SdwR//u0lC9StByiNbio5jUe2lwPGRwz/ZL7tp+lW1QAs9am5j
3kQ1Mcy5oucQ72kyfqMF4R6McGCQg30OREUTJZsKkVuV0RgXoJylndhNz+O9jdqYsHaVMmXtRMiF
i/TCPIrEchSm8bnC6c1VekSUdF8rJGUmJi4nKvF2/qDDxOB1rXMMUDCZJRnozj3Kcnpx5TO+/GCo
z4toWtRNju60+BeSKdVVPNDqlA28wwLpCRrTOS/iXYUr3vUMwX4krc1wfmV+h9BDh62cCpwWyVEr
QA2PYCAufaaBU4Cz07c9bTP252o2FvSLwiDc2r05sCCL9PvNQyj7cx1E9Fdu5Nx7O5tMDS7MpOEy
omB6JfD55NXi9aIp5nMrRldCF79wEuEmHDBiQLTW8H/5ex5MMilApdmZCw1iooT3rSTnexBFR7TR
IzJ8Nmiet4qfnNgAGzY3NepBygge9E6HIxWIuxy8AIo8HNLpbXux8lif1rhu+W/UzGmgJ1M9mWzi
3nDit2AAaBEoLO7PbZFfSgD4MEpIoDd83RZLJogV7dH2QqoUa/YyLRNtREpsZR9XKvMXZ3Kar+oX
f0dIELFYAspIxwfTQuuT3yJn4m+Gb4douCHXh9yaK2XoT5+VcbLpzxOVWPsU/j6YbaDlfk/ym7Yh
Z8fxLNv1GmJxxg1YTFyU0i77KW56v2OkyasfDUdPN/pfSZ1ZA8aTxFYd5Ix2WDHwD4KgEOIvWMy9
ZPrzEjjRio8nAsVtF7TTecfwXeZru2ix+AYRjMMX0yeyuMZmtlt17WCNEC/xIIkYXVYgSsgSjQk9
HECiYccnSP/Vzj1XI5FZJhh0B+85mXRUXfimhYomm1uNpuZHyejd7agWPPGYL91Va7Z1YqwcmjvO
hhuPKFA686C9EpvasS8AAoCcG1WRe/b9rDSvUuJDV6giQBBciXXq0/qWihy1QFzCWEJIU6G26qUK
JHcF5+6QFRo0iVL5uigC6+zfsgtwKxeRooUVeh5hi9M7ZkSzIQZGk9zU3NM9hGSn+eWjnWO85ruH
zQ+gUvn1UrOc5l7E2DVqKz0h7plZfmvjPw0Vzjqzr79j5yOb3RIgyWYlnO0J1kUkwf3v3g1lAKsJ
jdLkwMFL92ZrO+AN3SkUvzFzS1jVhzxuWLVbFABgY7P81PUI/2iEF82IV2F5oC0Bj2HYImx05afh
UZuF5JD9IuEsnNmeMSrAhis3hmM2JMYCxiTKJrvOpgyIkkrhUwwCc0UnhU88qF4osUebjMdtOHuN
m6nvwKSYT0gO9l/nn40K1Ks7K0m9jtKLWnB+ni/lls1hLSm00ciDn9+ozg1+jps7jtM2gwzetixe
/zHyqp69kwQGLVTohnc6dVUxSoJqoLv78fu/Axk7ssk6ezvRJHswUBnnre10PjQJrgtm6OJ1SkQp
APjJBvQr5Q3uM47vuNGSlSUkNVQTaf7V9L92Yfu/Hz6MJ/fz6pUhZAfmLfcuLSXcF7lPElLDsSVP
xbh5qZWHdOWtv7ugz9DM6G6O2vOpP1MTJfcLcFRGpl4dUgaL6FsCk5+kUU2NTVsS+hj7sg6symR6
qP3Db1ljDa7eN+T3geXCZQn48wXTEBsP40KlQBXHN4TPjfGwNj5RTYPExpRm9LW/e9rG+rKF7Ps0
A7UAhS9Ubw1+Ged6li1Xu2191WTQXR96yL+9nvktQ8bQz2F5VK9gp0SU0PC25ne2g387y++csMYB
hrwTP2lm4LF/cvIsb07JlMfcdGEAsNhe9ePjt9l7hORKwy0OyIqVpcRGnUvF6jowbPTps74vD+xy
3S4ZQvI4biARRkoyFbwJWtKeTjRSUN4FbepaueNWEZ3V8e71nCKDRyA9E9ShQx5BVKDhKdnqB6eI
v9HsbgQ8W2YTCkDbDds/3PvG69a/uGWk68bRCm04xN12v/+aRSrA47izGA62BY8gGqp1X7WBr+3u
3SRuQfPB49qz4cJ1alYNUpJj6M0wlXhMAm2EDER/Q5FXW8oofuamI5b/n9eqSvQOebRPjGk8Etkg
CxqLO2/OCKq/vOtHk9X7Zv0N1lm5KkXdeOuqqjMnbym8CXim8qcEcwts9p2jBY6b2ZXd8T26ps7Z
rJho1fqZY3STeUMwvjMKWOCqNLxhRyV2fgbDJpSDvlTtm9pPbMijHlAEYAUY4wEi7S+tOeMSUYPW
ievPg/qXqfddktsF2qbweJhpoI63Fd1p0yA4O8uWHy/+ABUt23vVkQ2pTQR+mYJds0cV54SzNG9v
u74LUxrBMVdFCoICNNw0R4Y4KPJVFuMyoATDLHV9Shy6L2blCPwlOfAILmX3aJyIdBkUgfgs/ldj
FGKeAuPcmoy9rg9Or5bDg/CHnzOl09xUq+Uuj9eUmLdgfYagfXIBV4l3R1bT9EoZv8v/oNua+/D8
MdfB7Dv8GJ28WbxPV1B+/qzh4gtM/2r8v9o6EUWLcR59BYZl26I3+s7BMwu5eDIVodq96YBuFCLg
DuyF8e17Srcb+l4ZWxHAUk3b9ZNK70aaYFLnxo3YdOO/UO5WbQxEBJ7O1qr8k+COaVQrINbSgBB5
gKGfmbhuujvAWyzqGJE+VE1lIz5T0xI+aD3mBq9AmAp3h5sME/kwofk/VZBqgWOPcD1AP9p/IT12
f26FHHIuvoC18S0ndQd+LYyeIldMULamvV1L9IB6RomODPvpfj2Dxw88P+j7aRwVlirMiHMQCZ5B
Bs4amf9txRYk1auD0MdXVEoydASEZG6gNt0xBsqH8PUXMVY7bKyLd9Cda+VwGyfKBdHqhHTTQ/Jf
9yn2WMSXaZcWWMd/2Y5ONi3cOXdQZhNrUppxrvKyO5cJak8uFDKFZpYtw3ey6fmATptQ8ahmc7r3
9BStwKfnCG1fWf6h8+FwQlUndTxf2YZjYJ87BWC0+44QaiD9eBUESzyvpuTpu5CItHNQp6tgY8pW
qyZPB1iu610Y3kR1/F3SmjF3n6nXKcYc1OUJCVeyZdcTDWBvaLvzCVKFeCVmJGopZjtQ4n4/Rg3w
aVAt36p7lIy9fzkytky4QRMY9yi+SRyDfguW+agZY3RFs8PN1T1e17j+X2OmNCqh3YhUkQQCilCs
+zx7gVazanP4kNgeqS8vVR1cav6NEtDEhqcuJyqpT8mqeWGGtoDLfqVG5WCPZ8tpOHtAyLBGlBWe
JkMfWw8KfEwQeXhFwyx5cYbeguzDm/xQR72gqpIDH1Bdf52DXA72nhj5uDh/+7K/VY0yUKjB+QyD
W+9vJiu7IbRLAJsS3jRVLQXuDYk3GTbBJaCGM1WW9JppUPy2QEmAoyf9n9yvYcqH/241620dq4q6
EqQOMhH7uTT8krzgV8l2+Dw0zhKJueyNYKRKePgXQyN90QCLUruodJ0tJIQhijOUNJreohHyqYW4
fK7ZpMWCBHHp+WVcNfccp8dm3ib2dX/AmxC20YiiuBFgX+B/7+DeiUrpZIfEM5Fr7DfzTiJui0k1
BT61IxSTFsh9kbsz8c0cDekHYq+P/EmxuCEzR/ZRKFroNhNSOeEGIwyxJA1KjScggKlyoRomztM+
FM+01smAbwg+NJVdVLlijIWGmwInNU4gsdl8hD//Ig8APKSbLAJh5JcPdyRUMHepVO3X3ucjabxF
KOPu7V1bduICwUjwnekgKta6OSYXRqu7d9VbAO8uxYs/cwJpkx6PFr9Lzcq4QT85qauXoKAa0H3f
VNyjJouDx1cqFi7jVwRTeJlvkyAGbeuQxML5Qi8Z8jBhBPlMIfxgiL/iWvvkueOFQ6zl6KkR1jWX
LlP/xLl7y+YTLYDXROzjweggGCs1NGH81gaiXyoLwk1Vicahn3QoEaaUxJoGb+glzr1Ssuoj/Clc
0kymUU5CClLOYRv6ab4CHwsfRVlLGBqoJ1hWtbeUVQW6TaDTJmDZL0953hTY3oRcyr3MXN+nfIah
m+v+bafD2kx/h8EXAtrFYRkK1/m8WAB5ERpLt0GxqQ17VM2b9OYu3YGKSCKRT/hp3kKBmS4BeusF
I8d9HwkWUx0XGiJuKkV8RZoNQLDUGbg/9YKGBHnk6zYXNDaHUjqECjWVhO0r48qIUDY8hpm6AqXD
e4fuXqMu4cAGMeWuZjneVGqJM7nBwYmkiVYMGvpaIyIuqC/UR/8dIKaZyiPAXdJYkWCGlys9BgM7
VF7C32DUZyUYD2GphOptOlFWzaJM68UXSctskdRJcxDhwE3e59SHcNpQSgkAldtBP3OK47XKzDyf
2CkMkVqYtTBqG7seinfbO3pWNRXHK3Ul4Q08LzlHwqA1SgdPmT/tpNHXHACiucMpvlip5cw/YpZQ
zpq6F76aEsm1WQt5W94TbycAemuWXeOwmDnmaFTRHzXrGcNnxm24/DlmVQfH6q3bSv7Dilhjjhxf
QR+s4s4wW9xh/8EnuflcDstnu36/pAi67eqiJ1GRd9zznRfxjVGHLL5bUjAMv5oH9tCDVjeBnVVG
NIHkpLsDwynxafnR2l0ua9hhcd+fXZUqcgEtvin4rorxhejUROdt1f6FiZGJBpJGktNIl3LmUhlw
O6No+3ehXAGe3Naj97OL28EJNNYvbyCqns3ePkFBuZEyhje8rAavRB9gAU7m5FGDNPUNzD0qK/a4
G8sy1D79mmBViweHnnrxTfA6eZIlQqrZ2Eg5vi1WSLcaJetPlQA0MTthEp05IHYmsyxVaXz0gFXY
bkrvzsptmUHkBe0kPOktHuo/ZCs5bKgX6n+VgavOCZkfjnolvn3ZptwWBq5OZNTerGl/cSDbdVZd
+tivwKBM1g9wYnpbq8E3zKwEZ7moFK2WfLuQ4nWZoluH+wjnVtslZuLVOx5OhNd5VlYMoWRCCLDu
KKyW/VBqBIYz3E2tdpO+ovo1z6X4K9NkqzcLzVA/tMP5+ClZ1MoX3+R73Oqk1R0HfxLP0bJ3IwvT
O2yfzz+CbAsOogk0FkneptMABOVr9izNn7mMLD18zU+ZnxHHom55q+j8YTW9R9VU+3iovFCNZlW6
vDqS2lVIMPk9Wchbg54WvjA293T5dpqaKlqhhg4TS52PYSF27PPwmxAs0SPGW2TW6LgIrVRmFZNN
afuGl7NaaKQdnXNWi+Dl1kObEJvVieBppBZ6igDu8EFaYcAb2YPh9X8WXdl/KhlCri7EXsPGYTFU
c2bl2pfQC4RRc2ktugCQEmBnzq6SsquhHwvAVzJK1qh7v78jVBx5dMl64xk8pgu4VmQ/0LgEXrBI
E5ECD6vVWaNwNgR2KCt8Ug3uvEqezUug9esgWgUOLflHAyknYCWWVJeFiJvotwmFJYBrYxYs6Y8u
9j2yS7JkcoUbvY5hSpgYRKQVL3g8V3MLYyqdw+OPG2T8I98tLjHxJQj7l5exIYiPtrF3CqOuYkf4
SwsNimG1gC5SJZ2sT+ftC/j5Ij56DEozuLnwuuUHjyjuiwxr1anuxQLA+PscxbhMceEep/lwUx7d
DiXxdfXVnpA6Df5QxoH693FXCILFcZOfypVT6X7gkfkegaA=
`protect end_protected
