`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
YwZPZQx69ZM03t6W2LBPkrTZmtXzx7BGOEJ82ciZJZybVQJzqtzXKfjTI3MfzS2HKJJYPQahLdjP
ANT4OdcTQ/oP3uKmSYCMawrWeVJbcrbrtt/AlSoULqr0I2/VghZeeqRkEQB+g++/V7ACji0Yc8i1
IIobi3tnDJxaK02y4TPfdaVx+tM+xBGZ6IYcX474ykuu53vta0USj+nbL/V6jdBfiJYx5NACzN/N
T15CtXcBMilJ6OtBU0CM5Pu22DA2FdC0AplBr3K5Adq6objnIBcIC63BJrGY7LHEOQcxqy3rRU+s
9/tLYEu6in0FDx4rRVKPpt0N+QCOoibv0ANUKGkUV59DOuuiOZumFsgDCnVmWIYtK3CAJ2BleTD3
w72qb68dYSuIw3FC1XySv8y8kTTbBdFGt5L7sn4riryMl12H70AFobYET1PEHE4jEFryHigZnNWt
kEDuUzcBVPG5GT9wlud9nMlcw4oRCxrDE+TEJ99sy4mOQt4drAPjKTGsV4LwvNouEX7SsgVOTWiv
Y3TWWJWnQpvV2rY6/T8NpyZ7PC/H0ZdaLvvxqa2/Y638RaTIciD6tAw2HadD8fqri0L8CjpsLjWB
arQI7m+7rstRrRPuEjPAwl2E2RI97L798t4ayvR8i9SbyQCNJFcWxh0l03+yjLAUjdIC80t1ldAt
Im9YOiiZ5TxY9N/GneMY7pB7IiQi64R76lqosqJMFfniBycJa+ibAKMjXNoq3bFrzK3wT6d4OaTS
Ooy9AB189Kd/AXtSfo71icCohwVk4oX0xTPxJ7b7/gIMDddVx7QLD+QrpkvjuToYd9v7bnh2H+Rf
dWg8tqzDmqOa6abE5G0eRoeJfnl5VOBV2wwsR2J/mk9BAtqcT3sx804fWzJq6Yja0XbqJ7xclsrE
GVx9MHcIf4j/8AHHZXVJwVOVqDmfsf18ApsAh8FADA5eCwU+/0S72TYIekR6Qhdqfo3ue717N4dc
IDc2asg1g7qsBpRxjuNeARdbr0GK4zcHO/+JxB8zHxcaEO3/mLfRJ4xfYb6Y0InBPg7680MWTLsp
za8HKL0BrBVxXPVaXYHt5nWT5k4fA8yYCfRRwmY2AgBYtHol047U3Mf+3Ni5jrsQSA0Oj6Hy70si
KenssWhR3rcjSx7mtd1yedFwxLSa2AN1xcbc79s4OAQESNrR3J/H86qYhGTECZNYws2Zo/n91sgT
dneBsVmj308q6TTfme8pYpXbHl93wGAgoHgEKme2uPztkOj1KGcEn/cgpNu0DSyyM/998cX+6c/R
VEHPau77LgVOeyowySMGzWCaxK1+XDouds+5HeH5WmniKYsGR7JwC/WBjgsgY6mgTUEZa+HteGKL
Os/PJRDwaco5ZmVjohxg+lKMhY4ncfFpbUex++hNYefthy5w3NpnW/ni/oC3pOa02/x9u1muWYlw
Awgo5jO8xqwOaF7QgeP92LOWfR/nKxPg2kqCXZRpNWRsiEEiuA6cx8qPEQ7T6f6Vl8F4wKE2iZSG
h65yAEfSyCasnATmqVGI4jro/nQN0fWq8nWCB7LZzULURD53d1Vn7NRN1LKy3b70sxo8uFGbAXoV
/aOjxgDcUWE0xPzJnobGrZ+g0DuVQQKc15+v6oBil3d7BRNyuwp5RTv9VnW/NB7lr18jnES6NBo6
O3PVrI84WA/V7kB4XSVrf7FCatyXpxhKe7mYPDR5BpU9AaOxBTxieIE3MHTIPhEY9VgdfQvgoskP
vQSsRzF96yRp8OevEr+kf7VK7n0UZdBnA06Nm+aPUKJ7j9fVaDMmo4IlYN/s6zyBdMUvin5ZzvP0
2RsKtANzXZNO/qiTPIyaUbF7unZYXOL4gl+lntVAeB4WAM2pz4cJfCFQc3XhvfsON4a2oAiyFmAt
dHWqe18VFUtiTeA/HxJBQb5yDovoIS3r8uAB+hqnJMP7TdqW3vN11VIfwuIPFvIxalkSqDxARI2w
TZJfPJ0EcdnzaxJkraEnApubOO66diHtMqPjm1z8M5oJ3NPFmuIJJ1BvKVKxbaX9z+5FIvSKaXfb
ktZTl7hJjqlXo54wpNrxW+2KU5iht5OPLl4q3cZuaZspiWW57vS397EYuGPYZPyxHfTQ+aAey05J
wglYmVWFcvXg6jhHYu5YBWjcazCRDS1IIBYDgLwOeitP5wHAyIshKqQiQFlr5z+oMkwAVAICntuY
TMFCHpZSQoeehcic5N+ZXcQeb+PSIyTUCF7diYnWVVBdxhoe28+6DVQYBFol3+RB1JRJiruBS0Mx
ZaqpsR/fwpM5nxbr8O4ewGUDiDk99kJDcfA92UQtZZRc2JWvWVQTpRrKPZSSpM9/hwjfAyrEWGNJ
xI+us+/nSSuLNZyiTEx9DD0dCNC+ckWUGN0urJy5ocnPHWof5zG9DY9b+0AGzEuQVNtOqTLeytSJ
H0+u5XVG09bZCnhhqpNeZO1+G3u8212oEiv6mHsy7zaU+l+1IadqgIwpUUOm3RghAcPZBQdQ11oJ
EfPtD3xVHUZcE2nLgRdh5BZQXmwNHTdRMMnm6PsiChrv3/nF+F5Est6MqNrT0uTiIH62i+RowTGy
DjU/JGC/vIv1vxweL86T1uB1JBOzTtml1KcbJ/sOMbwKk34SSFt04B2q+cXs2vvfjEZaDb8uXZOF
YjuD0wG5rurH+tvs1neq6vP/uqq6Bl6/kOamfJYHet7JSUAzWUV6csaZLuEU4BdUJKWTxXnJHFYt
uLRMlY2wYqKuBXXyW7rr18ED0/5tdHPGnD14HmDZFAgsTRnAOS+93lfAjXljiNFObbBBfzswQs+6
8JSIxDPAQSMy0o4AkSh2ROjWs512RlzzNdH7g2Liit67OWOLLRFZy3D+BeK2T3+zIg1/8fLqzvE8
1vlt3j6Z3MlYevmIUtZJKYDA2CRa/Ho1vGnVayfaQYdEWPO6Ma/voQY9iC3Hm8faRbnI5/YNfCCW
/6OjKujs3/ZDfCdlrXEECy+nd1HT8pbJPWT25wum/MD9hvc29Rbda3FkmU4OnxgGsN2atXOLg1uA
XIBKLjvWjdw0YcozC8lEMmAKyEtCu0BH6QmDFDsobqULW3NrORdh7mHs1ytEhI1BLcQIJSi35gTa
XQZQpWSUt1LNK3ewlLl9fdPDkiuPYlycNH798QnBrEd4/kaS8a0OVbh91++oqlmLjoaQzTkrhJAy
/jgzHRg0/brjuQxWlD02IOT9AKaz1tya4SuXuaI+wDAB4ech5UMjxfIwhp5jYECvu2zfqIRiRWq0
gXuxEx1tagZMn7vVpQDcWixfiISHmPi4eLY8iWGBHlYoIaECNB4NDOZ4shC8JDnfbUzwoIScwzfz
0Mtnrv6VyswqXzHTsXhNIb8RW32J4HjJ3sRMqnZ1IBulEKiPCV+laH5SH/JfceOZX7KoWLnzukJa
Q6NU2cPetKpBIKOAVL8cwUTFaNsuFN0ZrtAxNE2Li42tyPQDE9bk9ELek4X1iEUFhc7zBZTohZlf
eLjaOx6e6fACiS+tiYzclvlbki2c+OssV2ccmYhBCogd3RG8RQPccKZvOUW5ZEjHhh0o3/4KrRQd
aFW1K99FUIWtMpnLtCkHeHw80SVKqw9a3OJwLqezScbNYAG1m/Zwaqy58qy6BKDhdkPhVU0RFLZx
NIiNl3tneFH0STmjSmWYuC+cxnLIMj1D1Ecc7AAu2GNjfuvXA8FbP6zc2YoRyL3Tz004NOymQmUW
tUklJnr1R9BU9JkWfw6ErTo7dyYGfq2Y6XQ1ApD95X9IRWDm6ccRAowjsbpC0TqK9+TolvlruraU
tlvBOvMdH1aubacq7nwxqbz4arq4Cnrfsv23YV6bdWErpBQIloY4/fFU56mtsX3juzHTQsQAMl6g
Oc97bCG9zXXLOYvZ0Q7CFRojMlouvLHyDCVNemOVYI+YhNH3TOxF2LGGxV3MC708A0E9EZozrVum
7wdc6yOkTsm9iSt3Nij/4uRzhwybdBDKNedJ2Y+ROiZ7A/Z/QJWKnZ83HGHg3N/JNJxxUN+QH2zU
KELcFBGuR/G+z7KEsnAAgyOJxV9oeEnjQaNveJjD+KpJ9+DH2naEb5ahqEucAIGYcTH8psSaJHS6
4vYx97Jwory413OpPubMerJjZJn8vmffygomfbPyckYfD77CXNzQEPe1lUGGCrFftUXUNkrD+xwD
iKAB2t4Kbsrz6OHNa1uNfIMDB1V/Er/b7l9OvR+36szm3nRE9rt5mDAhG4nB4Cd646FFKEK94cwr
Wov/q3E/28WJJdsB/ZoacPUzHXLhI6K5zIDTQYZTCsdqlwWZXItgS9XKbT6fkc2u25jHjjOrbs5T
HksOAcn7ox8qGmeWDZV7J+iJF9PrEXyw32XAdpKTQ8gPQMnc88BHavyN8fda5UdHe72zuOwft/fu
dbqZWceR21Cr6OM/FU5ltzxgbwoJsqfR9jafaCEWRyKiuJbiUQ7y/8cRKsbYsXt9Q//WVtZdknFJ
L+MxWQeRsIRt/jUCg2xJ4MA9EIzjhYJSyA1yUaWI5OJ8qNF6vI2ISUAKkZDJEruFsyHZOp1Xo3VR
MVVwpApVhejWpc6BGAOqh1GhqqBsibccABUNOOfxuGm6FaMgiYda8VKjJsGrJ54rfCSMKrM5426B
v407XKpJ84ZoKT8LlvpSANyl/eQ64Lw/VJsKgQCGekAE+iPgsIbSL8zJEzUlgcXOl//DRY9VYWzj
7YDHRKGANdUIxnc+xEzqAwauGTUce/Lja0i2TNVpP16JQZotEZPk/VpvthrAaaGo7/oCri3EEcZp
/2vXX6jBNSz6jLSODOKGXLPHA+3ywxgZQR7E80+v8rCiePD9BiFetq2K+IIbZl2tUWPPJ5DAPk/A
ckqlyyLX8wPtcuxI85yMJXNuHI74jWPYWVycDwrpkz5TC2oGZkpgP2V3R7sSE5qpEHadBhkFRYfK
wd3+P0aRuM4bz3KXxWONZ4vErCeTEpTeYQww4WYGn96q8DvNOKDEkqt3ycqzBQJ9Act/mvx4mRu/
bzfL7Qddir+3EBD9jm3QGnxxU6tsD7qKt1gaDKKQAkR6Huvvx/YpJ+pa9tSCKaP0QV7bmS2SHpeT
kX+W2Sw0SBpew703IP2fpuu+rYhDefMvQeRdHoN8h4YWV7rsr5bbqgUlU7U2cz3rawQUDxspH5Ra
eyMapxeIlsrt5/1GIVIfDgklq6y62zcUZNAYD6Crrs2/dAZf3SD/yDbbyC2T0F/tgHBiCP5e+c3T
2ma8biy80UesvD9MoHwpA9aIf5QwwFA8EbL9jZotzfTnft+VjRhfvBvHiRuBibTD5BgzhuclSr5k
SeQckDO3arPwnB2MOazEsAEZ9cJx7xKaYa8U2htplxpC1EDhFWkUuXnVf3j63tNyVy8jyWnblYKl
9TCRa2bWuzHPmy7D9VnoerDG9Wd/2gNyDgUkRtF17JzxsTyqR6bs2ETXT/3u3ipTBwrlj+EhKyox
L919FKrxKsJQkLYI6nw3Ae8XtxlUAnhp4Dctx3Rmo5RoUmcOtTQH+AmwFeOtYeUoxifrQqnkrLQy
EKMQilMHC37HRu1LGa2LsrNS+wLkYhgksl9YOrysMVnSbpsLZXXW7zelfkJIxvdmFcx/SxwIzbBR
ED9ifDWPOxd5JTXJbjPYTXVFQhWDJWSJ0FR10bdnNQ4aca98lNvLGNs4XWeJ0hFLin9MI2PcX14b
F6GtZqjuwSrAAKhxpyM1cBkoe416OC3oIb3waasS5QBT3ul81I9gcAkmWX/8d3Ez8Ptw5tnHsN66
r5O+QLx/IMeGQHv3KokGpHCrMIXOmvZhPbRIfsQ9OvZ1wa+Da/RDiaHGsIX6f4H8Q8MLmnfA6x04
oB8voAhCg7bjKc27zPvWhdh029ovNxrVjOrjfl28MIXO4K0xPy5/EDGWkrxxf82ZliTOV5+CPNZ8
AAvd6cWag0tZzkhh/p2qgvTy07tap19J4uaUWqTPElknMgnxsiyc8epnClJ4xd9KftBavu3pyz6I
PEYZw0cKAiUmD5AIse50obN/KncECWZuKKoxotRRwjmxgbCP2BSI3iICXQNJb1Lz1XmnfKjKOay2
Q0F+4vvQce9R8ZenGf8vFHDcggd2mSO5tTbeJ5Ql3QzpqpFem8hcL1YmA4UNFI8rKPeHXEZW52Ta
5q62BRdBzHvn4GRcE42qPQD62WVjjjul0fS80xO7iAijiuVQBwJGaHOKcDy4tIo8KkbJj5Ntd7tm
WgLTCRinXH5jcPqnwhuRsM3bo6htse8fNVto5P9sVzmaQWt4V4u4Mz/Hj+r98DElmMWEVgKQ3vyc
aVo9AwUoXN6n+1gRvHvgfy6vxb2oVkNaaAivLAGvUlJcPX2EL/jcl1UuxrHATAUXDGLTTS+d9lZw
H2g3K1ZIw1GMn+C8JO9tTBYQqnjwnaBRZmt2obdGSH8xt2RmIRtsK0v+xtHNw7k+0oD1v1fu5jJh
ms14BMjHpul9h+AFH+8AwqJCuWMF7Mnv4WFcR0FAXCF8NStsVAjk2IjpZlu3CK+FeWDaU1xUoK+k
1diPlrKibA62unqmWRjSaRltXDgyLBzCqCKM2gAyb55PZTwoE7ZgSJlWJ4KhLHNPEN+q7kdkM0N8
mlWvsCAGrVVebxTdlpx5kfYiDKmxYYlOzWksdzGKix/FOLzM1CZ0MBdULHTF3BkUfnE1GUpa5cCg
DufAjQsfigZmYsZFUky/4yIdcFMTmP1wiKOBPLRr39rV1iWfdOZ4SAk1ucP9dc2IBklGQoZ0u1O4
oIp0akcDz2rd53O3Wo8/xXgngybhfkyqfGZJeVS+sZEki0gNHxzesKn2q39+8L350tvsdJAivJWH
dpWmm5X0jKghaBs2tcZbx4IyO+QxGMkt2zEbMZyAyUpVJwTwEMUmFbR/U2T71+x6FKFp9GOy6O1V
EUyLwBcxgr9tV5LiC+fsCmsrYjeH12o5GTeeKDw/71kYqkqspwXEKaJ0KQYeJxMW+tfREFPZORvk
N8fYleFJBf8LnLJFTP8jDQgw4rU1RblawrMpWaf3ePq2K04o56awk7lV60h6VLEdLv4E63/fno7y
zBDSS/p3xphToePWBsbmhkjtKlQsfiQQMgaN+7oRxpv68NhejcvankYj16HN6CY4K+j0if5u9SVI
Z9jIVEOEmpYYc8Oi8nZ5pUOWyuLqJ2DVIeZ9otS/yBARO6vLubx6ZlMv1ZLr7NEB5y8uxHsRPXo9
RLCsaucnj9RnCoOYseue7d+308qv0eLesSiJs0K/SUIDe5vMTO5rvTa5zaU5YkOXYZBLuK1J70YJ
FxiBvSJc67M6/dDMmbHFNQ1VhEiw+ZPh1+1NGiJKreOtyDpxjQpJTvzmycbe11UCb5LB6L39Klyz
BtuaLESgQ+/C2iyeGK6qUDXRncDISL3z4Lld1bCH8iCbltk12OkXcS12U8GICLMEhRW1+voEqTMQ
MeoWty/1fMarvO50W2hp93dlmvr89jySjtfNNTYDNlWzAj0hGlHDDPAt3UxGcePbxigiU/KFIFi0
+abvLFwqSLtvseWxgDJV1w4FlPe6/JeQ4p7MZxfDIu7p60CA0lpEIpBxjmdMaS+4QajBww00fOqm
tioUQLtgc9lCd5FVxTz0QSXcg6yI/jddJbDKLhkfY8H/yjvKpg0Xu34CkQrMC0yxcXDs+p+t5625
jRpACOf36qw/VbIZ3tmtBZCxyDnt7PgMaH5Vp7TvLFRcaOPl4RX/sBoJd8Yc2lAEBDI1mWNrI+za
RIDUYRO2xVrHGP78hV/tzWDOP6zfw2oj+IWUydIV0mzMo65kbzZj6SmZKcGJAlkUc6rnl3YlLZOx
spaRc9MkgvrrwqFGvuvMDgxzlQe+jofdx2neHGxIinmWxl82DtMo9LbHTAHWtkyl/Wt+0eLxeAcD
7YMr/nOvE796yl4EmkZn1l/JWUBfiwEEmn1aGTcJm9hGKfyqiMXpV0BOZPTclrK3EqDUVONoqCFf
AKqXdupi+/RxDuFyAn9Bh8ulRi7g6qjbwnJOtIa1FholC9hwpFAQ2ZLDAVMfgksHX8mQ9YofK7ZY
mwY5A2OGLGVgrIUOS0wdN/fQ0VU0+I5z9VW5M8wy6PJVLCnhVIRpCqV87DSBKyIe2h3uceCskidm
kzRPHPEIGPytH0f7I0qvMMVN8q1Q8E0M7bvea8vtjAk1QHo1cbDi8Zlj7mOhAJ8739y26HbWmUzG
8PwdzAZ9mug48bFM7/ONbl1HnThlWT/oia+lf90ouZVM9FuSQvreP1BFbrRAGIf9YXe7TsS3AgXJ
VDR/1Tx8KJbCIPJAx/K5p6fsDbeu0d+BKVzf2lUfRECsfTodaieJf+7WcdI2OHyBvFA0VM4rWJ1H
rb25GBgqt5oF5Xj5gG+o3GIgdrBfOCJvFs/fTsIjvWOs5ePP+yLSS6TK54O8WMdhDJcHNWPLoswv
StDOfC/ZXcdwU6p2LtWRPpCTEZBH6Xt67BxkgPWmPA2rQ1TMSu7eZF7IZANpCU16IlejVpPIXxtK
gahYoZiggz6YMX79mfGk3w==
`protect end_protected
