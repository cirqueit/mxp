��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Щ���GJ��%�����h�K?��"�J����;	�p�qy|���R)M�i(�����bQGc��z��%/"���s(sX���7�ߪ �#^ ��4�)�˩@��_!��LAU�$������G��1��ҫcDH��8�o�	�Eה��ޕ�X�%/+���^��9�zRC����\\��>RXt����)w���g���w��+xS�D^"Uj�|���=0�X���j�kﹷ�I.R�@���.= Ղ1p�@Y�0���:A����,0�$�K����)�My��Z����-1{^�a{�e��k�j�x	����@�O�:|MC���c`�)�=�M�����tJ�]�8�ݖ�j�R_j�e���x�A��4֭+��ڛѓp(��-	�[NYPt��P�hX8�CX�bV'e.̀�5V�vƖ��v��a�'�N�g��Z�o�(Y����G�qV���N���DY���'�_�P)[f���mC�g�*���;3��$��gC�����dY���v����V ��&_"um�/;��
o�<�$���.������9�1)a����� [������{��2n�̐�⚕
��I�-�B���t�H��E5�\q�&������)~33������J'���
����/3l��	�G�v0���X�^v��8C��Ǣ5�P%�ȉ��:ܽ��(�Z������1Ro�L��m�@AbP����գe���ipu���8%�z�^`��a���{l�({�^!1v�AР'^�<�X;���a��Mb>S�͑�Mzc)��CQv�=��d̙���}��f�!	8YD���5u���XH1����3��þ��H�{$ْ��`�a�ѝO\$���V̂Y }�X@+ߌI�Tc�9�cȑ��[�*濾&.Ȝd(�Ğx� W�q�af�"ۑ2���͡��ER6���oQMl�N�U�|\gݜ#+?\���>s'�j�>��� x���A ݁|�׃�֖����h*�QȒ��l�U:�byG�/��{������k|���ƙ�C+�2��~��Di���c�pI��Ұ�)v�d�$��=ˤe��?�G���N���-BE�]wCB��b�Jݭ�d ����
�P��Y�d�P���լ�}�	zO�i�2�i��_%�̺L2��G����e������6�,�X��n�b*+�Q��m!���GP{�)�c\9�a���Un S頙s@�z}���zf�Ah�~>J��<�����*u�<�:� ��X�����U�LN�Q[`Gk�����5z����ktcI5����Wk�(e�ӗWj/��XSi٘� .�^���lM��+Ֆ�}V|��t�	d[1.��P2�W�9��8�)��]-N�aQS�5�5x
E�n#j˭�i4#?��]�I�h��#q�覲����DV�8�_��8��D	����I�wv��������V��F��t��3���	2�iU���/{ԓ�P]�$���=~LE���քt�� R�>s���~�2�:��W�
���1�CN�ġ�+��w���o�