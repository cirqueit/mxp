`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
6my6mtFrVAsFldvBe6wQR+XWzz1uogfbgTfbvf0hShDegYC+BCcNmEXM+Lw+ALrMzZCmGfEINWk2
vONjK4y02W9NeUJNnci+dNU+aH5Nk3Z65tqqG+cen6k72jgjgj05xleoUHOIT7OqpkUVoxgvn0pU
UZWggZU2K8DzbpNh3Ndc/GTviH2L1vN6S7YPFs8ePzthmtyO+pX2luhp4VwAm79PB6yB8m6mVBaR
07kv3vxhZJOcu1m2gg4FL0p28v4SQBgM7GUB3+uZlS6szCpfz4HZs51V+RyFcRAaB8W8B8AX0EwH
sypuViMmCLP1oI9e5HVOG703EJSymxnor1zQpJvteXu5FH7hm3VZHceIVtN2EYfkTP3tY5aIVKcd
Bv6mR48KzFRX4Wl7RI74z3RvdF4ZipUYF5B6O2jjp4PU/NnhThlWI2s8Rwf1aSOvGN/zEG6z2NAb
DxNTzkGy8k+7eyiLMv+zsm5CGZZp6j1n19xwF4C+kESn69Bui0z9aJAO8Fmg0O/BtK7vZwSc8IrA
8hDSROZqD0H/VkzDgWLQ/DCPd0NzGgiWbdM5qW3bloIGa7BONEjoiy7Ok4FFiZpVxhSTlXT8BlIh
zZK1GzOSscRWIYzC5dJi1l5B79kNUBb1pE7PZ5aJ4O/H2Ve7NiEdLV/9bJqjJTYNlFug1zcylT5c
F6igem4wieroXxjZwgU5bcSyL9yN/zkXuFyo5roL1dfiTiK6YaivM2an0t0ZU49Alq/OJgyBLDHP
ml2isFPSHtwX+0dolKdPCGdiQjMqKHwIvSdmAqVyhd+7p1zcvOHhS0Bl83D/s0zHYXsYhBU5z5N3
qPLXe3I2ej6WW/x2N/j5rpg2NHRsKXZjvtde2QE6jxJkQn8JXhooR8vZ3KwXcJcbJfx20FQ38Jny
cGan6VAw9BgEczFhAI3JUdZEI5IE+KDZ8KUXVMlRdoc4lr6c7rk6upQgjQO9am7kgfKIl4HF32zb
gs4T8w2sRZYGN3WvvLCWxjdUktCUWQfQeHFfWS1GsbMW7q1qb2dompzTFdQnAaWOPY777ZmecJLb
FLvMVUrnRD0AbCJjQ0a/hSoKEbsLKp6O0ujxRoFg5FThrXE+Z3E1nJHT/Jz5HRzz00biKm/lN9mU
nG5kUmq7oscIkdmhvzUxdAesQLIeT3ro4qKQdgHU/eokKOTcEWI74DgVwJ8VyB47FhjbdHNgaJHh
qJIvGrV2fhgxGenvQeG++dpzcPabvfLB0mxdRXQIQdwSaz9E24msfw34VMm3g6oBcA12F3rgnV4s
6IXFa2X4Tm+KzpVZn2xj3+aRQDIk+V7uic3dvyoQ98Z2hcMFBx0ePPSAEfuaGRR3ngwSzyYoLqS5
APHcl1DR46JEwGdPssRcqynmrT5wWivIAu/XA3k5dhGBBj9PAkUcxtniX2jvGBXdJQ+whd3djCAD
SbUC3wNvUBTMzpixeE+Vqbak+8pEJfhCZxSQgiCGnmaqhlxjTql+7ENhw1Wo9hSJr2N9UUQfJpfH
xrFhZCIJe6I1I7ET5yq5HsDQ2EB75FLgKONGFjSWsMxnAI8Xj287MM6bYnT+h9aB5N/IuvqVIZ3L
emWik0DW32pV86yfBMCGoChc8snPM+u14paeNZWP7b1HuOk/v6fgxVJAMzlVwSllPmvZIGbdciY/
nvME0VNCajQyNlVWjDWlZeesKOQ7rURL9bRGcWBmOuWvby/rNCmJzk0wBnycvvaLj+CFgGkW08zr
Spbicy5CtNAnUyod9NqEcaLxZA5Wi9aiJU0pNgsZlXjchJr+Py397ZbNSuqLta7vBjajKeiTRZfn
23wGlHLCagioFJiOeCBSEz6UNAjFMdIJRpW5BLKRihWntVNqmL25a9I3HS4AQXRJ8167VGrIpofJ
lj/+QsIJSxQBtSRzSQHB1cQC6Ub2zBu64Lcp3QcEmUhnm8bcz5mQIhlJ7yMltVAyjyr1vjchGsXz
45JK2jb05LXdR21EebR0SCd2NS8tUUzP1Enm0nXZhookEVnDM4QdLUv63l3+drNyY++hq3H5xvAO
LvPkqTvHx0K2Kt+LotEY+1c2fSNpyDEcyqocCY3Avne5hIAxrATS6brHWlMbeo6vZFztrxZIvP8e
iLLBrSfZAmfF/3XM0/MQ9ze6BaLs/BCMa+4KiNm70nPtrfjrH0sWdmhUun1QBpTTnMXyDi90SdsP
N5Ll9pPHd+OdYf+H3PTzB4WclRmZyc5/E+fpeXCiT6DxtlvggrdCJLoZw6kjoI5FyrfSLDfiR6OU
29oH7DBCAudOFc2LiAhUjMpHLbuuzYFBU8m33uRfKJFCpqxBDT5/xJGnhL2i3Hf+Y2aQCR+SA6dy
NZhkZzMoIFl48/la6xuJ8u/ymge3R/SoP2tzpuatFLlSMn0kvzwLreBsWdvvj+CZDZi1jpctXKWp
M/54uibK9xCdX6d3d511MgQpvCksfXzKD96vbiMrbCArtQJN6wneslq7HI2IMFTB9iBRRcky92eP
+6F4fGwr413EWFzo8k+dW+0/pIInUyDoHD1hErvUtq2N+MN1H8wcnFhXLi5y+ykHU6IoObp+LiH8
hzchE7DUXuX1HUOAHVEZlibBN69cEJjrlCels8NZYaYDILQ/3vUyePoI86jhOlHBOtW6TLMOf3CS
dlzf7W2sWTisQdF/cehfvNcutSTeukHmTiweTG8NPpCBHMA7ORMbJ2qKPT3d99oM8Of2lkLOdAuR
lH5TFJpesPyGTmkwULZaw1fWEx1Yokqr97H+/yank6qtpXL/BwfoN5xBctrBhejWyRImYG5Gu4ZN
w5XfsOPNZyKSTEv8Cuk79XEyUaEBijAviFQfsnWaYIUQ7Zx72pTBFslmn0hDWJb6PiXmW17OMqlE
e2DNDSsWeduQq+4YWRiWb7nt4Ako7Wh99Cn2Y8JkyMtuZMXIv081xxs8DtywKNSGbKRnX1Bl+vsb
PfVA5Dj6o4E2xmdEnK2I8jQ2HyacSJAJE1iWRA6jKi8qR2f5b4XjDB8tx8kEArECj9MiFISIIuH0
zn8JLgAmUbOj4D3k9YgdzP2VL5jv4wOgp2pHtZy7dPPc7TNyJbRHokfqFB21lmNIO2XnlqBKAsGf
HoQf+n7W4aoUdhYZ6k6xnUTmww+Y876i6SGyXeniVi9quQwRMRN2YZotOB5T5Xm0J0rsHDv1QRUM
+7iEii18TJNDQmmK6aiurYHgDwA7SMLO4JSyI0FFHhSvj/K3qktBU/wA+5hW7R8mUMvZ+dkN/nJR
8GW+6gqOq0L9SK9I1cir4n6zOBeGuINQmFclorp0KgjlyEDtWM4jAYYyfLHE/jIVWOkLYBaNy3GQ
64jtRyOwjGo0557ERL3+EygeAuN/ZFOODdt9lhjLzEwRvQwEE1gLU+CGGseXGQgNmPY7MHLNs44J
rz2fx6CcJXckeQqhn6YfRLZd6Id1fWruII8VhqvV8debgD1CVgkm/7N4Q8YQy306n6QEaKEA3rOa
lGQG5P3eensBSNNJS/nOK3AWkS/Cbmwm7VhwPONic8ioofJfCvCktPah6Z4UnvusUGZA6/uJPsec
Hhw3YeOGNAcYKNht84NzWCmtDCs5VldNMVqoIoDep7QlJmBL7X567Tzrs/FNVhlPP8EH/SX33CN3
TaP8ofIJgfcza/YdEJM/BBBh2VuD4dbEFPpfws6ifrHSokRm9UVqFEwJCA1BClkMZUJyPVfnoCR5
EmdXu74Zww0S0MJ4Svq0UE6nyIyGKIY64p8cow3gooKna0ADF7wg4WGdEljmftXTgmsa2b5z6j1N
wT6uHawmE1SvukmUxTbQCJM55qG4/G0EUCsONXqUktZQ+xXnSkINnAyWFAhWivADMZ9OenG7caiG
jHa5+7zSUokG0B44H+W5U1tpUWNGg0oY57frb4Q7Yo+BpY3uIzw2QhbWifwoFmfdK1ngf7iHXz9m
aj1d/U2IrOqhNQi4wAIwATjDq0H6lVEi0LyB23PQVTyhDzFGt15h6iMmN7AR1C3gHlAJh6Rjo1R5
S6a0y61HrvnrQN7n/73DrBsU1MX0HFPnJRGoFDRYOIjuAkEVGhOq+0begb2UUupf4lQyI+YMWvKY
Oi4RZJ7rlew6LTykfAyKMKP2dqdmMFwci86RQzSlwY/nzrwD5qLLlKzpdzTWGZD9tVMf4VkKzjI3
hNVCRa/5j+a6E2x5HImVnLZPZEOTRhBCP0wCMX8TAnMD5Vlez+VP2TBO3efXasF5kZtkMUWQDbty
AGd6zD5PrzE28eqtwKlvts1LEvlfq2CW1uLPX+Lc2YoklR2Q4RNQM/uWGTDVQn/ZGXdWZmnMX0Jp
eVyWBFbqvvv3B4YaVyPmAoZ3kbe2BMkWKrZj24O+UJIe2siO7KHp2vPsBZn8B1+nuNYxqgiK26If
mQpaXygMopr4rmHVFhYPwqrt+D3yXjXjjEQt473VCMEJakPeKuS66VzWE78X8g7GGFknUdC5k7FZ
j+Dl+l4+8V9cvXKqq7d7GI13+P5aqAStp82z7wDhX8sAaIpdkBsobNLZ8PjJ3cNgla+rpWFHcDca
NLAAVTDb3kMlxG0W0DRc855yt5StIZn8qaut9rjduMKd5Rpr38YWq4ixPsUt33ilic9YVRn2Sdc7
tXUBtXZ4x9yKLKsj+bJdwscMMCuLup7kjzyS/uWCewFY1ol8ja9ERs47cGZRTz4AdWIXZnZ4QzG2
gnP01I0453HnAVEMKu65tH//AYM7aLOTMIwQyLp5nopY6guoNgIM9CjkaXVdLS4zeWzlIVV/TO4e
Ch8SK7j5D7KFrqndICFAZx/P9dxls0zbej8Db9ItHBGfZEnbw8QoBOV3yuYjyD0jtPzSg8H8b9Jb
OBtdGY1z+dyk3KNtBcFZcRKJHUI5WzbFgI1wxMtDKTpr0FG0LXnXE69owQAP3AwOmDTpN8VT5hLt
PGq/Rs1BBYASn8Pws/GiY9wQVTN6lmlOfN4By4Y5mjwhnQG1wzsGg+SBR2h4pBS6OV283XKz1Gll
uMuQN//f1N6qwf7t0nbvMFC0Bc2o7aQbfBZihVkZY2VuS4rq8iop4+gTlyrnD7mbsau/kOydAF7O
G4ekon8y6GolYIEzfwpkvE7NA8RoG2Z5WAidyfbZSsnBOr0GbsxxxwElFbZWuiYudKEwkmfC/Z5d
NbDhFhT0EUYlbA2MroC0gOlwEbMHWjHgukpz+WHhmJ4jVf/o8YB0pit9nRnm7WtZuXIaCcEf73NE
pTFIxFIRSlReDkD9xoZPPiKThP2OOWv1AJMDVjiotSQ566sMTiMiJoShswUOEv5sI4j0bFnnYvzD
ivcOK3udg+ndVL5BYHi4Bpal4t37Sgua4WYaorVsMFDnymiN35eMr23Lg7t+LvKPzpHsCn7Huo2p
MNpS5ok22TmxmeH/cjV3YDyGGEPymlL5uvWS9XnlJeX5kxguM1VqBcCYp/jgdFZbi4ZpjBKYtICi
rERiL80ZMmyqUqQHzYofHMdZX0bP5Zq3hn0UWQgPIItiiKntg2ZRH8ZhMiCIZ6EdhsimjhczWYTt
f5yFZP12gt5YtYjVnqWRo8ni+F6koaDYmCiGsJ5jDosvLlrj6oPQP8pFBWX9Xy2RiuucwE/LGm4N
xwZEBhTt8V91p48RSjI0C5ulCClcE3AI1RkaOSUKhUBueMVwWh/S3Pd/I3HRcU7nOX6J/J26U7IJ
HIoDVDOg4w+djYbMOajVkdwj9Kw3eESIZeo8TyjRb/bQLP2Xu76BTpQqLHu9AhU+oXHEEDkRgW5y
+Fo4PB8GhJYQt/Q4Sas1A70fD3uTdQohcCaWYUo5Y0bVandBnuF2EMcTXsiUG3ppDDpFb880y3r6
kQvkCsBlKSIJUj/zGi3qSG+zpIGBkkCo4h/Al1EKVtyHnVbotTKgcy3bp/HlWrDCpomLUB2TohpB
bqkLtb/Ring/AXCh/go2vNxGUMvb10REwwZew+y8oCBfcxIGu9oe/NQYPFbA4hoCYSvE+5n0LOFA
dcto8zY3cG0U3jGhtEmnr/CnadWOZPnG2ktEeKGNN7fQggT0pQ59NthsoCPvV1AJyDHe+9u0NN+F
/THqIfLAboBX5gRHBZ+ZXXLzwpi1NKLpZGaQuPlKqIHFLRDhxIoMUw32f6c0pGGvRh2ntJ9V9InZ
K1KfQWJAWVoKQdDdVb3ThXbyI/5l4kfEutbEhuVsmiyv2irKFVaWjV1gUK6aDofJ9NhsRrefhLnD
kVOl53CVlhRQ2rLcSL5bUG95DVygTVI2kqmzrLTo54UH4LBG2YhvrMzAEdskMRwEJg9wez+sOsZi
WFIEzNv9jH7w1mUDu8NWS8iFkCxFOGFLcD7W0ocSUWg8j7ZncTVbMRjFGqIVkRdYkIkiepNt8zpT
znZ4utNNxwAJN66/l1tSqvSDk73NzjqaStV1ouV4SqAU5YhbpaJVXLS5CGf/Wp4DlodbtB9mPLdj
iIsff7qAalN0JH65xJp+FI12Y2IAWIeMMJCCsmn3iNOUqsXqQgzGGyyX9C6GGSviOuZzPCvRqol1
yNJ9kQRHpVTIh3MWEc3DDG3bTBbxdIauZBervXQoVKQcbVHV/szBk/Ua3NuxvYvKL1wvmdciFCvS
x4Fly/+qkXXP4ojsLZ5MSvl5OXeCDGhDjuKvDXkPufgHWKaQ9kJ2oC+0L6jOx1qtg4i43WF7tgqB
1glgDV1P2gZ9igR3R1m8VUm4Rx0uFCPsQv0Bo1bxy3C+3yobFpGkTBFx08LYvjvyVUT0WCxM/s+f
wvuAMif8tK0XIGSZkQfO/E7L1avh8rCR64vNrQWUTz6e89KWGG9Qy4ZZGjbmGN3C6ClRzQulR16o
b2oxztdtNEjtFNIwKUBczrSI229afeQCMp6P9nvdl988f91L5CJfmvNJYh8w0IYr+qz+3UTVWAs8
GzxhR6i1mtaUvD2dH4nvZP3Jf3p9SlOU4xmD9Xg4eSwik6QlwKxTczJEiNN++pwcFBTKGvlHnUl3
ZenlBLvUefQ2nhyW0kZHiQwhKW4nw7IJG+MzwbIWt0xzX4LS81VZUFR3IhMBjZlHWqr2Q/vu3Whf
kmPFC33sTNbWVepUAET2nXOqspyZSYgx+b0a4mpA62KGznNWxAH83LpALJT5UVN55I0ehaW8krhI
+nX1clx7lPubzwlxq6yX4YjZFfAoidhabtbcoV639EF7eMug8lYMY/gySqnoYo01emuBTlk0p5ix
nHdLcTNQTaV187lGrVAwbx4y20SGoxk2PtsTTZ7hDykHWuysrv8O8uRvFikEr16fQy0VHAQy1COp
G2q2+JjjINvevhJUC7zBCrnv6/dq9Ydbx6j25G7ddRMLlEojPpuJLiB1QEgbOniw2kEF8N/t/P2U
ZoCK8rmz1OpPbVCqBTO2OGLSidFfxliQ5gVAq9xpbU2cVJRAp+y69nmgDRvuArccHze7ieE2G3vI
aZfL7oubtgLab3o/pIU3BUp2+euYfepgwpQuNhKtf0sWe4B4r1jMJuTwhUqz1dq4pUFQgaVFw1GV
MEA4YsVJ856ePjqJ9pMkgWwu2rt2I57iUHBaDKDbiy9d0WjdvIRMjVXM00xabcgW/BlGVUt+lkXo
2PsRdwlGn8b7/UoRq5R6qI0PjTE8fLgAoJigvkLWWCSG0D67jxBXpKVAdlVtjqu0ICksitGRueFq
0SAzeZpMWU6rZnZDVMaAj//06UbgJZZBE/nBp+tKfSyVJ1agzhXcrK+VvS50SR1NPs0AodQ+BjeK
/Y/7954otbT3OG8+x1Pv6s3y5Y/KYlg1sG//C7CdgwMn8zJY/gIpKO9PdCoHIShJfa6761fti4e5
ull6HtYr582bMVF/jTu38slZ0YcLXMoTQmNsbVm9+yjAIc0HnWzav/a98X/406pMpOn28yYlYJAn
58Ry6bs4G7yU/MNpLg3bLfaSorY0MbKGMg+oXDcFNZQFz7TDUVuICIGU3Kjmz+1UudbDZuOEm+9f
HFESe7Y80DiUxRCbefB2bkwNFBK+GHSeFW5gGmvki/g9136u2FFTyaSDIq/D7mgJBuiIEF4iDuoC
Iudpt+2aIHdnevIYpol2t6su4zBteU9QxvqA9YSW1M6Xyx7kCZEsMyC1U8RaNqLLBxAwzVGGf4hE
nsy+gDk/ON5uOzdRpCudWmKSYre/UplG3YZk4F00lCZDy/xE0c/9YJD/3NJkYbM8ofPbh13OuBfH
1i8hY5fB37LXdCfKezpAtrImrhTl3SvakBYGUqLsNE9/zDMUQFpkZcYtiCxRUgKfh4wsHh1LUlOQ
RPcdptrKlXRyy7XBI/Q3+Vh61p5YwmzcNRjeCfdHn4KA3vR+PVfyH3KkXcJKvgeHzvAIZ9CFGeBS
s5OzWHCCmQ95h6pSivew7PnreShp/mQZxB3cI6QQnfByv7ngqHszuKh/wbGAZzCHC8VprbH/A3cg
Dvq91bgIHJHYQ7Lv02HMKjQgNFWCfv3dCbvZibPw3/EeKYpdaQu49mn26gPvhIZnEDtgGC/eITWL
OQqeULSc931SDL3YFJPVaNAIm+OAtWSyCSzq9Hfp2rNkXb72L3sZ3qaVACmHPs75vWCeBfeNO8xu
F5JuLaZpk0t+/7oGAmOtLVgBzTHAKrT4rwHYbnRUL9X27PwWF1eHSdDpOdMJAVlHXcO3v1amBuxu
XsO845txCt46+jezsibMvYYprqeipoK3lfV5KLYY4aX7LD0SbDJ7js5Vvr0V8s5YNLkz2+YrdryY
9dJIYIOQhZAWZcSCr7OLqjwIGn6hoaz7Epznd+qpdx418h2iOTmf5wB4p+N7NYtsU88Rd/Li8fgR
Xy0OOemEnSskodMfYtBSmIUNnsHuBxHFOAIYhkVGOYMzBgIojBAxZmK+Hd8dqyVoZTfZBlOXL4Yn
q3DDzI1HMyMpiow+chE803Kr3J2k8bjWss1bjUYhRAX7TyjSLzHI5NJseAn55eVTFUAbMou0196f
3bBmNm1RaqWCTZOOM621bnM4haLfqiwMSlKRzy4AqvtFxFUvt+6W1ejSYGT3skYrcJ+0DgbdKSnh
Wvsumi0FVc2XYuqj0X91UcAUdwH/YmPppPGVH1CPCnAC4o4E5sSCYWQ3IqyzBlLEAxHIEmKHZY5q
wSjlJPeIxufLUX2AKTJtEgbm85+FqNAvN1vCkMaB6dEDIf8lqQE1rPWV3Fi/4Y0IlVTiwJSvNhjG
7C66ipMCCxkBMA68DXnztUo1qEUY/sE8Rz56LeXXwkMqR8s3xR110Ea9hs6P5srnDit81hXc06OO
MDx0Wmd+oyW5vqOyLNFc27sMRtC92Kf52fmGwhqYiaco4JR8AUMrn4Ra8j1U+bs9E8U+EZDNM2YC
/rKRN1wxrDJ9DhyuAWFX+XRN1d9HACkdv8KURZzXPMo0Kn5NAfx3zFjf+3xbYneckhmoTRNmopyV
7sdbNdLmRkYAqena2mDFRBGTq0uq2YAi/FiXRUbDA2w1HFnmzwHMMW/l7gwvUZOWRHyd9nSWNMXF
PqxooEP6bFapsLY8ZNwzS1AxkhGzaxvtTRnNL6hXWg8oM0QiA8+p8AMrIoXlLMaD6spgctNgz7EN
ooUmKsZ1RBupu/hFaa9MtkeQu4Ernzk0jBNXYUpKjDutrzR/7VXIE6trondE8mV/eGpNv+ekzwS0
5VNej0lf6fAbTn8kzt+MB4pbqkLBlK3N3vNoBXE/FfP8f2cfjje4K4SkLeF6llI34rHVgPiS26jz
LwG+m5M69kfEvSnPa1yAAz9qID2SOeONPobaKNqCi246Fg2mMk3hCY7uBen1pr2bQ0QUig7kWFby
7OAoFny26DE09pzPx7oLVHTnD135Y6qPA4jXJJCBKl67r5CS+9mk4fqiFZ0m6LrVbTYHzFU0Lm4r
gYHQw/6NQ6NqkDAuYcoDDY8SSa+gYQ+GAhDGSwsMaa7ZXDenoZ1YTHGH/VypLSEYHqyX/FKwEiC0
RnHkFe1+qopLUEmfgcZHrGuKNyMh9/7LJgq0lYmQ28m4pFtsknMIlUJPjaxVIxOZgW7eEu3RgHZ8
vvqBp6NfjVfKrv2aTgq8oP1QMjasjw2qTGu+KUHq8OGJtPZPpECGkKuNjTJfBJ5W4sCVrUTTxADo
fidsKNekqCfLb263tdu8dKZVa1vaBpvz4mDF4F37mmoe97gXPePJb8WnhipS6baXOOzG5LuAZj54
uLHY9TOQh6Qw9xp6N3zQ1Umr4oayE11HiZuT2kBbN6qiIKw/icF7TfpbwjnwNA/RmmjseYs085jS
sttOBIi3jiVDzQ3DMZALQXN+ulywg/Sht2dG8y+za0xzDjfB8KDiQKRxHNUZaUOeKeTlFKodT0Va
e4ibdkG1mHuYSKOXJQMnGky/Kahu4R03ek3UIGLpfwCvwJclKgIUhj2TBBLmW+DQdz8Okubxzw/+
h2hq71KfJTKUMLywqcjef+6CdJPjqIsqku80OzhkqffVT/UDQn5bJY7QBvR8YpndWNRTQmu/oNSq
Z/dzESVH1FrsbyIhtTryL6lw1vdV6UCvlr7P4d4HcQzHe15Lm6rSo02lOTR3qlP7XR1sJjazThxz
XwfIHVoc6JaRnzBsEuvAWBCwdLki5fKMOybenX4NosAFkrlOalpbgYwMhvwecpufwR4tRMypQf9G
aBx1UzhA8h2VT0gYzHvH4SU1//2TWzwmuToM15BwkCWupgDD+f+fKz9yCJYrLTpK9y934BEvs1Je
oq5GLxSCSH6rdjH6l0HTm8/L0dtzVenE6O7zi5lxQMorjClD9VDD6p7nQMK1GWxBQ66HleahiZyn
pnOiSoijDTjDFgTh2HhDiPH9SbdMFYwpWgf4x+E9zyZ7+y7fN67l6DdlSAa61yZwzn4ZJsozOjB3
jcvth82jaGhgXuozQvBoCNsxRounu1bqCJGAzS4Tvv2z3HiI4hvvp7+IKaENHMDaEzM1zB+mTAnL
4li7YV6/Utj3LzykrLGKtR+ggf9pUZbqUnfryEAPI7Yk8o59wFJr1xRzvut/0fU2NC91AtFhW6fO
Dmcr6IrMe/35qRhqx3CC/jfMt1FNUhzOkFrtrQXq6szTBqnAeCUhqOzniWNoKrKBF1mxJUoarnhh
mpE538uMgGSO9xYMfrCjfBZEOj/hEPlT5gvARvx0fiUuLZTPN9BOuHzJ38K4yJPMhD1Of5sJN5o9
G5raRINGzib+PDwWRR+TCB5ca4eCYKBlslcmes9UiuIjwlYba7jmJwY8tmzFtKVHBMA9Z2oqOPbb
ApLBOaH2VKQBzZ0uGkZ7MQq0E/bWQaWS0SQuLyQrJirHT6gJdiszT+gQTRX01ZwFchDyef+EEAwQ
ivSz6CzHw00PGLGSYxZixroyopjtLMPiL5IKrJ7xbln2+ipMjwXoMdfxUblYrRXH2H9XDhRxycbk
0Ntb8w1zrNvBp3Ox7BpXMlWGTM3RaQ7knFq+TQmY4t7vROIpNdKEB3LnjOcV+/CbhrEYOHupqqR/
gSIDCF27+1iAsNSX6fD8/ajbWWJ+ojy9hEFBH0/7luAWsd2I9yWG4cYdAl/Ui1M3TQ2Sn7Mjbwtr
snQwP0fQk4N/xoVGgKLtwlJ9ymtgLG3MZTbs40TBwoGmZ05REvO1tznTd+V8+oZtb6Y57VT1fEdc
vOo1vTfYMFcdB5ZuLJY5qwddbUH4r2w2oRkNyWUtj8uEEy1smOg844W8MWM7Em5li8WzaHkJvyxq
F40yNTFrE7h+LeEsIKARFbuK1hvWi15hSw+D7aQsrhxij/qfhJAT+r2AO4VP7szC0iNFj0tDOYKu
kKf7XWnbRBGCNs1uP2iMmdkGJiMl4I9vmYYlF2Ud2Cz1JWrn0otFO+7JrVTofpe5DVQ95o1mv0zr
Hn2Q8NEPQQGQa195EsAb/v1DeCV/m/fJdzQVktQuEFV/7AcQ0wjeBRqMjxv9QkhscnrQXJcQ5njx
mP265332/CPY6vUkqcvK6WdPhpqBgEkRNDUN8U13DNV3BANnryGSR2S5OBdEN5s4Bz4KGEJI6OlK
uGoStoxbwhlPKdnQIwsMZ3g9tFIb9fKd7co2qyhx4JdlUTsid4m4luYwA1APGhopFzUgR688iAUj
lekqL0cg1Uq5HiGESKtWx6WHnARVS7jAT8R+rCKm0j5TZmlzkryQRGH4CmRZp+HCP6qDQTIhCWFK
4NjtUtxtw2lFIt5r0YJ/MoXEvNsLC3kyXZd3RXs/R1d/167Bu3V6o5X1hKs85yu2wxaSuHrJ3N+E
4wVBGzBQhppZWhV0mlSvitB0w65xQfzBLvoNHlahPURLFIL5eddoL7FE8Ks2sIvcSgDbiFhS9Hyt
9Y1GSm+WB5I1I7b6qNZrsIuTWUvSZBlGWWQ2SGCnGu0acrzhih1lAqpCYzKP64yStfe6W0Ec5r8z
D/nq9HKQ/d77b6ZQJgIYG5rwsytqq3mv9C8syfqVgTTYEOzIihxxxaXJomCUmtOZ5GOxVHiinp19
YNjB2kQfi8YYootvfucbSJKW585rSpgFF0b97PSysL6G0Ho4YAFPSPXOqH+AKLFseh/QEzt3s7HC
Bj+Q102Kgne9DR89y1sHFmpJDpxGk/0/el1/wQYqQDBu+b8iMGgrWL6bSGCHBpYkCRTvclaIvhEJ
BF3LSQ4Nd6DcfaqhrGtmxNi3mOZZhKEgiViWASyGaBKj8HqY02PGwz0z9EZvCbA0bzZNHnReS7wz
vr5c3WwQ7gicMagDj01bbXcEpMHufybIMpBSEoll23Om7dTZm120qG8Zz9INw5hKx0u/+WII9qac
OWZE+1GOhAsEj0TykU3cbwyBy8rAeg1Sy50ornQGAuqD+B8fgeeA9JFNmV3z60uEqh0Vv5UKFJrw
yVo1ZJ/iYB6ifNjOZLOVRXqiODJPPsHq0QeErkkvicmBKpuapOYdKMLwnIuMWeAjbwoH2IdSP0HO
7sGfe2pIzW4zr8QRhOrg7UpKz/6KuKc7CVSjU4NfOLTmSe+47SUglIFfdvNIWDYXNvniJA3guvuD
YdDBxm1Ac3Lfcqb4xjE5EmiPoCsjrValOmb8BZv8YMGihVKx8NTsrGeM0S7z9RZvTmiOhAXvHMlp
knqOly9WxjhQfG9PamVv6uPfE8XquRwvihT9/yL7d2SP6bYKwBg4h0s6VqbAHtsE05yTcm8ORZCz
SGiPQcryPiffI47E/3dwiQv5ONijnK5aS4h1qOBCRa+vmDuV5tHvmnEgA03HV5z6xSuejx5LMyYs
RhNwdF1SLphKA9gNWWFBFUAI3a9OO1FKOC/5hq7qaVzLMxpf1P5lBMkooWPc6uN0uWXn5RibMl4O
M3AtJUVdt0DGxmUhyULDsa5VycS6/J1mOrlUc1kbKsIaw2AZNM1Wo++3OuR7ntCk8EtcjAf7rc9h
A0g/RFM2iphD2UjigxxFqgZ2C44SA0E9dH2IuA7+9smqQ14FvH3uX7Hz4Uf4NiD1e8sXjt5UZaIq
D21+O0LUSFo3ojXZ/EQ01dYKrrp9JsXfc0hwGA6qGRHFSIqBs5OAQrkQW4+xTz8H+aptOhJZyI0n
jaVirp+v63ndOB5fPDpkOHCb50cpIpqQIq2jiUi3DCaGRcb4vKt6gPxfFdj/va2ds2GpaLbHaUUq
qc2CfOFCE3JqZU5iSVVSH/HX3GbN6Vcvz8iRxrS/u5DAkcR8sW6k1L6Y57YlI5sBqy2o4TtEVq/7
57P/xdiiSNJ3+NSiIYdFOy3jetzQDvBXLzT+KWAjiS7aRFYVcb5xn5mY6UXLwN7K69v+6zJrqJBY
9EPm7lQo4Yy5f6J/AbhDsQAF43hel1nqh4CtJun9iLk6r+4gQJDERG2zC79vBrNwtPbf7r1osTqT
jmQNFneU6n6RPmrbrCHWx5cebeoA528SiwOkqTPcBlKzE5G0Da5PeN5/3/gtWdnDJQOioraDFNt2
1/qhBav6f7D4bsK7LOKYWGW6DPdXzaN/DIOuBA10IA6Re6vwL4FihGJSOdiPfvuEjqw1aHVyduoY
4+414nf+YniMi0CM8hpbAVopfgjBGMX5dnYnEwdvJ2VHv5qw2w5ApH4tn5Q+WtLL3pf71lBUFiTE
9eezIXhSQVxQUQQzCRWwlPEROHJFRfz3TXHzpw5GZGDwCSjtM/IX8qZ1i6ZDgR30/FLfGNXWztbU
XSWSbIi2v1tfE7bsGweJmVMgbj5nx4M0Rnr1NT4+NhX3/GdfN1A=
`protect end_protected
