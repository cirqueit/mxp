��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l���OLkr��K(��j¢d�m�iK�b!*��[��?��x{�SGb��5�My������kWu����!dα���������g�������w��
�W�GŃ7 2*�s���1���;�|�⓽��X��B�P�k1�"�� XH�Ñ�	n@�<�){�����}��J_9�ٖ�u2��>$0w?�"��Xʒ��=�7���>�r��b<�	9�ĳ�T�5,[��B�������3%f�%��-.�7|=Kk?y����e��%��2�n	��\h�O?�݋_;<[�1��3��K`�DtT��ԳcF�mQ��̻]P����X
��X��OP<B< H��U���m�6��l���?����/z�pe�;���.F؜����R7"U���L}b`_�Jօ��\�f�,����I����w#'!s�f�����oW͓�!Rj� �M�MV�3��IY��;�$L3�K<���,J鈆oMX�͌x%�7:Jkb�eyȸ�ă��γ�I�	���|FUN%ϚGW���B��>7L�t߮�͂���QG��-�,QQc�n�I�U_��R�oz�ڼ��xz$2����}Z��t���;��o�[Qw��k�u��j�S����A}�p3Y����lu�Za>�h{�?�ױQ�<,��}���n�\�� ��U��ݵ���e0�.3N�}!+`�br�/��K$$�0q�-�zgZK1�^��Sݷ��F���Jl��A�xE�k�lW�M������FJ�#�+�M������cێ���P��^O��P-<|f���;�m"��n���Q �sM�97�bߴ��DĐ�^s5�
FK���]+#(�E��I��};C1^��P73OY���W��.��5�dJ���|���"���K�H����}�� d��:����	��	�aWzc�,G5�������+���M����~��O���B�bj�������j�ԉ%|fr[��ӻ�?Up�G��YO�����a�I���t��N�̵]���E�/*5�S�
v<Gz�q(��9���˧-��Z��2{=����X5��>���v⢯��O��:P�%Ѷ�&�;�ۻ�".V�̚�;���k{Xl��+�~]��?��TOK�l ��Rf#d�:%A+ʹ�|k}�M�ӑ��Y�C:AK�tp�r����2`��-��cR������#���r�E��)ο'����|��.��Hf>��%�R*W�M��i�4�{��q���Ok�¬�4��-��[��q�V8���+���X�G��گ<���k���/A���Y9���e֦�����r>�|p(
�or�i�J(�'�%��o�����/M9�V��P�V·�����,2�C������4�R^-�d>���Xr�(�u�憤��-dʻ����~��C)���#"��0���˓�F�j売V6������gf�9���q�Z2U�h�i����*ϊ|�-Y�_�N�k�D5N,�1"���ϋ��O����=G)�j�Y W}^:0�>m�R��P_Y��j�W\ t�@Џ�f�|&�V5����hm�nP��R�T��ڜ��^5�O�I�N	��ϱ�m�t�Y�v=ɽ�K��<q��=��B�I��ڞ���T�"/��ܝ�
�bզ��GA�e�"�h��S�n�g����1��n^�)�h@2ol0A`��N���Ga�ebYŢ���zGcmŞ����ӺE�*M��OF��T/�Gwjt�F��*A���6o�LO��d�.�1�i���1�T@	��b�D���8(񝋦3.
��
�1.�Ŀv2�9�;��e�.��	2�y����8�[��o���.��,=t]q�w��5т#�j����}z�I�85;����!5�R��O����C�?[<=�UO�q��J�q(�	`�K�e� �!�[�����;J�W�H�a��j�����x�ǐZ�78��\u\��8��<�:W/�`hQ�L�żػ7���.�" �x�gr�TKtLdl!
�Џ�Lҹ���l_H|�%I���>����۪9LrvL �U<�<jǥ�M"!��&]/񒢟�4�MK��o���Z�f./_���	p�s��&G��2�C�,�t�툡�{�6g��j�o�~�睆�@UB}h�/�D
s���B�����E��
	�HCK�Y*GfR��"���a���&���J�k�(��b��л�0ZMga4k�H��ؤ�\�P�ε��0��GA@*�����1��o��i`BAՉ�eL�%��Է_�2ц���v�$'��$�����50�)Y`�6�@�8N/��L�X�>��j�}l����~�/5���2�Y�?��ね�]�-��G+4耨��}�~�<|���Í76�u��ֲ��7W����Yn���T���z{��w�ɶ�3!��a�l�n���*.L�h�������q�����M�0e/�b�'z�P/��� �g��xz�d���%2o�y!oi�ދ+id���M�2̱؃�~Y$-��p�b���f�L�O��)�B��VQ���Z�]k���Dw�1�([�^�e0�\�������jH�r�\r'�j��xҙ��=m���v�˛�!�H4O
�,�P��K��$�lW#ڶ����c[�^5�D��<��N��R��QU���V~���)?P�c:���S�+���+P������ˈ�^�e��ԓ1��.�-)'�<�?��!�G�-R�W���{ȣ�0r����8�m��s���t��J�q���^��p<�~��;�sqN�W��r�9^_Pl6�|�&� ixt��Q	Q�e5y�~ĵ�,�����Ȝ��oqvH���`���@CP����8ߙ2�Y��\n��ƁP3�J}�"䕱#AzÅ�c���p�?�n;"�Y{`ϰ�}�b�����i�Fc,Ӌ¾;d�l{|�S;R�W3V^���=_�:�i$�73?7Ҵ4n?�b%�j���5%�q�J�X��sE�"v��"��e`Oܸ8�$�";d�+����󋲘��
-`TY�	h�Ɏ׎�i ��\S��֭ܳ+P����W9|G]�N
��L�C*o�g��Ȓ_�ڧ�=�ق+k�%�����¿,����]�e\���(S�)�).U�㶷m�q�
����OB�{6\6�Q>�+�x��^)��rA�:���r3�l�bg�P��S�y��o4�r�{�D�0���Ϊ��/����7�-������t4��(�5�e��YR ��QQ�yVS��\�If�Vo#�?@��2���Y_q�fl�M��9dV�2��t�ʏ&7��<1�}܃��<VA�J��
r�%��i0���)�@�x�����E�i(������{69-`x��Ir����FҼ?����;h��haȨt��v���}�����V�=�g��o Ȋ�R�3�!�FK��2z�ݪ-FWg��u蜓9x�!W�z����K��n�7��{����_��E�f'L?�_�D�(J��N���:6�B��������n�݂�cȟ� :�a�Uq�����u������4�J�m�OC�n�ڼ6�Y��\�?��@�