`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12192)
`protect data_block
yOJMhS+Gge+TxEskTvRM2r9ZpEa8Ovh1o3nQJWPQCmiLXPOZJ67ft9Q+nT+HJCTJZkWNcTjDIsbI
PzB0PgSrOEe1eFLT3lOuugNmNYWMAYDhzWPeB7odYEk9Fw+48PLxwLuGeaqX9o8XXGBuQOyBFHm3
h1nAfM2XCEWSki2hY/2OJ5W3g7/q0GciyYFLHMJz/dhRAyWfM7eoABgdbKOlUI5uZu42p2xMl8sa
deGzjiRmFqB0HwYN9M56SsBWqI1Zn2dg5Nt6jiNcE0anjt7ABxq0QzPLMXS9ROTc8KiG6TmXvYo2
Kc1QWhY43PPmIjuD+PpFd4zvH7YZ5f3rS+X7gbioG/WQZPWG1gDDOmb4MnmuGp1PElxB7tYOp6gG
v3+TotcbQRGohruyUGhBZw/nrOUv8rUm8YKwTcPYWtrXDblqLoq8KSKOm9eBHYhUkg21lMMblKai
vjA4idoBeCHeCXNJNcYRXybvLP49olW8meYFL5KRcNP2vIoSPQ61CbTN8dHqlqmuDVL/h4yZrU0K
wOS1Ia2g2N/+c6ELBdrNI3JzMSPQtzaTn3lgM7tCgCPh4C2m2AcptQ5JkaTU02o+wJhJHK6javSJ
nVI/xVh7r5wm97qVjQwJpov3Sdp0bG7xuXmgyy5dSyCGs1Xq6bSIDGSWe93T9NYn68Lu4GKm+ZzW
sy5oJm5U3YqN2zCGzceQbRL/mYFz2jTxgNuRUMMPRC0ivuYzi1LA/c/TwT18tlWcaqiWl9aTSJui
m+iRBCdT6cNE3+LkVz8r0rMPmRMbvpzf8JR6oprmuUiyykxczz9Sm7kv6Bm1dFYGpJ6bPJO1vMw2
wBJJykiDkjtQRKLCq5jp5KW2mPjaE3n45IvXOHyCWje0TNw8WzjCOQyIUXe1q+Aiw/f/PT0zzSKr
fKgyw8TP7B8ki7d4AbnOz5J1WnFUd8dzJN/x6b1sOz2T+beS4Q/3G97GdlDRlwch1WdLXS9vtckE
nDuuviG9kXd1BNtnVFOgOvVOqWfoelF04ROUQsVWHy162EwA0q2YAZDV1SZCM9/D342t9rQJkUXO
E1ZF2QBi4yNUSHOMGEbFpOs/2AbysQuzfFZtpUh4acar/5uTseW7/T6c/zMVr8PsegVTdv7+NeZk
hioomEX52+tquOw4hhzR7pNbIc2dkVjhASzxvBo+8WCS9LefEqSKKnlRHQeDEevpgm/lzA3Ra+hN
stM0d9kuRTaMA0z41ygWnEsKB+ApQ9io9oFjZUc4jy5XQvzFBkgLNdvYwj9Q6TGUiQEUVxFm6M4X
F8IHnySiPdIZenEB0Gss9TzWv15xuCy83Q0b8Eq5zBzfA/iNPknc3UfcXmIwjUPfNjPR/xku6xcD
zyE+S9GROM3gBC9aFoJbViQt3EfUvNkBp0d04d20kdCv0k1eWGOohyTtHIKzHyMBvfzGUdD0JPEs
OtSSH5FllrfSa8swTd5BdlfRkEDVtl5Ie6dTx9llx/0x53e5HbNZ9PvAnwyMjfhAVC7/EaLkgS81
QAztyVCbuw3/0RkNc+hZtaEAHKERBLMlrJWnPD1xcCVxjhkusxJwe639MgjE9EHO1cpOESGcQ4Fq
FREVgaEhEwexCQ9EteuGQixY+8uNyjUIBExbhRAus1IRH74tg5lNOHqRXWtYSeiTHYPUZeRDP1yo
UpoHXhATTT0DQiCDsedi0ycZCPrG2ugedBSe5hI6Eu+Giyenw5Le3zGWD+3e8fHQxhX9uFQlmuaj
+CFNMS1XBdamxp4p8rrsj5SR/f+wESHRG6ggWdvlU47oBXvxbYW/ABrrPWof49s+6EFniqvWS0Y/
PhCl11UDL/mdGIWh+9BbvXg6aiaQx779YA2qXgYRzSOtO4K+g/SIMFk/oHshLBc+p/CBtrxhbkkp
DzaNaz8uLt94bm0E+ANH+jqlmkEE7PyJzojBjkio/Wg3NBH/dO0K6ReUryB5loAVaylYZwv7kKCx
pBA5PPaSLzyEL+xVz5xGl8ffF0rCI1bjMmplkMCsa/KkLgTqMGaBf2e1wLuszzLbgDBRHgjsX62n
26rOjloA+uciIMZ3ac2FOD2XLgCHwBy7ioQQJioOxyI9FTU6Whe9U+MbyqT7wzxtxCO/mrsJ9pVp
g448RXOmswhc4WiiTmH/5FuGewDjTudagPY6gHdLNyUl5UI0Q9l+RDwxZ1PrAzeysK1mtW6o5BN9
EJCBlnbou6ZEfXzxasbZVm89tcbig9hZrsajzUJhQ9SnAPCJt6oO1vBtfp82t1f9EBdUOJbVTGsS
hv3ZrecxLcX/NA8jtT+N+zJTBGRqKEcKg1GmCdWEQ0W2AGHs1MBmIrDL3ROvCiAiepJo7VEiuLuw
U1UGlrXHIE2JLriSE+NxDqRHqu7HNRPWIN2FkG+aLKvU/BgRoZDfZP+nrHwynIJRmF5CutdXSkcc
1yipdR7jUY4hsrj0U/SWc0g34orczMPwzCA/nVkysGFE6PcMFIB7OwCavG879mQsHYoIH9JHsFYH
cyRp3cXBYP6I4kquAP12ScRyiW9AN7gAzrv3/GwexMLQ+AfaHuP7/XKwJ+WHivRvx9ayrTLNLSbX
h8P0/e8u8KVXfXpaXwrQDtz0UV5oOCMckWgOjpmJy35lSOooedWpqhmZ6Y+SaeRA2z7ormX1i4v0
lQNEeztEUG6XpOi1RENc0gJqDoZCCQL3Mgv2ZWg4jmqheK+sJrruxetfE3t8rGoGXMOuYwzK/miJ
7cp1J/vojTDdfuj11nKWUv8R9Hw+1jhUWMt9vGC93G/vHoIqTaWM2FyqdsDz/Da0gIGk1Ae5HEKS
7OHQ6hjNdasUKDvDIb7rMPiimkBlAYxN1xQ/iNJxgGpOptDLqQeMRBHiZaVS3Tx6Hj6odelowIBh
oEw0Lc4a2MaVRQWHKSMa4KHQQjFSkCHZoGubTGIWyZISvE2azaOEgxECuSdZZWBGl9XtcvDBRPpD
KgYP47Bs3fyyJiB1mqZ3nmZWdVdw62eXx3gnzJCQogpaw7iB8pPpq9ktMMrurkKwFPk0d1dN1rHG
MmYBBuaQ6Ng3+4cGwSWxMecrWQmhzdCysK3poyb3yszloPn2ZJNt3voqeoqSDBEcFRZHf6WqUY0Z
RvbG7OrC0FzfLRcqKeYLRQ8rpma4oKnPpEfdT4jiWKfjxb0LUaVJHXVRcPnfmajefu97X9XSGe/i
jAqdYXZ6fnoi6kl34tsGsj1IqQHK9Y8AicYQv2kRr7CVEnJsz17KY4zeScHRZ+rJoU6A63bZWm6V
pMuxT6PFXDdavBwoe/qdsdloRDlOElkAZjg44b6WdcFJzlOG9Or1Txl5bs36gDHOzPLoaxPTWCF8
n7BufSwwrQX241QyKo2OBdMn6i5rv2RylamL4rZkUgCFcsNQNg+38k5+rQ5TWHvB3kh2TD25DhPB
Nr6E8FvUndNSg7oruMmjEMEPGeYpUAS2yi1eXGBSb7IYGoQDNB86nKHgCwmfnj8V9w2FzZ7HrLFF
eX3D0yUldSvTEoysaI6ECD2v+sr62K/4hQVtC/lTtr8VyGwVM8Nv4LRrTFOIjGqFXHmjnbpzkMRs
muZ7b1skSv80VHAUJZWmDrzNMUgMNTBfq/WpeGs173ubtDJW3Q2xcmPUTIifyz2xxO2vagwXel50
NQ/Wq0yhd95dr8YP6wJrjJ0eD+UEeTVkoWKu09O9YgU7uPXT8Vd3ss7whMbK4UEOKhFUKCEy32WM
AzDtLmCHyA7vloRGbqq6nvSAOs5Uf7IA1mPOVSaO+Epxwk5GRBg+4YRF8XN55Hjvtjq7ywIbg76I
/FxkD6sJ6cTGmxNV9gARmV2OIIt9FOLiqAxVuLrFKXKlHOdj9GwCekzJBTe3cWoa0JtysvGUe1jJ
lH9jC0gi0CjRcACii3TMuNz4ET4/ceE9kqOyOtW5Yu4CxkRqEPZrjWtRkDLBH0A3mZNHFrLJXIav
wXyjOHURYlMI2YSkE1zdTHHQHDqi+wMpH+N8G7LRZVIM7jXNxUugETZZcLjJoa2SY/heoOBC7rxX
tZNrNVrinUbr6ttRkZFyPIJMv/OerH3HKg7KtmOJPeDSPbLYRcdMwMuU2y+kQz7pwPUvvcqpcCuT
kuSNni7vOabqZWFET3bSxAObifqxZKxWFh7XdrzsLZMMWDy4yK+6diKnzDrhKT4ZU8wG7k2DDIhN
ONYPkEtt4ggmakAG0SwbgiA490iPoUAMU7vEx26arkEytqJ1kO3J2BPfPNwZ+aAhtSfgt64NMBkt
6swggxjAPxcwBrNiMIRVebDS92ChL5O064YjRdM0nj77zm/G48yQLHl5V2o6HjQ3TePrjCEOuShx
GsLXfaJdFyVhvE5o/HgOlL3CR8tSZWOozfnTyOQB5A4lfcmORp0GqK0XDr7h2/R4qUmw60woTcFo
OrSIjw1Ha/LJamwnu7bBcC1PMNu795PE/eSEckvIuRKQN/EX9d7Gfxiwm8vGmHvDuCBENVOQQnxc
UZCUG/Vc7rVeIQ3n7TRbNDfY0V3IDDuusbyd3ufZoh3BcYrw994VpiiTYxt+H7Fzw552c5tBkyWZ
YvBTCcE/PTarmL7Ref6b6NbUCAXtCjcvzRUZmoz2v0CivQil2Y+bDtsf4IY96mQ+iR1+UBqItQX2
JZoB+jI3U6qfPpWqMYxVGX0rJddLCW10VjkmPNODIA2GChtog/jm0i2n+RTSXnR0KSIOXhlJbPHo
5xgtikXEI1JzUgaFsCB0yDoXAcYo/p/jdSoHFAs4ulCkqslaGhZ1k3acjxpvzsheTu7I9wcGurDK
mpYKUI99JBV8qP2AFyYhfhGPqsxeo6hf3NxmyROAEvus+Y89L1YfGmuTh15wuH53nFkJOqslcuDX
dFQHRfcvZcvwCQNF2gkRuYuESkf0jgFDNOzBShvjt08AHqlac0B8tXGIgUJJoLEiSM27drwGynEW
Ad6md6VgcEjoK5lkgMxMGwBT5lp1FPb1WjscoPUOSN1EKOrlRMzFPvVfpEyjJjHBIcX2OTfgafVE
WibAtyzxsnDLogzTPS5dt6UFzB2buhonM5cN0dlJxzM+HxfZ4ezjsexzM0P3Bd9Pwy/pajIzv224
Ecn3WXoYNNyTVbq+AxUH6bemqPcPEhGvDf2TmJEk/DuF8q93DUXWZcO2Svv8owkZieUkTdAIkxJE
tqBcIHmOS+UbPqtrYr81cUW8Hp9wkXELkP57+5qOc85pABsNvr98kCx+IHELlZf3IJz94REfWo1M
D4eanMlrLjaVXfXB+VWBCV1hjQ2nHB6YE4V9Q5lHadu6OXFZrF8685I8QUEua1e4k8/GeJNFFMwB
y676GpdfRwWdJSUGMpgBbbhyP26dFrHE9u6RjzUFOwN/gumjhn9TrlxvCrN3mWVeBGLfV2khrBMQ
akVPIy2SGqa6OGtURhmlmnvN3oOdqc/WZ4RNO9wvAZ1prNGyoAdYEiLAMKs8LuLrazj3SLVu/Vpw
ylQ2uqhAtxnU0MVsZC2berS8cOngAETS1rAUQr1I/wE9TqeyU9oPeYlrUysVnb/XfOKkXt8B6hkk
+pEUuJCvz18fS579EHO1loYimLDBRxQI7Fk+HkgLx0Beq9OD13QCvaCBC25jcveoXEuWu2gHXK1s
/PmSe2UJC8juYKuXfK2UAk24+AMkPB02jSLHrZ/dnA9/vpERNc4I1aPfB8BND8Qe8ZXtz3sQKqgp
liYKXkAU0PzGVEb9lTN1xPbEbMCF0qN3lOjKoM+r29QixDtdxUfNCXG8MNMi68ewiRGB1Rc72Sjv
9cQXtlSpvVtOlke5hCiuzaKOx0yC9gwEhPJQtj5IKX6Kxj3AMbkUYI5yurNVfEW3G7TEZd3CFmjA
OXVkPucs/byCzMGlkQEV30RSyuQZ0EJBPmHJKCtiJgTfj+goiHTHEcCiJCIhyN87aymrrbZQKw8G
+XBFz5iI5KbaiAdrC6iJvHFiEM0M4Gl4EnoYApOI4gG+musDmoFet1mUWmEVxwBohsh9Xu3xpyCH
1cJUMeepxcCwr0AYRsbfrQV+4LLz4PhU6+IqvuD6UXtwFTJL3oX2heARaiaHS1exj5zc18aTeJSQ
sv/eBnSggA+z/frAQq+8Ph28EIA5r8DGVe6RUSnZ37Rs4OgwGdSwqtUMq8bnqf1yL7dxcwQNsQG9
aKM8jU1CYHGEQjXXcrowQCJxhIbVr0iuhr8yyMc7F50x2ev6L98Bg1RT2ZWMTj77ymWbsA+/Kvz4
FamhuL4dI4szlkk0TwvrFHinw5cRsSW5nlw6NItL7wFFxI6aIm/5KQjy5YuFcrg+/2tWpUvSbXfx
H5Mvjapnyasa6olXfttDIePgWqLsEMbtKZXFFIjRk5O46N/Bt4V2LQvuQIouWW26v/VGeFBe14iR
FLyD/EhkaTtXqQcYrKvquEVcDrvd0AMwr7hrBtjavhV6lRFQYF0a5PgRQi5nRJUQP0bWKMfRHnok
KqDE/f3mT1nTlaF+XYaAWWHD7HKuD36Yr/bKbRQ5cy09s6XcFk71sA8hZnOesgXHS0jAP0uphzqN
eeEoYdHmODlqD7Fr0Ew+hEuKGo4t2A+JO5rrspwfDAIcMBV7Daws6dm58nER6FTYjS+ltS9k4u0F
I9+sPeaSPpLs76jS4N++YHJHeI9ADkyYKcejWqvDXaAfCmA7U/Ax4F2gFBiN7+08HdeKJ5b0XR7+
BecIVulkx0E+w32Y9xQsHU7jyLXsnxY/Z80V4fUN4cYGIFA+bQ2kOEpU9wJC7fEULAdKqoQBaDWo
+dwee3qY/M1Rbtv1PTACdYnYRIDUnsYjGOiXPnHn05n5QYsCbeHILqYy8YiG1HPMpO07eqSyLWJK
dey+vHOkcn/9iQNUZkWHimXAgjgXO3siR8Fa6rK1dGCKWPvCUXe2yDixv6vCFeokY8TSEM4pW6O2
Jau9qG0RjeWWOM/PQ2sVQKuMu7TZxC4wHKgYoXvRRZt2JRtXKohqWLYVEjlBnRa6vQR+YiTM+gam
cuWdfl0KYFN6WAC3zqn2glnU2nxQC+akd45UQHHtNVTg5v9acTfItz/WgiBu2xX9jZx+mIjwFi2z
qiqmA2B8QTwltRpHUQla4rvaVsugFc1NDAo5WVnnokoEzoAWtm/3/+GKG9zV6M4zqvVwU01pNzvE
0IDNqlUisKBi/mwafJQJWyUouMrmVsJa3wVawHhr6l2BufEhi1KQxQQ3M8/+X3+wHT3Tb7zWO9JJ
T7EEsgY6yDO/u456P8i7YvNObGCAsDFNC/MTxrH5NSJzRxMv4ZxPeIHJOENniEu3VIvwOb+mN68D
14MLrFhZBokbSZnSue78MmyVvEnFnqwBv6UJ1gUnvfQhFM3IjZo0GMNOVo/A9XnTyUA6HKxn+UEV
miSLSQpbAM5NY8syDWMf53yJQ2ZQ99sMs2B9dMatd8a17pgC+L9DKRhp9SegrNvt/u4/HVqCTSCN
csKQpi4eRS5cD734pwNEut89CB/ZZZ39lqP74aN2+mgWatDibcf2zwMIrbVM26sgQH3bf5+Iy7J4
HKN++M2SdkBb5koiXiIF0CEtiIYPTnhXuseTgHRbBHuJ2lgzO0cwSkYM/AW8EvcORWSV4oxJELrt
ZLS+BWTj5e3MsHxLA3aPcD8Ctvai50ubeKCkaQ4tOMHCQSu266OMyN0bHhvx6NSD8p5B9Q2De8Dy
CSyL27tsx2hKXGlR5VgrbBXxwg04T3PcGctkPTBNk/1Ophs/JWPbryw5dPBXsEVSsyYJzutGHrXN
sm3UtKeImhnOqjxydt+7KVWm0PJDs0hOWLOEhdJvXMj0vlxB3uI93zn5GcvPjI3PiJh4mN/qFgXV
pTSHMAGA+raEdhky0j8Ngyh+MYejv4dSAnG0xZflwaCwhKs+KfhdnnR+j8KEdU7T5gWim2Z2qqzW
WJ593aa3I+zaYMHGmI5eRF9ijd7zIepwWxNoAI7arD6rKMMjJgE5qAVge44xyyb0Tj/OWsxrGR0K
0UI+JpB4NrnV3sq7tUvRNsclKJIO4dVSkLDbDkXj4LEUahIfsX8NXVdlpvq/+iGTBRvcTGXuvZfV
jxxwU1nnts8do7Pw336Ky0WTHB4X2ptsXrcGG7gli0hcuGZa+t/U0t1J5xDhC8YFe7jz43h8yn70
bCbjhrCz53VwCQOqyHMPxFrNQOldlvr+Z3UHv8fMriVaLFX7OTzwH77mcyfsUp5HdDkcYnY8Hw1L
d51r5fvlE8dt6CgCwou0I9jUF6vp9EcjbOo3Qkd+2vgMEuexVG1VZie6h1gxR90UFstzCgH0/FQa
tcQ4LagDFnjZNlPfFbqiTwwW3VqGo6AkZYjG2JHubS2CfvmP8LhxQDtEY0z8NEuA3044OXkQPaBV
USppfOMkaguKEF/nH7z36ZCvNY7VQ9eiY8t5pdjTGY26i4fzK2HrOTmjRiMRGTKS19oOyb7WzNbS
80l9vTx52GJj3KbUWVsnnGMUpQ5QPEPpqjlXYwcUCHnT6IcpiGVkzh0qh78sDfPyYOEqYFux+WS2
jVksOEsPWAOLs3jYdJhlY5jS47649vhC2+BBSBdIXIL//P8DSyXn/8jF0FOziJdiUJqpPjg2yrOX
PUa4bOcNBoo3w2p6WHr3gKGISuSVAQ/QzSNN++NaYnerNOdeUuk+pr6PTFF6datrjkka7eENsLIE
HgpHxPwRHyfO1an2Jct990dpyMW7ZaMiIJGFdA8PET/wNisPViUh5/P3gQxi3nAtuyNOzpy2gXid
xv6hun1fdoPKwZt3GBdFsBabghxXVkaDQYqTCvO053JRHdmsenaMDcIrg41DLfIDWVo4D7RoPlJD
B0zHkgchZt/Z0NNRN8B6scHI3o6KXC2izsKcVwcSVuE3tTahwZW0p7b9plVPwQ/gSIId1f5UYD2X
QPCnY0kLcbE/DP0VTmov6KktveJqQAAz9S/egEr9BwWqe1usJLyWUqHEREH8A2SnlqKgsJGyLKt6
WRkO//0MgVrYFidBlJuMRSZCGOlmQsgnZDS/vtyebntKxlBVe8u/1yeuZy2sQUOi0NDs+0IXG8Qb
uTo6avmwuX9+U2KzsIa03l0MZcVJ2Z/MBTk1YxKR8GFUjdkTa/4GHkvXRo3YUgd3PjVWQfADG+qM
KiY0yLdlpWeSB/Hu93E4/lM9JfrFl4w2Pozqhxd7WYq+jvw5QQGSk6kkuu3DvxNAYB02H9Yw0XZU
xxZ9ZlUGe062ii13rz5UtLNjmp1X7aYRuohzMU6I8f5lX3lmaoU8dC9q1RvroPy7esJLwU1SIWbV
Vl3RfqKfSG6atMczSuZnm5EenYYWChH4r4LswUd8CGI3ecYy3LTWcyHY3s34RusZn2GJ61A9cFrz
V8AyrXchhei3m6921slYemDA6BB9DxEc3d65OZETyaOSCOHGcYNXYOr5eKcXkwbDR4AoK6/77sni
3Gz5FHhgSWJA1b2w5i5o5G99qNidJvWq2dpyjBPkvHQdCWJL0nfW03tfRgzaNkDrC61rKnFUqRU4
2oAx2XY2Kyr0b7TpJcG73LM7/0HtbRKcuXLzMiNIZcUcZGMEVhqsy7W98h8XsYTrGcFbXqtiwXke
yu3usTJ55aj0goPcMWgoq6i6yIFiwQsICpiDKtZ1nkMihwyl3jVM34PQ1i/LQxURytLXUDGVt6ET
T2Ng5gN8JhRZyAePA3Hw3Dcr7s1ou9QOWtJC5eAtKVoBOhOvTa3xFGU3E39LmSrunTNNlZhpzCvx
QJ59DiXnWWP/v6LIrDvCK706orO08ZlksNmi6s4XCXJm27SwInwA8bBc3HVmXXoL87hKa/HDh6eN
QODac8OXdTBErPRxerI3kxVCQTc3iijmtWmPBh1RZmk/rKYymCsJ7CjLydRQkm+UtpJ74WdAbG2G
DMqr8Yko5+6xDjYVJtZQXSYi3qHAVUNcVfko8VwapclHDYDW5nu4bZnYynAxjHe7zrOuBugolnnk
QYamfRx88ies7V0Adk7SdtsGjEa+pklZiRYHSUeJKsdQ+QvTkfrpxc/beFJZDLOcsEgI8l4IDiM5
IACwltGGy+06PygIG5fg9Vvpxab3FsOM3k86h7D1V7t1C/cnQkPLDZ3cCxm9E/QCzAyRuy3rG2VK
LlXqMzeiagZ8ghTTUPMnVAElJnIjHmy5TuCTfs6rLo5Nw29kAFEHCFw2BLOixQQWJvdz5HSxclOm
NgrWGHSe2+mLClC3ArRkeO/18aI9ajcfueYl3QoLO1dZw7oAtuv0SQ7SOtIbLUEMfcLnZAc3+fMu
rc1zp1/ZMoBR98D4cIASoJ3wcUXsD/Tk7CP303+rE+fjoqTG9lTq0Wkbkc6GzyR365VLlPETsUbc
CYDKjSv4KgAXgdMoz/jUDXHDhrRgyqcx/Zoq1g2gXlxMhLkLcDtvY1Uq4H6JmhWw1kdjM+ACh2kp
spa5cb5ncdvcEnEZaoOFYKkbOJgYH2XEljoCPP7q/kgGisi1k2VaKgFPGVJBq2Vg6tyDcQTlJW0o
31/+tnDh4KHFTBqppLuFUB/q3YxCMGXlDgQtip0n3CFMLibKqv7+kSIP+9NLpSpimKCoV+7fFYjb
YxX1ypdtWGj0nyAf56CXl4foVRFWOcCBJYuf17rSmSdhzkLmrZlEfHHy98JngOnffUHqOR64K8cq
Vmd206K/TUL/LhcZoqPVw7MMCZ9MStUmD93lMmDsoRAOqdrMw7taJFPBLqLY5AYck+YhsaLZoJB6
ZDTS3TtiICnxK+nQNiLNH59LzD9E8vn061mxpqHWro+W9COjpJwLUtBFuh8IbhzuYbiikRZ+QOFg
NYdpDRpupLKRbWtTEgwP0nNoZZNzN+G9XmtjJJlIlVQv8sdbueGazILECs3Ob2QwSiTxlYOT76zk
StvAAa2u1XCAe79UubI2XT01E0a3URzDCJLKpoIQh0TI8nOaKRyixSQdwgH/a4pRyZYbuiWXTFKJ
+Ubx3xIT4AjyT5i9eSWugtnH5+kVH/qvdwewPLACsxGwAmL2AI+jU2r6IOYuXSWAm5BsfNOw6WYa
O/gJ2lrWjm38QFBM+i0d1oZG0YPOQWMPr8izrrjnTpQY/YH4xAgYiZ4tasvQZT28Tvr3PjpqHro5
ZtqRWUAW7zjCRlsSp1NJro1Sb2b1Eb4Tf+5Ve3rZJa/+hX2IcjiSmf5vm7h5XToFXJqwGcFK5FDZ
YZ7ltPgzThbD229m45tNSX3tZdL71utZFB/QVJYylETpOJAI8mKH0KUoInWkSnRvvgKlT7WP74jx
jnGPfeykMk6D0pcnLRoqqEnfr8Njf8/k+NmWAkJDbIuwW/4ZFjjlR1wEp0OKHuhegBxaYzzGu2Jj
iUG+dVqewzrgF8yhhA8EaA594vDw6U+Cilz4ycD8/cLKML3Fe3tY7mWmQPLVl266eCMWSRlp6uZk
hDyT0LjDhnnkyZHPXXNF+RdusJd9dZl6qNaWuS/UdmFf6e/TcMZXgyHUIvyU5ZF+S6cx4bM9UEnP
LkM16aquV6s0kxef1hUzXl/n7ami4UDzZqDjqlqtAMxvJ0x75ac6D0xrMrcVVkbMd5YGu4sJSq9L
X1Igz+Cp2xokAKw+XPKX/XFc35yMnYUjijCyiU3Bcg1eNmaZ0kTAUrGkyMaHadOmTPVTQL5t9/gu
sbSK4+vvIbYWsxoz8+UjPLLVxsRBF5JFI0T6UNqG0hLzC3+tOhPJd66/Bu+KCMXv2dxGq73BhfwF
tyQCaIlHdMY2GyN/g0cMqFv8QzMF5oWUOoZrg0rl1UG9a8XAvBdj6HZaQg6fht7TFAr6tpM0dVq9
ObXF+DPTe8bojb9TReX91/PkwAIbTwhY8dF0VZ6sDvw0oDFvSFwgD8+8fFb/MuAy0+nvobQzoBEv
OvImpa2DskyDWXcRzZ8kuuOSebqvK6Zvj3MXs6ekL3dnD1kjWbxjYwZkqj3L0AgyyAR9phhRG3tj
i9c1/e8rfzY7ectaVLkcQxMPba2JQj3JknFLBSD4hqaY/oE5V8bBvcBxRNR92d8LWcstVe8fa5Jf
YkGE8aCs1/fNW9dDRkvJRV1Ec63wKse8ShWELRmGCTse2Hiv29BD3c1mbjBRSTERtnrkjxfeSyMU
u8JRFRksk1SYsjLRISaWdXV1oy8pI50jguK+RYYqG3UqVGBlmqrGDYSdkBTKrBgmITXPGY4sE5SR
IOOwgNHQH8x3u8FNXTZCOvsFndJpAzo0JYcMHIDQlMyFdhliYql8WIX3v6ZomgPOD9h5EZOJtKtt
NDsG8hzqN1jheVk9wYIHYDknjoVIiSGp9oO5jRSVMVS6k+zfdjIodG1ChXHNZi+I5T6aolTFWViO
DGJgHgnGObx/hfPbf+faji9WduHYcCXlndiiEUwlhJ2llW7SN9wz93YKlWXvnCY5oru75EVOWu03
dl2jcF5190jXj7ObL77/ra4hTzZZzoj2QY7CnZmpQAjKX7WlmO4mhI5huAMfKo1r2VqHzLnndSw6
6BEIQb8Fr4NPfVLjqB7J/wbwuBaGsAGQieo/+iLw5rCVrmF17Hq97ATrYbfGlanv1RDC23I0TLa1
0EXNZlB6Zyz3MsChja/5SjoDfPjZB8xLzxXKZR4C46Ce6GkCMxu4+sbIjRCC0tRGLqxdcauvZTBK
HhWUFE94YRr/DAdCswSLKmSUlFQTXw5rfMzFFa9BEOl+efW8AgiTRGfM0GuVq4Aoc7DyNgwW3wEM
VX7yR2ZtZ94v1Dznmb2JTBwUL2s3UcgBxbPEdUAO7qMC35uflmFmulxZyD/fRoOGTXc/kfHopAxD
IeBLQbWJzNIzUSaViH2uX9VKbgigeFohR6cDr5wev6nvb9fWA5LtFl7pXuek/4IeTZBmAHClGj0H
iWnEWldj1ESevDt6tcGbqxcu8/1ii3y6AA2x0Kfcsv/lBWNWRFk65UEeEkGfsL5FT73b6z/K6lMn
0+qfG+JexA2uMoKfBahlPZJiE5AFk5FstJh9d2wp6LfaEPoQy4KClpOIXVOJ0zq79ikVoWDmKkDI
xPNF1MVnNSZo2jP29xx3CMRsP16qOv7m5kZrGajhZ/rwtNOw5RBlFO+yRAxausbOZaatFdn97FLb
XxiQPioo8QEbywygveQN5t6TYMDCV3IWplpjl+99SzPV6TZYlOBU15qU0aqWhH8Yvr2xqUVNTFKU
FfMiSlnHjSDkVo6Gq9hTdX3ismjMjTM4UqaTa4VlwODYPV87ElQv2efmktg0RQEI2Gf8FnM/PKDJ
98PVO/0pMek5zWgDxJJIJ1dXpVFUcJ5Rnigy7sB3/rsesb/4klUCB9A3KzsGkBgn9VayfvwDgZfA
REIb7H2li6Kud/zYsvJp/fk2XIBsg5dKOF+PRlJEOWwfeUmv2KjvFB8PxLA8S3zBqfNGBBo045I1
k5NKTu8gL9UQ98wB+5u/VLXoepfxfO/oewtOomrdIIu7g7X+PqC2Xevip8zpe1v7K1m0h33+DPhh
r/S6gOfBtRkPhOIXFTnwqzUU/GjuQ7oiR25v6bBmqq2JS1zEWeniQXUvfe7NfXy3q0R/WlV31e+l
D54Y1Cr0Agw02ySQWNxOkxS2mU/4gKq6Sq6jertIH7XhTORBD4y0LUeeQTMndYRGTF4PFsJVOn63
omeByOwIVDBKhqBtgvw7XNvcmHcMQk5CDD18FJFVwu0dBqbATaCWeCCPCLTBWQJGCwLCDu2nFvcp
fV0EsxfNUBGce2DvYxF/slEU9OWA8mmAEP/bPPpp6X+3z1GaUnxXApO2XtkPl3JuMMV7i6oV6QOf
782bHO31sJA8bMn1zPUWMXU1ZUoOGt4noiBOfMeHqzM2R/ynIrKtXQQv5vl+AkI8NqCb1VtBFOYr
Svzy9VQ1FpYSCmQu7Zmc5kBfBiv1Bs8EsfNjMdOiKG3DlLXEQuiQKr8JWwe9vxeRi3TtVqgZFFIx
T/XeHG542ojcSmL4hblRbC5cqYYOKuMcxHlUE9SsKsmmh9LYQHiDlakSi/U/1Ba59fDDuwjg2iaX
FKXrv91wTukx7z2rQsbWZWqdszFttOuF4pJux9blcR4Xoxb46wHbMDdq3IyKJT9iTkqbIrDM+xQP
tX2i2GnKDmbx/SApQvaihudbiggTMcXURAyY6hUmHcm6XHMHM9GDZm7v24ne0/eoGW3BhGS5onQ5
a9p5kVYa2W/nzBZ9RAJFQZUy8T0EMqsYUG2AV3q++HDI2KhjtG/e0DiYm72RtJfQAJrgZJK9mWEy
yK+mu4j5sGUWMLq7dyDNhK0uPM4FAO6PJYaz9cdlcDY09vH54QuD/Urgxw4zR0xFx2T2r4MRDwDN
jPFo0nWz73teafDx3N/BLcbHSgeVk9glnV6Bx8Cz+QxX6DDGAFtMZj8rcqJ/ugPCDS3Y0rThL00X
0igGgsxJ8/wWbHrRPc2BMeGzv8+qG+qe+hJDxFqRoPwQRpKlIj/lEUV+Bxo4UlFkvIwVrEnOF1QD
+aNeSNkFnW6pIof2SL+TI4yUzb6mO822Q1bmyJw0qzarW1SNMYfXpYZUd1ubyERRJTNemv7OJuav
q1tAB+wv5SVdDdJx+GOe75l/mxiTOrcEY1lQUpwynBOqpMBVsYmV9E6LzNuFTu5WcAQVX8WdWHso
dOQcfVx6mS9154Wq1qM6ztjh5vUwTPQ3Grg1iZ57XRXXcVa0AZy5k6TP4rZ9BOLdoKDthXPq4URY
+uUm3nWu398PnmUtZd5Rs7Gi29E0QrNoPByD5W4BaL7RdcowCTXx5YO4Ea62rsdLNzrbNszUpMaM
roxHXPLxg3h2OxNDI2WtiUNMCoDb5VE8qzyCFm0VlD2CgTJohS3moKQ8xSRHrT5huKI5Oe629I6K
EN0wIyzZpuQ6jjtVilAnOPpZ5Xgr0jB8lsrysoceacJcdlyEYyE7v3f4GPLjAU3fHgOwM2qnoUXd
NK0Vt6lLkQQnMvKFq780D8jMzQk0dyXFDwgT/1Z8+kbyBBqxkbmwZH7d/aH6lKNg+Wn5gAvlve27
ykqInLvOuOSD7WFFSMPY4wGIxvM092VUp9V+Pg3NNeXmlaCJ4L//Y6BzGrajAvzdXD3x0G07vqvE
vrO/EPGM6z6I+Rkmvga4adPqSYPjAF1ncKRxjswqP+E1ot0OTWHJAIcbzPBN6gbpDL3qchbkoPUE
hAFIczlZFoEo1vvwcXV5kZCgUyslWPITj0/ljhNjO54Q/02LVe+t7Ut1ufVM6mJNKXkBVs59re8c
gWQZ5l96c+p0G1GZuG+ObosE4Js4x+qtL0uGlXQpKS8kQsqzRZzIvmv/CQGzZNgXCpZrXE7oOn3S
XlNX22Lo21iE+S0EP5skVN5eLXvNNtC9qW4seSxNp6fpbhdThkn2pyjY6YM5fT4uITM2NLvMV8tl
lMfrBo0omrj+NITTkBf5Xc9gEskNDggMgstXVnMbXsEPExTBpYBRC3WMPc1qDqYepDWYe8IS9A7I
pYn31nHKeVlftZnd9tx77ZfGfyLGdjKWhl8wm6E05Ca6gRMbtCSqaJ8/WCtXoYXIi/mNLoLwFthY
ScqmJaqFl0ar+AqRfWz/lfj2PnKWo0zlVatlUakO3QlnI6FPnSKYZaM1z+yyrTIA9YTjcY7Boc9C
c4rfQ2iQIpy9l+1dKPAKI8es+BWEAPcf2/31Fk20HU20xKY8H5aLNWjM4ENF0pzTXDjzshvfePvC
Ez7VteF2gYJJl0Jay5f/Y8RcMg50F7c5gT/xErLnoP2pacl8rvggbuXskKKU/+5K0bs82NHSrEiO
PjgKI2PADWQSCum7aWFHSU+X23jir/QhPDg4jUz+MYsb44IXzSUg+lSYJfqi7qreqgdcUlsVH9Da
c5ZJ+G2L2Il5WKqD6+UNdsCdwM6v0RFgSRUD+63+aiYPVNmkEft1LnGAwIaJ8Y5Y1Cf0k15RgoGS
fZjs5AjxiWhEiPjxFDZe6NZ3MK2CyGhFaZUmQDjH4URSh7rPRvHEzE9VVT+ay+4WoYqmlaGbfKmk
U/U+OFuwYFQBdwvEpGykPXWJJphcrnf5nnCQo47HmTkuYudXvV2sbKNzkpOH2l5Yr4i6E+LZzTNA
/XPiBNzjClFQaTvljjbdJlmoI5vLWu2L7kyowYUbjYB9lGFFrjZw8Q8NVskTs+Oi43fIobKayPvg
3YjViFKS6MoK+TqTmphdlkX9/oBFw6lbphnucqM5EmKw/88RgPwGjTXlUUp+1LetdtN8uDYxAOZ6
qFvDgd3taYvGC8cDfyGtGcTLfWk0UhBTEsw94T+QrjoO6+8vefDOqqZ6bKv+laTalSWp
`protect end_protected
