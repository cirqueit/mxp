��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l��Н(^��9��j�-��]�ޖ���q<6�RYcW{d��fɯ��[��x�H��y۷Bԥ<�� p'S����hJ��F�@�n��U�j�U�:*lUI�o_��^�"#�?�c��~I���OUT�lq<3�s����4_*�5潇�TVq�%�Hzn�tX�#� -�Yю�v�2ԑ7��@�7mj��-+-��r�%7	I����&��Ͼc5 f�>p��;���낒�@`�#_���x�sC�� B�R@3�\B�&Fb�5�ѣJ���7ds���U`����A�3DFg	T�a�/=L��1ݲp�����	�� ��!x2�˅(9�u���w�P_O�N�fJ�z�'��3���In�7Q�^��驻k������_H�b��?�(�js�_5F��!�ݕ�|Znt9SR��4��0Q ����)%I}j�8 w������w�&�>i� %�k^�`��)Rm�o���-�z�v�g��~��N/Pڔ�$���V.J�ƌ];ߞ�ث9q�]���\���yAp|��q�ނ�/>[�3:~�~�q82�o`@%f/"@~���ү���
��R���SH�[4�Ⱦ1ge0�\-p'�ܿ>^a&i��H,3@bX�=��{�H	`�e�}���e`��6�k�Uw����x�f���>�g��5?�*�Z��o.�R�X�)t���\�����#mj�s�FɎ�]�|C0'7~
/�%�1C�2q��yr�}����k񲊗(�M4EVG�x��7�~�0�<��D�[��kG-���Q��b8u���5A �*����?2}�|��e���%���D�Ǚ�(Q�����05ĆY��A��U������Q�d�M��e�0@�K�!.�򤁭� ���􉥴C~+/�BR�0�:�K�a�m��>��5Br�r!4�5�2�9�&e�_�u�h�|�=�S��'f4B�N>�W|(�7%����5��H�ޭ���`u6�ҩ�-���7Ͼ1)�F�ZTuX� I�qu�͔ߠ��Ȿ��`���9`�����Lf݊��Gnu�v����/%�E�Uc�x�X����2�QV�z���/���s��<�ί�W��cO����[z�8s!g�ak��4Jn��I8�@��P��R���h\e��������3�\���&m��:_}�q��:���Ra��hj���帆7oG�wm��c�IbC�LN
�����~Zo���9�}�$��gۓ]׺���H�,�h�lXt�xcV��ZϤ��-��u�o��7vqC<�D�����i1�{�[�):�AښR�d�ԏg�RΓR��r�4�{bK.�;3����%۽v��ټ�s&v�
���y�*|;�D�K#w��K��JW��E�~a��L�oJ�!?nDA+�e�)\�⪇0Z��D�#�i��l��0Z
>k��j��2�2��\�oj,�j!< % �ܫ��Uom�R�	���:(��0�d��Y��Q�_�/@9bZ�,���(A��z6�>"Z!B��E��f�=�M%K��e5�v�~���0a�8CM`�V���	�;N�S�	�t�|�Q��b��f�j�aX�˚�?!�0�'�0@|=N��fxN+8�K��6��Bl��΂����5�y�#�?}(VENEt�$ah�t� A�(-RC��KO���S�
��P( ��`"^���a�|����f�Ƨ�(d�b	�W$��������C�maR�2��bl6󁳟��(�-��/�;�~勁���P�ρ�3�>mg�a��%0y�t���Ș�fK�wЦB��;������Nm#����eyz��[��E)�3;yJ�����(���sE��������)�+����L����no��2��i��[�����0�	P��hlƤ���F+�6=`�Êi飘���)�
�<f�H��oǱ�9�qC���(��4$�@U���.ˋT���9;E:u?���6sЌ�\��X&�Ll�j���C'ѱx4a���`ZT�@ۚ�'mR6��)�+C
Y;4`tG��ɻ�-;�
�����ts�mAk)��Ǉx6����I)-��W�=q��4/�����7Q�f���T�1f!B�D٤�U�^�r�����#T�1k��nׂ�'3�9�� �[ĞՈ˖s���B��셮���H�G�;i]x+ �I��`�v���3�(i�7m�U:C��:	PU�w~IP�%0/P?C�������:4˱���P,��H����=8�2�N�-$L����c���������^���U������Ϫ�C�%�=�_�@�	��|/H��V���s `��܃�ɡ��}���,�쪌���~�7k_ׯ��n?���$Uòi�:#wQ��K�-Z�˹#a����3�x�8�-���x����;�R2ƛ��ͳ=Us��m���&.�gS9��"�q��X�y��k����N	��-�nWE'�ub�mc�'z��/�[*a�|-/�ѹ��
�lo�Y��{� N=����0LN*9 ������NP�fCt�Hplc���2H�ESp���>�ꢽH;������
���'T�_:���
�N��l������FCbϕ��=	�3�JaF���:Ad�e۱/9���63F�7����5��5�t���!ޞ����N������ �8��'@GD��ГH�J{��9�ݽJ!z���/ '���(���<�g�2���ףRkJC�׈���~���_J�dAj@��C���c����"d��BC���+��"����ɂ�z��L��ݞ�2��ʈR�W���Wj�2�����R%�@<���>{-y��������i�ˎ�H}'�*��:"
ndL�
|k���0�d���Q-��=�u���:Y��^D9��8�A�&�Am���[S�$��,Ŭ'����B,���ҳr��!3)�dl�F/�n�}(hC-�jpΡ3l����bD�/�V���
���`+�6� 8�����ߪ)L-�]��t�_��9Ε���_0��'uC'��e�ɹԣDەCHA�sTe#G >���3XO]�.��-+��At_���U���a�7a�m&+���Z�Fo�V=�kW0�%ţ�ky��N��c�-C�r�?q�"U� /{K=4(,� ��g�<���J*K�OH�.o��K\*�qGm���P�0��C�rZ0'a�� ����E���ك^'-�������[�����C��J5ȇϗgp�vd�#8���a`�.��/*I��8D%��A�V*dD 	y��K�ŷ$Xc�a*TkT�_7�?IU^`�-��3�m��Ψ��ыh���gH$Գ�b�0���z�1:n4��iI��m��řU����o.�xGq����EFؿ�-}X�����J"R:����3�=�P�V ��ͻ2�<^��T��O.=��Ǯk�κ�k�\#�7��P�����B�a��AH�\tU[�LElH`<�TH�Y���ҤJX�u�)���O�(�v�>Q4�[���sj{-���nBn\5�{-'�murI�� �����tI�q�?�S���U�='f6@������:I�D.)O�V��#[�T�ր%�����V<yF}����\P91�1���������fn�"P.2"ԍ��K3`G������v��PS|�NG��1V�X��Q5�(��K��'�������P'�U�Ih#�5��y h��Qg���h6�\cd�0�y�d�?��9֟G5��/i�(6I������o����e!BX�r�6�%�m�1:��?jy
|�.��I�F�dr�F�G�̽�܎���o]M�F�oU<�:�T�jmϸ. rlh�*�y�� '�\��n�R��۟Leid^���;�<u3Da��(¨�Gy5�����_�������o�F��?eG�g�źuo�Dn�~B�Y8&Pvi8�L0%l���*�F^�4K�PU�3����Z-���c�?ֲ�Y�V9�!�����(�>WE�hYͺ�h�=���[<
>�I2|^�'�>�K������hg�"�2M����jQ����(�L6�~q��^�;� ��D���*�i�Ie�
�0�Vb�V�b��j�닓�QWm��1[�mXv*Ît��"�u��Rug��o���Nw5`�S\^=���u����^�+�؇4#��w$���`<�b��)��:k��4���yn }�l�}Uc%E��<u.���摂�(@O:��۲�͊����E�PK'z�P�68�y ׈ܷ9<`'&���	��lB,�J���'h`����E�8�2�!����E�(�E%5p�x�[�>�"�%��w�����J�PUx��w>ע�~
m��?�����ob�;g�(o��H�a�_���ë��'������v����aӪ�N����_�K4ک��Y�kɿr��b��(e<���ɑ�%�{̋�Mj�/��DT�f���]�5��T�`�ge���m2,�����w�[���͍��"��S�3���:"$�d}�������'��9���ϲ���1��'��Y;g���m��:Aʘ&�2��f���ڱ�;%I��,�X����pX�|3��7!x�� ;�X��~0�g7���l��ˊ&�tzhO�����z��.�<}�a|g#�X�s�4, ���ME����W�kDt�ٹ�'�
�t��w�A���=%�-���%�X�4�e�a���d5	�_i7'�:�=����{��. Ē&�P��Z��M4�؞�)|U�#�d�,_#F�q��չ�P�@��y�d�º�sn
�ܫ�(5�	V�%��۰��J�"������	A�__��%T�Y�Z���_�rSA��!h���۫'%i�n)V�Z�p��63fr��qzrQ� ���R�c 7���*�}����s��j�."��K�Ǆ���pP��\��q�(��Wߠ�tv��o��q/�Ƨ���a<�X��Ľ�Ŭc~���;���3LR�$-�=ɧ a�-��_�u?������:*X�{3L~fy��@���C��yi�E���'c�<��t*W7��p)@���y��q����}"�����j���I����m���@�9'��prk c�.JOK��βS��<�}l���S;�R1�3��tHѷK5�OYMh�{�>����gCv���xr3	�V� �!�5��&�S�o�6�3yjB���*���h�{��so�2���yt(R�o��@@}'���-���E{I�pH�N��O�z�<S�Y*}���g08���'l�z߇a����j�^"ͮ|�/Zn�տX������q�w��9H�0}�PȬ���iQ�xN�&M������d�{��S�;t�;�쀏��L�u��n��!�?����Oց{�����eo7�b1dV�KEM�4��s+��=W���k.�@�و�kFSx���~�g�Ep�K�slR���}3hx�-21U����
�$R��S���vQ)Y��~Ume��>�4 ���c�dG�`^B�*=�8h��,���C�mL\D�O4�����p�&�
��q�/����oy8��=Vb�Ѫ��(��e���Þ��-M��؀�y�G>$@��dR4�vm9�[�NT�u�79n�l�;�� sq\�sp�`��װa���jh-!�F5�Jh��ւ��(+_���F��z��>A�H�3ӧP�
�
��e�A(Jk��tbѽ�gm`1.!�'H��9���I�(��ч}Y�K�J��� �q_@E�[��u�i��sKb��EM�����'��W6v��З1X?)xN��$�ś�� r�q\mIL�i�0���D��ղ�M'���pш�*�t���}4��{���^H��qUaF��5,�{��~|��x��B��G���H��Y����\��`g���� �]��7S"T���6T�D�fHυ`HSt�=ˏ�Rqf�x{"���IRK%���3�t�(���(ػ�'~!�����݁&���zK����6��v��-�^em��|��Q��ubSݜ�?��c������Xbi��3 r���(ݛl��0�p��a ��&=����w+�VF%7�'Q�b��NzO������CV�i���L����ـ�(��BC��>�ڽAV����l�����14�5B�҃�Ű_ْ���Q��{���S���T*P}%�2��x��1��>��2�������*����"ы��R��h���Z} �� �|n�����o!T�������@w<��8