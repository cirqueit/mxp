`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3840)
`protect data_block
QuYqVIhaZJULLMKCJcbmjmrusxwa0giD2io6U96MSs9UXbt6B+sPA3reT8v1D0LOXuBSNcWfuWGA
tgPsu5iOqZl7ulBC+oMTRfv4ENwpmxB6gWzVsZ7QNa/O94ddgUebiOR8HyJCR7whx5JlTTA94yZR
TCJ+XEAL5k5A25lkOEvs+tCt3fWo6s84DbzKwdp4o26onb1LDnAqFhTA1WLjMduEbGrgf2m2b7js
alGFi6ZEcydFri1KHcJVq57hCaGpW+lxi0fIY5zCmFJTXHk0bN2HMQ91fqC30UChlsQfAW584SKN
juPAaQ18ILEP50nhEL1clDQZ58lfWs1ERDdsy7A1knaTV4p6vmPs/v/92dGXJUv8gVkbCUxulHPi
gbSbRgUPk8ApqBjZn1lvV2yVd+bieDUALCOTga/q6qh1BZkybZ7kSOkDkRak+nEk1HfwjEss3YgA
vWEtslBNCBsBC99RHpNVQIeUAF4O3LOei8ug/9C59IpGOVFXscLB3M0oZ6fJWiPhvG8wQtJUyJLo
PeJT9iHfA7UZpx5zOjlo3sv3Izz3Pcb+jWNHjLaF8rn+eNpJvIhwp7A2Npfounamt8zrVGezoAHh
ZGh0pdZxR6kJz2Bp44NeTPE29/SstQza1OtiaGXxiS0D/zsZHN6gWVnWme/o8NAc9Z7On0ry+8FX
O7fteKVZQzkxWpIlPpz9xkGw58YXXR3Be9cZcaftylkGsFqab935q94uSdLSlKYEFyPzylfCU4hB
haxCDGSYgmn/UoTHqZ1eMypttqj+YRTLml0XqEYdMBGWOmAtb3vMQS2NLRMD2jQ0lTfLiy9a86gw
EMlIp9P2Yhmnc6nAQ+QY8r9CyMNmb/dVYHQA8RShGouNw0zdWkGD0oq8IHo/waciA5hayUE9uKY1
gp96PXwcKQG6wOZs7mpXjOkyEfi672DMaLiN1MGqDUznRvOUrliKOJyu97baFvZPY2OF2ZneCa0T
65t3WbNfXH2WNwISvF79WSpOF4v4sR7y/aYB1pMXpEbTdL4Ox7tVs46lprT2eFKTSjGQM9XFySx/
VyNSWFKw1cWgQo4mIKojl8uupJZcfgFEuCezpaCPSr4CHTETP9dIfPZ8iwaJ7qmmOvTsbjdKQLsG
Wd+MmEEi5w64Rdx2vEU4RIfQjSqX4ackzkoT5P9M8pvC4jzZYzkX2kpPdFYdbIpuT6/g/Z66bzjS
u7aF6qUKPwHR9Z53lPFf1Ifd+H2CY2NVnNpZiTAyN+NdbxPnCihULD5exE/lcVcrpZYQMikdypM9
/GXOKgc5SRkQhtl18TOaChP4+p3wSiDL/RfY/Y2JpCiMkmnE/mZTIIsfVvXOpKJZ2VjLPsRnikTV
1BjPeHoba/CoI6+npoWxlXbdI9YzB8wS9D/u8gYzYbbOaqCuj+ZaswaJqXS5NbrQbvq98RbKZj6Z
EpBeVpKaUTlRseT5QzDxUKMqyopuCgqmtbNeKblX55Izxr3VBPSNu9wjQTzYApUbiJl05bTM5VUr
XDsDPeYmh4fL/3+4IHbSyjnv5pUCB1M0SVal9t3sdet7+KBr8XH1AKJ1ON00nOUW6gR+gFgFdSHA
MxxWilU4cK/7qhyLYuMNKmZaQzGZiIY6kJIAmNn61oeY/vd/auA3f0KQuuJQCNDYQD31MexZrot5
o08LN4wclgaCae0Qwl49BgaEcN3vtuIiSk+QwfEiB4V14Rfs0vvVyL6IBJpZkixwfKczhVrUCONl
p9Z+4aizmQGAP4R8DgEz/yV9/id6a6gw0rwje2TzJ51OvIa+7zb7Xl+NqGVTRhmpi9YUKGWx6RU+
WWSPmmSc9GUvVuqjjwXoJJz3FpbFysWsTGAWYhv4dQxDYZTmAl149xlHmWGkeiGfD2yxi+WWv/lD
1xdK3asslHWNuHfQ8heEoOSaYy4Q8OCyRBQr61WaE7hiLBuRsOdXcr8JOjYWJ6aVZs/ZvAlLAOG3
5MBdDR1ukRgohiFC5ssH736SQPU/KJyOOSL4iD5jIuq98y8/CdTYyLOitNR6zn/0Bhb1/ISxmulK
j6xyzml1VrXCRZx1UNi6mOQj49+eWg9r5YXqiLT6JidI0qyTU30eraeXE8icAPNYRh+IJV9hhAoX
erQnL79B/fyGzi4ZU469Pzs1bynWrWqQHfSikDqAV87ovG0HJ+YtdQkcTqCFgh+q4yPCcahKVSxX
FqtJ5oQn6okDuxB/JSzUYFnW8GJvIr2wmrjXRgrEKCxYxjyeqR++Mb5gzjLYgbU+o6+7XZAVulXj
ix/EFXEUEXN4Eje15/5yH4OkC7CsSSBNgE8CsZ/0zh8wsjcFgQ5y5pN9WgxSxcywhUsAzkh9TuzL
+YTkaOMXI79hIr1Vo69jeZVOT77t8jm0x7xoF43BXpJWeP40XME4ti/kjlqBvBMklDWd05K9fpNl
xRDwM0mH+OPE79lYXpldsxQKejVZiKWlHSd43YLwSw4YhpfjzcCTus0meuDkCOYqXL751d/KYGbF
CFwzZ2YvqUx+u2kiFWQzVqa4nCoYFuh1Rg7jGvsO3Wai6YU6iP0a7i0Xl3rfiy05woJMb1ik6eE4
9PEUuKFWfQV+RMGk2etj9ecbRsmQdtpVJlHBllrQmljNAJWluMMlRal6nF1NnTBHCXFr/vX0bXZi
ZQyqJVkWQRYBYP7ZSveR8J7G8DKkYb3C43iDhmPM7vgiI4ee94OPB5BCKv5mp2ML8Re3yYVtQ15l
sEPQXOZ49YJo8N7L+RRG+wgsF7WI+fnk9KCK98EdVTTZQaoqrVkAswKeGN951Y0UiCh+lyfDL6kS
1HR02/XjINNJVl69iP4EL1vZaRMU7yEI37/2vDR6fNJbIGW55MYVO7nmFgkk7W4q6a0+r1DcDNqp
c+saBCDFbvgRRY2MHiWN64w1HXA7a9euOy35ZxNsDMKNXeuN4MfrFuTPrbTxUR/2x1bu40xeEoCK
MJ1OMvn6rfOKgYcRymjgpHbjTbaOWvc7wSxVV1eGibr5Pm6R2EnXYd1R4d9Q3dEU95N0WN5fofkp
XZC1qw0IBE6rt3UQ4X4JTh7CwoCGC0ZHOPHRiE66BsN7cqjCTrFZ0AL5Rpm9mlbcqbwmHPyb0mw1
LqFfStX3FcI7E2XtCWRlLD6q/LA/8ogUvELl7osSESydHgxZEfxaAkcxsToUd/T/+6EGdEQCsZDl
ufasqJQo41vCmAcsTe8eWaBWdKu6T6shwh6fbFhsb+eS0flmZETMjj3RMlzp+23XIFNQ/TZgtCc6
lDvM203gZLJSL6njieyugTTnr5Mui0fOiRHFrJ1Vc9QC17MuWNR6d1T2xlDxpHcMejO0eIRhz4IV
zOWFJ+Tj0EbS1xdyo6hLprIsaYExLa8CT4lE2mhk16WOg8WWixyuJ9QPKswwfMgld6em4OmaZ7VB
Np4oDb03Sop9uj0YcqBDazPHXNMqf1X7iFZA2JrNqOkCDwXdx20VUZWMc1WMZNp5TA9Hemo2wJRb
dkGqllF6lHCeukY8pRZWeh4NqhEqRlNv9vSdwXHj98TIhqLdB0Wwoc7v0obAVud8Jv4lKC+zBt35
E6A2w7YEgkS5KpUskdF9/x6LYTrg4XaRxIUCSznLrid50tTitZJnIu0+SR2Zfllb/TJE4vlGdDl8
swvxv/W35O67AEI/w/I9pq4GNaxo+gXsvTR6H4ySAdWsFGv7y3bjb0X86g2e/NKK2zk1GSJTFDMZ
vp9fOAJ+xuFlsIuxdznIi/qEhRh2qLftJhqiLPfhlWb8FhZhmuKJosO2nRA9LejWRbhQr/69+HP/
0OkPh5Oxsbni72uup1SdwpZFTunD6xpPf+PgHzJBUlPC1arjD3l9P+68wcdccyPsOaM9namA8Nod
FwaNE31l+pa3eoNkq2HkCcomqkN+DeBLF/hc6BFCwq/Xzzl2lEclbV/NLUPh4cabQlZJxYAZy48y
VUY5wJlNWyA5gvMV3pZ20WG24sxUnIXOML+4mLPuLOKPpKCfsXxyhCmz9VO1Ayalddm7kqnfcway
xs2v+fYREiFBmpKHVKeP5FPf+InmcUsjnqSVPt7DQf4iQlsfwcdlvIhRV7ePVGrW/PM7A3pbunxD
S0/g72bVBoDmNw8gSyb3CJPm2yDLQmRgOER660RNGbdmQojp+vzCUol0hZB/QIVv1Sr2kLNNJGQL
1Y2j7ITVowzNQKTcZQahM+TiZx2OcOo0O0j/rI+TzjqF9e+shBG19mEvWnTUqmn8lp7tRlNTctM/
xHbjyVdFEJ6lMYPFshPPTlicao9sizbKCW03gc8axBkk73fzJocL4ngh5HbB9+bCX+7nl8yUKOH2
0tcMHYKwp9uVkWNDlusSfo5v3YDS3bReJlLmTefUY7xTG+twHeIxI7pZNYEFM7s97js8p6MwC+Tt
CuqWp8jTUNAzEH4MeEAsD6m9GU53L0O4WgVMrHnqgEMDraxVRQggNYYYvo5rWG7yfiv8rKpKlkUH
+I3AB44yBj5VHloZZKOLJI83Lg+muYiVCl684KepK0N4r15qUOpFcgV8wv2SVnlzANJmV8RyvqlR
KuXKSswVtKEdmQWrcc3fPpYFWyM9PmXw/Brf4pPa3cL1ZmJkwOHXUnGvWPvGdAlRInTx4068riJU
rCMrcMb7Kp1JC6hFHhPKfZeFyWIzTpleAWEvitAc3D8IySH7b9MEjgVwFociMk/PiFEp/OS1QCeV
RvU3pJOWR1Bgr0DQSi8bqJE7JwMwifHgKSrEvBNF685xWeHQvifBpTgvI8fZ/rF7+5GVcpCGeIGz
qd0BItgwpQqINA3vgy6xRFEkwQAHiysKIBf0odeNunApdK8qXa+FiWtKqsEMc1KJSmqzx4iuF8xE
aNbBsOJRV3uLfy8fEUpGl3awu3SctKXd9VKGDIfT09+TSg4HoQuqBHn381mOnFNvlPCpSqxCoKHR
0wpjvA/rlmBfnuVuRLfQTmOUQ6Dkli2VPbxcJB5BioJJI1/WqT1X/xiPXeNYeFfW7Q46glSjrGB2
5OzJwWj7nu/OQceR47l4xPikZNgd41dfXf9gi0mYn/mK+sYchcEWTk/CVEoWmI/cpJMLeHJUcZa2
ZgQKSpdn0E3x8Te4nsD24+aTAxkc
`protect end_protected
