`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25696)
`protect data_block
enwBiMYwG8WLbyHLKpu5sETxtpnRYQdTdZEDNl2vKRMB1sz71WMYkIk/efL8k1nny7xL4ZUVD3QD
0gXjQAxM38s78WSzC0ujDsrcuWZP9/wk3PnY3e0u3bqNwuer0lYQexe1gbu2QoSJNf984M4mgFdm
9PVaKq0/00OBp63N9w3kI3rROkQ4bx49fVyVPgtbVGac+1ULMObCAzDXPFB/ReOWGvza7o/LYgP3
ujutZzt9IFmJ4/1SV9HHUYbCd6+xDYtwV+Ag9IYssa2vUasD9xmvy0/pLiMp2g2oroWTxcbqOPmb
BWMJvXGLDo1BDRC7xzrzcPzCjUTaNs1F27AIvKtWjaVwEgWsZaWYyBd9+6i+jiOSoqElxFnD6IXw
AQwVXuU51N7CH8gi1FIowxZqBS/EqxYuFLS941SX1QrWR1dP7SlfAOGt6c98EUNpr9sMp3/bQ0QH
65BSjAYbyK564SzXOBnrY8btT6UUYDqRHILisViLB6XFzJaXvZVEmXVFsFGbM06zKv8T4/eto5SN
sP0IrRj2hk+T++VsyOHCQm507w9hB18yNU2smqdh7+xzCy9w5ZhVlaTdeh4FFQ8eL4Xjwy+JRRDS
T8xf9YF+wA6XHBBCNMn3OjsHAcWdmO5Brn5fV11F6WOTZeQNQVtNQtbasmSTcr+9+rorc43RN1h1
y/LkPXFaK+suhm+i2/7i5YKXplVDzuDT96kPhsfydA0eUOgkDucDOMRfsywGjlJWbs4xHT0zAmve
M4GLj3CLYPkzyuiOyrNiFz45tiJhmbd1jL4evzQ8E2VmRMao51miLGUylr2aJmW0qh/VW2wjPiS4
R2NNKIVR2PU6Xnwx8p6LZ4q9OjWf437uxnF8vUFMjlDhptMs6YpsyoiLoCNZKq5BwkYRYZWfDHrE
1qY7Y8fdzVO1tGlNGAOHkoRljEYGS5f5KiP0TlNs038rPZX2vsqdtlvgVINpbMU5Mc+YTPnnt0TL
yDKLiO+AlWgSd3IJ4QKzFH6R24erSrav8U2ZBQcmbwYCo+vLvpF/PQWM7Eahtu9SL6UTEciRxz4f
OrcXUI06ILwSMNzV3UQB5eTgys8UOKjTXxqyYo0wry3oyLKZQe0ZOPK6j1bpz2iWdtjxDtBcuozD
nf6V6a+buYgf0d1DOD8RDhdI6PlKSc/lKJFKAaSA4DlACc7x4W8igIjCD3OXqzMng7dWqPLpOQsu
P56hjlL5tnkjgx0qLvIex0z60NA1ax4HxCZcyacqi+V8DVbBj5V+j+Fe77+Hv5/bj+6oAsqKsy0u
nJ9iNuoImMtbAgjjn+kqbnOpp2QVbz/NrPK7QsSeFgplW6/fVAjy48GNVnkbq4yE8gysboXTxNaa
Ijv43ryBPW4ZeyiCHu2BDtyuYxadneT5nvC1O2Uzhr99e59+nkRB+UTBg/j0GkexfGwuFzvsBBPa
nq1gy8NB8vNAsQr/x+SbSVrBH8l9e2Up8VOpKjXPEGDQc5k1jox9Kb8c3vvnjiAPNoc6eKrd3FmC
ZylMafl101kkGMsTsIN5J1DucOS0j/Fx8QXXlQpC4II/KkW8D+cf7IJIEibkKpUq32emc9XfjP/Z
zPV/hS1IR5dYC6Tlt89L3w1mcQS5yN+EP8T+c1ya/TVlmd/FXkbABosNdeUNToYo4KFx5Lxbbekd
BybFWAFj5JLG4FI7KCE2FkXcucKMr8hZu3bMPXZMhi+LRSSpLC9IU5PXlj2lqx8IAus2sW8xJYR3
H/0MNqovNTUUIzMP3Jhx7FwcCNlgRWPdm7bHMgA7XD9N0bg0h7qsD2ZXBe60XUeuav29JpdMaO0V
yoxG2fRluOl/PvPf6iXDRoj3ZylWZ49GZsXF1nfK4+XcXsk4IYm/7ANXiITlFkubyPGprzYcLc9c
xnnLj1c+GFB1Rae8zAtRdtw7qXOyA3UrpIbNWKn3LyNIWtmIPeFvX6FlK6bmGubkwp7wsFc2Eqc2
GX90n3/ZOlByBAjs2H+THg4XcpjgUj0TgHjfwa4LO1Rx//KWbL5tzo0vIRLQpbQ+5HkveO7RtOWN
Alp+W67kjQB0lCh9kmURoHcWPkvJNC0Qb8o0iT57X2D3u87BVehZZFEBH9wiFVfZvlsqymrLRwia
6sY9hXVyelyzhJoDiaPHiqDt5EKnPF4PQGdsHef215BollUWPSY4kr98rI5ETjGzdm02aohdGxZU
FfRLwqFQbroi3ie7LbXaE4N1S15G3wv+7IYEZm+VhUjk1VlponjFNyWNYdwRNWQETUh/i3YB61LN
od/zMsBt9ZlhtFt4cqykPKvyrFMDHvxra2VRlfr1lp05TuWBiurpAZbkdlE48G/TWuxWTBfrPjx7
Metxl24QMWqcpfZijREP0IQPwJd7rCwI8XD63Boo2q9GDxhnkqanBTNw6TfJyM2POE8R8bep9ui8
xYTqbf78qvxbfdbOzgijGTCPhoFOAMonLmQlmtIIO/kawvLdz3WglOlHJwXTDkmQZOsp1Zqbw1cm
6MrOd3n1XZ0HVd8FhXeH2ug/twI6+nCNvl5lNEBFvIbNtI34rIcLSdbw8eWA+WSPfIqtcGel/3+e
O8P6MzAL35JEtNL3286kE8bQvLJdqr7LYohsPLsbIB7gUeQe01dtD6hx4MeDUWMOobAdbnEOHL+O
bDrAW9CnYrWEqcCL8mOAz4yjiO4nTfX+6MZbKQEQ87VkV3I+b+4pGxNw4uxShyy1GdJ3mGG631WM
dAD2x4RZdZicvWhtey9TRj1U5kMJ1tUCESkD/VSSExGIORkaIviIXdt5YvPOTg6nEK+OaSrcssNg
yHpkfzB7c+yHvcJhGoPQb8IpFjM1LDRA6Ah+/z6IT73WIIM20VsKr2pqeQkgpRlMTa7TS9JXJvGj
61tDZ7+3BCuNsjz4LhSa4hDYHPPikc3fLiPnyXeztAk0HMFhEjzMWBdDT5Y2O0EVhs/SFRSNO0aO
2x0YqtdPdGcJXzAhM0ijKnGk+8IJM7Tix/GYSh0boj1PGHI8V+gWKwhclaq1hugzQ/Lc5IC4QRct
nsUlhyqxVgEGoVzCpQ+5lKfH3uvDCkLRRB84cQf8OXXidbG9m9Etkmp0RFCD/kq5ZYS9Nyj0FX6+
gWnvmVhOXwlpfnAhQrJPjK+PnRMkKfnAFaTEw4IJVZcjtu8CypVDuybtD23jMzrULigzuw62Hxck
Rf8Q/LoTEPhhZimD3KUtcQntPxGxfkGDfLsq3uCdg/n6D+pYiRp/Z4RpzqVVukO2rUwzZKCKLrGI
K0RDtQXPxYBoQ3Bh5VB8IG4WCKjqOLZG8fhApqxbP4pZKP1RXFOZK7AVFj0JTh8JnTQajUvzNLrc
aVfkLatYw2MQsRUD+yaQcwcfq+0DxmvOlEylH6nJ4TxsLez7hngS4PBWJtswlOoKzdMgiBQ9TK0+
+/gduFPLDR+11uaBfTKnwg/TFoHvZqAVzgbfORMbt/tH5WKdqMSNbCPs204LFmqPHYf8PScKFkWS
QzJqnnWuOHM5T/U0g98fe5VlOwqKTJGxXJPHA9tZjApiog3Y0iKhFF4yoHj7qlm2TCGJ0ubpBDkp
MKgp+kP+ke/tWjmmQfQ6Dzi1ImLbgjkafu1Zmfqd8t3PRK6Pio+b9+8ymtcp4u1NDJw8cLQf3jto
RwLgY/k4TSydPxMNdtNZIf/h5s0WOLXCZScCX4s3ukTzVPb6dWEP1/WaAaEToX6QjJTWoNqjM+vs
5wzIy7cb5OGvVhsGQ7PqFMe4eb6V7K1AB3DBs74bBz6RZAPGiZQnu5O8P9tOLCpwMnhx9iOuXRlm
kpKfcmnm6wCoDrlmSZn7xjIr79C2Jdm7pOhV2DQ4P+0cUVQcvmckBYkqUnlenglqr0YlHSrHcPmh
uq7PXuikdD+XXUCGvjAtiMKoWS3yFrySrFGrWHi/3LKQgshQqkZ0Hp4qaMbyZOo0Svz57VDDVNYg
Hbg6UmTeNrrvMurJ17izE/wOcZb9lP5nUuiBZ84rsxsGlXarHoYa/kX0wG4IdcKvxB2zszofY+z8
5Kk9dBlkjuzUrNwSK+OJg7RXJaXvTyuY3hOChebMz82Bx0PHFEB/CiX8YDY+GuM0tDg/Q8xwQhvl
4TJXErF621/kSDS7RV9UTbeoNzotcujWpFLIfROhcH5WKVHaqfavMKPXGRwALg0AEBtCHTaWQhWp
GX15XoPnxSClMZOQG4X4YsWXOnqrqEu2CHDkcfu22Q29vTb7AoSZmdKznPmN/bZNVbua2PjoSaDW
cSniDEbKRKm3AoykURP0E8Ds2KfqHch35aOToqtvF5C/SYtxtwu6WDmGKvFvMLoJWTXzfH1i2eYp
aSOwVPFexgu067+IntmaoQOOgIa2krBRfrAcXGWXgsEzseE44FDQ++JuExzS/vrT3zNLELXweaq1
/yjgydYCDDWmYKlgvAYUChxvO3Q4j1oS337kee0KO9HR3cRKHn86unRw32jmyrTYEsGTl2LlIv62
wdlbYgUV9kD5BJByvVWil18PJlDzBO/wWj6ydLmrhJc958fvDjvSMnhsE9MJ7w/O1/sCfe5hncfm
VRknEqG1k/UNIewY1sGoZn2WmBg2kqtWhV4cLcySeiVgUgFR6LLsc4lIa7fULe93cIvXjSuiifWG
32TIaVocV1PeBXjfDC+UoZ3LrUfJHT9tiaHNpxPl2ugGDef/m/ppEo1h9s493TeCE9Jd6y4dn+gn
tLhBxL/PJzqqs7wX+OigcL7ED6DNqqb2UYNsJz1teQ7NbDAFMKtdyabkeEX4/jBIAbM2rvwWnylc
YgdyRVsd13YEXtWTGVUi/R/JSzRvEvAn61adGynvGRilJw8l6yH+8tkHfPq0oYFlwJ0l5CoF4iwI
C47txb7/b80tIgEVUzZ7X6g5qzgOSJW3Z4UtXpLP9yjsPmxn0jp8TqVR5htB3aLx9l/4k3ANVUqP
qtBn8R0EgYZTb0c8d2sKcOLSu2F13eqeESKqvnwBIJzoT0Nb8zARnyvgB43Scghd7lRMOjnd2G0J
QvsEV9pC1d03dDqdJIdMsamRJT63NudIrtyHqTaX71ASe06VZgwDWlNn6ooUWyPmlLbrjWFF/O8h
g334eAhFqW5g257iSwfXhK/F+0xc8l8Ek0Y1Fy8ofn4hXUU8cQxrZw/7e8aZvhyAN+qwMlXMesUs
5qklMA8Gjt44c+Uu4sX8gVHbwkrETTVFOY+Fi2vYEksvjueUab1mUNuNrBYAZz2FlVgKdp8jchIr
OOVmtQaRkYOIu20Bn9LR9PMcvkkUaY+DNBLTPEF5EZNujphsO3X2nRimSMzEtBUIqbxn+OUcGk4e
cIAfhQl2/if0gRAIbCOpLeiw4c3TLw6EEmlyxenwvm5Wh61BIaAzY7wZRPIH4cNV9jtLTMUtbz0w
weIr34PYcQXE6b+esrR6AkVclU1/d4jW+J1SgBHDQF8xfuHNiPYOCxupPnBRcS/ZMSpLuZOnLtEU
Nob5KM1Bh+Y9ILulpusEIgc9ebMR6FZkPKwM5SZb0wyH5t21z5+6nWLd+BGBvLn8vMitJ2mjvh4e
9qMCsPWdhp5dj7jXR1V8s6nkOcQBZUoS6AcEWQT/+Y4uWX+lK5n44wWkloaJ+XLOTd6O2DVzsfBT
AKxi5BC8r+Fk/wr+v08GWVDOZBrpn6xGw71nuvz93GF4p5nXnhT8Ly3lpAInxocabdJMVR4AWIrt
0XhCg/PIcSm+X1YCkzCaYoMPkhkdAS4z0RG6z9UgWHl8O3Mv/zVZ21DOd1uEGHAjg5woRgZKf66J
U8pZsD7Ujo7k7wStDMwEqruCf4vbD0zDp7IzWAYyqEGonvQxUmIEqeUvjw2wnkQ7X1qmt0pDKNPi
0hrJ882h7iiab5cnoMogTyucc+eYilcrLv3p+lkQfJMLW2eJPVGQXvEzGU5AElhN2uqyGxjF9X97
3VJUu6MQGYlbv9EsooZi55nw8CaK00NBJiYpgv4DXENQ8cpkD0l9vfu5Khc+/9cZjVmO4jmrlXPI
ftcg795ML6Vm5bghU2fzLuwnm4Ihvg+T+xSivE4r4BHsMIcNlithbXuaYzQKknRTB0fKQCRz25dQ
TI9cwKKw1C49+stpy87aqaS76wSG/TnXHn+u3AUGetIdEt06nEdIMPHVV9+AsEQPc7+xmv1JBjFZ
W5bsvKW2gphYbb1vd6GRhPyW/Y1M+kKE2REq5c43gMLh/CMr9D4ouF9vO1IQ7SE9UWAsjINCFPn+
frHjLWRGNP6TAo+M8NjEA80NbcSBc6hfk5qVXyEGdZuRgOZlMSsZ/bK2A9fq8fBVic+zvCCI9ADi
d7tFXfzhRJvxvswgPR6i1D5YVy1yeYWTB5qe6643NwpU/0mpH6RriaVfqAtF9zHimv4dDErQU9I8
dy0jACx2RMbBdkEkBYqzTyOU9HL52XWSbnoZYDTmiETt5Ocmn1HhUGlvvxRa9qL6IPSLXQD+dtoB
WTEsjQlEK12uIcfKe5CqMQMKcCx2N7KiIxYYjGG5gAMAZJ96TeCS2hf2gpnm7eTaeZZn+dsgFS/S
Q+k15rBK9UBWbrIRPdI+59lw80GXcC2yXxNCx/ZuPgv0LgAKXnolCUI4IM+rFlyCdC46kbzFOx+h
0+C2epU6HrXU7tKxkFL54k+BQJVuytWPUCgNlAwhixb8HmnK6R6+pPiocIffiNOgYxtY8damBARZ
46LMVW7NE+sosQ1KlyzzvsS8nZnebKH5S3kcvfKRcQ9mfZVUBqFOc5dgJcvT1qnQTmiSNfDxabVy
Rb91lku2JK5kAoUiOZmudeM2SUC7d1hpaN7EurC91mZCHMnv+6JEWJKu/vsSRrKuV1e9dZOeCSGj
Nl5YmEqfYsdEl+F7F6sNG/A2CpJjcezBLpHp+420t1UVWPfrJCst6ULFsn8v/RNITX0kswCQmEQ9
zYsQLogRu+u3A33+lRE/lbmJNjFZgzSVbaSnbG3/GQeDrgX0JA9pzQVPycifL6I72OC8evTPh/XD
dPTD2gV7ABSi1qFiZ0DV5vbzfrRXR141YOr7Vonu9i2TDPtcWfig0VbwHVS5HNp9d653GTNXdrMm
zb3PzswBzly8jnY6FphXioiTzHCeDcjL5JOsNZv7SspKkv9NIMSL69MLl7P6QpNqFl6VXqJhrAUR
BKJ+hHnCXLWcWH7lYvDE0ewFvYaWjWUM3vA2b4AkOVyBo4PiJObw4wLo9APm3QSGfSAPfmk6in24
js3PgsfNoO9p6f1m0d8mDzZVstUsLn4OKszcowF8kKKZv5ZymTdsIRHPRxvjvZHaivYbwiywgq3S
eX2XAhMsfSUpYXGVqM4kFuR6b9x3tnFVUT8i2SD/qRHobiAjlhoymNKNwAuOEsKs/f7rG0Ejm93Q
aNAKgQitxtDI5Remx3luXkwtw5eR4C+vmwHmqOixO71+su251QDMl6m73Pw8Zar9JlsI9QS0iHe7
dzIRtLxpQXML6eMP1PDEip+xKGFZIdXqmDmzsjk8G7BP/Ibfr1G+lhaamkQuM7Lfww479gquys1j
vuDapcZ2i/eeE0rHHp3E5MmLH5K7MpMGMtQlBv5RTDO2itQg9Q2tkoeAQ1Lfe7tvXr6DKzIX/yhp
RgbWpBn1XpQ2cxTU06eWjuW7LSCZYW3bVK7PJ3WItsw+XMVqWbh1ZSvG6bfBjLrsQS/jir0DNSsC
VlSbbkXV8iQx3VpNidFxEsrifj9G6Uw+Hi2cPI0oR9jRkmbb4BOH+pkCcp+QpFlNTMMNudQ4QP+K
K7j7qqCHT2qk6SPL4R6HBp3R7swH/RdTi8m+ZqLoRKG/q2grYX7xHs1cy4q1ZShTI625f11wccie
7TEzdxRNxjQOKwMeLHAuQRhBqPOlljUGT1BT2HD3/xBQccuHJiQ6p39PIesCkhjJ1ITWyd0HVGft
hDwpRXYlY/AckIJstVn5zidzvQqJVpI3D3QlHRVK5zmgDrF5PE6nRilN+YFfyND+H7EQYHhF+UvG
DE7QaHxRO7jWhMydZJsManiOTGABuMRESumEF9UXs+bb9tBU1ZyzS7rQBobMbzRSOGtDGeH4WO7/
VJuWoPOqqDbJ5AjNpoRPi6ygmA1gbj+xZX1MFSM37nswVgSbsvzVkqmizFDOwJSnSFDGWMljsMeF
lEYrK5FDGBZCOqvd2NDZ/dW1gUt4ZTn1n59F/S0A4HByf4++EYJWzdazl/nJTpr2ei6Wz8aHaswk
sp7utuTL91oa/3jDPamQufBNM1kMvWp5Db++YBXcyYX5zXFk/CP6qyizE+JnsrppgAhnbxK2ONiz
dcM084qLRDJG7GIxjF6IT4xmI2j7lSU0up3HcM7zfSOQ7cPWjvQ9XOEdBfIWXFnpXS9keDwRsE8r
4Gku4+oh+EuGuJ3VETPsMKENLP6zT0oD7HNUqQNAF1Fze1MGMjd7h/ZRssS6B5qlWgrmREf5WFSa
+qf4kqI/+pWKH5Z/qsnDTLhgB6trE8bVSv+Vn9jE7BAn3DttT+vEPZYNVSDVVziewtwTo1jTEa7Q
PnlOWZyNQeg2bjmX+kn2ZfUhsDse0rftdetxHNEd+wE+2kBGhHGg7lErU+0TraLZ4n/PflAqCXYc
Q3C5OUIZOnpQI2fYbIDzdkaewKObz3GrkHbN7z6PCaJVhN0R9FN8nDaydZ7L6e4q7e3DJF6JCFB7
Upx0Udw611rhzqaC728NGZEsHptYH9t8D6R6ejhuHKmWrOeApCGnnF2QCkiqwiCG4sVDLKsJga69
uOnJUocJaqzvvlkZfob9xXgSnHHSntxKR+cBgLcD2lFHGf5Ui/VuVieLTz3RXIO3/o+bmBdqWSZX
HrijSj1s8UdYIdhXzbc4a1zoG/6SO2zCpUcZ2MPKPZyVV5UIKQn10AYRFVO0NCCKGFZJi2aa8Xs0
Xa9rrG+thekrfn3LrGGX5Yp9mo4pBVEwqREKqH/e2I40IHTyOw3zT27RtINlkOpbn2ZCriBHPfSS
arVPvU4t4IVn32QsTaF4HO4xdVAb9MCN1EeVQRsXYUEie3JtHzmjZmXPG0QxGqjNk0qgw7xv3TT/
ks4mHOoDNL3my6jCoKrynmbjVR83ZkiMAK/LJHaxRCv7BAXlJHLBs+EgovpBYkoSj44FElip1pLj
eNQ/lalHLN+qemhLA08W6jevYany1G9k1rP2ygk1jtKyf8WnWGJwTAFhSJa6YGsh7N1gfKY42oAp
9v9NmVKPtXLNFuJDOMoDOCaZ9p4OpCnMreLPdWfflplCQYSEDZZCP3TzXyKpd/q15kyCHTfJNY0g
cV4iFsuo6xzjqOSYz6vBhKxaCWY2e4+k4PpooNB/cYWXjdJ1TRI9kduo0t9owbjFjBplvYKkdaF7
Kiqs4gMvYWC9/K6TkZTZ7UgJlEUat8cwxvLaWZnXbqDq7Nmx+G02Oo4UY03C/Rxbk6GhsXjnQXf6
FhCFucDPXKXp0BvBEI1u8bSxVFk2Wr+yAEaXevJzSfwByzRZyBkbm8gRGhYjKOkNxpSBVyvftizE
YjbnlYEGiYbB3EutdXqdLr1xQM/2J3G8lQYKt/x96Mz1CmvsITOiYlbapGY2tLGc4HMUvP+fuUQX
1hRmCCbJIG+vUham8pwN1YzBCgMDegIoalInkHUEPSSlDQ5uSV/upsXLzGHRnA+WMvbpW7b57FZo
y6oN1cKsHSnJUpAFzuU7KjP+oDXrb/Y4IbEwHDeyENX2oSTlWrDfl38XuN8vzkc5Eya/sWoioYcJ
N+l5X0w2HGKDibH1pcNsqFdQR1NYeHGooIwx8IR82zYlVCAC4CHH4nxgfM8I+C/3A9mCCPMb3/vI
Yn3tC4OIwes+ePMevAZgzzjhTX73g6motipQh3RUawFNKAEpb1wuaEztlp9r4dDVnx/7qNWIBzBT
8qlDA0qSuH0P+vQM3tTZ9rCWOooTPR5skAhc8AJZ0ytVoqQzADrz0BiXhFWHuMI7OIZsXjfUnth9
T1jY4Q+QWTsLcmI4ZOOmUU3sZzNUhzHJEiAfUtS267pkor7O4NOtUH9WK7oDDXMXMyhGiIOt9Qo+
eBq+Bt4v8PwWCvvmEvwhG81H3ZZ6hKVj+2Ze096nqjtKMhyHZXpNkyog+QDSB8zfY9e41ZedGkbB
ttCG0M7Ixr9luRvh7sGTXJ6yDVoPGcIdm5QGDBrVMUuCLaSkK6QFUVMPjYA5wBjzSLBctDdkSopU
F8sKWaIngENVQCSDj4GtEI76Ki9A+RUFTuXJVoL4jSMBIW/86P7rUnr19OCbIiMzTzS+p5F0H1aB
7t0SbSE4vTt23LzjALb0H14unEae/ebOivK5RCWGPNXzYo30FGz00etSctpZCFNUM+2cNq8dgRVK
1+2vSFxUm6m3qEBJ8vnzhnmtAERP21lp3tlb5+bJtUpazmZLrDSEhKoZPsf4kiTjzu57OB4whH41
8wBse71e2I3VGGb1IMepdU83J6DX9IVKTRhkRQuKAbNjgM3j00NY2DhEXqnJ8OTiAJB1dGwdt2DP
4zXAZ7VMDVQS/XMBY+Eduphn0HgMeGyiY773zwMLt8BCMimD6mdZ+XCVJgSropwvOUPjfvtXfvmx
yVMZs3kQH/E3/AIdJJLWWVsIZe0LVk4bXoJkVhctvingRw76xZ7vmNcU8HhZSMedyyvMeiCfbTlG
bJl7hQwrLUPtiEO2PUI5LwioNj6N7MiCqwEB8ouxpU9PxeikM5+6wOBFm0DVhuS3s9c5xcsBmoao
BGGRq2eMrCI2r4yknEIMWo/ftkwyNmsnwBc3ljV5imHLu5rgylsW5Fg4nLICxEbwIS0mJphfIVhF
dwQi3pKlTnZi9QX34ZhRCbt7/1JCwOoS13q5xdgyho46wtTB4bv0GtGfig28qZZM7/4domGa/lvJ
C72Jy8ZeLNe8uOO+SEHzK4VAJnEyUyx11ZUbZ3C9gqwP9femYNwzLIxcPMk4nxfWu+bHM4lk2JY1
tHcADC+dhDAcMeemI9OfRNX6YIfye3knTyQv2xmKNOa2DKunCiTk9hFBr6Joac/cgB0nmCS1lbas
XHrjP0M4A8CcwNu86ZgSUqRmsHM6Zuos7dYgQOMBOnGgzKKuVUUNRh0/SWJK6kSb7ZGPYxlIe3Ye
KmZsPjaASLff9mh6zDJbV9O5eaddaAiynnIjE5PpkfumbS7wFWJGCUdJe666AGfomjSHa8Go6g4v
ahXYfZsQyfc39h+KbZS0/o5vnsDp8YeVcIheF4Tvt1LlzL73ZczJIsfk10s8DBLs4SJ/IDm5JHDa
w5CfephdDgV7I2IkXqmRuN/mPe8PEPlzbPX+LClSDbdYJ3QY7AUnzSEZpU+YAit9Lx9Uduqr/9w8
2R7HrpsdRCijyOeycKu8kALVX5ivwMOEGVFArY1P2DxXYiEGTwMAnYvKLnF1M052BU2jMgGnAieA
IqaKsXuz5HSvL7byb8jeqKTEvkCS8ScREEXQMAy+ebPJXztpG1PS9Uy6niY8Fi6zrLYdqCIaPqBn
B9qUMlzIm1sDDu08zkFmXBFAmBLhOAX+kyKIJ5fRG+5SR035dWR9iuG8Rn5j0tfXO4mw0rxB069z
VOT10Ccdud5HA3EtrJzwLhficl3EvJhysNAw89Ed7rqD80GfUJjQOjkcSgyyIkF0vN/+NPBiaLDq
P2YDZOUuM87NZib+2pyVhmmyjPtWkiK2QI9PXvnLT1Oix2s9N4sotTplaw7JigDG7bzQoZiXa7W6
ldUMbidakMd0AcpslKJkF53jPnVGpQfYyHqz08z5Mv3/0cqWJJ6uTXl9rWneY65TWTgNm2ZCzAyU
xa8JDlxCe72pD0m27HxuMqQj4454s3PgBTKINusqHpsISUmB+/Sd1+1MWrCc2oGeEj5iS7Y8jGb0
VHIPMEukj6ANAHyZ99VNH1VOqJdJ0ybzP3wsaD8qyyfliREzWCQOfFd62NO3MWxdZ09djWGNN/HX
W2ybnmek9SqsykCfZNqdJ/fFZ948JEPt2GAx0KfISA3v6hiSBPlNU02pvSthHe5QOFWvYQO+BEi2
ygcu/cCNwBxslsK0fk2zTWJWxz4PWgVxWfi3+caNyb2o3xyT4QzFcsk/uJ+t84ebhrvqc+40gSdu
jHSThXiDz0G3CMq6IHy6eUUfqSjLpl5bwHbdLf5jjKftQe0wqRpBVfREGUXJd4GT+rV+hNoCp4od
9dv+9v0FytOBEX2XHbAN/4UakbhlmY72KVo2HG7MLCpugBLqb9mc6fqdD4eDFZKBHyHS0zs4IL+8
7wceYXt0MjdIQ67qJsYuCDs+B91ubZeGnuwGiBQlyRXDf4+TrEn12ahrozTLqD3qU1gXDZ4qtBXZ
LBQO95RADhpWN5QVD7aNb7nJNs7eOhYFBKJVADMPJSU6ZRqcJ2jkRtqNOOKy+5ybL5anWdhHgDE7
5g5QEIYTuvPUyBgqse7kSNp08ADGd9vD+bMkZML4r7mVJmEsnqo+uhwHkY+nyEzDDvBo7A3uYSn1
VDHzLhRFptMv7XhcFcsxo6GoAiGPZuLHVp+NPeyndsjro5pru+3s0/ZHnLy350aa2InkqFcjZKjy
RkplPsDJIX8knDz9VtRMTEnEUX5y8TPtzj5jgrkRvsNCqln5UuY+a7RFKzROdG7fwMAsaCIzIctC
SSb+KOA3siXNl9tOcpQZ5dW6qfLnZbEljkHzBj/GitZj+YiFFzXNyvNLI4N3UMH6WeTaU2hsjFSa
BcUeZomhL7aVdhhrU/iUEy7KKOJw/7E7yNWjYIxwSYnHhkylAeKCrsIWepoLnp08SDW+4+xJ3KPF
D20PRM1yTy3fU4ZOMNe4gdQwFD1B/bkYrX4q8Od4nQ2FH5gWuR+JwP3INhGAYmAk6Z6djVifOKoB
shtQq3tNJFp3lEbDwSorXbvKGFNPuoy8ctMJceIHrl3Zwqli/pDOhBdf+70LmEem0K4oztrPlZc9
6nzj86AzkG8c/dIEGhBWjSaCB0wXQokfXAL5LIHlFbU8ktns2RnsklrbZz2olC1Je2a5WsdG5pjQ
oYWZJ4FZwb1DmhtyQ5b3LIjK6n98wG6tdbOrD/O4YnbgWyXBb2+2tIwFinQjXCTcqA2THNG5HVQa
/sO9WYb7zTpD+sw5so/7Jpv/ICtslbStvRe+2Qq9GCD92WyrbAwdJgd9yf7Gf+teU+52OKU/gOFC
N+ppRZdxdRTZEWfiSvYkJ5dOsCWWWcojObRVGdfvBFqwlrXrhM/ojIXCmGGcFzv4p+HyhWeKODak
RXFjzvS83G1CtgMIJzmxAKaL2ysBVd0dRSfLKhRkmJsN8PMTTvrRnTzF7NeP25rn0f6cw7Ct2z7U
JM2Dv+jJpeef1x3f2Jc1BT6QLta3/vdPcb2NARSaAv0WnMknMYLeGTD3oAPNYnYGwplXIFB5+DG8
f+T2s4c19UokISiSpNftsZyY0Aw//onEmVbksNKO5i+tT3dfLOI8SfJtphG/qK5EjjbjvjtrHSMI
jIKUS3H4i17Ia853D8CsYs4LaB3L4Vg5HdBg/A6/0IavuAhX+LmRAhn4RcUr9VMw0y+qcHL9kk5g
eXbNkL8XSe6k5oadHxai8hWxcIA4g6KieUYVO5pkjK7EE4PHxyO8YP5phaSvYkVWjmR9b/ZAyDm/
v33xfO03pcEcvmFOA9GxDcitIJVLR4hTxb3+lSXg32gnXTz3BASjXXLD6f8SQB36BRaQKoI71iEm
GIKPXOYYLaT3OLLeWTxmqR3mt79sz3TR6xvb42kjNBVVY4UYzD3EBDuMkRBuwgKkT1zXkIPagvRn
F9U39uETb11uCV8Q5jEZiwPJHBrL4g57Liexf8OZiGZRCqMDLseBnQIcGNuecgYmbeNt62fQtP8v
/keC1T7Stc32qDrv7+Tzud+YfwAMBmHhFTPzsDGgvZP35LVEgXMgQ7Szu3bxxHkcnjyjZ5YnZQQX
798ZdQIwNIlurxKayFcMzZ2E/3D+BzpZ6I8CCuwa6W4zzWNq4SIKluqEfdV2QcdHmM9O3K0YJHNr
5jOp0IbVoAqCKKqEYuYtuHl+vBxcq/Hi6Bllo+gLafM0gKZZ0FPTqeiv2WWoZauVqaSMnt0vm35a
hcpSv/U4JbmdnaPkneUcrAjNQaWEs7PrPMn3dzb/RTwun/K5x1a2TIryqyuClweYcAVJDX/j3JDt
BJjGhMrMxPMh3Tq9s4g5ZkLL2DCA/QPP0ySWW/jUtPZCGaG1vWQatf5QU9/W5uLnWbSFDlMN41d1
//GNC2Fcwezjt36Zxq/JUCzYh/YbhkuhdRTDpXXgEtvXpvFj1Sp5jflYsMp6jiH/Ps5DoufDT2Se
5PQbLmVwXGL6Zr+nk7Xy3LWbID1HgW3hfCVd2AYguJHwFK89q6LsavyxANVEgZqDXoo1pouQDnCE
WhPcmgfdNI+vAdY+RuiQyM4UK1VN5+N76/IRmecOH1BE9jnPW0JoS6SdQG3W9BkcX4bXIydn+4RI
c8iayLAWEwVmXwlipEmLjDhFkWga1/5fkdmCu5VdmqjTsT3GRy2DC3/8EC9uHVk0zYPzca3WpxUa
KPGZuKNkyu87cuaQkxNYtTBV02hvh+4QlEuOA5F6q/Tm2wtma5u4mad4Z4p5yEQb6gRZxKdtS1VN
Q3pgepMm9nV2Ih10yh3ZMBP28/5BaXtzZ3X+Tj8aJdzymrRTDC80i20Kv2PpeZijTLgZYoBt0xcd
1l+1NPYTCKfFv8BP7VQdI8ye5+1MP/bGRMJxKz8xRDzDCJDOYGuyHHecZa5jvCX9YATBP8XOczHa
3fYfp1WvdjrUzjJlLQzCItiK1nNICnumb4krnSCyjx0AwmZkmI/5KZu1+lstUZHD6deKdk0BjgpJ
OZ8l8pbroOQCWTx38r5zXcAyG/mBDvUJ11CFpqM0cLdu1zt3TpMPFAZoSBEpzsMPBMw3kyWC+eXf
lRguvNdlpWLZpUYWhQXERE+bs3mFXcCVuMO1KX7Bl5cNvBGZVYsYeU3+d238ijOKoavrM3tB0ccB
Ttcy91HP3aZKWiNZ0SyH/hbXW8Drn+QvHOKgJk1Bn+YCzc6J1riDdl5dVG5118y1Mb8ej2hfmyUy
HMAa6OK9vL28Q736qeWgfeVtSP50f0IoXAYMMJXbvaX7H7PSZNvwZMe0idqoRTh6FzQytuDtVxAO
hXVk9fJGL3UC49cmGAiYhSEiLehXpWJYfk6Ms75v98LuxR0s39rSG3qjxL17GLuQY6Yf3XP0ByF8
O/jxpJf48Ke0jHdPeHX7yTnT8cDxmqqQWxmICrGx8obGe1OclLTOEJvZwO3egps+cFI0oWqf44Yw
7KAbDG7AvciajPQ2Li5vOfqkdqSj8lmhtFT7kP8Lp7DSMcrgHvmyb5Pap+964j2Rpp+Swz16i5O2
g4/+em0kJrtZbYvR723BrKLCRotrem+5TMSTsWj6wwnOVXM1LwTOKSkC86As864HbximVzXJOnsk
fA7QOdV+3z7LBPYDWfxOz9x8Mz9VtYUl86fPUSaaAXCsxUVaMWc8emTlMGRX1uTlmwRqLFvWoowm
iXLL5GlILZkSgrnqmSkz8PwRKGlDP9Q+M+n6m+fpz7WT6vYzGNW16W8Y8oz5xQxBPQltTIyVieFf
ddyRyLdFxLdqHZwokGN5Ul7Qqdu+iuS6K2sM4lgdRYm7HfAGrWvnXvNEDQfU2Ny5HvFmvPADokIo
/VJQ2relAjmQ/CXgLlVh+ucmMwpoOI51DYlQgTq/ozygjxJzHhDVdBS+wN9J4wlPfs94YfFLoVTZ
Mu/GlLFUbqBSnUX+tZvgcp0w0iS60aaxyG7ztoz+718DgWNv/eUroDLVDObG8w37qlVhtxTB1zZV
eLGH+x9+RDAvKYB9zuhvZoxgw9VKyjIR4zSZwzWjAfYajcHD05ytAwB+dk+Vxsp7VWIjLq+nITzD
frodbCDE5xsMs+skVGLvMaMGYiXdpXfa5Wejz54WhiF0mHx7WWHng4c/mM9HYwyC9FdKdPCiU14t
n3maMER4Lpbp+nvOZuN6kk3+yt9uDXRhbL6Li1mKKzjN2QD09YASd6z456IzcVQxGFkC1Cc0TqyP
tEmmUzXS2+7Rm66eHGBBfu3b64Xl2TOupqtdRcZUKVliw34Evt5RU1ToxcnhsfRF7lrdrzSIoIy5
2FwvKnxq9T2VkcztDqdDAtkowgwKGOU8L4YJucrzjq8rBwKL9l969fwro6tKVJez+sS76mRtai1C
M28P4VZA4Ljla3qRWo7Rs/N3xRNhWISn4tYp26LeCQpYr36yIk+BE6A6AdyJ7s4JdLDU6NPBjYUh
nk56jUzO6KyylT8kcP2UkGsrNjCVuh3E/hpHgyOR3dvJltiYPTe+IaiPTVi9kRZCZdQIDwyw3lEJ
GkAug3sfYv9vBebq5DNiJB9IMA80lv78KPAL3v9bdWoppAwJhErJmcUAoqmeHuifRdCXzL2E7iZk
8w6yeCJv1MUrlgbImdfIRbU3E5ZveeTXAGuS9LlvKAr90OZXCs0qwA9q0F3wDze/WybfxY5dFuFt
84B1RNSVmW5wwxInL2/TydFv5WWaQQbWViFpN9QN3ZTZe48LGDmDJsR4dNRPdBSWVozTPxk/YoeV
31OiPyU6Ojmp7p9DQtFiQfmX8uA2oYtHQZnwmV7dkjFbzbT6mFWaNPrGAsYUxMld1D3fFJjTHeZQ
XjHVWJuqPL2KwUhahrIYIzmJ/xXYDyzl3r8y0+PCpFSKjYHdB29YRZSHu4CFptx2PYNKMNVwF+k7
LbpBb7oAP6kPb5asq04W0zQaFTTdzV7huhBIZZIM9KYn1bSD6/3DJKYKgTeOelgXQEeIAO514HSH
6Vj5EVmu6Uz4TkAS6UvqJ166eVZ+6P5QCg1SzUqfhq/MFcCDKSNTA5RBKbXC9k6BL+TLPeapkfei
6dfYmC2/uVV1G/2ZzQOEpP2anm1Emz3ZCTiqb9HRPl1JTjXuQj6ZIXlYQIN0J/pMSDpx/JsEj7Yr
etJqiqQx4b/UdsM8DmZ5BGGuMsduagMKbNNw78igjsVTvu+UL63cVvrcu5TKU0CV9m+4sunhZgG0
kdze5UuIJyEmSnIeurjIKUqPNs+2Mtm4ewWw3Fph78YglTVMgLHVQkCzDRVDhcLA5ap8jiCJUfrG
vSyvrOwU4IJNQU7ti1+0BjtTdRp5uGFKkkxNcCw6gMKmDOa3V0ONyO4hnjpqkZIklv/L2uJqNRpx
I/mjfW10/DWKNt7CrIg/MTG4BHdEybr4A0/VazJzksx5GZGeFO1L+Ekm7Gdi5ttTeRvyKvogEXT7
ZyYWrNiNO8aCj2skqN6zDV+a4ppfm8x47mzNpTQ7qPE8l637csGiCPNS7ctGyYGyjcu504/a0KYx
smpqqaO6L6vpnF9g7iJwIvy5JxWcwUj9MD6YCmw6qV4d/D+eEnKT4ZbuClAUrv34eSRtjxmLltZF
szZtEpKH1zvMnEH4oi0VxPKvRm/uNHxJYDrBL1KFo51zCz4uroChNdIlpDHjD0lNkTY1GZYIJ3BF
JNo5Cfu7oNtRsprczqkl/LEuFk8FhGup7Y6sYW3dfp5meObOLY5KYz6neuWjJCwE49u5meY8colI
p+2YiBgRKKMzh8hIfPHkXBw2SzW2DvaANr+WU7MjMlG8F6++FByDT4Bwiod2M/p//kdf0nK9MT0d
Rq0Qx9FIxfyIRMsqQIymfvO5IXDA3BC0zWZJierY051s5yQRQTPx2Gg4dRHybuhAnihhoROa1qsj
WJloNMvdfiBn8m3f4zA7mj1FLvMC/D7iQ8SofLjMfqO9jsqsp83CAJIGubbmtaDnMtaVAv373fA/
iMquHhGGEdlj36FFmaVdoK7kQDQDcn0jUC3Mk2HuvCzs75/wzxozh+kHPQ3HGU0/fhxVl5ejLxZ/
yp2eqCOfS999AO1CYb6+NyfOucJuJ7K3a1i+ruXfjH2m8ezZfx3KZxHYRXGjKiYa++yjunzArIMr
HZsxSyLq0ZYdswjaLJY18f+/O4+CvKjJA5wnqvvG8H3S2cDpOas5JVGbCNGm9a6RwXtgZ2/VBAjr
O+EYWRvvAi7W9v+NAskfvk9tmadj2vRoGvm4GxsjSjb7hisU4V8giSG918F+pvVNpEOr10iDHXJ0
uPNHezHPqtrYFFhj0cbElsFO0ajabEIt6Am3Mm9JjL2iPyw4TFERUhbZSaxRkKCrFyfABYDEd0zO
ia1Dl/NKlyOQ7tB90QPat038umOt6R8MURcff/oqiqOBnQBAj/O2XfRu89eN9u4e5aOrw6A7kU6x
z63wFi+6qj102SajFkuQDhGLkI37lhutwiSLJYF4V0+Du1IkIr0jA2+t0WSGq7ScxWjCnbCrFAgP
vuh5WfWmqFrL/gDK9uYsMd/j7cznS1F7k9zo3OmfsKbOpmgS3DQaWZ2H07FBhklFvLbc79DoxodM
/Ofjl+VOBV/KhdOGLywf8dbCP6QVHLjzwcRwfLdH/NhzGkxxHd3YecvVqAxroBBrnCG7ldH+F+M3
vsVNksvlN9u6xvggONkq2c/JKcphxPfASNBCGewcWYpOChMc/FCRwrbrGnkWjqF6Z9/oM2/k3IiC
D7NAcvZ4V4y9b+3Ak9fDQ86OBJMtP3GR9jYVskjbq+7fOjTV/APDJtqdDql0IP3pxt2K3niMZEJ3
c81uKZMuIqBq5wEmS6ms5zAEsiMWDz3SU/x1ISHkcKeBZy+YBiM7goZpwpp7Z7La6qKQM9ufL9Gg
Yf2WkzE4DTrJ6H+yKtmUR5BSyeydGxFWABdQTXS/ZjZtd2isRM1hfb5LkYrzs51FWWBQmbKD9gHf
N+qekcoG0Dhsmryhuf/gK+4ExPDtCTJGtqK3n8lKoKoYGvxqsbBQFWogCGxDOkz/CXFc4RJtnt/V
vhkEP7lVmx0EFlhwka2sX95iq5KeUZ6wKfPa0L24kP60hAHLw+rBmnTCsXdURQOvvMEH4uL+fE6W
ZdHJ84whPLE9rvL7B6rI4wtfaIKUUpqLZzTUy9DmTnNR3/4ooNkh3scZOhbEP2CdMY2pDhQD/F9i
+s5kdizZMCbhEPyS4dz/O0eO9MMrado5VgJWkabPU6EW6h+xh0yc6/wjWFt5OLzUV7FZu/ouQHHO
eHNow0hz+TZ5dS9Zy+PU9QFCpPDPM4qIIRUEYtAERC6+oW0iLMBBajzXmlPwdNJOf93GWpNuo0rp
tqkEfLxQ+p7oQLCk7hEbuwyNhJ0RAk8E3WP+hWqh4K8jPI/g0cCUSiAC5l6XZRoPl8dZ5UsuilQT
T37TEl23zCNTkzSrSFXHlWjwqM2h/UYQiSqzL7tgfsSwpddkvUWXAoUnWM4KUlgrPNqKDVeIX1jT
aoA+zUEAP+hqkzX8H5J6yS0mVMHq4lj8hC+OfVVHvFqE/L3IqFOOrSDl52TEDuFAELywzUagRK6t
pkeuQy2gJybQ7qTRrHhv+xM4WCT5Arj1Fr56m2w++Uir3AuSMnJd+FCl0Rtkz+aIMAG1Fa/ESugQ
ftrTfWe5BtkzQzykShakuQSpXFY1qX1MUw4pN9rXv+MqNk004hmiNMh0m95VeS3LgZuIdFYA91PW
QVDwdWmkxWcw3VNpqvUjgZ4dWMimtKSoExHbP6AMowE4YE0vcAJX4719TOZrV8C51xaIVV9Dhlhu
0iXVXsV3hiPKsV5y5504QB4Nr2U74SE+9HfA7jML2Q40C2plks0rS5GyXLkFVg+jVPMOUZ/QT9GV
ehZeBE5DIFaXxYe+78xWnt0R/A351dBARPg8r2VHBnS1f2wI3XYQ83rwQpfVCstqAyIqpqjc0ZhX
iApL7+bZ1/yUg4UBHkbUca3QJnd/nQZ2TXgbW/p+bTYY8Pm5bA+t4xUEClwegJL0Rm/9ivBCNVQI
Y142Yr9dtirZJEY5drdTod7MUb4lTQjhEqkp/h2ljH6v4UJo9wmtOzwxvFpbVp8h+DEhjQlpjvGe
PtgMFfKCho5O2K0P2GGeyZNiA0/lWHREfxAJTeTTrNdVluiSAyP6gB2SNI2VTqcoU4RkbBhtgRz9
hQfcvGtEm4S+grjoVmHJIe41ApuuI852eWimCEOsxube7MfcCzgjodvQrNh1VDfQI72flIhenUz2
X0Iv8ZzFETosP1Qdx5POBzn9qW6kJtownmVM0qJQWVAMG0E7xdADTpiDtbjuszG10OXGfKtmmjSI
MDGEBBAZ5aCF46LuEN6l8BdgZR5ZOgaU/RWM86HCHtjDhDq34YXOqBJshxY3+24LYUkQPnbUYqfn
1XH9zq/2WiwsTiYxpLTPrJggnHyEo8Lp2r4rt3DtRn4fTs61oJ1XKSS9v1h8+5cpXzBjJ3OOa80U
Tml6h0Kbw0xOAK8+AZmMEAcsQa9Tx1Rad1DtwjfmtggA6mtNGsJyqFfXHnkYiWTRT/KjWytqYVEX
mbqp/1HEsKZqS1yDZ1GiRC2tKPq+teY96J72hVGGcXTVyoByRdDXgOwbegYS/4ij+UXz9VEew9P8
ocEX9rDEsr9JaezGECT7XIhgl89BhV9szjoOUiEJvPH10HsX90B8vNWm2L7qRP19fHepRcq0lUg9
HdIcqALnko2AdsZTII6b2u03hkznHz3BCb4oYqN90CC3yVSSPh0ahflwzrlk2MgwrNML33rKBa5Z
Seko7g6NLiqVgSPJPE+/G+ciknYSwwQbFMXWrvbZTajnsw/1AYycfxJTLeFwdSZY6FJfXTh787OB
Y25vGZu3uo627/4OeuVkn4CS2I5m5KuSQoCPz20auzbqZIivlv5/YFIzQNdJTqvjKscgB7c/WL7v
1WyqhHTxC014KVn45wGFc6mYbFOJShx3oPgwM+A7PND7DXAcJa8U7ZtS8VtIHhi0UgJg/pi9rkOV
ydyV0sLMHwgYLf5PReN3cRe4bzP7Jtu51BDvOd1HD22r8WAdTV3V3aOOj8NHwC7rG6smZizO8dnn
NolyrcB35/uFtRBWgnTpYrEWWWCJLkEabHO83MbayE6X8dwkAhqZQm5x22QL7ihQi2DSl/XESYXQ
BcVTUKuX/bxGBSFTVAHvDqC/3BPo6LbUyAhtHyCdcDTIvsogdiuDgeN0LPYq4kxprKuP/LBgjTNQ
W9l1fD8sZxpRie/IqW4GRv4sDSEft5HhP3OszsZevS3kQf21dtlIEPIal0AIGrB1d3TW01zys4Xr
JgJNFiWfsA0rF7VTPbRnGJUWPOTWsWv4N0RiiBCPEhN8Xxjes8Rmg6xgN9sLKJAGEZfJQ7Xzfq1U
r8pR6taNVYIraUNWt40XtMQbazvCshyK36Uy96p0zshajDzf5pmWCSjBpz8CY4psgz4ayCsDrrfr
bg9TCM1kEkgRXnn1ljoJORa3grQs4kExulbtKv2q7+mxmqt8MvQcVbcWNKWHaumTjK9Zr1m+fkVN
OuBDIxli3FnP3ZjSd72C2mmEhSJvZl7FNeVNL3vP/pRUfNJ6Px141SCjJ19YGn/KD2CoNKBPTTa3
7lk6OpeTwLTuFNyviSSUKA+p9OLHvrMekBmwRLdic3TSmnsOb/WqNcAJV7qH24czQBoyHc2BkG6X
mYuj2XadUlFNJI8dRLHkmZQgsLmMBKg4ytAlCLwEWW3lMR/E6T0f+Vwo8dbg9FnozOl5wTCB+vuG
H2WBtS7GOKEG8wEbonSZwHf2L7bHb8EguD1q0A0VAa/PPeI4VyYGlYbzWH7EGKLInL4JKfKzmC+H
TlCkNHxg+4vgsmFeLU92aBgEoslVuG/9feK1Mwe9MkZtNwBOjtHGuVO+0S9eESgxqBP8GLnMcdne
Z/0o+zmcufI/SVOkqQU7aKFJiSpm1DVComdgAYqdPuQgoG1grdz/5u9X8QmHGDpt0CzNiiVmVB3b
6cTxMpRw5Xj2Y6uDRz0xtVNjMoPr1izFoKaqptU0JidSpEBByZwfUDJA4duevAAgcHfOvxAn5l1f
40mqHHrqtQt7W/v1KK8anSnMxwU4aSn9AaiXM6T0677AYVbp/qtMUlo9nhBwRXI+qcEusgfiYQkw
fhJIU1vHbo7R88mFjZBQLhI5VdnDADqXOgrLgvDe6wwML95hZAc+QCJtLIO2da5BPSjT1sh6nyy5
AxoazSykgOFCisaMBu4RJzo4MmeT85s+nk0IcB00bGrktnFu8VYuAQ/SEDgpydXscFkB0vFWHRbF
gbxFKbll4xIp2yKqX6gjsD8yoH5Px/ZeoQ17jTa57oIGVfuZgEFTprsmECsspBxUgOyjLhB4J+uF
KHztR8rdj6oprQ433IPV0QM1IgSHLnKQ9ECZO1jt3L4c0E28fXYngN09jIWfbKAtc50N2WiKGO6U
ja3SdMVbkB+NcCDx/BBgFHmRsNeWIJ8P1KK8gB89H4OHwLoSWBYDKytSaQYaB2mfYQHFk6Yn6Ech
kghQtSTtm6sEL4U5Y1bEdYYkQXfG9YVm1MovOFjoCJRc49QoZ6rKsSYUAA4vivK2rwnx4GRlN86U
8jVXFmoEm1z20pKvx9Lf5+s+4AfNMhdLB7r8PcQbgagkZycObPxN0cSkUkdsKWRKSrwAWnTYOMR6
vwJxhe1TW5qVhqFcSS/cFXzFPwwmhmi8qL5r+qUgfwvQQfzYqIbtcnr3NJg1qAjRDQZfY6M4WAOA
qLda/fl7UpDlwrALIZWFIszpmYA2vA0FNPiNfscp8tZAb6wkk/aQ+9e10WkhxTwjljFOGp7o3SIb
spEjJtabMyRBwdAeZ0hdFuHi7UO5zxLNa1wODt1d7C5Olx2n9FMQlu5XBt7owdUtl3bIEenMERmv
/T7+Kx06o18V/wSk6jRHr7A6cwA9GH0OdA7p9NJB6D5AZ6agdTRWtYWExaOapJa0Ar6Q9dLEuHgF
8cdQQMFRKNikoGrXalEqBiJnJOujXiWD8BSuPWnjLt52RvBFY2vTYKYU4ihCTBNLdAndpV86HObf
as3sGNWW9gXxN95vmaoBiL9yvqg5oe/kV6hHAlaSSFd3OccBJ2H96jv9EwXx/SWL6S4SqbDqUrhA
UGQnf6vHRidcAUkCEE/IZOGVShmh62s2aw+nBuK/UFplOqHEqNOCZWww1GSiLDfOoyGC1yriuFv3
llzSL0H+aBPZZ7bXeyq98KICjDucBPKQjL0ZHhbtPKkKIm6uFfY4E0aKVvWaMzV0bKAUp8CjkJ0e
827xtcwzWmVQik7oYuRlqwavOQZrBShOdnf6pqN1bf3d5tsEjNyJtI/FNpvJUaopYjCQHu+81sTS
79UBut4ljrnsMPlGzR3HhksFRnP3+GotHhOI7lkBS1UYaDNwC2NSjqEJCNfJmV0q0t/qLdjT5KNA
yPRz9aFVZRUjm14Pt6pxL+8GB6FobBo2OH84mOuZl2jsd2Z3CfMo1vdV0dsuyrxuBlbja+z+ZL/b
r9AWlApUa0w3xFEQ0yxiCHIwfGjM8rHBbvJoOr0nMhPm6J7BaGXzsHrNg/5vNC+fv6bdLzeTaJuZ
ajNSIuX0UAFLFaytMAupk486Q7ja4qRY27Yg3CdVMJ3UZBPhxrum+4iZkaeSbEvJzgcCPz/g+E7O
ad7KWsqN0chb1PKCM5Cg3f5t+bIZxApPz/zirv7v9ichoaY+Sbo038ay2zYvIgBF92mwefcaYIOu
wPdazHlWCSnNCNNekUoOhqPfGBU2xDss+wwMRIt4o/WeJQqXVLRNDtjNqD3FCsYFUMuzBueEBvYY
vYgVAesUVxBa4rF3D0RuualfSFtlajpYUN6ByDPf+Fnh3OdKm+tmgZgF6gkS/eOS+isD9q7ECXSu
vrT8G5houxQDDT5VBWNGkL4XQ9VOIARGbEEm4MdKrG/9bwLHjE5VOak6j4IyjujwXVfA4nXzL3mV
L+BF+23wr8ggVbNJmDz1RP9FIZXx1hp0p6fJSzyz0B2N9oCK/tPKsmRYOKE9aBOwKSDSPLDeyTI+
TwEu1vVFNHi4aFT94VEEF0Xlqi+o11aHzr59LJ7v/IMZCrfw1Z39HZtRujDctNOL88U/TVpwumRj
ATmUVzZoilPShRw3W0ABgZ62L1voHsUMh6AYyWYXX0VBFldYujTZ2/bw46Z9Pt9Iuj8tv3GdAX8J
Ebbj3E//+OHGlUoLclkX8UHPL5km0dcdh8lQKhkCF09wbxgwNGWz8eLPoKltrfKzJ/6h+USZERjG
0wiwym4l2yS/8W3fyd6qmTl+fxUe3E5Xz2WzJjwx/Y0EshOVcpMl2h1aTk9tbLAvk8cO58QiSxRi
LaavjvG1OoGfXkR01rxa/8NJHQzt1c8s7W+IqooyRXGoX743f9SHWr2hrZy+nRxXW8q82DBwkWE8
08KrqedwzsW6+2OWQ+ESnur6F6FHWQsLC2pt/ZQcMdajn1aPPqsCfGUby24pt37mEZDg28ZELbtV
6TwCN5aLLpmJDzgD6109VGpTQv7EODAOtdRsDdpreTP77+ShxSM/HPCG2ap9Rl8SKZR80GPqaqRO
NJfh//fJ/pKslDG/hgxl4Bp6F/f0FVcs5H3qJji1+5Fk137kJfG7GC4bSHF52XZoEVFpEmJNxcER
ShYFc0kQ5XC1QLjB3kvZf3xA70/W1anb/QDDe6PoWx4WNKIdCiAD75BXmkXwBStAiOVQj7Qx+Dyy
Caoya8k4Pi1jg3eqMR4zBqyZW+P7N1zNzMhjNQmojjl8XJnKs0/vFT5OrolDFrNLniKPK8eqqJhZ
WlbjjEiaKrR8W98kJgI9xh5HIE6NzYQpQPlBAEejtfG4APd3WGIKB/vttGA5lPrv5Q+PTEIOBdHz
hA0iV7CYzQq0mLASj7+j5uvxj+vF6QxJ4Jay9Ok/Ise8w8z2OsH9mFoRYjCRuDfhcqOWf5WPHFrT
aaYVwrtp+BbtG+IC+panBijfccqoubgoyXcNEKu0wxYTx+M793aSPBUZbh4JEjHPVdrd2h2CJy4a
+lgoBwyJ0Fy2i0OY4ZmyOMcAnMXQnblK+xBjTWIXhUnREi/DNHx/RvjyFMrcFMdGrkDL9HaNeEbP
ORYujUZceMze+qZaeQpAO0FUTVWKiqfr8Mly181XUZkGK/N1E2NNb/GOcmUZ4hIuKpjNsZ+X/J3Y
EXLYltK36d51+8c4HR91AwARS68yeYiRWl74+SHHyb5iuCMiiXR2wakl5mgo0QwrKBSujkoXKuTx
UGj/REaLKJQt+YlSTMVqC8UbtIcQdvxTEiHm8AzE625eveBw5Y1sv3PqdJq2c1IjO9xqmQW8vkdT
eaiApt1UsYYh0e+HJYhRWKntVCGQLY3JkMYazS+1jz9BnjhucdDj1r3uI4hkf/94PEgYB5AcU9V0
zPJqGwtfk797Cue3Mcp4klw38ZODXv6ZCPLFEWbWYITC7MV+1BS7XdlhzUoB2j4WTnTrx1zu+Q3y
qPe+6tRGiR8jmvUtRLk/UP1RttVGkRDWl2OH0KCHdAMYsE2mx8k0l4T1cCMATeY4VUudgD3gLaJ7
K6GNPG+Pc6Suwm9Is839KN2Q8jNEkZB9jA0vUfYas9aa3KNufyxpUX06AEoj8LD97k41Nbe+AYEi
QQ7QSuBn7+uu+xlD20VtRUAa5/nHKzBn6D0c3Py46PvR7PJRTb0jM/8As1DEsRJT0vndGQ7qefeQ
sbjy43tPbBNMzbf5e1ngcSM9xTiZFduFd6xOCJHfS093evVlnZeSuprYcuK636rUFeekuL7ScL3/
VmFT9gm4HO/vPup8Y5KZE+yZsLwwlqQQ3g/9jGOIv2bW8qjgoLQ0ywRgSaJSttzt7GPNFoBozMFg
ow/Y/7G50Aa+3M4CvlAOknnuD2XAdP8YjEwmCd6Wj4+LSlls471DQuvrQDdAVEyiVQ7GGedWKeOc
8EBorGg4ergAtv79jwCEANcdsnCMM+5SM1CB+lvVsX0Et2oR+CpV3qeD6vqanj9bpDG1zB8ev4Nj
8yb4i/B3fhNC10pKNLEoxTfdGOd2HnsPWsjqQnN/Leep6KmWl/jrZHCLAQteLyWxD26neLudiTJN
374MzdaAJffsnwU2zWOkL+isBSdhbaqR7NiTPgdIJsQu023ZhF3+dLUPZ8iUH4tJtsQB6+NhKGnu
IXJOGUuZKyZOep1A7zHX6YD/4Lr+zXdQ57KuSTRfjOBgvW63B6l+UxYUDaX6IAHaG+wF8z6TF5Hu
kzFox6oYTMf3BUhZKDyteZekH7NruToHhHcNoaEQZuRkDAosqUTjdcDT+poTZLJt7ml8M4xqYnD/
Vq4VAVKt3/TdUrMOumvjVNiAXBLtzohac5Ge14Rk8AWkrHnTZZLxpP1tDjj0OhpbLT9LpDfe9ud7
BiLq5ePoAcS2/pPbhwvg/z//N0i7zgeNIt1xeapmjOCFAEu3NV+BoKL6cIWC7gwWTe1q/Ahn03Z2
My/j0c4/YRAnYhZ5Jma1E48c6Ijyy9BF3HlT5bOhMEZjIxEAaMrmVnY+Jy0TyPwSdeeN88yc1pmR
ZYE0LqmC+C1nZPvBdPA3lPtrbDAUI8Uzs/BEhUo2pD05jAcT1RGJtDyKvdubuDiEGcP+6RiRpEtG
9XJNaPe+AelIRP3sMgqIqMmmCULaG2FA5kBEYqdzSIpAVLJTzPOIMkTwij+xtIwglSfOYUaluTAQ
9Zg4wKRGbiihvvSWS5LyCThJavrnzrDY1qYTY6N7FezXVQtvePbUrhYDz4cfVl2KNGT69Vn7YReQ
zjJPVGA0VXvCRCKtsEouTnF0Yw0i2M2NVVXtl4mawrU7AGzWhcxUQQXnmTuRWX0A5Ldisl6wrEb9
LXNLb0UJJ8RX0SemXdapvh17y4DY1cCCwIBMTZa9SU2mHnJgkMg/GHJeD+aHbx7PKtlOUBYfY4nc
UJfjAXZd41mVIOjeo4LZWbgG1ag2rhHQehdi8e6wDFYDin1zfvYJd2P+frGxPaTm/EwPeafOCZJL
ZAJEIvqXS7SiHLuQT9lnZQ/rbIxq5qmyYj1a1s6iHZgK0wbOJD60e+gTwF1fbZ1PsIcLBN+XiBqK
Ewlp0vTfn1WfGyE104zR/bffP7bjrEwKQKIsXE3+ADNJdK4CLwS/SoJP5uYnZrbVAbUCb5yql4t8
dtaKPpQLWZakIB984zUoc+IjDgiZXaLZ+iaifpxvjFxVEJ+z5+UDeNuFCX3r8Gtkqc1EeojbMXYa
C5Sxk01vAxt6k2aurZwSPLjx8BuOQY4OAmHFB4AL3wflG7MkNbF1Um7rbOOSNL+2vjR8bX6TWDTa
GS73c76ym4GJXIN4k7DgTZ8+//ga92BndB82faf+9EgYEyZPSfehwgwdAkybni8CwYzX1d5RAEi8
cephKy4vGZbNWjblRiAZSAaO3tocdJy44cwEBwWnvqYl/ZeUfQL6D9U4re7CzhmO8ZtawqQkf49f
nCYA4KgTjpAZVs9MUSCVYz6jYDVhr5LO+MfSFKh334rsB+WeDnVISGLc1H0xoLyDpbOv+g9gyOqm
VK8zzohGGhNpIlSlUCntD+658og7ZTPC4Lbvdf/x7r4l9gNS2kUSwFLEz7xuXn0hhCgQprUfsHsL
IRCnQZatv3q2qx1s5DXj2l07It9Paz9ZDL6WPE4BvK45v31DKY+iaQ8uZnbdOMWMN90NdqPipoIj
01WvqunF/hqnha3ZUMfVhQ9hphOMQD4c6NfJrCVBGWW+dt4MdEkA1gXHrNYcATZvjkbMBdLm7x3u
r2QTXio/Mx5ivEyUEvJ7BDwGp7Czg7P3XIs3P+9vowlPUrGXbFUSDX2eVkxniNOy+MKmtF4dK+Vf
Dx/OKY+RTE8o0TNgpTCN/LTp/cYjTKEwUH8R8saDjUQfyEehu7/0+iipoR9PLKtY729v1cRarmyo
jAfG1lxqiMzTImGVKPwx2epcWdjt7lljPFG4tCs5pOEp2sYlFimeMeMLJ5dpyiX3kltgLLnGOeKG
wQtFSYHNrKQrggScesYQ4jQtaoQoFhK0CqXF9hMDVC0FVh5s716V3/PzzyyeIGSG8Tsq1xVl/gkN
qQbSP1kFUC8TUktbgGjKdXOr6p6DjApoqnsy8uuN/qw8tf9g2+a8X+j9jpsPdUo2yRQp+Dq7v+GH
ywz809l0jWt9WtQYVKNKsZTn5WGjlWyHRtUXtL+SxucxWkUKbdpfw1JMuq63ePA893YYA1TUevbi
CUZBtL6WNXIKEIVoGUBiYkPmUI/1+ZlNDqzLcnKoEqghzWxeAOHSGt76AVyL8sRoKEvdMrKfjzYj
kZZ+ul690DpALngocfAlMRe9pgrinPUyZMruFpoygMGgYGnLNwNzyRG4qMFBRjYCsaoLuTxBum7k
YzGeyB9XkRDGScPKqd42CsVYviJF64/oXt3C4wle1plVbERfCOUydXufeEzJoAS5U/Dd2/nopAW+
tHeRw5TZ/3IuaPkdqKMp8Sos8CNEml0KvTHfCDq0v991KzqtaTJxtGCary9ME2x7o2TeCvjkXp+9
p7eZJefJt6mZ12cbuqgm4JWwJHWXLdY3dxEQfCNE+aV0CSTzV68hRbfqy5PO8qWUECkGyxbRYAJC
pFMLRamluw3bUmXx7bNCykIsTSmQgb+gtEPfm5T9SEGXRt4nOzD+F1iCW9GvWNQNu+OYX7QMC3+v
ENxiH1htF7c0+EH11nSQN33tGN5uP7O7/wyxsozoxXyIRyQW6waGlubaWLpyFFQRuIsumITX0kSw
JD2tv/eWHIWchVmiUBbN23PMm2P0gB40JrDbcirWDNXEus+yE4WBjZkm0qTo9Y25llyxp8KHRsaV
2SFCgrME/6o19lZJ/qQlRvbJEdagTvayI+rVse+WLPj1qIWbl0cfFBcyd9/64LiTo+jPZ3AFGrM9
TUGJTL4JovTGtiZuWHHCDjT375gx105+413E5dSLA/zopeuRiw5PtU+FzkBdpQrb8PcLio70knOX
uZRZWIOirvAnSCSwneI5AMS4lC6WMQUyCl9U0R6mwTvY8LcfAIhV0MfJ3uJlWug0vi1KGy7TRW63
dATOibeU3YPNYaGb4dI1JdTv/CGnhptrf8HhktFqWkflkuohn3tvd34FY6Wr/WDST0NJKW+G+yvO
IErfGRFr43UKQuZl7xpv8XIwhkEKda74C01hBOucWcjQUFIh3IqFqaDf/YYNVIp9vfth9HlsVIfH
EthO3+/2XNcJaAJKc1eK3bJ/gyMu7wndEx8UksKafZp4S9YF9H3tVsIu6c/1Yo5wzrftSGI+id96
LLpj/Pp0iEcKPytkAA9SzioyYE/vq6XaTKqtZWeNCXNVCnJk4qOX7IyLD0mqt6INgh+t81GEMvoZ
VR8Ypt7dKyK2622N9GX24TKE38KG6+4BT1qpWw6RW0P9czLjDAgHdgRAlweHIpnTD34fIVeeeQha
0U6Se2BdnSi2Qx0lHZdSfpPtocfhCGnil9EPxlopiBa1EgKxqLn68bS9vySXnZ/9/LfbRLWXTzfn
Uwdj7l/3kxeMc1o7kDFCi6C7VxwldJFSs/IEIHoMtvtWs31RoxCsC9MfcnQvjJB+cnLGWb30JdJI
VXwG9HIxwtde25Owqb0C74ZPuIfkoYFdURIhkOedExsUwlp1s33kOhYebLoxBUerNmffiQKni1tl
pV7gat9gYqxKBYVrWPCUoFZjZWXPyrj+N2JoK7QpftRZWTB2vqSrDctaCSm3dyq63Ucf+Fjfahgb
sF21qTQ0qwA9ibFa7Vt3JbElSEoaUD9UplsIs2zhdvqhnhKBJgVLh4RAl1ZFv4/bnoT9Zx33YSer
/7fKp3ZqAge8Ik53qG0l6HSDN+IJqdjMIXsM5sONmPIH6avlGKXHUcy5VAMynS5mk7VxHtanzWuw
NoBHaVYkdIwZ7R9UTowIetfbpUPf0mebXLQmguI38n3z8cst0cqdvVQYXepMuZj8WjydBNLGG0mz
uVVEDdJJd1QfPAQCPLuE4SECyiB493MSW+y/6hKwYytcFuI5roe9/AV47I4bkyr4yT/8fC4EXRRb
ussbzA2FKgQ1uSZfScJnNMFOFefdNCIAWOAzdeKmI+aq1JAEmeHdt6hkmEKfqLhhE/XwIaFne0AT
u4sqGLU/bG5Rl0wEVpriLXwG9jh2iKtZwbspMi0bU99Q1rvuD8KnlipFdYst9kIAHxc5qOgKLgiM
VCL9T9wiVH85P2N0ZIBgj8quLEta32Cqzs1MHVQFUMf4S5TdohtDeLkRca1FNr0yE+IHRQDL87mo
XPC3ecVhqhKlomj/BcVT/NDoOco8OXZASjXHTW/ERIXeebNmNqYJySrGs1OAkqhSaNklWRiuNQmq
WURtBBUo5KO0ukOjqqFQhsDb8c8l6rx6yiLlj2K+EHDxOSK1IYEDJjWFKf/TPq70GgAq2DwIy8sP
nvdQLKwA21EsPCNTCnKDOlDxqboCF5UYYmZtXq2RxewwCLUL586MguFZ+MNs6ZyW2GWMcenLjUGJ
Kg4Uhy+zwgpTR06HRJggrg+7m6K1gNF6EVDYEcGgYmMRmtQFE7S2lo4+zIlfxVd1OKQEQy2hX/eF
G4P4KAtlIgZ2xx9NDfIyx/w9Er1xZVex2lXgt2p6GUXjEzHi8cZ6x5acggu6Txwjkl93IJL5ptg3
LAJwjJ1YnRKWWkjJRFJeCvW1qoQP7DpGKGng7O72p4CGw0IkZNTqq5KYZLf8OFTDEm3g8/IeZrqc
PSad9DpJiP2jFRPKvPzfenb6l/lgbRXt5NEwocdHCKPWQak1XhWvEMNlyJiyW/F7NJTlcafqe5P3
fuS1Cnz8Wil9zcvkb1QqnC7fH8udYGK5fIdVEqieq2A6YYZsp9V1GOiETYP+nC7x6wlIHDbsFfl+
UPlxiV7I6qxZp0QVSo+aKUuC3eCoy/Sibn4+qD00991ZpRUpahIzGnG0woiQ3N9GYRGyMjhnZPzi
7Rw7ZUfZQtIFmV+foHcbIqbZzzPiRAeS2oZEI3CFhE/XVvPhd6DVwr1Hr+ITV/A+pN/0Ubuyizj/
VYBNJvyO6HIrwli0Z0Y66u/CleKlgPmtwplo1mO6l4UMfzEFiQxQPwCIklumP5DAdc2E3qRx0Jgj
GnNad/RBjTAVdS0HAsh5KQ2V6wCD87JD5nHvKuY72IaJs7EvyU7xdmVbM3gD7Sy0/wficu0KywpA
r60uD2siJMRQUwm2CNzL4GvRIV+xXv43T/xm+vYFiEllhMfOHpGdA5cC5+ztbfYXlPVJsZQ3ayt+
KhLYEbM8nuGYR+hx6zeeIZIKlRV1bjLD54Uk+R+Po9iTXrU/PEZTfGTBzkjSAwlCCGWA7wkIHIOs
++Ul30vJeL7E7o4Rlj0S1UQ7mkIKK5pV59hPUd1rXSutYyB0/2v2vYm9heJkWjS9vZR191VpXIVq
zwoOzG0O4LaE/RYROMKYe7k5FsTmEWySa0g/5cAWtRLnGTLBR1J0s+1MVMzH0aSuophciJfscU5i
AQ+Q0cNFKh1hwmG3qSgq84NpdQxsA51TXT9bxz4oACcvEGkPCyrFvxMaoTuPWapo7qZ02oNKDnj6
DkCkH7h0+ZIvwJkSmFaixAxySk1tzvm1lZx0UXJqtQCcaKkXVBkOh83fxxrUNBegxg3utkNXzA75
Qv4VMoTOq5YskbhQi6qkMbI2pxsDLFlxEIaVI+wtGDdVO2Ax3G6deW7yxzESUn4OSUVwj7n9HtSX
UTUDpZh+F7HbLkqWxCBGEBB6k+38GfgKIXfGfdUSocBMV5GB31Gwr4zMo13LLOnqKzR/1kBf+wJa
DeAnGa+a17Il4ZLSJz0KpkBJtpNhyxjUc99JvIDH66GDWVCfOn8wioudim9dtAugXargfZzBW+jb
xU2A9PqCu6aIVh6oe/JC9xopqsWj4xI+U6PjqaHMwFy3Iayglt3If4GcYBtvahwzUSyzON/w1g3v
iuvM7rjg4T98r0gJAPPv2hnfRqkA5ymv6nNeYij1rRWwUWMOk/kmPlYSrnFmi/9w0r2Nd03Th5Df
bE2nk76kX8UH91nhsPXq1v2kajFSLgOj+Y2KJqh/Sx1D4CvX0Ugv7fmKSt67VluTh7Z2sw5a31Lf
5CRiJOIIRNcG6f9LdDmN3Mx5NNA/zt+RROE8VmCZZLLRcVXtGYzVTUMhu5SGUMTTbQbJwwWk8Ev7
TLpKlPBIWzs7DHGtMMJeoL+ElWWLqRdCON4pnmfcVspZV0fiBtxdvmTV12e1NSJJvzv1SSgWce30
ZXW7pZayMwowatNbR0+VaFY/j/RUt0XlxiC9qYLRqo1VsHQziB2PaaRTybw7jQbjrosYTf39bhSW
V04CBGF0nHnzy0htra3olSo6IBLy6EayrwiJlZ9ikQRBGQoxh8S0hB5Zii4ImyHqCE95ii8gnzPn
5y+lU2jfsxDvOFXK2M6BCQ4SDBVllPFpZAHg46iKKJSVhixpIYN+Rduv+loB2augHtkgXYslA1eo
e1SqGFgamoebuUCybK1NmU/FocONO9GX3xB/CavWine0q0fcGP/IDSB5tyAsZTpm9F5JPOFny07g
Mt4nWA5xCBOkFrjiGUIyMUQLNDjVMu92mDomR7tUJa+rVLACJf2QOotqkkaoGDPN6JNtA7bC5FDu
VWeU0pEFIJsBvaje4puMOPz8ffEEPDiUUzPQRxfr+XpHQLl0U+seoA2MfEkbtclMVFWQGE4YzRGz
jWCC6Yu4gt8B8DT1v209vLtDJAA6cz1C/2MfRLpyFgbpJt31LAYXHyz93+T8HOasOPcOGmHu7K6N
14XsWCoxqWxpAxkLOoQo/QlVgxkAooet0yq3eOuECmzzP90hILG3BYrxFHoTNgfgxYDELx/1ch69
SOz5ngj3z9IaZiu7l6mRYiIRTrTiUK1azWKzd2teHC5oQ0ST+v2myqwrQtCjHb3Fe8IOpLqUZ9Fe
XFX4czHFkU1dBqSqZyii8OvKJ4iTZuPs8tbsT2RE35Hz/S6qTjgQGtlMXjxgk/356qFDQhfWO7Q8
G4h1WNzYQ21B3Ea0IdD1yPf9VUnzVGnanW90HO2pJKo4t2R1Y8HoC0lZmQdsVb+0mj6yYFaMq3Jy
giqKmSWz5F2Y0U+TSPzJTtsXaQfK6+iF3k6ivSO/50AvJ6GgMYBS6e64Rjs17J57eEhRxmlTjYTa
LZW3ZTCKC7oe/q2g2N6hClgqYJEwUJN+snGJzO2fzuVL9llJBnXYK5QQNWoAfl55lWioGB+uj/Wx
WGb/ykHexDeyfRp+7KpHkxBiPMdmTV2pfF+VkrbZNWbkPCxuaFp/FNmJ7VBvc6EdI4s5eIhVr/pC
RrJ0S2J8lMKJano0UUhge6pl/0cWhuZHBDbjAT6vw6rBhKc/IPUb5+FcUMM79Yn7Io08OzXyJ0Q0
mQq41h9njMuDC/Iiqdr+EJwiM8N09Mr5f1U03/zM8tQAwaE0OL5pV29yC8Mx+q0zEuoEWG7eVMKm
OBAJq1JqpkdS/9o6JvlI8RHhstHm5cDBu0QaOB4bQ73btGFP4t56PH7gQBCp6FMR0kfm86xc01sI
86kA4/WfNIbBsRBW2aPjzhVJeR96DrB6jsiMyd2U4OTPu+XBPksL6Axt8QMCiTgVUYoV0E1epshk
hVVoiNDXMuOOg2rjC+t5hw/oVsOVU6W4l1hagDWQP2tIamDyfIR7qPbI33fxh7bfqMpmEYKJHMM1
VkShAsYZ9hdfsGnNiLqS/fj8RGrDrpH/Cl2SF0MyJH7jXetB9yN0laCLVp0y629czMJCoKIzKppZ
has3y3AlkYmWyWrU83/mOYRNwVslPWG19a3Faw5VokaOFNy/OvQhjgWm4GdZzQSlyTsmUnFyY4ds
YXmMAT1Nn/BgA6O28eF8fNV9fbQi906GMo6z2uBuPYILXB9Rz5LAhGhePv1RsyWw8h9WpQgukcmX
pe5fCgGCeGS5CECtco72Ta5AKtEZalLFt36TDyVI9Z5q4pQAwymF1HiXUsBgwFBMderOThJYchs3
sgnXoxG1AOdVSP+1Ap9iATHgkWhQ6tllANbu/pnUU7Xo4E6FU4s54wTQ8lg6p8BO8TJVRBBX1zkc
1IUhsCZb1EiwUAweHyxjaq9Q95LOMKQwhQ3MqqVd4AHun5GrbfJ2skoaFeEtsFAwStZYa1+4mGTS
JhJuixXzNehVY3HhS+gL31LQs41hvMs0qVZ+QThkVxXZfqUuDztyLY6iq1Zgdx/279RBKfxfqJLk
KHRCul3FYWbsq6lfzNEcp74zCz9qo3qFIIKpKpi8AUQ3JCYSOpzZ2mzoMNrRHCx6crxYbx1mtPwJ
4GP7yfAg0YQHjTtpHm8sCPiXqFO1Wa+k7XPWLm431q3gtKjjArsc9dADJYU6MHBieyXKhJe4NWMS
oV2oaoDj9AQEVR1xtG1g3wA3HJqc4eWBIF+rYz93HTaQ/lSNOMUdYfizTOsnGA==
`protect end_protected
