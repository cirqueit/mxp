`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13920)
`protect data_block
SpwP8jaf1OcWJFtTaGLxccTSKMvc87pr666Zn+GXrmuvI8VMl0bIZO73lELNYcgibcWlbI6UhO8a
oQiXdW5jrffDJPCF4EcGC82cyPqYkLAUFvv9Qu4G4GuyjlMszN7Y97vKhKdSDJxmK05VApLcFFRp
FpRv5iOXieIDG0d+KpA6deGaGv8gxKnyI7qFV2t78gop8brYhGw7AfWXA6ociJsj/YuUB3BSOTpE
j2tA9panmvZkCBphRDE/IwKEf0YRQwAHkG4RY0R62o2nwm8SOyUETcZdNko7a88odLp7knWb8+GI
lne1AcQ5XmIM8WAxxDOhjm60gixEAAm0jY8ON7FbmcEJ4G/HW1ccAeUijP43ioYrMKIQ2qZ5cuXz
p1lJApIkOmDcl/G7XEWU7Ivp0ZAo9WWQ5KnOkFj/cqmoiQT1qsgjvZ0gJj1lSdt6hf/Tt/DeXnMQ
s7DUM/HJuS4v9RGvs4tHTpyLYXD5d6Gaq0DNWpZhRnsEq4aTxSIvKDmkYjOs1srmxIWnVojKxsR1
8dsUnieivPem/grCjpqxG6t/1i32gmOVVIZeSKmadDxxOB/xhqBxu1wQCmuGQhFyIsU9vPwg5YN4
BFYSNZveQFQZ+YNgtQHdDXRNOrwfgJFEzJn7iudBdaMAucX/Vw0CaEU6tW1u84ZJQANR6LZYWrld
AEpw4WUqtSUmh/PFa5Tv3e5jbldsMMhWujoGXb1VqpTwhrIba8+BtflKJf2N8+4JX/4SZ6LqkRCR
mlXidKbiKAG/C6Jrip0mVk4q1lmdfCt1qUb+ltaA7JXi65RI9m2tpiSbtUkX79b2RlEXQps68N0c
Z8eL+ph6rxsrIh+tYVhvo2VSQFz+Lc/ZwuwC5hoXYJZAfjl2GFTOy4FY7C8lBo3EmI8Vwy6T6wNi
0Dir0aug1WF41zjIGa+CaWTQQ/Lp4kFMk0jxspcgvGbzh8cwIYlrWkuYwiaXnDUluZcIgL3E3wJs
bF5V04liO3MZXTZOnuIrr3iLNBWX1jyZ3e96Hw01oYOzGNE/ZIO8Y1xZn/YQdWRBpHrA8GuAkavQ
57SGIAB5Dk0SDM12rw1F/1S70hP/KdKp8gSYht0PnRJ5h3C2yy59K9Q9kWC8iLPsAMGRamZK+Jwy
Cob6I35gHWVmdKGwVSZSPHGeDM2Un9NFaMivIXOyvk5dNIYmE9wP1N9Hx8sgilJ2A0GMsPLCUiRd
aDRcHo1G1qERJuEDNYyJJf/3c0fIDjp8EiE8IaORBkVlBpd10StR6KKDXpERiX5CCtBpIrYIcADd
lMICfGCxaPpQEsaICeGdsaw9zoNCPldXJI838VheOi62SaU+CkDiICAZ8/BZJvwLDOWzKEXj8qnV
iTqAh/dKV5UtJqutnrHMzo4/WmxYap6WKfGwpuQiJcTBw2aWweG6/lwjRTOBsa4EtGx++fGCg/Q2
aK9mKXrjW457F1ujG+tMXzm8uCxPeyvVBuwKZJh9z4HTdn3lfIo3EahNhJ9OdekB5QXHDzaXzsE4
mvspD+DfUmWjul/3BeIiR11TSmuFU3F5J5xjBhHV3Ag3qNOKbHriji0XenPNVa+t1/oLQOGUlJ78
mChaA6xSNrttXlCjZqs6Innl5EUW/S6Dc5/7PF3VAmo7AMbrNRVi8BCaDLaFjo9bPd09/pSPl0Fr
VLI4/40p04UL38inDZ0lPFCepL6Q7uPkPTpvRU+dgXlrMa7QiTjeax2EmMs0a7FK13PMCzXx6OTo
i8pMF1hXi7WwhTa2qoBMkQpFFe3ks7jje2IaRpMWQ6M85/XyGRl3fKwnhJrk4V5A+wC0UPBv0LWl
JKn4n9pBvMXxqefV259GLL+G3HcS7Ddw2YE5/2jTQK0hnHzCSvuhn0uzMIfHxnNuO1fP3xMrlhar
0mcFJyqcY4dyiRKtfs0jrxVN6GmBZyxMNu+Rry1RMvYdnASoV7qR6EYUAtB9yCX85Yr0BV4vsc8v
G/dbcjvtTMfp3ELXlst2fhlE7yNNFfUrV3uaGQrF0wzynK/0ja72L2zl3YMR8R9zktFkoVpsoh1B
/s7yGNzxKPSaos/NJCRBuDaY1jsTN4To2mmG2NbHcwtTr3NcY0G1pGC6u9yXCg1P081O/t9ks+Ap
a6Udy6WQk5rN2AeIscPOzbzq/SZxZ0o5HqdBMfAqg6Xyj04zz62Qu16sa5CmPIHCy7CooqgpKcgd
kpluSvmQuArqXf1ioqYmIQIPmnd6nDSGv1782n9KWG6F0xteL7qaasqhb+l0IhppLm6FUaNgOOTG
B+8coz6UklxXZKzO0Q0RGRjhN+I+6EKMN48KYepPT1iPaUFKvwQCFVsyyNhAp/e8rMGvz0e32E+C
Mlslqs8YVxIg7i89xl5YBXtapALYfOqGJOfQJWAvpp1wzA51myWOCjXEOcdW4A11aYTgueDm88m9
clWb0jQUOF9Sbgfw5xHi44NKjufoQ2kQaX/GxPaEVhVuzm4wVrTtqFHHENgvsAvwQYQwLppVplDp
uoRmYq9PjyVGjdGA83vJeaJMeXigVisieQdpW+Ac2hnX4OHoGjK5nXDE47Y5s5Cw8xHUu36814ps
sl3xsYeVQqk2evqTYkKBHG3+qkkHmPM70x9mIsyilEj4+o9615itJuaN8o6lijtmtBuMir8WpSii
+CgYc+NO7JLO15yvoOY81H416XD8xIE/G1caUrIZrCM9+gQSSUZH2e9XmiwFog+7Zg2bVrI/tn1q
GIo8UMeh2mUGZ5hqfH+msuwBwi2RKQph0B/7JBnBwq3LvjTzapDUZUQKf+y0YKyQBdXlPh2j3H4Z
mRT9Me2bc1eBWCgnz5MWwKE0dG8e8sunj0EQ9Xd4EC6jOk5roAIiw/0ZboZ1R2CuDM81Gb5bKWxO
O+ekrEVcuNBZPJGsdYFKbeXyPGlWUmF1BcpUYVTLn8lqPKr6VgsaKuWWHN1cOAjKd7snFflVSTUd
5urV05+qi33ZkfLNplRgZyPegCPyTWVuyC0QWgUgS/PbinzEnqrzPopj2sdprQ7SotId892ArKJ2
3Qk+uS8ROC1R52PObNamEOCK7VAsnSkis+vb+Xd1Bwq7DhvOGNdDbogQadgJYqB9rU/wsmKrCOnY
l5nr93sAKdAOrxJ/Fd1kvx6ks9Ms0OmpDon5fz12IDoQBjKusCEaw45s7xRp3jJ0gsUSADrbFXlK
rScVrRjvVZQCcjyDToHFfIS+DL547ZaVbfDk34iLPYoX0P0S/xDzeJZc3KQjNryYhK5HyMNVrA+i
tFhevnpGfYWOHs+DL1iGHJYsac6eJv8qRihp8L/K8HTKrDJTX+2WWyveHZGsn5tZmAzJKg7QMhFN
pmY5fv6ig1qtiYFK5P2nNy0BbbtaHDpiBAbBV/0LwsF18Yu/HFAitUQjoSh5/nvtQd1Ni2JENk4Z
oma88pHyQPo7KBEw/9f8fbPfoAhrq9eUUvUkMRt68JlWAS9h3lhneCfhu0E1a8Gd2YWkSAGK5Xbg
UzzWjitT117m5V+6F4DtIWNJr5dJBr8k1SciHYk35mGc6zYsPVXU2hX5MjFKlo4DKipTuCVlM6rz
HA4LQDpCBSWGsCkS2Azn33CoxWvzE33OmQk2d7Y1aL765GIrIz0rFjRtBWnXJ3yrOE+pviEKv2W0
4YbnvaGdfYnqfwOJpquYfnzMUGA2MlUnwQb0XRgLC3DDJ9SrgrBoQGW7FKnvbQ1skFnCKYDbQZm+
0zOvwOP8ImqKsUsTIT3/sm5Gl7PasNDtaGLBduCmrwJbrpKnL1AkCfCu4hfY/u4yyrYYpvUzwqPY
Vd98FeBFccNsXPPo0naABZNc5lecV3+OkdClnURdhSyFodnPpaXjB4T0He32Viu00RcvLf8dGtX2
uuclT8IoQxGNvTyReM6wmxS7A3q+Z4GmlwNeJoyJqJ+RgaQ3d4hMdFlx+q2CkPpR0Ar3sbb850b/
B5znW8kkf6oRl4L+OGpvP/kJCIVlI/DC1CpWrsCWbTdZk/d6B2Ru/zZd1tEWb2zVtxiyajs4AiYb
EHuuIKJS2O6WyHkhSc0PqF8zUm233JA58IjE3CWQVAmm9hPSCEcyFWqGRcEUCEu7dBLbO3h45/CL
2yIOCdtOlbu/LJBosogFQsISMjH7z0HpL+fEnjy7neTZYRHs7ggOTIQDV6sP/l3N84wm3logVt9F
hT31W2x1BeCaEpfw5UlA4UfX/FrMyzt2BP4lNVlTv8P15vtHsFYnvmeHqYme0R7sgDaiAWjcBcx1
/rWet6MAD7bL+AbjKr46v0H+pkEfcsOKrJ8uswFY5p57mIZgdXacstA8mB3fVGwB6CrfObgkACQj
+ozS369Hju42k79t/86f+FgPO/YtuAOVuzupEWKJMVgWdRiZqBXm3XCm0+UD56IZmSI8lszUln4O
UnTHEB5rGbeabMcnNWE7+mQGbLR+0PkboDrgrlIGZuLTQpfW7u8zsuHMtn16rUaMF7a8ENmZ2GoG
gaWx/vd0mALw3YdO3/XRBF/O6baH8Mf+OPKbEave3kzlOLIfspVcg1xmVa78rZHmroWEy06lsa7z
/EjO3lqLSzX73XCkk07swoTAqfSgyZtplj1LNYpl4H+TVWA4JmoNAJsGRDXTOL3BkZT4vV3n61u3
IsMlzZUTpudm2qI3sPO3ncxmznadmIcLMskJSMQvo1fBr9N9UxYUexL4mRTDmkqNh5oeFqrjuXbW
msKo4IzdHH/ev1hY80E1xR/BuKbWvDquoZYSDL5mGO2i0UTmVGZNxmxlEi09LMc2bFtCmSIax/ZI
Xx784sN6bUOE1E5eCQvNBEE0l7NLiszKf2d8ojgJi0WTvZxt/Ucuk3cZrb1+GAhePqFbr5v157SM
tUDrRPCXQY5zs3U3KUER3LzlA2QEyFVaRi9T/eZ5P/rOAWRatrWVQiSq+BBWBkeDEOettKIYMuxV
PaFJ41g9v+nFl4IxQvdmfeU8SUKNnxwlcLK+phIQsVEoXwyME3Wu6U6x1lFm+aFuP5Q/cWTiNMaC
yNvnJV3WoEd8FXX292iISZu6nubEHDEy15v1Xp01x3n/NP+uzvpYvXzlhgIO9Nvzw24Wi4Ur/Rv9
vmAF02n5Cl/uDJ/0Rty4hScduu4c/SxC06cmLzX28gR9X3niFVeT8OtWLh2WBGqTqZcucYqWUmU9
OW/PjbL7YsjeEkD8bLd6oBQwvFBjSm4BZZEJCTbha6isFjB/hHKBm+K2yHuzfqc0nMb71Q+WtgTx
/8YCBj0qDrGh4Ssi+CE+XRJjDxkHT+apB5VPnIfc9KCBe4dPjn0BRJS46i5EO7+7Odl3GNktGkXS
MD4Df9OxZeKFQ1AiXSjvcRPUvRz3/BjuYaAKBVK5nIDwIyTMjXOXce1RQCgy7GVR1X0ZL23bLJtB
h5h/bHn1eMJ/fcyTTNOQmN+U4cmXtC4wgnhG0WEkYziO7HkN0gRcMzWQlIHh8JnBITJn8xmTewa0
iuWvXASOf1McJM6pzCtgINmPnjb0FinMCR7tDswOrleFMdrg51nWShCqXOTF2HOa78imvoyGPnWs
7vKCRUoKfBlYzlzLeXvgI08X0K0yZmxYrCNkNa75FrhLTQNGbMz0fLy3EWAKbBftxw/M1nFh+La5
8z7CW/k6NqUFw8vUAnGMIG4/yewK5K0nhksjolZfv2HhVTMPYhBqC2RfZtuOeiXY+ElFJ2b89HmO
qfEIf7ClF1TsCclJAoVXadD7AwaGrX5B7yQ7RtujunyxxoNbPsNZacJmUJN+YxnOO8gX7WH7bFGB
J11UmmZgclHMh7K5xM2gxc9b0fa248xpJ+gaLDHhlJmNTwdK07KTsHlxQkLR+ugPU0ypJK1qf5Wl
pRNCdaUyED8Z3DCUpP8z/MOh/0P1EW/1TzLYQZ6ErvlPmbTA0taYoDNV5fC69XJlghgBnmTustrm
x5tNDzxyR9IRcJwID1ON6xkj0Y875lQCIm0MoJ+WUiaSIenh51Jz7aYlbd+FR1vijGo08waTdEtN
1t0Gz6N3/ZfJ4nvhHlf8YmQOD8JiWFSTqDQtJ0bNhz692O2evAUvqJtbdu+FTcD8xFllDNGzvF03
bvWtqbAS5uvCX7/ixBVuSqCipdPLC59DCiHIEghVEc/g3jdpWoJ1QKMMHD5wOf30veIv7zdu44nX
86nb3KXnpW8/fc6ddJICVlbTC1FX/4/WRqbAcVItpMAgPbMbJO1CsptqYw1QDxrxuNNW6cDYNlNs
SJ0L96fe9oXteHQDQStQB2F9M2XaRrPJnJ5aAp0S0IvahLTdLKlDgi8huddRTowWNLUciMsqMCYk
gbg7Hcef3amEtKMftcTLcvTaQua1zoMUSFAxF/7Jg22rQfgtm1X1JzAeLoKeNYPKhCNSkQgYDVgJ
8qfqssLefLeDHjshLoH61BKbqbPzmusdZ2PW9oLaR08ggsoUx0Rxn6ZxeHqMAYsHsKMw4z22xp/b
/dR6XTCMb8CjXiij0G4GBg3vPfluXoKS2e17hRvNwAuzKwtUv7ULoUslsU6R5XnWi4vUWwVfTME8
0sCkeX+/QfC916EQvAaLrIBH1M99la9IRroG3ro5OO8zYV6gDpRGP68JKI/zCxlnn9pPDsLXJiso
dFKWQJyhI1aOole1JtrDnnayFK/t4ZWwYo0lFMAqGLM8NdA9iiBXZ39WontN7j5gY+je3LL+hfsl
DkaJKXOf4ZZpAJwiaruH7VBfPcLTKUUDKF7sOxhaCnjn6rjejCrVugOZotUE5rALy3/o1sSRW4KY
emPEAmM25iwDgKbVO2vevoKcyf7RbYqo07Ee8G1GCL1iBjJHg2j9EE92jKJH5bFY4ZSPiIMrjjXh
Dwfc8UUgidL9PvFe8QzVPW1q1o9tKCtZX02VVW+abUUkx0UswHJh+BR/89RKuOMzxVUYkuj9F4PN
LT1zOtRUYI+oCK6Ed8yoCfB6dB1eSfplqIpJnS82fceUCY+0d5e+N3JgFfBNv7bXwW43VHNdE/6D
O6BhATFGeKWRMCF7vOQGnwyL9Wzl1kILa4SMSh7Jdqr6WdXVnDWlVA9UCtwPLQ0myDp+x1ub/Feq
1ZbKzaMvbRaUitvBsG0afyRASFroEgWXeguM6Kjgl9VLj9Wz4ufu+Odwz5j2+7FNGJjY3718dVSo
rYSgY7gfyiCHL/Nn8SPA0CWIahdVbVffu0UwP+ptddKmkSwY5QMxg0RW0+XGSl1k/Cj16cudD7o/
DMWg3GxV7iBEv4PtmQcF8SLA2k0V/y5XQvov4R44DsgMZsnir6SYPcw4DiiK72LANvO+XxGkBT4M
O9Z/AmnN3mlxYdDrwB65SId7vPBMTHg8zHPNaa99nYA5K2//ZPL/WawEL2fVoyXojuMmeTk0W+Qd
DKjujiotuVnP/a9qHWcy8nND0Ibbx46nI590Tdo1Vd0KAJSZNlHj00MqVHFsdl6EIVf1aEHFacHx
/YOqZ2saJ5mEIerTMpcxxtnSt7gUQDjYlNzWzyUzlJ2tgfeZCXJjN4lmRIRSJfbNVHiLy5HO2iJD
+ywEBXEFdjzFLktIvKsx96PLy89Gl/Son912Hii/G/12aBYZN9JmiUH4OGg1sPVQqUPE7CGo+E5k
6Mnw0zawCy0PkiBzq/EI7ySlzq8SvX5bb9otil04WuwbJnOEJbfu5R78u+WJj3yZqey0ypjTvDP6
Mb9Smz4ZL030RprWcpixG15SvJUxhkvGJ4D7nXUffdVpAqRwSq0qv2jKWyjmy/0xwQeWDynKNKA+
nibZO2kMPfuhtMWtI+s6GAM8CsPbNdafr8Z1mz17Ax72M+XdkyUEF+4W32VD/bfKS6qmhX5s26ca
mZNgvlsAA6eaLTBchzb378DPAHYxdQNBMKT+Zt0iP1GUGuqP5anNCyaWG0zFalmR1yY+GzC8Kq22
OyqSNbSXlC4vY0AYmoYCqCdzKWt5y+E+ynpbYB3Dx46PFJMYTZvhUgfabu+59R6jRVSCuqr6QlVQ
tZs2w4gK6zxqmoFMHeCiuTmKWqTMGyOqVE7uiwZBPnQuOVL3dc+9x7WcK5qX49vB6+sHPEcTy/fl
uw34BvuW7gK4VMQm65BWkSNhCbOWe6KHSFQGd79QJQYxBr70XbiKV+mcm622qnHa46S3LHdf3xqv
gufyTW1F0OWCrBk6gUYS0EAliwth5vMQmtuAWL1njbZPekM6fuHegsQ0G/sCNdJz0qySTGnmQMjW
57Qcn78xaEa4G+pfTcQYy9Z3ZPSSEGu4hGhixgYXcOsrNriKHY5GIiA8QbqIIc+NXeGxCecFbSAD
6lz5sceogKPX0acFB2LuxDU+5j1d+qU3FdQ3AAcfFvcIJ1xmrcFZJD5s1EIFoOkcItV6eXzD5iQg
qgN6yH6SXYlIzch9a+Sdlp9MKnRA+8elJx7/YOCRrHbZAp/Cu0IzN4UN19RPRdsZkcef2WzRlh8Y
uD4aE/6u1dfOWN3lv+XDgr/PPT00qqPCWcwhJXTXNAVKjqa4A7HXChJ9UCefZSYQ5LrEc8DHQ5xA
xKvzB91A9h67V2Nn6djX6u0HRPr/ggETBGhzNuTU79TRLg9uhymFQJzS4nu22u2wKyLZvHL56S+y
cB4IlKID7r92STq7UM5BBYfaIbO0DAuDIgBylZl9uxItt0jgKNxb7B7/zbSSlyxMknI54PBujKse
N8Xc/MvuUDKAbwx8J7Q0btgXKn8OhXuDlC+8tXRAn4XDtBoBCLUp9fpSYvnWijo7A4r3fFNDKHaP
wDswqDFCTxRu4nDr4zBEz98J4pSZAG1gRxrusgDiA6s7Gj6b0LLzUN9wlMY3JtK9LPDFfbwAKybO
Yc6R8gV1wbT6PiU0FVGlH2NVvWDN9+QQj672LQju0kXhfBjZ5fL8PeaLZl19K5+SaFUbm6UdyrO+
UotOOMedQZZU8PUiuMV6YerMRg4L0YGcVZcXTAQOfziTOgEouDr+u80XbiSZ0DBC6KjOR7br/D9S
GNkjLc1JVgaENsx4QIh0ufdxtnJNmBtlv3fjHuh9Bc6QTalIAHoCQ/rPIasj28oXbqHJgEdiZ7p3
IZUv0pl3DK75j95/5XNzFAdgwgRj3ZKu2Up2qqJPUR3mXBYifbWwaXVekiw54ephs+SJC+cnHCBD
/IMD+0DZIf8VFlLSzSDYtleSMvOXNHC1gcwh8bf+EyI9AYMLvJoeCBKsQzKyQnv4r6BaXzeMS1Em
Yv157YCuGO9DCq69kxKYPZc7um4WV6aU1l0r41JMFWC4cemEvD/onTOt8ezNyqLzytXGGXGRZxz+
kf8Ag8CkAKNGHTo1pbN92Xp1IAhhqmOVLatGxoXhlYgPQn8Q2hv2DyRQxo5UV4hVsKHOO0fy8rDq
qzhRaVaIVh/gQBncmBz48bZKfGpYcg1keINgcK33/4CZ44G/f8PtCW79oFdhoTPRWUYzwmzEBc0o
5lb+mzxB28i6OTZ3JTN5InLQm69pYB3ggDg7OZX44GodpXc6xiyVroRUKlyAJg4wZSFnfp8OEeTP
t1wQnzNd7XDShNsnWI/LBITfuhmCWtbDJyHrmMoc3ivtpCAJ2ybvmyDqbXzLGGoUioQ1FlmkpJKR
Fkrxl5sriFJaSZpfMkTCiUTz+E4I4WzpQQzNt2bsZdKGZ0mCLG3ft4HWyZt+EcjPp+53l9ajk7Im
BXIfaNCiVFGjTNfw1MEDnuXfEZLZ/3pabrhImaXec4o5MwHMoRtJBkmYj2wFrUR8P0d9GjCcrx+J
AaIPBtAPkKqMnm4ca/QtCXG/+kUVmyTRz3qRfKeIB+L3zyf9/TRGBu+/sPq19QnbVx2HXm8+QYfE
/UJFKQ27azetXAas/Z1rrr9DDKaiRvvWc9VXumoK7UX3vGc4qEZr3AaJUlqHUPibmBsX9KxPwcO7
fIHgZ+Xw5fmaqe8oXhv1LfOKmaG2nLBplp0qk05xNJnDXd/Tw/j9A2HmZ2vw1YkubhDwihj3rNbF
zEXy8L32YcX9HV1HLHC60BDtnayN2MxKlQrdMTrS1FdZ3z3rk7P1DHyedyLN0Wg4vk5ZmX5zpNAS
ZJr0jQXcz6MPDcuEuZKUYlil8epUgTBTtfqNK1XKzIxfnKWJNlQ3Kkq+l/NiapgAUxrV5peiQGnl
0ZsrB3p3lJMQHCmcjn9YADzAhO9Vopg0/hLJMTHQtvj6E5wVhhBPkgvAazBNXqa53sDykAL2Q0Uk
FaW239V1w9FXIT+zBK2izw9O9KL/k9ZUKOXnfO0F5b6IE6wmX2NAUL7tQNJS45EXSjJ0Sq1Ct6qM
89bQfiMv5125/AjpveSB4CtZ5CnBnviykBv9zPL68ZB1Dw56Zy2i+tcta0/fulR/v9TO9ZMqKJdL
pcb+S7wfmNUnb4jVmyz2a9XdBdy8PO8SiUBrciXzuUJm4zc6S6HNXz5wkaAgQ/LWLNbobfM0zMZB
l4uOW8qkOh0L2eveYPgNHjzveZSgZSRk/w+EKMEXegBEZo0CqmKbRS9KDTO91metPnatUsx9Ntpm
i6tbdZbF+gd3ywHgdRf+LZtzdrILJB36AreLPj/y4wX9FW5i00n9s+kEgXwtGxmsPTJqkpw3MNu2
AOA/WeHVsQhDs1sxkEU0rqKFpRdZY4P6cjtLBITNDMFl3HWUOUSgl2Ijz7cbKTGI9PxEMh5zbG5C
g215L792Sd6pAur8NjQ1qJuqcXvMDbzrwH83tUSgPDAS/CCsyBR3ytJ4Qb9WVnSq30DJODQO5HpN
oWWdwIeREikdtEVIu8iwv9raPhoTlRkHOeFKLeT8qxvApoDw4PmpcBu68J7/IbdlEfaV+XVJyQ3E
ob4WVLgr17ODpGHGXBYSm7e/SW3cUx+BzvrFE9ZBd3Y6kwr4GckixuhhAF7kmoC9ileAAg7gKHVO
ks43W2V9JxPBQAi6b76Q9AS3ewmoIFxbTTANmlGD+IDafnNtJmTATN4Xkl1s2EccF0WPb4fBYCiM
6MJi6wzcoIaNcZ7a5NV1dUnzaLkagbsVkE23xxr2EnmKYO3w02Ksuu2/7vWMcMmN3WuC6s3rB/PK
hOrsX2618+X0NVkml11gT9F5/mipsBzFbsGjgJcWy+gmXrGMEfprmgvlTq/ulunF0RG898PS5OL2
t4p+F51ZgluI8i/jaQX42ghHRN3XzlPiXyUVUod2aBY8oF07Wwi+nUjaLlGuP4/tlAaxg4mADe57
ZStUoKfpxVYZ0MKiMNQHE0zoY/zK8vdH7A7LAqcyLXcZ062O+pM7i8g8VHlF3xldfO//MaNHWxRV
yBURnEjE7S/rGxrxIIiHBlm3zcTH7zV9mp+IGWFH/UKIIlvcWO4T25pAyQcx/1D44zceK1tAbOdb
Jn4q86UtdACyh5ohQb8L++rU7ebc5pHMnArtb0sGzEQIcaEATN4Qz6Stcv/+6KnTbksrqaZT9gGR
8y+6Jf5Wz8UA7H3MBuMl3eZ34vyr7QabZEMJGIEO9h2PuFfBPXRCA+s5pVR/lZQDuxFiZNeDVSY+
+m1v8Jmywim0RWiQFhTkf8P0BHnJ76hRA4cnGBNYjOXr2DrmMfd8hCq2ZCIOpRiAAwjgtV7zECgH
8eFm4tNWIAHaH9dRlNsaMRw8y3ZFTjTFVmrUAo+AgSa+aIn6L4JEgAcyyW9cK0PjdSCa/E537o1T
W3IZ+lkJle9c7MkDnO1bFz76x1+VO21deLCLy9CA2iF850orVVt2YgCSknw+YsxHtClVqv1rPj0f
omOdi+bROwLUcvIXjxI7Ig2UFFOcntv61A1IsCv3FPu3405jkDBDlRHkw+3FKfdjnkPUmUPUQ9MZ
OXsEV598OkGxVyGWKOWIkOWA1idU3b/WcWlV1XKAftFFjpGuD/KpHrFjg3FA+RPedWysHn8HqC1E
AwiQJ6qcT91hgIYzUK4i4FmWQoEW2tJjgtLWc9m12rHgS9wZ2jjHlR6miZG8M+cAhWj4CThPu1WA
VkL7Ls5XM46w6CZNNzfECLwgCfCBNku8xzr8zRsshSKOhZnbEwQD/IoUG6/Dnl3C5AMR+1qrdMgF
MydTsMEItuJwNs8vdTkFBaOjK64deJT7cgW46ohnXsutJ83cFWrHbKLYU+4fGUFtbDbqSTcc16B6
PwmMkEM49j/juuP4lF95OR09ozn15fEM0CJPXdaI+goK3Py4BfslAgzxMBe6WXQtVestD/t9X8eQ
5P++Ww+cglFDNjnB84DjMyok9hkTs74RX9Ef6yTGclsNWIGibA03TBz39inf9b1mfBCKdFpT6LhZ
5vYn7l2wIxifyewkY37ghGjLbgsN1f29i3DGqjPtpxDC2PnhPtVoTD2953mVknrg+4qq9cXUniN0
zOHUEdoNWsUmL6Y91l6vFlxKuJ62uocfsxE+Tzp+DBl2VIma1sdUpuKmm2TVQ2shLpW6IZHd9B8I
LnhkCoSbgO2TSAOSi7l5ZgPMzm+WXWp3Km+erAEAGYy8ZVq0+EjBunoNFFafTky3jTUYFBMiDI0y
PbhlUYhabcEUsLVZN+kzpey/cnjTX8veR2FYSgbJ2KhcFMEOLw3dyMpxIgodi8B8V49H4BFsOGAR
55CrelTPAULvpJzjOOj5duWsgyzwHjo2nubcbz+u71Dm+0ouYBu//5J0ttkOau/kZDLhW8EfvfHQ
okmrk3ocRtfeRs3S/faSFufR5Nf1reKvD9LmTQixTn+nnndKAPRBlXP1kic+P6T0xmY9lywKmRIk
ReuuSNnI+AR6BJ3T2z/VX/ziwuFcpn8/TE0whiW7OGX9IJ+p6kLBbSdWnK6YnaDxaFg7HxTWK664
R0E8U+ONUE7aGTbUQNAGFrAu5AptvyCDEH5J7/STF9xpQhYTOd77wXdQxcNi6PQmnFgwF1GZ14Bd
0h7pwbwo+cLBhRoCpWFs3V1NyhAOLEkHdOLtk/5fnND8XncWCOKeO6khw5B72I/W70FuwzUMaF5b
STn5Tx2ryfCOaBVESsoB0lXzqt9f0cU+U3rUpLadgUN1ngVnYIJVu+nqw3raJA46O9kAd6dbVff6
6LFGQ+9VsNnmkF+7CgOnVWCsR1CEchCkvJEsbRHygufGMsYNQ4IdQX6QqSHic+8ekdcmXuRx2Mlw
d/B5Rpt9m3UOyKuARsnBlvWESqtnozK+bDOv05eFyVFZOqJt5w3an034QAy+v+UjrpAPsBE/u3Fy
2pJAkB2qg30033uKvsRo6T9Yaeym6rGGXrTFSF6W/oXrpb8W1aqI3J39joSYFGhAloP3m0obkq9y
mLk4STLmIZv5qSWz2QACigHo/vXllmSkGPH1/kDzhyYq9RQ17GzxYJewpic73yGSwU4h/NLXvxUJ
CCYd3uX4RdASMmv1j2MJma3PdOlbTfnh2E9GMkcRSsc8ehTxLx6uITJDDyD/NQfylaqmsMNMw9CT
lcEvO4l2mHnWRaApASXP8Dybs6/oOEXfuTP1CEWB60lxY/ng0ky9ArAWlRmJvdtst8LA7lQkHEhA
WqO0fszf49ri2zLmUati5pB3GDxFhQFWPdWe+iaCyQj2lVVWhss5XXLJgzO/ZkW+5LYYtkdrQ0dj
j8NmgQ3WGi2CRhZb5CDVqpMiOUbbO+XSZDPjFyegVMDRnxg0hseRTQhEIu5R4R27mCSVjJHMWByx
xJYwzw1ed9H8UHsDfc3YioZ/8xu9+KIn3YCL62/QGVF72sfO9Kju62WDUwkZFPJbwC9WzC0BhSC8
N9iuh6/Cc5I2skGPRe+zO6JiCZ6YqWH3j/tMIN4zSZtIod9XqkabHN6QY8rQt6V1rIVdyoRpQ0Bf
mFO2dQQJTCvwaZ9s6E3sknMPmV+cFofxGt9LIygPIVSMoXm0GVKGBkrXzaC12xt/rsDiLFi+9j/u
17SuvD1MF801wWySv9MnCLsyb57CTfDPkRdrtKCdyNtykVX+Y9jnf5JaH2vR8nEWLqck2Hz9k4Dd
AKRXCSnmiNSOmC6TbtwW20iYrg5qxK/mcKkMNzR33csq4TBpeUobiBF0wpNWtxwYVNtWWgrBckHu
EJxk3Z3qYQ1ggkc5fvw4ihVIWnj2j26PYilxL5BG30rAzE6xCdMPupIi9Fb7y0WUNcPf6vKLlqSg
0pxhIQHP1zHJpYMnfh03tAvRTNGSeobIP44XtducYXRdGASf47M3jXM4chfUxa535j3DYAHekT/u
7BgI/9LdDACm3BiBWHa64cmYbbwYfNkAMJwb0vb5wB9z0sgrefy52gwOUBkgcHVxuHujaOdN6gSR
qRTEkO2nMO2pfNWE7i4bvceIH5V6n4TT25/HxNNlhNLfU7DYmNezS21oPtw0fQLFFylQmEXm1B/O
nxK6dt4QDIcJv1UcXcFNT5nK6B2jZVQ6fQ6tkAA/wPvM6aQQVvkLxxmdiGNF8NqvOtPvtOcjRcJE
zmR+CwkLPLGhX062IYoCD/+L/vVilDXG/816b5lKYYwmxtHCfvSaoMQKoAeBf5G7/QX18APDjO2/
yFPnF/89v81kBzw0bSZJTwBrJENpo4Ql8wvKpCr7Cjuz5gHF/ud0mSM4w7UhhO9kprbO4nRsasTn
Y148CVgQ3RwBcEJye4F7ONp2m0ogLXdg5XRIEglr2/f6mPM/Vj6wM9Dwa9ZcLznsmdnIooqA+2+d
rTFeL4n2LTu2Yey7aY9UcwVNNPyVw4gRqHdJF4BB9QVYbGrp9GqEl/z7tOygaEMsDovC9jzfEZCY
CohoJCLifDM+Ps5TUGYV6x5GgfBkgtnrGNqU5bR8+H3z1o30FsoBxNJKnSv533aW+MlBv+ywAKAE
BIU/fxCw6bgP8ukfFcW4ccS2RZSl99jS+9CS74O+Ig6fwHbs34Lxy/RWEBhxGDeSL8vEHjpEAn/X
EjdhRmBiSuqJkarpvxhS7tG3zEYm81j62xzucQ2jzvcadyakH19/+mxljOBoB1IRhbtPzbLMs5O5
YYaIgXRblpc/xIvKjOQ70fzPtXmjkJvFaJCrMpmGDk8/sXW0uP0d7ijhwrdolvjrOzFOihshW7ry
ChxeL08nbkkKCy4tVQGZnJrveLI+asi9OU/HsgLBwlWi2wTBkLDulPIwT+j4zRkf2ou6S0QGGdMP
1B+p6waGQj4J7S5x0e6bVfo1mqFYHhm42OhG3IEEodRCGIH7ajsD7NOJDKinfTkH+PUKlX86a8JL
wWuyeXqYsNgV8SAlRRY+U2cq0YnKwHWfJk96ky3LhGEtMznVDFNFtaKr9C3M3MAjjZcCPOBGSCmE
4xt1j7XnLqD/mMppbuOiPFaEE797Wfm2DAc/tq8mPZaUGoVumWngWpMUZHH+si4pv7j1I+O9DGi4
/nYSZwIqwtJ6MuKVIt47ze7eCmourCNzMKtz/Q3K5pPG1PhhEwNlyxjQz/rIWOl+/njr3AjLN32e
hlaAthScElkDjub5ZvHtMQjjdqDZQ6wL59sESRo9q0p2++TifsLjEJMnBxcVg/PK4avPNWk+Axbn
cbxcJ5S/8D+rbD0jTdPeKurx1FRNVnteMRxzdSeieMkSHFvzgUw+JezeV+aMzDRTV8RFzrG8tP3g
Id4a6nGqu7mxbpWhC2kbpJh8YKeFadVNra33bZ7HbdbEGnQhrhA37GahzRBBYcX1MEuXw9QwlutW
p7t1wRFwQvYVmYr4Iqh07tVWlqtJRlkyghW530ykxbtp7wZcXpld+/WiZ+H4c906YaxQ8clkVNar
KdyWNE5OAjHcHdb0yKjsQHxupEhjW+/rrjZoltUpgx0sdJgd9vD5cmLBKL/mynFjbb0oT0TTWyKn
Z8L8Hy6O9+jroHInzXlcJIU3NDbO5wtI3JI8REqofTquqn06epUPGYT6a+S5gQHKPAVVIyjpT8BR
Pz/GOUNqCm4+JxHQ3HbRkC1GaLSppW0sn5O4qxDkfc3kyBySk8TW/6Qo6TIkogcChEDVrKsaw1VA
4Wow6Bt2BbS5LahT/K8Z9vgFovuzsa8jDdT8Qfb+nvLzf96Cguusi0RV05b1xOhdUZpVWxR/VxV8
eAEWAXrktBWMmk/+zL2ldDyU3elDQ5P8O7anYz+/k0q26Lreja30L2AAefFlLXVo7c15ZZhC+xwE
ZvRPMkPVClxtCweJ7pRswbPq7OQJv93f0gVRIvkNcw9aPoUNd3+UjvSjPJ0SqMEwoFfYsuZBz3Dx
D40GdnbKH/x5c8GtypAhJGyYzT3I6HLrMTd7w/OJVnIYdYxcfPpSVP4DeB9CmrLcdVl+e+U4yLiy
fQVQCYlYUM2IyyK6nEMyjTnQ9Qz3ajRPDjF2farT3LJUxzI9hMJcub1y9TblZDedxEGZCLbSVpHT
D20eY49KZFs0Ni7vBEeWWUFdWnJFBC2K0vJbLTvqzPk5hxNP+dVNG3UzpJV+fVkdwM7MBHIqnd31
jQ2eAkeOh5S0NC7N8K9KttTnFTNzedLxl+2wzpYg2AX5Whfr/jfySVUSxuwR8qCorKak2KarCpxS
py+s0KwG2wWGa/JUUzRJjH8XkFZKH4MfvzjEXsn2LA1XqoviYtttqVzxXqZssd/OiJR45plCZ59t
mrFpg19AEXXJGLf4u9q79Zt+u7WV+4J4yGqHQPyF2V14u0QILcmnwxddodsQfoRcL41niXV1QuKL
1AB8cikqYiWo73c6rY7Woj6XMJd4VrWFGy/Q8OQqnOwbYzExH1frSeJnHotsvvQtLJ6t7D8AneGl
GbsdMC79G7Yj3fR3RgDX6rJAygMXQfPgLXIKmSweD6cNoQ7yjxJAI0IjxwdBQ7frsacc6BdqjWJ/
qwzU6HJtr419XbST170iRBghMJeE0YsHv2NrmBYekupFl07/7g43+z33yLfyXcsspG5e0j8CWP57
i/lj+QOOca96Yy8UOllgXK8RLZVc25trCrd9la1qdWzKoyJ5zeszCmOC3M2skTz7n+DzETxssLZA
ox5sj6wqIzHcju5frqAEqg6zXy6dov7M6/U5McvHiR9HGX6oBJ18YJ30tLGAymis2KTx/Ml0/HT4
dOXTyx0oP9aD2b5vU9nawuAt59DJL+11uA+iqWyz8qvtXss6gn/AuATTkVxfIFp6I5bIB395OipU
L7V5aHoBO3aQ5VhHW1xBiv1XU0vmyGWOh9zmyMYdJK0q3RUrVvZ1TAV/IeGrHf0TGaxAok5eqo0J
9Bd2uhS6JIYOCpEYWxNc5Y5dZq//VtWv+xGAJux8UcwYj8StfaXUVCs9C5ULz2igLOS6NpArUcjL
LTR0beAXBXzlcwL4r8oLfTK13D90KJxRqJfRKrAHlWsoQsk6946CdvuqFV6o9qoncQWLo23sbrIA
xhM6HpmvznEZkFbvC99uHfZt4kdRMqXVpscY9BOVcWaMCUPVouQNd/aVllIu18LT9sFutPU7ZtKn
Y31hvKZsHzYq9GaJRJLWWoHcoUJmnsQJSZK3nAt0LQrz1XWldFFP7M2mJgzcDZpA1VbaETuq/dws
alAUfNLrPezzONmRQuO/peb1liNSUsQs3w254/cE8xh8Qqp5V8C9t8WdjGHwUMLONiBStgUF4rx0
XnQ/0txNBkyjJD6/HtjcRljshva4N4sXH4xP27gwRtzwhhYs4gRxAEZ2D5F5cf2Q5dvDlqvbKgCQ
/QT3j20XQoT6lpnV+cgI/6KDxMeOn6ESnhIOn8KRiQodfUj7lvuqeGqSvuxUWuS5vq5992wRSXZ2
IeDXRREk3C7CblKXCFJ593wcaGjsvvFSVybQ/JT8/p8TjNcPQT6+UtXpuWeL6xIWaHWz6cSo0kQP
3ZdGNBoVnl0iCDZGn7VDkCh8KrVeDhguzstpzfW6/ml42+Ds1ETUgfYwaWnTm+45GUse7h5y0bH8
1fMJ7yfP1t+cRC0l9qxBelwCJQWz92EfxYBauSg8SwTisVeZrT/UbZGEW4cT8TSBuusXop9qJwLK
+ncIBWE2XBMIEdxNpFXqxPlZQdhMgfz5EoskbozW9xKsv1Q4aJG9smd5yX5yI+EL2gIjsPZcykgs
0JPqOoDrzWgY7LakLk2nwR9/HDGuys7w7+KBpdODwPrSYta5pSr5fHzv5iuOxA32kgQlWPCGQS52
Zm4srYSCuMj6A6y2vAhlSWhU+u/Y1xnou5szgHvXRJDesBX44yuwbj9GoXWnx2VfUyLwIRbBICoT
SU9qPgalNijZopV3knNgq0lZZ6bc4QqsZgvHhZGdz9sLe1CghLrPx7dhCThBOsJ5Cz00FuISjRcy
HEO+03pBzuSdO3yRavGDdTwDQqidRl2MFulxHSutFD7EfHU5FbC8bm/C1UmeTbZHzek9zefsucce
h9lwTYQKyoXUU/2ceMXgMYdrgTXiNvl9AZcATb4pTanx8VEKQsutnwHnNpUofskwaK447uHPr2DC
uyqZtxBJdBixJFAHzjQH2UrsHrIQCKunikqnzTSNH00Iop2J7ufFb9RR5GVM4BZnu+dOn0pb57x8
Snni0FzLQJDGcQbO8vy7INHmEc0RBWPRbFcHho6yq3oAnppscEwYU6NLSDdLjWqzCM6v1L/csPE/
mKHFjp2+Vazq+0z/fSdZcDs8v9MTLNbjK6SwlK2mRSbquwLuAInZLH+iPCmW2fTSH+yHlWisPQzi
Ap5ec7UgzdwuVsVr
`protect end_protected
