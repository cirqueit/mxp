XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"a�_��_�/G�b��!���)����c97mݤ.��nL��:TGzBo�q��-E�D
�R����C��S�����ELr�ٛ�B�z�D�w�G� �/��̃��ʢ����7�T��#E�0ٿf��
�!�k�k�y�ZiNC{����M��(�X�L�M�S�SoE/"���F�6��=���q]�k`.�b�f=�E��Éte���Q����mZ�2mg��r���#wŝ�>�ì�b㽗����	����\{���y��89�Y��n�?N.ԭ޺�`j-(q��ȿjm�b�YT��K�@���Y�I�W"3�#Z���Ɖ���а��`�0�%��hоn�p�@<�%<� ���l����ш�����L��KH:�U��'����hf��躇F�T@v�!����|S5$A��[N��;RD!>O���-�o��x��<��8U9z�mJ�?���C,��ʼ}�%�y�Q��>���"a�҈ @��w�̬�;�。������ݣ]]����q6u��3@A��/ph�_��^^�Q��|u�.��D�.Uέ�*?��/ᗞ��{�ƮP[�ĵ.^$V̧O�Љ/T�i��8}/N5�O��6&T|T�^J�	���N�N�]�:	Jn �"�B��%�+�)M��W{�����d}o2>,p�����Fř�ޤY�B\M��߆�ꏙ�1s{�B�u����59z{I ɮkm�}%�2>U����v�b~J�$��تR�XlxVHYEB     400     1a0*��:�(�;���^�uFߘ��A1)��)x�ѷ��Rv����e�@)�50��Eq���zr�V��$+V��^4� �#|�&��"���C#�v�Xr�SP���-����!'�[�(p�j*���n����~���tfm�D�qؘ��\(+���L�@�  Lx�tɬԊ�Et�(��TT��k3���;RJ.����!��,�ϑ�2��X"�Z�lp���{�H˚nO��{��*q�2���-�W���"���A��6æ��x4�`��8ؾq;�j4��*_�� ��+�)F�L?����&W���^��_5��b�`��x�k�p*NgC�����N�+"��}N>M[NJ/]��+�_���9�e��.�I��Eƹ�C59j�$��N�٣HCaHም�SXlxVHYEB     400     1b0��� ��-�{�1mn_(����
O��^�'��_d+^f޻�Z�=�!\��s��!��Ԣ�~�ԛ��H���u����r@���M�dD���҂���7 *�s�U�3F�	8�]�&����0�W��3�*���<]V�g����1��r�p߃�
�������Ia�,�`��M�4�躀���/Ң[���0A_�tRD�2
�B��k��&\*}�/fv2 �l�\��BN���H���!Sd0/#F-��������_h"�@Tv_G��XF�ݓG�Ui�2=c�iBU�t�a	'�d%�{��w�4㄃�DsBu��ZVQ���E[�?�1џ�u���N�dpA�,N�������#(�iK\ڦs?���x-�?&n�@��6���8��(���(�`{
?�A xhɜ���t��V���I�v0b�2�XlxVHYEB     3f5     1308�wR
w��7K�~=�}m��q++�\����[zi���E��"��PWA���@���y�5�7�v\S�@vY	�KYMKZ���{���m_��K�ܚ{�==�!-���/~��z���ݱ���v��Ŀ��e�g�T��i�ι�"\�X�j���-��-�^���ʾ�I�܇M(��W.�IlTo�-d8�B��<�J��0��/5�G�����_S2ؕ���>@�W��]��3�<���0���=2��W_t֮���]�-��UZ��N0��K�2�����S���㪊