`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5alaGn0eBHRiM7FruWOzKvie85M4aSdRh24y/N/jrynJKfrP6QSg8JhOBxEiRHgjNZr01kBEq4n
Ele8oJQC+ChAOHCtNm9RMukMhNEdiSDPw6+4lvxOM8DtylRAoRnJT6vHikjyeuEP2F3tzl1G3Ylh
qV2DPvWLULwzDngmmowX9UP1NhkkgFjVW+zK4SF69DWOWUUJ0Abut5R3cCDelAKhjn1A97KkWZFS
qwKCDmH/83WR6TubnCS8IFERYBdsk05hFgX/KsSP6f0CKrm/GJp9srPkkm2CBwczTt7LOAy4QUb9
kbF4xk2KqowiStfCGRx9JGKi4ASZkzP0R13oCg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`protect data_block
EXaHNFqxO/mj9pEfkghGZMK/5gkOSKqUqK2B7387R/eLVgLQrXiL25TBWyUnNAw4yF/qd/OoBLIb
6S0yHNiTwpww13PYWk1Dkye1EAmrvCQQ/rtPRTpbstPbpq1A5NhfsAEXq3C18QxRVlbYMfAwJ8Q0
d0X1577J5BJ4jgdOGyc9Q4WzE3yzF9aYEIObMOXZ/nTsc74vBql6MrWmVQxhKw7klzZVyVRqTBx2
rXygb4BM4rjtV9+OsJ6eRAZWbQ2b3Hu/oqH7qwVfblFN5aiD4ONXEdn7LwLdhaY0v1d2R85uhg0H
ktITS79CGQxdIREvqKiToNL8Pg2NztAt0/6FZwPxweYe4+7MDB9LYtaFkV9JpniQcERJvpCeOa+I
NURfOuUIQa6HNxR0Vd4cMwSE5VhfYMjeDYYwSfkyl+hfZfb7c1Kqtq2PMLCGHKXhXT09Id+3KyiN
RBW/1haIrhRnKEg63bDSv8DQUFPd5tZLqUdO5KeXdWesLHhymOEcpOlQMthyl2rHbXGR/nBZyfaJ
O0dzcOTaSaRkF8IKNPsYobNXleY9TVl0PwZ6tIBHkb8XviG1iX+WAncBZdWe7fgx4ufOZoivNxXY
tpXC2tMpb1xTBPm95CgAkOuzmnYWy1MVVuvr6F78W3Uu0B+dNSr7hJeBDe9SezLhlUuelWWS6mEs
8LxSEIzSmsC5EMkvTw8ran7yv/f9HQDJRbAdLq8oHQmt4O6J/A4XJoiGPmnIgPJrNo1czNXBRQWW
WiadXzJ1OtR7dLWYYnagrl5BpCDNTL3H5gMbYmk94HxiXNYP8KX4kEOHSsq9P1zTt4UxGMFzCKu0
MRD8gQaDlDI+wbkua5O0gUmKKA6t/SyAnw5vVNpvQCIewX6VRZHjp5E4QFEGdwppdU4q7QXlVeXO
K3m0F7AXSN+bUlLPgxZZYN0xyWSNzUePKDkCEwyxlAnge0glWEvruWWgBuQVISvDnWXsX3oVwvom
I/uGAYmJPQyNgM1ACTVRe6kE1JbG97tPNBPHKRqt/sHhgxZg7mgB7JG+7NKhWw06ZymihEFijuRN
a93S+AqE3Li9ZYXMxRK9S9pKt4b0l49n9EDt5GRA1IGLMro62wDUxBnZO6V2+DjQbUmy59mc2FBW
6N30cf9dbx0wKvie9i0PURnIwVYDC01AXlQjkY1xnEAsMtAHrKR+gIbltAE99rC7K1f+PXQZo85z
leiUUYqEFVCvHiGAj+6VP/YkZj6Bc+CdHVjGEuyHsYcQFfzKVkJOt8epxq1ThX4FKt5+BlV4Ps6B
5UwZLSI41K4ZROTpYxMRCCJJmwHcq4SMiECjvoXK8ib2bbUIs2KO7empli4z1n3kma56A+n/XrgC
v/zFPGGYLEZKk6sxImysTtuYN7gyL+Hmo9DKu819ZLPrBXwXBNvSp3PYU1ewFrJW0+AFePGD9zNW
hitokupZmCA3uDy8QNX71hW57hIwcA5PGoMMtQu5mC3eeijBjw==
`protect end_protected
