XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����y�yv�OM�Q@�)��j.M[�]�{���>K	��&��#��?��d�Ce��"o.���Ѡa�k�2�R> ݺ?y�X�=�4M���(��X�,�)�J��Ӻ0t��[{�>���1]@o�	�JtY���kmf�/�e�}_��m�
����ڛz<r����Z���܎B.�������t�X�'B�`sC9���E�9JQ{���] rf�q%CZ�!�(�,*,b 䁁5��h��ic �+
aQ2�s�f=&S{-����+�)vr"o�W�ե�f0@����H�S��̸�@�0���U�cd�O��Y\�d��^3�3��$|VĪ2��i�iV�8@F��,�|(o���i���=ŗ'9a�Һn�'���Ыx����ctݻ	I�)#3�������OE�<��!�(�ٰP�n��}����_� ��"���
R[Dl�̙�k2�=�Ì��}��w�x��^�"5���$X
�S��,�����́�+�T�
�����@�)�ap����t�� _��4]o�������@C9���}=�>�G��S>a�J&�d�A<㟈�5ĉ������Sb�r��pЃ����]�Dh���������fc�_6U�I߃[[�_3Y	��T(���)��N��yԟuU2K��
j�2�~ o߷I�NK����{�� �.�H�F�K_$�Qonv�"��
C/�����U� ac��B��՘�K"\�׋����x����^��� _ƸU�b5�d�F[
��԰��$P
�q��0XlxVHYEB     400     190b���Z��6����UҼ֢�T��+7�-<1����-����s�<����&ٺ	��V>��� "+��i��5Ș�cm�g+�g6O���	9�7�\h�s�Z��p/��S�%��W��Vs�{C�eSI�?ii��w�k�0uI47�_��?Y3�.:�jr�bn\��QB�cN1	�,��; 7	U�^���F須�j��������� ��B//�h���"�E��b%�3"�dI.PB&z�� .��67���t�����Zg�lR�A�����|4�L�H����b��+�_+f 6��tlf��$�#M�Q뱥�1C}��-Ln�\R�<���e�6�^N��B�ϴ�=�Rw|MPY�$D�������s��UP��A(�[n@G�����O�JXlxVHYEB     400     140	Ð�~��z���0<W�E��Ds.�<�k�m��i�_��=�;�S�c�Z0%;�qV#�Z�*�Ce�	�O-�]F�wLv�r�	�쯒��?`Cm�����6I!7S��L���E���:�6
oQt���[�~��H:���ѡ�I�D���|6�1l��]@a�,��G6%�$������)�+��{�F��kp�e4�U�.Q����ֲ�W����Ӽ� �waꧻ���Io%��:���]M���|���55��bct�jPwҹ�A�.�Qx6J.�y���ɟt�+]�\���yuMI���$N�����AXlxVHYEB     400     130yo�Ű��z���J�}�O�TH�J��[K� na�b�����	���}t���"�m�C�����ZSRK�q��<+�/- �w�#��q��)4=x-+y�h������\n�?��-[*���r?9`{����t��;<���5�@0̉7��q�%i���!�3�)���
�)��y[�M2i	,���^����/z����ɯ6x��7�������'#MK�P>3��s�]��
��-
U�%��cTU�<'FL�ݝ�wb���9�5᧟[���V�9�����J��X����������gXlxVHYEB     232     110X����z�\��2�����Z�r1~��Խ!=
Ĝ?�d\ft�E3�Pa[3��`p�c�{U�!����Y>F��hX�DM�����	HN����ՁO����c��Jc��mp�[q�����M�q��eFe��	��_�����G����#�PRo%VҰ�;�ɨd,d��h_?�c�)�`��d_ҪB#2�w�mX�C7���d�����--��&��T!��;d�B�$9md���	���qp7��~�J�"�� ~�$=������s���{k