XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���]�4L-�mƿfi���U��%B��]����D�H�~p[���&:>�uh���*$�@����X�������d� \k�TrD��x3�.�2$�b�GTg"4�6!rC���Ozʗ|0��߃�5U3fT3���~��!.��<ni�R �.���*��~�M�x�_�-�a���vv���;���%�ܔ��wJ��շ*ǘg�y+:f�[M)�bZT��u�����I��fr�{��R�s�2���ğ�U-��y�1�t�M ߕ7���iƔ�d��AnC���qi�lJ<J�����L˾!1j�m'������tsb�P�Ne���+8KR���q~؛s�&����*9�U5���������dp9��?2�ZAK���W������̝4*�ٺf�����:W8c:�خĿ<At�V[Ar^�d���͉��(�ʤ!���I�I��u��)�!RZ@_����G~�3�����k�.g�o��C���̢��d]�,C�RG�w�>��;��%2��|LQm�I����&�B�����"������� "Ņ}��Q��k��J��@Y�l��b3��r�Y��8V�=�����UN'��=�v�MS�G��1I�v��>���D�o"]L4SuK't=�.�q��߅��F2�U@J�v�	�U��f��8[q��_*Ƅ�W�ܦ�
����4��Dc���0+C�������s��]��O�m��iu3�t8���V4C�B�x�M'�S@�XlxVHYEB     400     1e0A�u^5Dj#0�丕6Ǝ�;3~�Ty��.P&,�'�����3)��bp�F,� vq*�����yޏ�olcB���*^&�<�x[�UͶ���v�lr#B�aD:2���x�'�%ڂ���XT3L��z9�-�(�F{�%�[�)T=��2�[ A;��ٕ��`{S\	��]!���e��+�u��\rK��7��H��ߘ���s���)ɛ"hm7p'�Dk\��!�i)~���;<�%��b�ĸ��l6�M���lLT��ІU����u/7�<I���a���qz��Xi��4,	��.Zr�p2E���g�u�@������t��Q�NOƹ����~ᓏ(�&�8���پi�8	d�`.}��U"��#F��� cy��W�Hޘ4�i�0�82�ϋG�g���[&UW����
xa��Ћ�-�N���!�1���W��J5��
`�
O_o����:��\������/	UܷWXlxVHYEB     400     1a09�֞�uu��A�M��h��3Л�k>�^���#����^�m��x<��e�$,0��+SBoz3�c@�,��2�-�� p�-ZIA��PX�Ր���w5��C�✧�x<�:����(o�R���B��?�[��t��m�K^69��C~��쌚��^�ޮ�I����d|�b��7�
:��U���Q8(H/wJ�7�	2��f~�dyd8
U��]�p�^/d��n���IOt�H��ݹ=�V�ڂ|�^hv�n5˚ MZ�څ+�u���م���]+�?#�t�k��m�b(���]�U�~�],��'���U��a���$�}
g��҇t��W������0KL	k�񈓜t��g��:�}�Exױ��$�U�l�s�((�]G{S��ס��&�;�0DOI��Wf�&���:XlxVHYEB     400     130�K��b��N���!�����IA���J�:tUK=�y3��Qa#��BZ����?><������x壖�S�4��}�%����I�y ��ugnĹ&}����/��gJ$�dc�#�}�����ժ�N�Ɩ���!�8=�B`�c����2�!^>�Q�DM/6E���GT�	�	��r��tH��2��1rR�CU
�\���RUN��\{/V�Dľ~G΁�mE~d��K.o�@��qN��59ueh΋�J�]���"I�6�U��p�3���{��s䢀D��G��n�ǾM_��*��D�&�иXlxVHYEB     400     150:�5l�R,C��*˥���W'M�a{c�g��M!}j��_fN����A[,f��t��?��O��� ���(�.�-9�.���g���<�E������,�/^:��A'�}�����ɕ;ݴ�o"��Dthȼ�hX!���jq��迃�8qy�"z��K蓛;�V�ۓ�l;y�]>e���TP��;��F�"�s�`5���9��R�2�s+�&�GH3��k#�\)����C�n�Ǡ{�'`�l�"�#�u�Q{��|����#�c��-�bFu��������H����_����$S���{�:��r"�a���<+�'�K\}ڡ�ҫ7 �͵iB�XlxVHYEB     400     1a0��\�ޙ)'��w��/}Dl<���[��܁T@���L����(#��Қ��y���A+�k�Y���i�A�m)�y#a[��S%^���e��֬h�]R̜t߫�3�_k����
�sl�iQg,���t��;�@q�wUP�'a������Y@��d3�J�D��gK�Q��"�`(�q�f���^��8a?�E$��r<��&3� ��]����2b-��j�a�D:����28y�U�mH�'6�P�m���q7m� �)��u���<��4��gM'��� NǾ��X�A�s�'Hݣ;��kΨ����;�b��?���'������x=Pv�]�BL��4ye�хE�����u(��9t=`�!�q[�8H"^aw�{l�eſ�{��bö�^�Q�Y��u_��7�N��.�㺔ZXlxVHYEB     400     1806�-ݗ7�1/�s42�&��!~^��ެ��X�i�^�<�����G�몳^_��ҨNY�s���5��������=Ћ��`�.[g���+jP9J����+p��h��&z���� �=��!� �2�W�kI����{5�b�����I}�5I����r)C�q!�:!�I��d�/T�%?��!0�B����貅�@� P
�>v��d�C_[*�kz��xӰZ������3����Gi4�Io������Hx���U�����k�bt?���C�<|����=c��;���29�Y��1׸۸�E�fr��9P1�3�ז�p�!ǞY�0��N����+M�-�w �g����r9[E��R)Ru�vQ�H�%M>XlxVHYEB     3a0     170�u�7U�a�����K)����E?Z�Z�xS��5�:�M�~-$o���^X�.�1@�P�Ss!�������P.�w���Խ�]꽦� �)ێ��g�*�M���76(� E�\�C%:�����6�.�8�fD����\�����&��:�$�s�-�?����.)���~�l����F�D>�`�����3=��^&���cI(��"��,�}��'�d����꿔8�E�P_���>��:��*�8�^�ݛ*����nҗ�AYI�h��ur��H�?�S���,��%I��ZA8�|�b�V'_���O&���f����R���u�e��j���ä�!�m��U[��OkO;�X�Y~N
�����(