`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17056)
`protect data_block
7po5fNOXjoGTFqnLAm8m8YSA+tvT1L0JMCRL4qOV8dWryoK/UE8OnYadwl8LiEspp/TbPhdk2y4V
DeRMdTQI3wyyvNdB8n+Bm5ESj3t9R/QqHlSD/RsRAXbGrfUzdH0/aUX6j8LcdBJtMJQsHe66ZCZ8
PF3B4fXAwZwOGrzaUVt45scxAhPttCf2z5TNvHw9TqY2v95nuCODoTS7jdUn9BNyODxu1jnZ3ids
BXVxOGC2X7zAMMRP+Tk/ndc90BecMOD0IoKureMoM9VqHG9fc9KrPV3dZ5V9mxYSAA+68M29APtx
xPztbiykLmj7ZdCCY5I9Fk6Y7zJkhdoMWV5uWzY3sEw96yfJx2uzKsWDjbdjbZAUxp7zY5774+XO
NCm9v38+yszs2FMo8h+vQ1W0Nfl0URvayvHyv1qAlghGwWxngZ9vaecuh5HCNm5sQ1wejrcVJSq4
XOeibgtc2kjwSAOvpuPN6uyqtgGg7iwXrFSbQjIZ8NWIMDPWAJyTdvQQrEEOgEMz0KLE75sAulFk
nQbnG4H02jlHYYm0fWhUYQ3+w2qj2pKpt6zECUNmp3zkxKKKmSDeZMs31avXGY6Xe0D/PNbZSl+0
ibwM3fVF/WFp0kHmKMR1IwnAaw35VfsvJI5NElSnZaZkcJZD1Gj2VRfs3WnbcNpNjAHHmeX3RYLZ
Q+FUjjt+Sit3/4EidXe60Mna58BH9y1H3mvddQdUrCzzZPEbhAHTfOri7mWy6G8yG9FVN1+bn7Xs
MUwIdpYgx+O9s9xnh6o+MR5qOGzRy78IaZEaK77UeJ0RqmayfR+yrx5tTxK9GrLirR5fxB+G6A+j
NIP6M69v3mVdBJBEaYss0C9JyCla/251vPPBrP4nwsjooIXFrFYIcyMSBCT9Zjgj8WtkW+vAGc3y
QvYl6TKe4aLWpoLRi/f83xJEETWMBebb7ibhhP5Mrbu5o1drxeHEimWecMNY4QsQtSd+IL5QStAH
KybiSslf41VXpm6quZqTKsd/sdWMAckaEbb659bVjgdYN52MQlX8XaKbyXoSewmTZe/7sDhzuB61
tKqGQBVD/IhrtlE4Ua/c2wyUGP4luOtHwHYg188k9qWikq35t7cuuCkCISaOr80+Yh87FVYLlD9t
dmCe4xxIhAGMNTLNuESCCHUTxNpgf7GoELVnVLB+WUEFn1O5SFNn0GiwJHhmU3i88aIyuwsPgHdJ
bBf3Fw4NEtVyZIb4XlRpHnP2mXmWr52ChGsx3bwV0zpG7KN0XgXfUzRxe4VuGlKISyp2VtmPo8Cf
wCpTl0eQMlQLMmWPdWCrnEAbsSh59j3MdQ0/bxmEEs2cxukLccV0oMPwtlZ3O9D4DCugtLcw/qtX
veYnvMmR6B+nwtdVNhaxzUnytEm50+7jrvEVKAbn5Y8/mOwVtRhYLMJlU2VBrHaUw8NnBgH1bIZ2
+C20J5z44u+ZAaHAY8qrf6Tn62TZ/WiWp/SsNcqTDKb8w+1Wplg7LAZnF3Du43bitDP1xjMFAcNP
Hy2IPp1weuNn78NLYJss5rmiCKjsfJG/WfviY3no+4PPoRK5qnNqF03Ut8QTKdnPQEPKTaSvz3A8
kaD/qTYx2NuCVqPHbVl2Ckqze+NlH/MDTqy+ClzmaxxraipGfmNev/H2eNzmg0XFEIiyPBMo3/R4
LxzT4Nm2cBQ86iW7nBJzV7SXWHUiZcUtUR3/nBletJXJnI7t3OoHyRSbDlzPRJDJrIGjx1qMvZ+s
140bBLBa+szfgAX8ARLHIF5P5fB5qBQrYv4/7Zkf1diYN+7f07n9TqbSh7meavtC/sYgieaVS79w
umAlGxPLRDWS6qwcoscakH9D4eKAYf5WJiMmhXS8M+10nH5mAkRRpJcKU86VeJqo8aCxWPJu5BIk
+6cJZS2B3S6SFnRQ6lHItLkxU/rrcZhChm+E9EGZ+gPCK2xAENvAJd86N4BzwLn15NzBE1Mm8rx7
PFw14Pf01Vy2g2VdgT3N8pW/DSuPFoMbude8YDvsW89ZwYQpO5rMS4hz7zhgWFKDXtzGASxMd4Hi
jpbI0ObN4eYGFli53hOY8UYFfeEHUTJWteQlRS9A8mxOCjhqhgZZbSaUzDkg9olIBQtzJgwJ7UCZ
KIzRp6LiZJO4IUAUX3iy2aZ/DZBBbphncMkAJp4Rtgr/5ie7AuW+5muB1AB5MT/EprnsYKkq2EpS
2B9ofO7TF/AOWWxZI1LAaNniiU8/KMGD9a5jtagxdhywgsH+pg1SaBW3IGcPrBsMEesoTohOUC9R
1YGm0gdAMlGKoSESeRw7orTQb+GonwuLyhbBRDJSrG0Ya+2w9RMrK3XRuNe0Hg4TBwalRJkld8lJ
FSKHGXDFBGGlAgrhZoDj2tpskoe230g6XMyYc8UyEY8P3pMMgClYdPqQhR6X7GF4o0QLan4pBfLr
gX6sghooskbHb1dgs8j6unqx0fKMPUYRXDsWfOt1uz8PnJSjv+MK1pYSCaHVvO/3+MP0WabpL/53
fWMCoz8dnAwhqkpL6eFEcT09FFD/hkPbt+k7nwwDVzXgCqR4kDLHnrtPtoHDEWpy5fCrh8CZZqea
rT3cu0Xwyz/uYMFEGbsgRii5kuScQHXx2bssO9XF8FCdQuB88dq6orzZgfiuFQadnaBfkodtVDY2
3aMvsU1f/rhDslbwJho5y1mB1ghBOh97BL29MJReeV5l6yyYLz1odp1HNs5sEVUHFbgn6bL22HGY
CZ4nsgMnpZkfkI7uF/5KOlHZ0fHRlXUn2RItAmtFJV+SqCVXQvgf9O1b5MfdGVlEdobFaF/MJqrp
IKHiyGpQZf//1iDd0C6j1F+tT/sR7fDrAsNgCKWd6h7RX1it3pnLQseh974FPCJDTbqoA58WrvCG
4augHTyQxN/e/u9NORJNJ5d5rxwOQo2wev4tMN6ZQyc1Izjdq5Pcm3j2qL7071vOf/2APKyqLBDF
8Rkcnmm0W8gXIMDuWWz64/0eqHVne9Z/3m/7OOjtWXqLTmyJm+wTyHl1vI4K84p/Iufa8+mPM3V9
uLrkrn5WX9cTux8cM5OvIuOV817xuyMFh7kHTbrbGZDxyP5sIjK7QN+1lhyn87gB1EZ2LDrHqr5a
Q8GHbDatPgoxvKemU2GxHepvPTh7M1Zog6uobwkpJmZkboWczPbRPTXwOcV4tzTMUiU6RA0jZIEV
qYjUZUxDwcvA/KQs/tBNdr2JyqEev9PtVFS+496xDjLMm9C6pTz3nZQwvVrLI1vtndu71K1/OY76
6ufeHY57AjsFRyLcA+UBSE1Ukk10MKuxSD6ppt7/X4P82EsOKel+JRKXf41SgC+vRVnRhujj+3HU
/SP4wI8tmW4piL5jbVNrrOKz0xYMx/0v648IdHz3jH8mYgCAjDKxAp4cZwOGoeYj0wgIr+4wPkYt
dlN5VLPp7jOvY2SDXP3qwUcNoLkNdjIiCIi1MwjpgtXks4KaQO8g4eJ97wEQ80z6sl/3SVbPPgmM
GY/EqPVYaJrdGY+5NWoxqN22NZ57IwanFRqlPbRyXe0PVJalXAiFEh6A0EFxcpjLoN2D1AFJO90r
OtAU4jgfPFOnPTVjCNYfv6VNNg07zKhLkWda7xPagdAdd+yGWsW6BQKzZZBJ7xqlyGOoe4qYJJe8
O7mmW54yISraW4pf495wJt0A6g4w86oeK9QDk06xXVE/cSSTMH/VgWl29grggV5Nc9MuI6gSO2Bg
DfWT7V4qjQ5cm5noocG8T130EmaLwjIse1pLS/ownLoPVLBFNyQqjlr6A7WGj6YoYmpe5vqJIPNM
6lPFPhfyCYNiUpf1aBW1hiuyRJdUS+Q3af4aCx95ufyBtDBnAjFelcT1Jas/zK0JwBcIs0bybkw+
6iTe7poB+185nN+z/g6oyPVPDqCAu1qTt2DYRZt8uUxpUPnXuWphBciAh4D9gMzJlwo0hIWUuxkX
DXo8M1Z9DQ1Lid9RBzcALg15E2GZxKxZH6rAVLJ2cVev2iJB8MH3yOJqnMSvqEQON3OmSaeNVIcr
j9TFpOIFrqrZ4dKH+6c7PQClpnHDf01znRbTkE3awtWZ3eHFfkQyUGBdWUVrzV2g4uNSQDhnr/UQ
EHDoXAqfo0s7ltlbUTdjijvU1CEBYuCL17QZlvf5jzP417HaXPrzLxRb37m1g+WeYKvOcZXmz4gp
lnT+ginQyl6VfnlmSOJrdL1u0ZFpvx19GUpxbiKgJE3Sdesx6GPqiDEwy6sLBoEdGFDNUcT9cCcp
H0NC/bInRIkPaJuyTuGSHaRxaXQYXOUD65jRHWnKSHw7y+CUwE8aftC18G80S+56rhPE3XhCknXB
RIfcy4Z9uic+QrQpBuZ8cwgbA+ixJx7it944PTlZNAFs8NTpWPE+Yam9MKa7iboha2lcJMPQ1zfL
WD6EYFGK5eC47yZP8m8utu63/5M2x5/U9k9qQBXCZsjNMIGfd6XlsRY24GI+63G8FuMBqYpxmeTw
8ABxEzlAQNfjQUFtLwjejtag36CFUKEuo0GAVHsoJtgbiewZLnJYfWXUHkpXg5h8RkWNT8VGJR7e
+e8irqpJC9ueP+K5Pnvxte94awwFddK0GlzpM7jftT4yUA3OVEPJhL5Mai5v9RBwFk1tOY6XEXVF
A4sbfMIcUnZd28pDU+llUTysFX/4uCJdluaOaDdMnzFMQUG4J2p539L8vjhh458yWbMd78R0r0nX
UPTZH5idOb5liNSepG+ACs4cUfnQajBZvmU5Car09n8+o6rsTRR40hf+HDTVqcRAyPjR2wlfxVeq
VG1QuCTEHJHHOqxVyYzEAovk8je+N1AAITUu3DjyEPnBqTsV7SyybqOsABFUl+7vbU5xHHDGGLtL
0xVfmTCaEq5iLVLYdQiJgJAcvVTIIyNamnZagGrmFf1scTvgG6+/5uUHgR4oA0t1DWGGbrGKgb1n
AxDWJZTcY80Fzij5/e6ef6eS4i/JLhQA/dREvtODfqs8PpJ2AEpueG/dy3+ZkHgqq3iDH95GF6Sw
3h7p0jYjdxKxP6T00dUEhRihSve9QS+0usKOeTdMvMEAfIVoSdIR7yloKt9JosWr7TV1Qj5Nvkst
R0Nzcin9D6Ob5QFE4GM+P0IsGV7DjWXrDkDwDQc96dx+LYX6VNK/oczIfirKKQLfZWIETWFz7gkj
SRqy0BTJN1RP4mAbNqQtTo8V3lBXJwuCHAt04FVh2UwkTowQ2OuDOZgnjusS29k09DZSqJ16shze
+fG6rNrTEPYVHj+P2q2GRh2/BBmMXcWgIARwU9I/JuymSFOOWWO0/TpkVZQFVX+Rf8Gez9soVvCt
Ptwa6RjCww2COrMAzyRPyUbWb2QSFQmZcPcQ2Zfy1/p5qiCAb4oR8R6h6ey+nzru/u4lITPBtPZP
PAX4ri31JQgne8GT0PsbBrCHTUKzxYtcnyjL4n7VEYwfNMVnem2M95PboCoRjF+RUOn852qqRBdO
TFIVpzGChru69yDM86z36dbJttjKI/MpsEMhT7wY19zNyY+EHt6cH8CapfcH0UOLRp4msxA3WufK
zbS3EYGuOvQ1TtWAVkFh1HsaesFAnJxxgmfstZI3I/PLvfaAHNwdiAIpUcNZZqfEBhM8p70yzsGD
w/79EM23n/vC6oRBv4kdX4fCOjoEutvfLKjg7+9jtOV8QqF+L1boRh4r9H9i//5/vlCMcL81p0k+
W1mkUlVWx0HLVMVfNqjHVAyFrfOjJGnbYkrUBspZb58OKSpKy2Gu+SvhL6XttcdaloJebbuU2KI8
2yjxIjbFJl1fo3ZmIZg3R98DsmghjB/ZMK725D0yvP+I/VrJo0XeUZ6O5+KXkmpnheRxHfEgN2KR
5uRGATi6wiT10RI70RbenV6UHc4RCxeIEhpiR8wPdEzL3y2W2hE240vrBylW3eYRi6uabHMbZ2/+
BhlVuY2HG8jmhQe5NTE86CJokId+OYNiULQ5zH/rV7ybdPEvbZGNVQM2usWzSijpLCzvspzDlWoL
yH42/8Cncb5UJo1MOiHAElFJE9lAGtpbLebV6MhAAQ6HOVNxUkpo42DRJRESnarTGVKAbqaxrWaO
lFcmlPTGyXF8slP5G0UBgaMcVAy1q+wg7EnpKa6DKH9EJKaf5IebOCEKQNLmVMkpV0Icm5wqOxEB
lkExXkIkTZjF12f1WSZ2fZfZM8vq863GNlKwa8zSeS+6pSGhQ0Uq2GPT/M9NDBO8nGExqdw6hIuQ
KLieILR17OYyMy/yjaa8iPAOlE2Rfk1upfXOyWxipZ/T2+dIpn5AcrIfOyAiiFlTj43i16G5L2Yl
cqhUcq1vLlkcyzxAOIcn2zB5FzNsK7sGNM2lZIh5jn9KzONCYqQP7PZKxPTOOa5R/WqAU8TxMzc5
NhNZ32mszm39BrwMoFNypLwd0V1dzt2TLZxXZIby7Ye04BJcvmUxlAfK+HrycHkEF1IZ5ey6CbSt
fB6CTacJ+HXHjbg6pyifF7lCquYdTyDh/CiBwaMrMXBEpVeQiSadcfun3J0jAvJvxjkqKfK/Zm9G
DenZBUaiyqVxcIdoovO3G2WJTG+bAivfevN5P/XlSdsNSEUfVWL5/8q0W6yQ+DzmWRGUe+iWOzfW
QByXp6FOkETquQ0UYVThaWCv8x27333zH3x13j7HV8b/WjkmzyCjfntms5zji3RO0lTErhPx/mqw
+M/wtA4o7Z0AuWOQWXA4hytTdJzHk4HJrGF/FzU5ZaBtSsBwXU5w7VeFRGjuoWdNdW6sgKG4P9ly
34LVL0IKSkd2db9NIRzyhKkjg91jTGhhMsB9EFDHKDHAycyLRWhP28k82UzkOK7HFZm+NvOE9xeg
6n+/7ELwdewHhi6Ikno06loCU8I4xZa7+dWij5lHz04dXhYGb9T79R94GOAqJXl18v58Kg+M74U3
eBHXZLyJNtKc2rfW5kUj7Fa0AwlVPmt2juxpr+sMOe7LpFppOnrhJHDEWqA6orDcHavKQZetcdrT
ZSqsNJBfwcJsfRHYclA8PWl8jqQWBm+zT8GGI/xGpQgplUysDDK1utQzSoiTNaQKhO8MwkNhG/oo
Hmw3WwRJquOEfEV2eC7CLCRzW6Ut22fsPdinkVUUxQn2z0UE1sw6TbcLhGkyNcHEP4lg3iWgO9Y1
ItXrQPKShXHm79UpcYpKJ8TzqoHkogPeQ4O6H3tVrcKsTT65NvwnrUNw61fkJuri5w74fle38PIQ
gvJMdjrrvjhGkDhO2SuHn/q6j/5Q9kfEIgvrnQVOLAW/6aDLrTPtYFu7zsA5SsXMsuwl3S/9jZdo
u0ilvkdtscon1kUat4oUVoizvIOyDqN77HNUYTJMqbud4hrplZpRCTfopGzQqoV0PzcWiMxeoXvq
Oxr1SEIXHs8aTmcT3JFxlcI0c7K1Kk6aMvVUAHA2ngNCr3TVnC85Nx0M3yEbbOkLrMcqBOKqD6Zc
c9C4ti4uSXntsXFXkF6IFsme/g4Gu0SaomyOfPNPulpZaIK+qnHfkRYUihtm69O922ei/DNdQHML
/05b8y0RKeKA2OzW8R6n1PJBxivDAMOatWdU/ucQU3cn/yQeDqaGXVfJZP4vUO1dCcq+Lis2euzR
jhN7k4hlvtmKcc5FukdQFQw/f+6eOBdf2NBnRru8vCOviP5uBYghQmJdb5v/0D03XMZhPFUUXfUx
2Y9daQKNEHL4Vxi4CnwvpmSek9Jjc+FCX0w8csDfzAVeI/2P0Uq5hVJ/q0m87LNJgdfV3TCbrHEV
XWXH1LTIZrxaAUWQ7EYOoXEkcQHxufrUG1H6ENV9vfT9NPkl+l4/LkH72et107k/PDEgb/xf9nND
V8tT73qhuH7X3VQJJPsjZOHqXs5bJddDO7pRF39S9uL7yX54BIOS9nxNVu6NZzLe0YrEe/IUUgYi
HaHR+K4loWqKywEHcZn5AboKYt1ozuz1LF8DWaCIZ6MMzwU7VTyS3ZzgFtmrtzzmrc1/lJPEAj4v
6ug+0NAcq8Cx9FyUMsBmXg0Kvsp8+yhVmY2IBlIRFr00qzI6kMXCDkIECH/UgTcRTaavsngCVK01
pW/0Zqh1fvzg1VORFuABKQ/LYBXpgWJJxda43lmvWeAcrZbJprXnq+MBldDJf78d3nUZa+T9UqWh
X5H06DiduKLNeDYAvL21XPKd955b//a9gbBhOL4Nz5k1suGtV/h9g6LqHDno39TxhxttZKeQ6wbt
dcA/bhJaewhFLle4Ym1DZ9frA/m7G8MT3YoMp7a6viYLp/iMnmVDifKgg/PTMLsWL52JyXNMCBy1
+s5QgN+lA78ggXzJeMV9RNd1bQSBXLHH9IymVWBZCr7ciTG68vEO970rbfp2P1E8WTlLKRW0z4Yp
xzYoAdiZROmreJAZKgepMZ/QI7xCfknh/IfuMCfKOdcYAOofd8EjBZzFoprfntkGekcRlWrpQlWo
WV9hpzEII5BsMEwUTmAkyrd87jOsEa9EwYp9SPwgAJTGssWrG/2j6iEEgOF9DfjCUlDVGiTV0YSn
d4saYj/CQiKveylLbcLP6V7k3pdZ3jt3TUtkwgnkkiTp3BgooXlzfrZAi3G9jfOp21LA2irRwCvV
HohIDPqNFSD6fE/JW/nBmiiGfL2/6AHP528+nrufhaSuVmHylkIgc2iPLB60Fcsw2nt+6PiapkQt
fCaB4W5aUqoVYEamdQDEfWmZjZh0nn5aDMM7FkAt9Y0q+p5+ygsJbKKXUGg8CGnliZKEK7nrtw1H
Jtomb1ndhG5A3ECxEzlr1ytUby4TMbWFhnVXR/dmhNHgoLwf6N7AYUmesjnRYcEGrBch2BIy80EN
DE4Gf0W4FNSc67DfCZWOvfmc1DH9hNzC14HqyJIz0whupbRUx6Tmu3JLcCzRmtM/tsV+1waBbtUo
V56xrZJjkLgJOfvi7p8X8vtgZq9vD8iZh+mjC0fV28f5KBj+gq51/U/DXapc+0uamBEKOLncYRZ0
/zzA4mR0vJXOLt63gs+EdWD9AcfGicsl5pNS9GXMBTn1blfBYl8KxqCVYggkl87AMTxA4zq3wAcQ
hF6awwJEG4f8FsmV6CnUlru1UrEXW+436YRJ5u7P1jR/hcVJsISAXznO2k3O4phOWd4m9NZMFufg
+eIwD7C1+OXr9hCR9zw7rZcs9toe+oKSWZaY9ea//qoiFF2EclMvoD/6uojOEayR0SW15UAoocQ3
4ecc6QF+HTgIqkQMAMu78rkSFcYa+aCBdLGyTWxuVicGyqRqVHwkEQP3xDCK5n0KgDWDrrDt4FUc
mk1A2OmeeJcQVo5z8gl/vWkiEFvUfW8u7ONDhSYBGe3BDJjmUevhEOnnpz0AectzaZaJp3RC8qsq
thu/nCnuxjglQy0bK3sCHVuJCPZg6kHJ7+g7Uh/ZgT5A4zp7mpRkaqnIRlVCSKdJWzZcaFCUkPLU
q0IcpAsYQh6eKZplIfd7TELwpn5yznYss4XP1fdKoZTx9WpG4bpKwzIQUVj6clpBcm9lrhu2BzEX
pgOcLInMXZlfWlRxEbqBvOb8DSFzNYsld7ggUNNO5or+uvmSeaGl955AQ5CoSNLUH9GOopsFcARk
PJ4fquqR3MB38nHYdMJawWWmnGxP9ojVhtm7RHcwHAf8wDGwQi2I3/1loA+iomi6zcJMWCkRQdDn
cmzgziv28ZELVqwTEgq9K6PQVFWujTo9pVuxCLlNvSLNn5mF7TjJALYmzLxHNJPBIjewsboLGAAl
zBYRJqBuFzzK6r2uoT7V5YFoJQJQUN/KVgIkdlz0goOOp9rV69bRHKQCJ5fGrht1z5CxM0JU4aBy
N3S5GVhItd/VRFG1y52Jk653q0Ty2IEBpf0xObxc2ef6rnq7EHURm9NGD52wwyateEG9nyr/9ZJM
7+alwrQcHVtMUzoyFL/3UWkMhCpQ65Pnt3hskpOMb0S1J7f1j3T9F5IlnZWtGS5GGpeJxwepnYDS
u3HOBaDpLXdyaFhue+dO6VAFYFJa7nBymYWo+bagfGHA4dWB1tAKgjpGcCFf4jPCbij8Jmeb3B2j
FCp+N1BMeLp1vJg5fV8roo4nJD+JkIpW4iET0F4N/mDc2TldfiXlVWTHXy+yeHY6d8LfFsM881dm
0pQgKKOjTRToBqBwTL6iOuIQ8Ycc/mD67xeflKSc2gAs4IwDFDQFpUxrAgGzqPOV9V1HQXCGMKSS
P/WFHUrClcgjYFTdSHI3grDxJ9P+RpPDKkRcS8YO1hDsv5ZYZvH8R8S6SW8FMbhQdmAYq7XYaNXB
69dnr9IP1r7hI10j88xcgTogOMXYPDzUCz5WfJQZ8QNZaE3oS82Wz5OlwyPFWreDY0kZT9FkLwcx
IMFTNOFrzNSOUqZ9bC41upit3cZ6pBd+bp+04zk/QiaxC1TE5QOh0V2s0uc0AmzfvcNgBvKMaywm
LDCmJqhYF4SG9FWAG4iE+5muVrMAqMmqLcLQqbCbcBGyqD3VMxzRblPFrs4/CvK33/ISs5LKvk1/
Lx7SJN7I91nem7BCayJHuffIFwRPElTQ4+RyipLiGd1YA+KstgvNfz0aDMnq5nsBVlazajTIvxKg
U+py1PmstpdiEIs9Vms2lJHK5VmZS1A1Qyq5opASX0aaLkRzXYau74sGbkZfuDWjYZitmTWzx4h4
skxricyb9PTGkqwq8wuf2rj6DXzcn9oedJhnDqxZzO15HO59QpBRDyOnOJSUvNGi3ApKai6jSn6f
poDtiTdwR7si/sV3z5JTVUI34iSr8d9D+QwBJzfQsnZOTIMTBeFluNvrDyCiMHIODumI5eDeHmej
x3pA67E/cC6kzV1lHE2F3W42fPKYqnwg707TcM6X+WKvoVx4iAlR9RzJKjdEA/WgdrcESQQ7bt5b
4nxhz/tEMCKWuj4UyWQISV1oO2M8C/lwuesK0eKxhXET2EQmcKyGGo15EYztc3dNTcJFY+OabrSG
zDVtaCpvtBKLiddWnP+x97ScqIW7Jj3E9jlXSornJUFsQFckPNZUkxteS/E5m+OwxliDgeC1d5bB
dCqiSjhj812S5SoQQPyGeqO/GtcvtBnf3CLIvp/zF2VdhHdWbyYhMdG2EbMvcQ9rpXMkSPE586jR
xMczmG3Yi9O7QS622lg4rcstEFwbqLDLY1XtkO84rkb5t/sC5/i78t1pC0YykkbRhYsvFbmqhLn0
0bZpolALkWMXlpgphUFvm1vAbBnOp/8wIfIVRS6uW/lWkRewkJH128DUrxjz+VRBgNQbnJrWWsJ1
nTMWzv2BsQ+SLccupcvRePPpf5zFQ6cw72PQzxRGKpmdNdeoytKrzyJNWN28nZs52Amhjo4dZj5G
c7KD73XAbNcc14QNvxMEyD3umtARQ05in+9xMr2W52uPbMH6Gtz7OILITAcsnkSLpJ9TplG6DSFe
v3UQgJpCNiwL8rjwKFeyxquUU6PoVc0wqCJncC8zMFj2NlwEsC/T0B5OWyXIOwnhIB/Z1NtzfgOz
9KmXB3YV2CZizbq5c0ebAI60g9L5UGQcnslh5+XOWQ8PAHjWawymuoLuiHzmgeeB4Nwz3BTUsYNp
naawWhPSDfWUkt9KfrcAPTrAiVvHKfVkLh933BmzBe0AEcAKoeRSeKbjjc0ua54GKI3UM/NtlvyQ
6MLxOU7t4rSvYHiWme6ZA9u2YNSHtbl/hrbIFrinU4qFflWy0IUB7+Q9giYc/m158ZIUPgMh48jY
SyW7NoESyHFA6bbtr1gFnTOsA9nJk6Y08CSzVqdR7TF/9DXea/57/EeNFn8QcbjAbqnTklMPbOVQ
HPDoLc6kd/4K5Zy1zdjMizRIvv5MWAMiRKITem4pZCCbdZGaiUrKp/u4NLJwgBldvIMMZyEZEIlj
vPuyppJJ/ictHGEFjVVsFHzVeu3D7C3YTwBk00pN6gn4ywT8EUG5f4+Z2aOnFWAdi6k5IEDIYSoB
8Ic+PvShgbnTebSycWbbZorGg7KzFh/7XqT1YtSx/7eJs6OL04toRTQvyjp2uK5/TYmKHD9SYOS/
nBdLHGXRSfDmMzOTYK6raV+S3VvzodB/KCXXtzmLZk3bEshPgdfVoHdpPB1WC2iYC8ste4fzxs24
qWNIAdjdNlA+2ISH5iw5TQB1Y+GiJrDwrG/b8OUI5S4I2fysMDmVqnkk7Hyl3h3cAobS8YW8TBtE
bKg2Ppx6OgCOuldxuaGdhwweTzyVPo4adlm5CdnIudFZ43cxrtUcYSjz/Om0grKMfH0rCxeEJpF9
CmmZdUtTS9AQay4te/1iN6PK6wqyX0f8eWeXWuGxmdzThbTlpNlepjXk4ki2e2uCndn6lGK1kVVb
58e9kNVhR84GI6JPDkSgGunWFFM+m//Qd5ZFB+zM0HGvriPIO3IM5vgRnnlzTRfBsd38zKbjIBwu
fRElb4CUia4qSseRBhrWZi2kLeB0CUAc6Xu7386G/B5rWUrQc3Rryglk/crikOCXHENcO13oIc9D
Pshw2o/eP2YG+0bkhG5W2SRndo2sLwzEOvq6EsTZC0Y0ueCzuO0kaa0hSAJ6exyha3NeSvc2Oqw1
QRsORA3Qs4d8wIdMv+dqiyNfdLWzSj1yA1mZFUbK94LYZZGq5wKoP/z2O8+uFrHp2kPf5pX3T4X7
wnxI7pwlmneavmZphhBlkOBPM6XXt4iL63LvOAwYDm8HRfA4PsOyMnwgisCyq7befGpBYsYdmQjr
UXl8R9kXtEv+UOykQthcn65U9nIpmTaL61o1xooo2qh6pQ8kNv6/lKMnR2lZr95NDN/EofaWd0dA
X/r8OWVTrLNmdACXmI/LAjYSLr6bIdGZyae5NEwghegwKNY8iG+nOX4nuV0i82hA4RsquD4fQaKd
zmgWbJRucrYPov0SE45znOmij20jK/XqptxAlSGr6omb/4J+i9/bAWE+CTtIQoEK784Gwx4OBctu
F2A3HQYPEdqEx17PmdBsmZXQg1TZz1QCeZ3W1qQ/VcLt7d8Sj6ZcdwHvFp67D35AUqKPbvoPsT34
T/AUOpija4+yMRsvjDDw9j6K9+oBwVdzmlQTOvlrWPP/XINhavs4bhrBPamdkKMpH8Orj6gIEAtd
CiQ0kPDqFXMfEBSu4xTzqHoG5cSgWwDAGUNcywNZAB366jlcykWAcKEA9QHacdkV4zba9v0OuVyx
/l4AEu8OkUcXIfauwaQbw5hmxOdBaYGK6pJW8Z8M3Tku0G9jyce6G4+wLgP6IQb+LNUNgHmZwZgV
lBJqM6VMcT3b6VfFxGIeSSPBQAN+IW4iGe6irMsR1DaF6eIhcdAvqweJWsBrAf+AgojkCEIsJsBI
8p499aThuiv+23rFEtMI63YJbNfvZbuMC5FOvDziR3mKmv0Gx95Fu4MgtCLierwkW4xV76VbEd2k
rtzo72PxgTx5zgIZBlfC3HazTHagKCScoHy2OGfb2BBxczRNOS0XmM6L/cD3uKJCjDVf0SwVwyER
Nvgf+kTa8ymCfQU/aPMZcL/3gGAi2ZbL8jWlFn3AYMxbBnkS9FW9leOuQ06Tc6lh9FIfSg32PuFc
oOKHSJgoVFrf3Q8x+8KvYPhJdTGfQ0sZD4fShyhlAXq8+/1dQo7n1ZOrZKu+B3jG9SNK5K2gsfpY
nWL14IonYNkLa3jxQbAHtKUcuqSCAFnTEB8eXVML8KJz0PafQpDOEw60EEQUrly848MZo1OdOtRc
OHCqb8GiREBqqXMOuA2jueydvqQoAgeU0GuxnwqL4Q/yRjJt4pvqkQ1ThWB5+Bf1l59/NTF7+oJV
N0x6d0k48yMhIJ6FRL3+t4l1gwggBUqBdnwB+G6qO1WfCqYydJDHY2xsFnXfQfrKnEv0X4hfqWVa
Q2whMOgf2zw/+TXOgRxblZGuduKdLhJjeTobWcwUPvDaDkzkyl+Ds7n0aQbC3LQPTzLPipwiAQD8
az24nmO80s1czp9fx4YEM6UA6UHIOqp/vRwZOqh76TNviwts6703+PxjQ8FeAAVBcBfImWYAeMqf
rS13JB14f7zNP0EGS/tOFc0TZzPo5bs1CTjXvC6/aoJ9zYo8jU1UxTzoMI9Fyd1BPg0LZaZPJga9
J4+kSjPHp+ZlRWh7EjFjmCJaAIIbO+FHnOfuT/M3llheYnMD2568glqG8qhjPwrZ6gf9dtx5JOSF
av4bkxLYoQfJRTD5wbYWh1cEAUNTTd2Qm5kkDg+eWc4JjD9pPegpkAq9MTJtqYJYN0h34cAD1V0l
BwDm8yfnIvvs/I9vwHNUlnk8KU/TWs/I3A8ZN/KcOGvevNC5YoBtWWKwK+77ROTAbKwp+TIfT4L5
yhGD+PtvZcFBxuHVbxmJNEWdzY9EYszB+gbcqSx/Ju0xWyr6wLj6AnNpZYFA/KXSuHRPmqYSSi0N
DOLhq0c69p5ptkgJVoLN9R5Z+qoiVVVjUuQ/6JNZyErfHfqV5yiAAHFiszEe7aB/kZ55UrSDmXVA
0Ky28jGhwM+qvk+2TcLMuB6wqG4e8PUFbwIFoT+AXM8drPGpuo/T9j7KUl88plRVhkVeaQ39Bebk
kh7P1F7gJwO7K2zCAceP56y36RgYhP4n/B5Eegp+iA0Cfunv7HJXNVTq7Dfe3IGqyCr3eSRf5Bh5
C9lZj65jlKBmZCvf2v8YRQ3WysLFzwEZxVcesn7OEiCp6gK6aVnG580C/4b8oPSqwHEOIOEYZ/2q
IyrZpoMfIsHgFVJR2G3+xMrtHolvM20J9UKJHBa2lNyyaoG2kIoIpasfdoPdoY/qOQT263katpTM
0zwawnDxYX+WVpfsCdOptjZQWJjNW1WjLDv5xPkXz8N4SMG2nVf99PilEO3EPyJVTmEJGirWxH/w
VHnBvyURQTA2aS2gf6MNwzzK5ptzcZrDtk8KxnejrnqopPQldLkLC9kxIaYWEeD0+CQ8HAVveNUb
awCw9i3Aia3xV2Yj+TPM9JT+wDeHR861iRBOc01NNw/l2CsaZiOFnApyjOBOiHXaxfp0TDc/ufd6
jubHtSbwepeIOtY22jy6HzFEv0LSDEFcyPYkgXvWb3fmMKHCEOD6l1P6WZVMa9+vx464p78KXDEq
1z2ZC1Wb5VGPVKVVWrF5QVmaWLIlpv7dmoEGcRIkzsNsprOwYbAKwe5rS3j0UVW9zjLbVVv4FNIb
2Eeu4HxPwFsxXFCogJuRTk3MiS8tHk9aGAlgCvTMS/DZNMyb32TFszpiVvr1jq/6hymYCRqPzEIO
KAkkc7gsdfWPuUXdM/sU+Ax5bfz1Ip/fVhfrEgbBv/j4OVhJ47E3VhJaORR5oAV28ZK7YMoCB1io
y/yY29srhtQmboN6ygJJ5brvc3FotBk3MKV6eXJeVFxYroVVE1mRI2Hsvl4rKxdk8hLR0kYoI/72
kdqK/I595YjZ06vXbXoexBJy4ic9/Ij9J6OTfl4FVtsaqWEvxKSsKvxR/X6sJzVR6GbBU8OrwKHQ
juRfcQvmPyDlsIYU8w7b9w5tv3Eot/ZnFE/lo/B1ntXoXOYhX/jGVJxm2AxRJsToPpCqj1Wzq1mt
ygkCEC4y+h1QkbpXk4JfOuJpPO+c41l+WkD/XHRRR1nKkoiPC8uM1uwX8FY77o8yPc8u7svDEXOo
nyans518peOuciP7Ied66skKU8+thfVdbxbO8VTCwq6ag/6Jf2cZtd9A26a2iRiFsOHiwLW4fX+l
I9Pw3f+7/3ZQlz7Uyu2JQs2LBkXK3osxp8Cxw33m8LPoxb0vzo0iaDgxDMHCXfe82Oet4YJuW7CE
YATHr8bxrBWmgpdTq0nkhh6hObJPh20nMiDGaM8TC8QdvKY4AWZI3v617tc/1ZhcaKp4/pGJ20Q6
52ClCGgGH4XQJXktzBCJ4YHH98kPcfsdgEPJChpZoK3+5SI08WArimfLF+WBEHIQrmU3VOA8CoTe
MVY/I3Dqv4mfdO7MlsVnuVHCDSiGwAsIiJ8gfxkTJus+KFc/FWacuRLCYR8U3uCrqd75z3skZu8e
8kWmpDEMme7Ab1404eD7BLtFtqPvtG9XvccPWr1FCHVNVVk1kD9Mwb6RYi7Vpre5Y1lFu2PxWsr7
RsWY2lE7QLh6NK4HBm5TNyv7wRvAtfh92buZdgFcqF7VcR/yCdIoGLy4L2CM8Xr3es8b1EA5XllT
qjkKlHmWNZy0Mw6KTLP2kVvR0Me5D3qo9+oHAtF4o2zLUgBMwwpIyVZBJUZG959T6mov5t9kNvyx
xaA38E3y9eCLGkdWQ9cain2IfCW5ViytCpD47ItgOpXnOJ5RLal2fC4pDK12Ua9Z+qF2wrxKjKW7
ZeENO4f6Si8haBNX8ziDfZOTNRiZDB6AmTI4gdw4X8wQlCXI5JP7y8he0WqdY4Tup4oa7wvWYHNb
xOOS4BwB2ELRPCaUoebQa6Ys2czHWCOmuSAaEAzj2iYeKA1vGCUW4rCgxZi+n0vGku93DzBB9+sA
zEdo07Thl0MnvCu27ibFxHngWAM3bm4qwWvWoCMFRVCKibxkTNkc8j5Eiq5jWY3w0IRzKHloA9Qu
jIAV32VMXAb/6fsRXiuobAO3VrzUGPcRzRs61JZZzjTa2iMA+0xf+mIpm3N1tRD9QWakemfrciPm
0RaVlZoLNmXSCNjvvCKdLQIpH1i5I0mhoTgU9H4ygPS9bQrUAqjj5Btm1Sw6kFXujh/HXSeyyzQY
qcrJS4hy0SdPV1h4fDUbsJWwVZvdLidaIot2fsdGvmWXUygfQRVrVfo8TPtlkAFGWbcD2cmBkGiZ
grL5yinc5+rkh+87jaZQMktpJvHNyldHz5UEixISBSNZHU7pgbTkoMsXWqFGmiikW/DQDPsFkQ7F
EdLwWi+kVFCcmMSKju0J58xEqrbipQeLRBq0cDKdABOQe4GBVn+LlcvKVX9MH8PLsjZUXm6X2df/
aDTpTVxwQ7KvwK8nG8+nDWHtqn37wvDp99MfKCx4ixPxtKYMDGPofuOpDpfB/Y+K/e4ztXyq5qLx
MmotZrJd3j7c6c4zOTa93pf5NbB/32Rx74sCsVFU1ky7+iYN19r1FXJS2kzxbpdqnDdyjdlMgjWQ
bKAmngwM2h06WnChycnOK7Dee2d5fT6sFrDLkeBPHG/7FYcx7E/vKkAvoWv0ITupTUkZTf7zLsEl
NHS8YQUEb3kECBkNlfU0irdat0eBnHnZAk3Kj8GAVRPtEHfC5KhVEOoMtTNofx4FuvaDH+d5uwcH
V2bjJJqCnd29VKDAaK+wkFq7muGxvVAR/cckiUY3T/bBKmjv14Nj/fry919u5pvaFAv5ZCKCsnqd
MrjT3KMA1kwSEkMPtzr9EboMxioIGY2pasTkvHxc1LnTWYP/3ovdLdzXD/ocob8aRf05k+pePmfm
2R9MOlPumEm+iJt9PvgmxJcwDR779t21MaXSSPRRRNgJq7++UIZppxsZ/TE/7TW86A+1QZtzyO1S
y/ECTt73xREST87nAoS+FbYViDkD8wT7AWtfi7lpCkpXNlwiYBFteqdsyteTWZ/VlJOpzwSWUhjU
h9F8KS6geO2TAbawLQMEgrPqXWL5J6TmMiLkD/mx3+3a//VKWhBL+FU1Q54Zwyz/7aa0oSBELCBB
Tx0xCYV79Uzsg3mcjdxX/NDOvDAEnj1YPiB3l5vYRCW8OueZs5W+/3B0W/GAngWSWS/sWQAlX8tT
wNCIr9+zim1ilOnBLb5c5ADYAHABdxCXJwTI5amXx4p7PtQl2BtZPrk7gngW5YzpaKByDsNWvQgd
tMS0XViZNNwvqUofIL7Wvzr+zmJg14GKQSModdFPIaoKwWyDln2BYu5kYP8y2Wa8goSKPhnBYUW+
xMJ34jxYjtI2Vluwmd/DZQ9TIgVXZza0JBTKZQ614Cb9HDcHu8EdmQjPjYv/qxTE2CdJyjbXWFAb
h9osrWZnL8Zky2uBYnP1TTtR9SVw8JDcqxP3/CM2W76kPUVJSys5nKMXXVEFNMeVK/Rkbr6pKg57
PKbgzWCS3/WGfoKmy+SzJ1VL73gLjR6e681PnPGjbnel2bl6r2vb5y2EPBqWVrzYRHOniDHxiKKl
87hwEprWOj3B/c8tyoVTRutW70fAf9FPLIit78eMApifnhYL9V/nyto/Y3TGRr8yu3OSarQ/gibB
pHUnutM9Uhc3fRsQHKkxyCQIghrbprBV4dvHuF1NDnUpkqeR6nQtHZzmWEfYSBnL6DnFG4Bm1VAx
WsM8a1C8CU6t1e/kvGFMTpW2s3kvdfKyifCkvOIjicNRhIwYxhiLLZGRm6IHHK1KYS0zf9VZycMa
D4EYBdgHFHBw0C59tQHLecIA/z/c4PKw8BaFAS1tWjAjWeNZp8qNTrNlYgukvtUSWLZj9t2pYCtm
QLAzy53cPsagruVLv5RQUjWUhdmTb8BQNK9nZ8/8WGpUeSQEpvnQKONJ1pw3ktcsFNt+BjqF1CPL
JgneHEdFzJGBoapSG+ENPJ52aizoc8ax2KigMKWvW4GHfMl8JOKkEa5s2kUi6p8O+WZkXdxpywhY
OJuPaXrJcnw8cv8M0nGBlBAqpl+D5fjhP2Z3uWLp7oajqngKFIsjDUk1jQQ4iXz8A4i8nE5Yemwl
lK5y+Eq8Uam3ZQmbXlCz4Khco+4cQh9u0tDMOchzpIKNaiCmmve2xmiPEm7eaB0xIQcwjO7w85eF
7md2fDB6Y9CLTILQ+oFVfSh5Qs6xOKqeU+AppPm6+N3MtRqP5PS8USt8OxIpwpD2o4JgwxnD8+Bh
iL6DuGv+khjyeMpj2MyCJWrR7xk+t2MtoIZrt2TrTNAFtCVHk9pCge49h/4/efTpLG6MraOTGXKq
nALVVbd0K7crz1SNPL5EU4ZQlJrqhSTP1kJxHhPUT8NyECAjxMKYssM8H86XN9ACR2EZpt1m+1Kf
n9NvPmzymvUVRwnCBzWQ0rB7B5bFpwR3/wD8QI9uHEwFe3y2VkHdvXxiId9iXHMpEw40A5dkRj02
QifgETyJ2ne3ONG/D4ZBvsgO33BE4x4pfpwb1QIH17NSS1TSLWrXR5Da2hpj6pg0A0NKzVKAnZXo
1KrxVQxGW0Z/iegmmr2zhjfz7QNeNs+sWU8FYyWX/WejTYk/JG/dGuzy2Hcsbv5OwZI+MlcRZr11
1SlB6Vcsh09dMx32FM4IT3NKWk6NpdO2mLpXGx5E52eMXZQVjBreYT48dNdeOFTsNkdG+4h/7jmk
x4F97dMwzx/9DzFF3cCap681YLJcHsS0RLJO0LbV5Owm3NOKgPhXLTIiqVfKnS7O2BwkVpRrQD6Q
n3TpionQNqTRosh0unFCCLdh0qkHZnGzdzJvOQ36Qhexo8Ws2g5JCBzXWoKAGDFHGnG8wiAhT+i3
7cw2w63VpB2Gq7SAkaU88QTK9PNL14muRwaHDAH1DjY8bVlDI89MARvgLDsbGLCmv9EXg2UNUTwn
ViQIKc4nZgmnD+TxCt6OcUAdiYTc+lzdPLpcbbr0O0ealJLhSITW/4+b6JwJz45PYBQFa5Wi+3bF
woNRwgFou6mFTY8EXXxck9PN6ia4GakGMBgPlEbZmA78mmgNvKtie5iuiWZldCuJNxFf12fRzPda
NVlJmw6T0v07sNzfRuiq5m3tVwfZKC5MceuiPmt5zWUQS+C+/IT25tUOajvKpcJdOc6w36V9t9a7
sSj9WfCGD9r7V9kL3zecSnPzZbjz8B5yhWj/kPeYoM39NdZnduHY/9Npsat8MxYtFJTvZA4RXqSz
M0v5JBq42WTGTUDoUuUk3yh1kWyEe8i27iTuNpy24Mis2dMqWKK2sA+Z+Gw3uPprSTT4igxpYg0N
ZzvW4YMyUHmiMbQJN9dvRibPcNqxRphV2vvrHUVYbqK+F6WpSoazxnFlBaM0zdOMpAPta30haChT
RiSuREg0RtFLxn/qLODOtcwt1gX3bvLvQt83dIILTRDJPIH0h+pwgF2Q7jhcZ7eVPvNbqe/Iglcn
bxdNcSs83a8RdLS1j4PrdSbq302xS9BO+FY2wYe0bB9Tr7yAd9xC9TvNca8WrOuJHj4MrAwQthXP
ZKKxuYgTwFQC+KMSw2uLwb9SPgRvoIP+BvApyHdOcpUBrnxjXmJ7IUAsX6Q0wLPEg1/RbSgskYPT
oUxzpm0CmT278x8ymf4A3vnvI2CmHYTe7nk+rbiJC8l6XCxUdAQ4V6EORwtfejo5oufeaUBao5AT
HOg4R2TUmaONyPASLQYhVY2pC1bLMA2tFX377I9+Ywjz9iCp5I5czV6rb6ddH1kSap1E6tEZS31w
36XStgYq7XZlacmAUI6SFsM2ejEgCDrdqsfFoGVfBLI0JfUcM4Y+jH3aQg6V3krSa4EKn/rxcmYg
GRlINT0XBcVdKqBJsMGgtmDSPc1ME/co1tI73/X8WCwOTqp3A7NQg6JNSQaC1Sy8HwPX84r5+CJM
td7TqO3g2GhCaWx1ugWGACJczDgtrro+DYwajOXjENEQys/Efmj1QtFvmvu6ndWoqi1TVa0duQey
Gmz83Hm4LyCGmmcEUZdBjZdH13/O+zaNP04uX7c3K7Q/Tu0r/W7ZbkG9SfqJgpqNcRyrFpH3NEz5
mz4TReZ8WwcgmIeH7+dkOReq/EixQ/LK0BYiHCalEfT4KWi2EwWnPI25MzBmF8D5TUKvxTaOc+D9
2rt8fNyJfuu1XEX/Lieq5cAqE82I/Qrl4a0J7R6QekTDrEOfmOa/5BNHoP1inEFgHwNjS9pvQpF9
2a8xaf6kwtjV+BK+PkGBDqFf1/ZqKXDHOdyPHuBVDltVX95M5XSr8TVl9qY6580WJtYJ4UVcqVkx
LFF7qxRSHXayCIyC0FK4L2CzyU72O0DMn0C+51dSdZBKAXONPtBh3l9b5sjznRtQfgk1g2yKZgn/
KGfSUHvALVOcXnxldE+Sls0bQ3r+rjGrnTnao1D5d56nvi/C1MFg+BaczVwtNe1Rb6snEgNKLSJ+
jUSdcTwAZt8aYguhYBsISDZdiNFudNms2AJrYruBm9QBeeCXaBob/ltvEqVSb8zbUt54EzTdEuS3
1O9Vgw7vJJt3rFiDH2siehjFN4f8v1GWaekoiuEbN2s9aO9BggpL5X1lcElQOOOp9Ww2vAequDig
0cGufh9AdWD/oqM9eFlKJFgWL4U/c0fyh2KwGsjlTt1g6kM1KlN4+oLwFkhhsdRV+aSaGpI3nKmS
jElvaNSBForcKFXddcLSXR+XNwa21m9cD6acL+0U1wzVQKHzwFclyu27ePi6m1msTUg7sA38kbVI
/SQOkYzV4p9+qxqTlkYVwtEIL9Hbk+VMklxY9PXFTEn3aWIIa2Hr4x40lr9PHMdKLICzRDlm16cO
qPir+A7F2IyJVlhdAvBg5oqr+SLLNpMoxVS0fX7XfgIrvaYcU8aazFvpN9PEuIKoDwR5zp8puHPH
A3oh8hLDXVjMMNrhF5C1CSJ+h6GXmzZY3OB1k2WvypgSxes3m7Lsu0Vkv3y0BNYUcFAwaKmwd6wR
e2Rw2I4dQLpOIlFf4wHd3DdvCwI+W5C1rDcypxNq7wlgQAWu6aFFOsV+inIm6DwW3ZjWIpEAAjtg
z2yFHkOZ67T/GvBObsZyP1Yn2XWtuC55JJc+PT4edacPw7J6cAnFz8frU07/gOepiUJwJL5kHvLP
i0h8GRCgiWds7xDIBt/cYoRDWjLG6WVTXiOCHKUxgPgdthL828hKlwmsfAeZhxY3eZv2tqiCtGv0
VIrk96maL7EjNPNZkL0DdjBdwAK5pIIKb696fIYiri8MqRq2OYQloSs6Yej29eGe7Jlgh2SiLEhl
kyXCGc8IC9XK5IN+Vcp5HKLcS5y0TiQtLcxKk4Zx4aTzHPLRDes790xs8BIDDJ2EEyXQg0Dwy46o
VGZibcKXsQnoo+avsn83F3RTyZryCmr/zmNth29oS1rff7/A22rHSacNZYoAI5/qYwyKmtnDuWFa
ynIGD71MrwmliA1i7QWseEe9fZ0ZfdzP3oEjHWN6UWV4NrTj2bKUjRY6Lk1YSL6hGKUzCxooY/GD
UtY/zDcPwCS/NwXiHPi0ld/bsiGJSZ0XENHcBzZNVOAfSMV1z5E9zmEBqEGL8fEuimQXS19GkjAz
J0QaicUbUx3qLS0BSzzEPPvrrYJPJjrd2orjsnDLObrCUUFufDeIx6QRDe+WeUFc9SobyB+61D4R
gGiZT63LESsH4sAIM1tYeZszir6z/MXkJGLxgQPZooeQnbnPcSnt+4m+FdJWfjByEoE7F6jHqNS7
SV95C0UovDlw01ytyTkF7ofYpKP0uyK7Fz0T5KKWUKj9G1Z/61WeaCl41b7PpjIo2zSr3xN3XorH
4C7JLHJsHLWlCfmkBsy5Nle/ECmBXi0MP+GYYJ9ojnnG2P2d4BtU7m2bi/iichIHM808wBvafpo8
R/VH5eES6kZjZYff+r18HmIN5Fzenl2pHfCT1HzfvDjwKStwL2SxsgjGppjYyluhVrqqZALmR4AD
XgPi5Ulgew5IwUI9TuQ1fy+GQCT1aFdsPu+fJSgW+oeBFes5ICas55z3NBgkvnE/s9YbrnEPo4to
nzHbvk/KqbfTW5QwZg7EYkzdIMNJm7qP5+k2P2N0qJAAZ/86TKMqYmmpS4Ggk8d0F2JjJnpYzzns
gVOy9itKegFjCHKXF16epS8rywGVhZcxPOvpvUWApOAoiUxiWCR6hjrE06NBFDzJl/N92cAnVvEC
SidYViexCRamuo+WhurUOEiOqeuNTGirP/cHH2PjmJdYa83CQtuCS1LlUtw8DF/I/6cVow9Zjw3j
eTHL5qSEoYVwpyWhLg==
`protect end_protected
