`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wluEddR4Xhts8EEuwgjKb8cuZK2y+RrD7cAzSTBxYGwhi5tcX8szZgGz/6K1QvJbbflicZXEOiDx
GGWTAbtkUqJCoNnXTJYtx2HOcH30WbUR7sZfhg9CClWXaBmSYvtOKyK1a3MbbM50R6vWgR/vlKlf
hq01RFyADZ8qNhwS5s6pednZmt44qMcWHIujBPCd6I37HQYnpOSbeZn7DgUNvhGbVNVNyg5PWWWV
O/0fAFsGDPw1Xv3oHrnDMG2wGKOKI1sDFR2eEnd17HrmawnFNihjr9/AHOrvXRj4BfqYWHtqUxUk
EPzabuh2NgpnPK210zifjm1pvI11LEWlS7gRiQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`protect data_block
NUnuRKwDOiMsykNOnP2Ddj+MU4xmoOMI2RU/49aWxxkIqtIkOik+NY3gYh3rxnfJo++ypYEqjF+i
l73CRZ3AuoiCnla8vZgrhaf2APIGbfVFYHG9vdYa/8DcLS9PxrZcvHm5PO1McfBU/AOzfbse5i4y
qvlFkwF57NC/RVZnuhnj3izUacRpjUbTYrgy7mBXTOu7MhFxA1qbijtVFCKosKPEbrIr6tTL6+Af
3DsFQrG8XE3urWC7xODUqTU+TePZoJa0rMnpbL2I6FbziFIPp9pCw9rTrr0Afi31jxw/qFNM/gMQ
CbPC2vEJEWTFZ1hDaed9FtpN7uPV6ZnSbr40EGDTGoT0kYGY9xBBoMgX0GAfEZFLsedEtunv+sec
c+PnEBbm4xOWPl/4LZyQZ9jzq2NPeNdSLYdQKr0HaFVZi4cUJhgQVs3ztZURYNcZukZWrjvkLEzX
z2Vw2rGYYjpLVvjscPmg1yDIDU572xnyo+XTMo8kbe6Bm/Agx0/O5C7iozDy8f9IC4X+X82fD3dZ
MfM1ZXj6oaP8fV9jaRlBdDQMNBSOH5XCTPTtymhlwRPMsHYICcqzb+zTNb2euOJqO4v5E86fqNTM
Tjr9vV4YMluM4VZ4NLNpmh+JEWJ0HMw5bfWAiNmCz0F3qx2PDupjY/YhWFnzDJE+R03N4sclyKdg
/xR6mfSPg58uEetf/FXu1vBYj/Io/fBHgxpjwsKiqwVGaTXN9dhuY4AlHZ0kawkOtgiGycsg9BnL
t8z1dxWrwh/kiMNe1Jidthx2WB2XrbNzaPbxNiMngcL/JttQ2+zwWnVJXxvKrXnhcNtzG4sr3H1A
le0S2ipEZCx7j2Rlj0IzRqhzQ8Wu6SyAPMZaJSh9Pd6t+0iPfv/yiTz67IQIM13CoDgXXgYZX8xf
qdX60VOcKuyZRPRU18hDRCsQuEg+IZr5B4St/onkYkz3La0EXpnnHofTmcwZITGrEOadl1X7KWaC
yMBtgrC63DoL8Rnrjjx3A4O+mnAmVivJGt2uEPG/T4YIU2nmlDK8I0iA+JwfEVsfm6pm0Wu5Z5IB
dD7yoK9BGCuropYYUBxGFwzMGjMcNBoQkcrFzGVeq8OAQv5LO+z1yvyvI4vQ4/qIY972q7bXG9N7
VYKNpncKsQj/rMCFSxTeJihhscdEVNHw6AA0zC7nlKplKSlZCcoJbh6wG9Lj0TGL/J9vuPboyMaM
z0dpGc7sWWNBPU5SJKZ7oKVwO+cclzM4FPqgS8A96NTt7M4ja4R4AAv7rUbJbZZ9igoF+dc02KkJ
cv9OdlaI6cJ2ZJ6YZ4PVwRV/E+kyQG6KbSnDhvN3EIguCdKYSt5B2JnpSL9d48IPgjx6CDYAP/bw
WYe1+TVqJEoKeER7znAuH5wmbWERxxotWfN4OlhbzVCnQYyHzUEgg88V+P7ljrev30uI9P3FqVXB
WoX7JKAFgcJZ1Edf8rcm+qMA1Hg50dtKEPqG0uNUnAxyDtE8URGNbf9VPYilNFW8zVpBY262Yhbh
oYnxjp6hmWm+7AUOZsD7Xt0zrgM9H9qVgQ7OVi6ZQwNNgfM2I9VVU439h8oyGEPgDUZOE/dknftY
gev+jGy2RWGIcXv0xmqjWrekN5OFTzJvGvA505Wl28RAyICMmhf3BcA/32JOvQnUmHdeeJ7XsI0R
kcYN7PEhLSCMt8UakBBDTrdR9LgwQWhsAhsk4KP2cpkhYQF2sMNBzaY3vGH7HQQgldXVANtEqrQN
fk+vO059jg5l3rarlsgwCVbd8zvcX5vkyDX9x/ng8vgaxE14jZcexmONq0l4YWa5I8a0HkYm0Rse
BRQZU8UPgaqk5CWd6gbsv5PnMpTbPORm/5+BY8eS71TqZoQRfLO82r6hlGVos5fTf8jGKeoxFug7
/mofktOGPsziSC2ny3pcbyJZPcenTML5BHMbzwLesXENy9bgMw3fqVcqK3uSku7nrCtpNT6EOu8C
6qqRrpjwUNsDOQOCO/yrwxex5KpDodUyQeU+5pgwQgDll94wBuGNHnDZ3j5W9/FxionbOmlCD+m4
v/u7VIqtukA4/gQDNbgtAerv2CoxFstRRftSWOv3OekJDPU62k5KQ4SKtS8Yv6Hz770gZJWhU7Cl
axNJBrCqjXCwdnoBgmnVUfWfbezcwFcOdb0qGKfC60+1Pq2oVAVpjry88IJO8HgN0LVdf6eqq5uN
MTyJhpOcM3EZK5qv8u6hDcG4+fLrvGw+vzfsxCduPOWm0gn8seywg8OfglTR3AvI83yqxfwG+V0v
DdsELQ/w4OTCzjWdxnG38d8ffWetlQmW6OqoiSs1VM2AXlLgdLyBz1xzvV2NjmDx360dPePlHA7a
s4vBkfE3k03ZqGLKk+xaY3cYiPAecOTXWvYW+2F1kq5dF5X9GfhDSwEEe4dg++zvTmn+EgSXXe5F
tzZg9/xFKGK/luMCAUSQbyZSlUQI6qfW8a/SKyKqMu4LoIUl6XFoEiRPCrp6qo9hQgCMGfa6/10u
FREChtWdrH0LJcMEq/iBd3cU3d2afu5zuUKX9gbcZdU/TBAABcayd/GhHpzvpiwHU1dyw1xjiuBk
BRfhiMsEQY669vw3bAeOZR3hLCI1tErl/bEGPFT2u7Ie4DDt+gGGj15EGB6JwBeaKwBYfc2tZ9p8
3nrOYXgkO/XyMMWB7adw6sUNc2eNqqWO3zSrd9j0X9O17ykbSU/hxEfQRnRQMMBod4aYiTEW5OjV
2mtBaMcsN6HpcAwF6/KI/mGewiYjtcLBLj325B0lPVQNgs6ooIzBOByHEUY/QLXEqT4o1zWa+vUU
BppLANEfNEd11cTlsQgRCb+3cbKH2UsdTSQOZ8gu946NV2Kef4qEwf98zrGSaBow5IKa6cB+zWsf
N9LBAiGgfbfgv+0nLsbozJEPZ1Xs6kdCTUTi7Gn1L6kRVai//2grRbbjGlbTgEbyWcPtunRDbHhc
DxhfOQ+1Q4vC8dzGjLLmFhogyogbadZExyzMTZTWbuni5ZPUWSWWt23wp8SxGRyDta7H2OFx2ZzR
xy0HlvNXOJUHFzm6FctmfLv10vnxFp0AHlYT+zDbywE4BSiaeduyuxzVa5q4mYCCbYamQ2vBlZV6
sm73GPQkbtQJ4P483MhTkyFvbJEejDs+mL/u576aVBmwcvHKHBgYWmHj6dmWVeYLmim90Gi4YYMn
lDTcYlYdGx1rF0pWhy3NWLDAKBSN5EFYsjwrP+VmRGsFIMpNHHO5zGhA8wsxU+quGw4wN258bJQo
Gsg+mFS1iHDJlcuLmy+UXK3NfJt80ToPs5dKhhbKebL3g+rvYSEIzipobEEfXP5hEaF0rff0ACGe
jPrZ5wgjUfqgfEfqN1D+yE06tlxPV5E7EmMcypJjtDR64tDJsLiNaJk8sP1/vgtFdEr6B/Rw1LzA
nbE5ftfOy43xKzCmhXB1CblUEVmXH6Z/x/cILyrv4y26ZPMr5bv/H6PnuaQceeCi7pvMy+eWHhnJ
6/YwovidWChvNgvPrTD9ZUP01kAOuIA2hBYBIbse671Wt5LN4w4Kgt+u3LfMQwSCIzzMCKtb11aK
/wZWivZuqid4JODLhoxtX2qQvXPdjI0WgvjgQOmpj2734auQgHwUJ8yzISLBihA2oPovbKVneCkU
c4loqe/dGWa9SXDMD5GCVl5zF3etnL99W29OTntklfKgkIFs2znOd2G9EX7q9jf1mR38rDQUXcZm
iFRjPMNdRWhItFE5TQhCyR9VLeINSbg+Yn17Kun5+O4ivoUnYHfeRw6OohSFxQj1x8SAAiWE5bMn
VuN8Dq2/FftGUShnJKsVwIzGazIsN11UQp9FB695lCadCTawAYtva5UiQJvFiXq3ae9ZgX+XuuV0
SEXmc30fDNOJbxdSLXBDfumjV9NT7sSaXHcb19LvgoluM8ZTWxzj/ljmSfgxLbp+kjkRnbHgb1Ly
y0vwX2GfVZZtyfPRWv+541S/X28hbWod6latCqjyDTdceSehHeijdPap+jNfkn9FbB8GppHtQfmY
NGp9n9DiGN0rPvKySEycdMk88/QOeV7VwccnquzfWBxKwAYYGndrIkZeHZIE1AAcj6Y51bcJj01n
kBbmJctz0yTllLmak58ALJMNV2UoPmxBOefkCCeye8m/bk0nkiO6m/jQUJ6mTTxMAFZ65TB3XUmt
cQr+pFslCrM3//2QmvnQ+x98hxyAHjvErhZCOVUk/e/hhidTkhhcdmM9rzb87tglalJP4RyntqMq
/93xa/i/iyRmDIAbQ3s++hhCpHZsyamy5g6HPwZ8VJdPeQyAWRqoGmy274432286gODWV7Ji9D11
TOKX5OA0NicUZjeRlf0QiuXJal1BMD4Qh1ZzR/fTpk6vamsS2uQa3FEFz74idvj0S8eAdddWK8tV
SFumY0labHOODDlb0JWCxOqkftvPCGym5e4w0BpgXrhRWVcJKuTrZ6p9R22h3Oj/GTx1yLtir9xX
2AMw39cI5XzunNo/qI3StfBJI/OHeTg4qkZ/laVxu1cjq0B1dXC4GkY0JxvoAY0nY3uvyLlDJHxi
IOeSnNoLo0aX8BAK9uZzbSLPgHbJHnUOpWfyKvKCwAzFVzZ6dMt+fsHQWMgvZPWcogoVV7g6i5Ac
CLYxmxs3/8shGtY=
`protect end_protected
