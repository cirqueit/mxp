XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]x.7�<�l��!������bm�,,!�[nϻs>'�ވ�r���Z���&���3oF�k��U!��Bs4��v�V�_~(�T) ���ԕ'�h0$��9I!�C^ac��#��P1\+�io�Y&�x�7.��'�����	�3Tw�[+�~tcҪn�א&�^�g3����Q�\�<�;�a�H�ī������	����+�-е���_<���ͻJ��x(=x$�Փ��B2��&>�쨶���=�s��|p��f�U_�����O�q��&DܿEU���l&��.���+�R�D��������j�;��,���'�C�?�b��;�f �$�_�kfƝ������;�W���@�l2o�� w�A���d��)|�*o]�-d��oN����
�ѹ��-����/^�¬D0�?N�L�wŦ���kD4���a���^�EL���i�j��N�<Xa�	#w��$�.�'�.Fih�y>V������1�.Ҫx�����)��bF=>7ȼ���2lB���<��V-rmz='��^��'9"�z?��6�&Q�>����=���E�����`6Ot��RYY�Lx��"��(�j���O!�������ٿ��6>X�܄�:�6A�ՙ�u��Z��!:���^�c������q%�7o�6
����xW2W֛���H�oSG%�o�"4��k/���uD5�j=3�8��\{bƼGgԆ�vLL��h>� ����N���V��:�\�2�}������ѝ�K��L�XlxVHYEB     400     1d0��� �m��@m�}�]<�ztɸ��&���p�ո��޵D3O�C�l���'�ƚ&Y9=<�'_w�?n��@ſ*Z"�[�*�G8g�� k�O��t��I_��m!�.�������ͽ[Fi�\TF�=VtOH��.��tތa.P�Ec����hha/UY`0-�X������0�Jƕ�wl�ZfT��,xTeΰ4V�w�����1��B�t�z�DLP�﬿&'����DÇ���rM=�^OX�c6�}�W�嗨m�����Bn��1�dƲB,��s�	:�it<����KPP�"�<+�"Ռ�����8���Pt^-������T5��C_��4���k"XS���NkX����"��W�q����Rq��6�ڗf������^8��k�>	G�Iʼy]��c�mҏ�-���d�9���4�ܥ%6����4KE�o��1+�Kf�۹�XlxVHYEB     400     110���-*b�m[�[1�ݠv�{��c-��uF��&�owu��?b��y��&yJț���I����z+Y��Z^U�k�����I=�S!?�A����������&��w-�6��~��P��њ?\���n�O]�(/☟.�'d�b�~�Z��J7����)�)���kdM�{��/A�ΓP��$UnD�|�]n�X3:f��kZ��l��R8�Ŀ�~2cX�4��W՝Jg}�K��� �H�3����|��IgF����"	2���D�8i�E��٤TXlxVHYEB     400      f0*�H�� V1.�kFK;Û;�Z�p����yZW�l�Ԍ�qn_��F�������T�?m.���8k�Jz~��y&��r�$��bT��BV��U�7�PN\(��OF�/VE%JC,р�S��2~����<�7�R�Wq�|/��8S���}+΢�^�5$�2�ܑ{�-�w9�I�h��nyw.����ք1/�1�X��cC���/iC3�
PXe�y\�����#�V+6�Tq����n�Q[XlxVHYEB     400      b0���+$`
-���zN��(�v�j�RsC
�I�^1�'�׃1�tx
eƆa���R�7�;-�����?*��U�����M��6�a�5w�x���%�ʌ�v����Z����[K/$�=�$s��z��M{���������-A��TP���7�-m����/�bq��	&�XlxVHYEB     400      d0�I�3�R��Z��<#Z�Dۛ1K{!^u10D>��ձ�u_b˷��F$�9Gv#\2m՜�AB)$rA3��U����pg;--��OӠ�]5o36����=]��p��Wsw�����}Wrk�!�7%��G��8�����s�Z�V�9B6���
�ih k
_Xp,ZDO%y�t~ޚ�,�Ӫ:<� t!�I�8�r\]4o�l���XlxVHYEB     400      d0 2i�5�����;,IC��\\	�B���2���%���3ͬ����V`v�����I����86/���	�阩f`�F�?<|�5d��-��}G���Up��
/���\Ԅ��rlz�m��^� G�t�E ���~��6��)��h�@f��O1���<����G��o,[�9�>�`PPV�G�(4�\_CB2tw&�оLU��8��XlxVHYEB     400     120N�`b���/���uU�}C3f4��I8� b��f*̹�{?�Z�ٞ��^�P��ن������`��:f>en��`�����8 �/���#Y���]N�z8�UL��*���Q�Cٔ;d�e�����q�N����T��WG�9g��!v�$�'��b�.I��u;(:��%�DaJ�vZ!;zBh`w��rLWƅrJ��k1m�V��ί�AL,�Tǫ�6<aD�Bc��/��z7�b�5�,R�������C���q�����&�FD�%3�=z5N���%�LgXlxVHYEB     400      b04bo�k�����.F��֏�a,�#�� ���
�;]
�졽c����Ɨ��	�b ��2R�^�?Ȋ�R�pK��g.�E����/�h�̬��ۤR%G7/Ge�)��6��,�+p��T.�l � ����g(֔������F۲�i=�9BE羽"j��3����,7�XlxVHYEB     400      a0iM��.>Ge��P�2�| m����"^�D�����q�l%r�"���+�q�w�2G��9ɠ�SYXp�j�RZ����LA/5�U1���ޚ���&}�r��K��j#�;l����
Ky?	��D��v")�����#���O���4wc��XlxVHYEB     400      d0�_Z`��-nw�&V�`h�ǈ�(T��E������O�3i���T2gֿ�!�況IңTs\k���b���/V��5�	�]�AD���:�&�TH5; �e���1�aX�M�v��̈a�IVL*1��i"ߧ��LЉ�!����C���^��B٠/���GJ���5!��z�G�O�hФ^���2�H�}W� ]O��Hy�䒗=�Tt~XlxVHYEB     400     180ѢH���J�?�rkRq���G�`d��d$�՚�!DX��%lu�����A8>T��`p�Nhu9��Ť�6�yc�I-�G�A��3&�	��۹h���B���)�i�����)	�����S6�W̄�~j�8ͮ���=��$^��Ѭ��
��:��I�� �H)o��YX��:�{���/��s���6˷r[��3��|!$��U�g�2L�yyd��,N�I�TȼGi,2×Ä���u��Ê���!l�>^�Q���t~�� �T#��Θ�^d���F_��=�M��ym�=��§�6���x�����ޘ��_�XUwcBpy�����=�:��/X��$�&�3�zd���:���u�� X)�G�]����XlxVHYEB     400     130�A ��3fOs��W��74��/QZ�C[�	An�� �D����J���֭D���1T)VMG����#�Mi��Ͳ�S�/�hz�@;���f�y����*���m=�R&v�`�r�*�CB�a�������e�f���7t�(>smk�d��@d�n��D��
�g�VB��m���R�f�Պ��<�?u�떪L'a��O7X�Ӻ��f��m	"��ghhNM�Q�r/F�����8 3o��+�@��%�.�%b������A@]���\>B��i����
y�9�G4�D��C]�E��.mN����XlxVHYEB     400     110���ȗ�ǲ�������YI��>ؒA�j�֝ŀV��y�^n��u�\#+*ҩW �)�<�Sf�_��������{՛�a�cɎ>F�I�W��ԢX���f�s;�_]Ք#����ė:aga_F��T9U�;D��nDt�v^��{-f~��37%���1�u��@ʵ�W��^�XJ���ׯ����}C)���Jl� 2��=T%��5-5�����U�;H��:�d�����^: |�A̴����� w����@��Xmn�|��ԑFXlxVHYEB     400     190�m���=hI���ߞ�I����7�����)��G�\��邺��V���Y����|l�����_��;uϊ��çhl�CcVz�]=�S�I���M^��wŲĨ��e%ڣ��N,i�d~-�*v<� w�z+]��SYNǉE'B=x����	v��y��[���~rR"�$v������@0zp�8�� ��*�4A����\5qs],�W�	�
30d�+�k>�n���ё}�c��e@����HlC~��o~�-xY�j������"���U�����Hz�=_�\�aH0�X�ql/w��2�	EX��&��k�:j��EJ�f�9G���Я�	��#a���`}�E~�����?.�2���'��+~��8�<����	���אXlxVHYEB     400     110O\jz����T(��P&S��IK���K?>��ʹ ���N�cF#Թ&C�#�\�a�s�Y|�z3TUi�CrT��ǐ��%1���/��C̟C�`:���lE@���_O(�гZț��pV��3߅������r���=��v
t%�eF��u}r���X ��ݠ�T:l޹.��1�r=Ԋ
	�e6ټ�������i�;�<��R�6��Pr��O���[�U�5\��ۭ�$,\ �C�ϝ�R���b�u��F�I_uXlxVHYEB     400     110�� |�B2��������W��ؙi�2��!&�3��H�n��@s$/��ѩk.�5����2�
+eD|����4����������
����7�4A�}h��_Ô���Pa�2����=[谤~�.aG�1A�Z3��X
��{�<��&
�����x �oA&h��G�ra�I���O��2|is�h�vZ/���0[m��[Г4��VD��@�?�Z�s�����;�{\���o���o����6�J߬?6Gg~$��'���xeQ����XlxVHYEB     400     110#��ګ�^���8^����e��H�c �-_V����5��g�G�ޠSO7y�T�-�����y7� ޔ���>�y�/ӏ8k�$%2����p�)ϯ��Т5VRɥ�M�r�A���kJ��h�T]>���s�*˺E]��@��ËZ���15&�Nߌ�'���`�oflH{��Fkς(�j?�{�I>��-��_��������P�;w~��EBM���R�e �*Ӄ�q�e0�5��"\��}�����������ha�{	U�O�XlxVHYEB     400     100��MK���K�����!Q�����[�zH2��;�hm4T�J5��������x�`_�+r����An0���xZ>��&ly4v��glM_ۙ1��7�<����^s�%���@ڽrT��̣>�
P��+��,5����+�(��|�t]��>֣��=&��LՃ�Pd�n��/�M���-��ĺQl�)�[s�К����A���}�4��4�׊١��J����,~X����������RXlxVHYEB     400      d0����v��f��Ł���e�����"���Xt6ƳZ�.S�H���]�ӛ�" ��;����9hB+-3)��?Ї7R'Ib�Ҝ&@'b��Նq&�6�1'P��~`v\��N7�ʡ�OU3�=��V5f�]��Щ�8"q����?¦�l��T0ME�dP�:�p@l��q1�ŧ��Ҭf�ڠ�z�%	�Z++�Ċ���s��։XlxVHYEB     400      d0>����yR[yL���(e�6i�)���������v~9p�3���[b����������'��}N,Q����u��?�s^IHC�%�`p�ssLt4�A����^8���;��.�âD1b5�N��wo<�Mk0��w�����Y��f.p��
�iX�L���5�\�loغ�:& �θ��2i۷������XlxVHYEB     400      f0lķ�x��øL���yڊ����C�k�gUxGE�0��3�l�2+�9]����^L帬f:�ID�Oc��"����������þ^�S�A��
���.qi�SUF	�o#�A�=t�	�7�)��#S���c��̈��E>�m�;S.�\^�E!�]]TP�L��i�v��4��G�^���x+J�7�1x/3S�_��zN%�F����;6�B^@���9 ��*�$�/F;g�\y�XlxVHYEB     400     160bx��}�rcÀ�8J�<���
c�c�y��WCl�������aI�`��#��;�u@��b�	7���x4X���C��X`L�Rcc]yo-<��A��6,t�||C��q������w9�3����3\J�������@$��{(u�e����G�K�jY��;���������sF+c�C%H�tt;��)җ�5������휘�����D���M::Ę�F
��<C�Nr��V��+����Gǚ��]�v3c������^l��t��/4�M4�U=��)`!�8��W;C��$�n����ě�DN�/g�Q�hg�LB��aԦ�6��3�[4�Վ7B�b	�@XlxVHYEB     400     150����Q��,)�Se
Ï�ߑ83{�U� d�9�F�ba���0�bR'ύ�����+~����	'�EK:rPr+D�l
n@�o���N`j~�g��9mz��K�-��P]����eCyO��Mܪ���4���tôe��=(�/��Xї#+e�?�z�Cs|ټ#|�����`�r��^h�3Ӝ�[�l?hj�d�2�u�\���S&�ljv8A�#f�����(7 '��̥?�2]/�0N��~��o�;��EA�OR[�����9�u��X<����H�**��S"�X�L��]M�:���и�I��� ���M������`�E�[�ʯ?{��;!���XlxVHYEB     400     100߃��ɓ�8S�
*5	�S��ۋ�)Q0^�+����e����P�u�����:���2�W��[(��^�ٗ�𻿰��4-�D$I�w�?t$L%+z�3P_1X����O��?�c�z�I��wӬ�p^�x
�p��n2���)0�G������0����Le�2"Y�c'F�P+�Z޼Çm��E���_B|���>�R#pq����$�����|*<�I΢�h$ׇV���6�q����G�Q�k�XlxVHYEB     400     140�ֽq���O�s���s��Hu��s�p�հ�`3���7��|�`�s�@E�hWѣs0���D��\�͌�a�|�$X�����73�n�O"H;Ū�z�gpa0�m!S+�.-���Y�UvB&Bo�|�������/��[&eʄpƼ�Z�.4Ǉ�\׫�%��Rφ.W�����t��NHWHU2�&�b�2Ip��>\�C$&��*��7�&�#�+�ǵ-�_�C�Z�7+�!�!�.��ܬ�>`�8�F)��A���zz���QDG���Hc %��rH\"�{d�P[f, ۢ$C�$�V�5�/��XdP#���DXlxVHYEB     400     140��Y��򳉈�]>:�y���c�䇅j4 b�F�[=m�R�l�5>�Y_�"梬�%�X�MeFX�;q���䂍�#n�TZ����9��J���`����w�h{H��Ǒr+۩�Y�ʦ��o����JxZ�0'��O@�N�� ��PQ�����,K<��~��+�w\�L�.��ϡ�w���s|0÷chq8>���O!5NL�������F񚓰P팀V-�-+�$�'��&�P���3�����ԡm���rH�׉Gq1���0w$W_��|L]˜ICOf���K�@1� Ӎ���(N��)��)�XlxVHYEB     400     130��D�?�phrcw�vP�WFP!���&��*y�#��Ք��Մ��J�O�vr�/��{s��u=���:D�qc����]�G�Vpmx+BcF65���6�,2<m���ʔ�� �P}t�9c��)�9�(f����6�A!�>��a�?x+F��B�&e}�X�(I��r��gȈv���~��s��WC��hh����C����]��"�چ�E��`Ѭ{�� d[�l>AO�s�.G��b�;m��ڏN�="_AF�׼̷�Q/V"z�u�f�����ZƔ���BF��cE�[���RE��&���a�XlxVHYEB     400     120���m�P�KPSv��u#��q�7;���@  ��
�8���v�Y�^cD+*�_�D_�� %)O��~%7�M)���X���W�%j��Y��&e�;��v���Z#�N�:O(ٝΦ6:�u;3��ø޽�'�UL%p%�i	he�]�BD�+���e\�d-��>LW��:���G��ϸ%B��yW�~Nb�W�%���5�"'�OB��ƙ�r���C��2k�������ٮ$l�|����K����0B�u�nIA-�x�W'�B��N0^�:,XlxVHYEB     400      c0<��\]����$;�R��$>�$�1�Np�P��(޵�
�a��,s�-�ke2M�s���-�*�o���Aug*t�1�`�"��cG�1���4�����p|8�\Ҋ@�$uS>�$Z��:uH��,������*%u��9o'$�&1&�-b
\2P�Z�ٷY Ď"���J(��C�XϏ�~�{q�XlxVHYEB     400     120ye��Ж�$�\�E���Qغ唶��IKZM�9H�_܌��M�@g�����^��ZM�@lc�>⧅�D��ODU�S�Tc"eEa�m����$>�d-��b�*�-�5+�ז��g�8���m��$M;x�/��T�G�'q�ɷ�
��~@�'�@�j�����Fj*��W-���R��2�NP�@�І?xJ�f�R:�<�mli\���ak�kLc�Ҁ1���>����Z�w���9�GP/�m�j�ל� iG����B����=����xh&� �b��>��XlxVHYEB     400     120��Y<j?�����Z�h�:���B�.���>�wB�5Mﯪ�nG�:�
�*�__�,o� !�[R�<*sZ�*a�<z��5��&�UL������R�����e�%��Z��i���Ӟ�,��@R�z𛾒!t(��R]�P�����{(��c4��L�w:o���i���zj[���99x�r��u?��#M?'�r hkCfF�K�Cr��8���vg�Ey%���a��9�#R0�ϙ���g��Y�0纩���#3L35���c&���֨�׊,�BN��>eXlxVHYEB     400      c0��"��-��U�[�B__�7��b*&��*��ے/�Q���2��
_�1kۤ���� ����c�iP�[6���]���u㎙{/}~�g�F�O�X�Bo59�C����}%a�tڊ�u�-��Z�>��AVpy�(Z�i)/q$'P��gw�`�n��,��̎+��F͗�3'b&��Ӽ�NK����/A����߆�_XlxVHYEB     400     120��,W}i���ƿ�g`��o���C[M"��[R�%�LV\i�o�>,�ذ8�(a6g�zg�ߴѩ�S��J$�D�#"naf��72�]����D3�;����	:b�+� 5�1,*�K��A��D&E�_y�gؽ߲��Wj6qH���Kh�΄�!H���#CZ��f(!h����2r��v�Z�¨�^�\5�$ @ �����Ma���R'��'���L��ZGd�����m���@�Bm����		�	�'^�57�$����]�֎uu}�!�k)���(߀��XlxVHYEB     400      f0���=.ۜ�[�� �!�T_ 2P�DD�xl)����b
%�L��҄~g����󷮢M"|~�q��?�!��_is�M��Y�^/?S�%bw������p5!.�)�X�"d{�ݩ7�� �� �am�mM*H3iP{�����*� ��`E�+�T޷W�,�y��QR��*�I�/�3v"�Gm^*WrTd�����l�.'z��r���[E��Oq=�1XK�XXlxVHYEB     400     110.�\��DNqup���{яNp�i��#�:��M��&�trW=&b��{�y۸�Kr�����������veoZ�e숢�7d4�g��H�ZӞX+>�ؙ�;�����:�0�?@Bn�{�#�(?�_9���������� =�����Xƴ�����;��X�:��2eiqR�Z��D&�JgR݃��6m�2����$F�:�A�GmB��3��:H��5p73���|#�=�g諢�Q��fa���%� �T�A��O�`�J�XlxVHYEB     400     120�Y���7��0�w�t�� "�w�Yz�XF4^� ��&��Py_0��L=��ϱ�
�b�����&�r����FH����z�R[ߥ�>�|z���
x4[@3��N�jŹ�f�6�_1��T��ei?������`���0�*������=�e��CB.�+j�K֓g�}����2�L�jh�t�~�I�H���ZB<ZcH��3���A��(�V#�nȰ%P=S�R:B���1ޒ:�۬w�4�7rGN�j�%��^��]ēMAC��U���w�M.B�!h1y�XlxVHYEB     400     120^�{xJt9O!��s6��!6��?�^%��`mW?������[a�m,�!��Е����gb(�q����2����� �n��g��Y�i�+X(bV���ˮ4��M�K�s�Y2H�hޢ9�����K�Z���١�p���8�؟Q*�
��zE�ĝtYp���dHt���"��\��9��c��*�	$i\V�&���tʓ��ol����|�n�	
\~r��UX�:�o����������~ �E۠��UH�vm�=Cb0F��{y�y����/\
e�c5^a^׆�XlxVHYEB     400      f0���s�O����}#޻�<�k�Ȱ$ݠ����������@W[���!ca�\^�>i�3 ����!��?�#����(�d��?�
^O��1M?��$��[G��8���W����#}�p!N�t���L��Ր��5m����<j_�E,:p6$�J�m�A�\�h�p�����H��gݎ2�,U1İ��@p�Sn�J��1�saV��P���jJd*��-|�v�{D*�^i��u�NXlxVHYEB     400     130�x@#+AM/\ufo����x��"���pa�K�hR� ���}������yy-5��y�»J��,���y��
�U�!vk0Lv�R�����1H��3t9B�F`J9�9�KH��������7���z�M"55H��@��o�ٹ�|涘S:RSb�@*1�TCi�m>��?��'0�"��d�2ކ�*������oT�6�":�P4�7s� �mҥnp��:V�c<��)�iF�MZ�ƂEq͚�hIX=gI {��@�<J6�B�F�D�R��+��^��z8B��d�XlxVHYEB     400      f0��z+��J�YL!c��&���KZ�?����o��$U�����Y��!)���@k�u`>�;)�Z��ө&(v�I';�h4��Cy(K��6wW��3�7�������:�H��:�9#n���.�6����G����.�Uh׊���=�qM�G`:'	6�7^!�H��e�0'���̿��wQ�]�&�[��p�b~vĞo�;�CYwa��|�Q�V��ů��9�G��@bf;(��XlxVHYEB     400     150$"�\��.:U��;`� �,	A?�~YfG���/���V=?HSz�I�=Z�( j��X�X���;`��^�������.	��^�?�7c���7��ߙ�*.�t# ���p(@ Mi�n�EnC��N�(9�|<�yJ*�L��?I*R�x��8������u���n��;i�Z�~�i��y����i�^�c�Y�(�c��Q���\���2���b\V�-� �Q�f���e}A��;��;t[%��z�`Zm�J<�ac^���[���U��'4�йd��qD��iurܨ'8X1��R�ʰ�w��t�|KN$R��<[�wg���A���O��4V�PS�Z��L7XlxVHYEB     400      c0�+�V�R+6���h������F,ղ.���u7PJ�vۯu�MB����u�`kKLM�UF��j���o߭oS�^s�?`�>\���JJ�`b��tCB�Bt-ʊ�t4p_�U��N��=׀	]�`�}���0�w�
+�Gzs.�C����a �G�[2��kVM��X���?Hs������)�O���zW�&�GXlxVHYEB     400     150 s��;����^�0Z�	�U}�Hta=����	S����(�aR���oSN�ݸ�O���O�c��xN�0�
$T��a��C���:�!
/�ݞ��q�f��;��;� �RN��P^�k��L��^I�Ӿġ
v�aoV�X3H��O�������yb��XOL��0���@Mb��L!����?[�y_ʏX{�c���i6d�>�a�ĸ��}8�)�M*)8)S{A��m�az����)'6��E�+A}���P �0xZg� ��]��(���U�jz�;�+�o�y�ؑ�d�E��ߟ�?d�A�y�?�	��Ig��bA���/���OC:�XlxVHYEB     400     140,J�S�'|@Y�1rPk< �]#N��FR��{J�i>z��gƛo�8��ޚ��(�z��zfx[���Z��fEq�K���ɯ3q"dl/���4lܵB4B�m�}�#�D�z��8�Ç���)v
��`^7�/��hP���:�+{�7���(bz��G.ze���aL�eӯ�;����`]��'�l�}e�ͻ���R�}a�`l�6ʚC�}\�^;~]�V��i���	���zf�k7�?6�g�r��V-}j� �܎��zRxeF!� O;'	I���(;�R��/�����V�/�OŖC�x=�g��%�x/��nXlxVHYEB     400     100z�iC- ���6���̦<���ڵ�P�,F(����	�m]Y�;�.�gQ٣������}�
��b�٧Ƽ��T*�o�Z9��>�3>�.hE惊�&�C����a?�Ř���)��\7װ�]�:� @����#����~h�t�/|�A��
N����޾��'(�gB���A�0t>徽>x#�[��gtN�iw��wt6��8��L��o^拡���2���M�Z�v�N]�����.Ą�n�XlxVHYEB     400      c0��KF��n�. O+i��!FG��	r�8��1J�h�NTX��	��Z�T�KO�F��j�طPGD�@86��?�[ڹp@�{��U:�
,�9j��$.t�2�����p�����*��l��e��2)��e�����-�Hjx�~2�����2�H3 ߯�����FF�xi���rҦŸd��z��]XlxVHYEB     400     100��1�c޾�+\�A�J^�jK��xi�;���?�s5�w	&Kܶ����Te��뤭/w��7��zA�3��W��q�eZ��9/[����= �
���=y���=�Z��)��l�8>������+�8�Π|Z1�˞5<��g�>}�eZTJ�!nqܹ���r]���v��ʛ�r��ae�3���H�����mX���D2���l�uIL�#�gy���^	2�=��o��#^�B��u
��}G�fXlxVHYEB     400     110�2�q(`u�滑>�����&˓�&L���sdD��Y�����J|C+g����l"��q��5 3@����ILV��ii�{xS����d���9��b��N���1�<��wg�c���C���FQ��i`6���Mi�&��W�������%�+�l̴�>�!���ZS�� ����p��t��6�6�%@AmV$�0�?��|����
%����s}�N�6�FA$��d�~�$'%0����Vڽ��1�JF����(Ƶ����XlxVHYEB     400      a0cSk��2�N��r��HE�L�Wnm(�R;3�b�{mڕ	�C�Ytqΰ�v{�.W����I?I��q|Aqb�!�P�[|��>"�mh�l�)��ڽ�D�eܽ�c�}x��þ�s�I����C��Dv�^�90�!��R��������I���Ȳ;XlxVHYEB     400      e0'�O���)B?���� Ml������#�!�=�'D����;���Cgh"@(=���r˧�cy��If6 �+c�}&u�)c����W�I4`d�쑊���-��g���H.�8[�ǎ�h�^�\ǺTu�T-�"�a( �?*W���W}9��B��]���_m���tj^����W���m7����-\�a��0�S`75��f�ZE�4���o�XlxVHYEB     400     1a0����u��v��_���� � �"���Iv�F�cs|�e0`N��D�,�k�9��y	^^Ќ�r3��%��� �V�#8�2�j�^<<0�`]�p�� 3?2瀩��6#{zЯgF���J5��&8R������������MƶFl��f���������^P�6�Y���}���߀m���&�NMĀ��Sڌ��!���r4
K���Х.�r�+��o�#v[}CX��q��y����y�`X����T�]��� ~V�<'�=�)��Ǽ@Cmk%D�GYn�ޚ>#��U$�Yk��`�X��9���rk��p�hc��9:i V�a����V)�#HSh��6ϵ��Xk��b��Z���7�Xahd�>P3J�)=!�g�Xra�7#5<K����6ԟ�t���\XlxVHYEB     400     150��?K�TT ���Lb��tm�"`c���6�^gGm��O�#���k%��S��'�o��a�:;�d��.�Ϛ�j�}��H��D�Y�R&��������$R]Q�.d�T�8y�lz�H̀�D�,0��[LB1��a��]#ߢ}\�e������-˄�T��B��Z5+��';hm��~�����T����>P�N��l���$٦�;��H��}���<�sg�dp7l��a�Mp�/�f���vh���v���.��P�L=*n�qM����g�#�ǡ���I�v�oI
�E�����~��A�����gUmmS>��l�v=�0��XlxVHYEB     400     120���v�ֺp�4]���Xkr�-��,1 "�'�]��s�U+�����?5�������7D"bE�y�=/���	g��D#����.�b��ۂ䛡��t�?`���G��.9��Ri��蝍6璉�
IM�+��Z��2ft~�Q�F�s2�chN����6�Qz�Ͽ^ �,��N��-WG���{�2�0�Y9������U�if���)a1�L%ҞA2.���+����������$�CpY1�f}EN|�Ӧ��U�yv�����E�"��J^@XlxVHYEB     400     1d0�W��c�	�Ħ�>�X�{o�h��0�_�	�����USH ��]��	D�AZ���x=�2��B�t2�ᵢ[m��I�#hY�dM`R�EȘ����<1�������Q0Y�ɞs����qj���O��t\�p��UW ���pX�~����x<� UjZ#W1Z�@IX������� �E?��%�%����Rs�#P����Ӆ/E���p�B���H� 4MeR������;��6��[�����H�N�O��@\@���L�ب`�q-��5��]������o���uT��xcq��\�v�Ĥˉ�l��˫n;a�!hٛǝz��
�s8T��en�����2ؔ��G1�ȋNP�˄���yH=g���^/ǜV��iY�u�L� c'|�),��͒�X-�EP`�ݴ\�PtP�rgM��w~Y#a�n�J#��aH���������6XlxVHYEB     400     120��&�c.W����r�CAY�S֑R��筯*F����gyJx��0n��T
���Dcy�~��8\$��c���̭�I��0��4��l�Iz��D��3�Uj�҇Ӵ�-�t�e��	��,����h�u��%��V	�ĕ��H��<�hBj�*�7m�wbS5B#�m�$-�U�5ڏ{��4��OgO면�����S�Xމg�)=}��^���z)�f�N�CK�M�W�Ν�}���<4��1+���q�TW��7�6XA�1s�ٙ$��}�Da�%�d�_Ώ�V(�XlxVHYEB     400     100u��s<� q���f�)� ��gdc����J�b����-���z!`l	�@�:#��k>�0���YB��.4� ��p��<�_]��˭p�Qz��P]S~}X[�y����5�i.=�UIU
�������_"z��L�����Ĝ�X��>#t��������=�T�N/�y�X@�/���Ř��F�=frp��aq�'?!Z2K�v�1w���G~C4#L��v(��HlBߤnh+�K7j��\9���m�XlxVHYEB     400     110� ]���� R�ӏk�<9vۤ6�#2R��"&	s�u�4�{��?y�[^����g@��Oiщ�60̀��,��N:�
��X6c���.�Y_v�d�7w�BlvrU��x�Vm��|f�-�o6�c�i�o����+�>F��`A�uh!mU�v�l�O�\�����u'x {F���çf�m%Ĩۢ�2�@�!���}C��*�C������T-�x5H�?���}��"I�h��Ն\@D72/Y���Bz[ D��o+tYP��a�����XlxVHYEB     400      d0d$sԩ��*C� �_@C)��B�����4������jxAon0M�c#B��o:	�Y �"j2,�m�|c���Y��>v?Ѹ[
�;��^ߖ%���Ѕm������H¡�F�u	,@��R�x�y�B��t�*,��ȝ�%�s2���{��֡�	x̔o�|�b�(Jup'o��/��&������3��5�6�%o�@XlxVHYEB     400     100Lq�@�`���vpG���R�	��%aD=���jd1'-����<"��+����M�!�I�KI�ssʭ���������#'^�u,��s/<�b@b��o`A]�Ź�&��)��UqE&s��E�ʬj.A���}�E!��D���d��5�)���DE#�)��#?�4u����1?�Q�@Z1h`���^=��NZ@%�fq
I�b.:�}���f�|�lOC{���ȉ��m T��cߺSgU?G4�Z��A�@AkXlxVHYEB     400     130��̾Y��׉�ƙh&.D_�C�[rU5�MZ��c�<���-�N 5���3T�CM����8���*C��ԧ�D�kMH�������4!'4�q�*,�*�
���5�����E��8��
�ş��l:�+�i����
�f�AV��|�ˉ+�ɠfM��Y'�����h	A��g>��M�����b�	=-�!W�-��/כ�!r4 *jڻsQ�Ǿ���1%��t��*�J3�FRJ[\#�d�ֈ4����{՛�n�^�_RO?�U!��cNò���<���i���ݬ��cUy<3��XlxVHYEB     400     120ߵ��M��[�<=wr�����|��D��'�y8wy6w�%�y�9��{k�E�ȕ9�ֿE�Q�|��CG�t_K�򷺼�w�t�ۋ_���%1O[|灑@�nu�.�q��~�+� ��w&hB>���F8��
'ߦx���p4�]8w�v���hugp9R� }4��/'{,���|�Yی�=�c\A�ѧC��_T1��	�������`��ʲk���݋�U��۽
Ľm�>@�z��Eٯ �ؿ
��q��¯L���Á����uߕ�
"�]����z$>F�mXlxVHYEB     400     150ʮ��0&B�C���To�Q��j!-1��]W�j�f�f�,wH��]�q]P������CֺX�
��Ez�a����ۻ��m�g[�}[	7x�e�Q�߱א�
u?Sc�b���e�4Q����:��(���<��N"Fێ^�T�t� V>��]î��$G������*���\�yo���ˆ�1�ڸ
�AP,����#Ӫ��t��X��]
�S9�(+5� �Xg���|���ߏ�����yS��Z	Rpd�n5�wI�q}Ɇ�����	�'��לU����1���å���E�Ln�I$��n>�kR�[�0N�`n�з��ڨQ�����؛�8IXlxVHYEB     400     110��R�4^4�I����F���w�|,��`���ֽ�jY�S�jU>,}l����R*y����K�J��U�4�H՛X� ����,�) G�E���{�'�;� ��!l~]�T��3l��v0ٔ��p�fX ���rh��J	 �I�r�>ϕ}��1zX|����3�[�7����r u��Z;��\	��"e!��16
�E�%��(�]sPEI�e嵪�n�uـ|r d�
�S��g�	�3`B�k,��p������)��'�N���]/XlxVHYEB     400     110�L�?TAU��L 7Ӂ_�	^�s�����zx=͂T��J�6Qh�&��I�L�z�6E�mT�luH~.F��=�Ԝm����7�4��`�
[��'#���kI_��yn�B�I�}�ż:;��_���%�7�v��޻�ˌ�x�5��no�tү�¡��r'^���~�!����~P���(������}�UN���UP!�ǠV�sK�*W��)�qi_�'���i���V���uHMT+=f��]D��P��\����C@�7�ӯ0�%���̑XlxVHYEB     400     120���}����\�tG��"���-T�6�TX6$b��@�'4�Ɠؐ�QC�`.r��c�зM44>��E}h��������v��RT`�91589�څ�n������&Ɛ*�mUnlMz�Hy��Q�j�(�t����P���ID)�pL��7��7X����h����yw��[��$h44�"���!á�B �j���8��7��}���x�������F�*8��z]�w®M�v��M+FE�]�|):DD�_m�>�+�3�CZ�u�����r(���ҧ*FXlxVHYEB     400     100�&���H�	v��dO�E���4�[��������Ѷ�Z�{�k9K�u(���d\zh�!�$y�2�R��Z��y6���C�Q	��9Eh�&���n�$"Tt�X$0��=:+k�9�jb=)�d�)Nm!����k��YO�}��[�>���&uNU:|Hi����6�Is�['�̢��2���ㅠ3�+�^�Au韊�g$ǳ�;-7�:�wK*3��������E"�q���}/���1�U�XlxVHYEB     400      f0X��8�Y�w�1�64�Q�U[N���&�����H�d����!�50)!-*olJI<��P�d�լ��2��6c��3C�z��
Η�%q0N�,�a�GV�KE�Z\���Rd��jP5ס�J���\츦m�h	Te���`����Kα%�iXx]6�O ��=�M��%�{�$�!���n]׏�m�W��M�#3���k�5ľ,=��ûW�J��:��p�Xpq<��#0XlxVHYEB     400     120#	�m]e8흏n�z@�� &Cޢ+<�<'U)��вZ�Y/?���8��
3��2<r>�7�e�����9��	�Tea&�φ5���_=;@�Em��Fօ����H���9�ʨ;�_�������\O�u�u�pD�!m
-ס�{�j@fF�#��V(�/�X́Q!� 7\�B�
�o]ؿ�K%{�'m{�S�cҚ�"X�)�,<���[�u{c~Q�cn	~����^����û	SQ������Xt�ئnf[�pݫ��	U�P�
�~B��\^�XlxVHYEB     400     110�����3"5#��_��f 9���#
*g:hh`q^ڦ��D�f�a���z~�5t��/[��I�i�G�5��*��T������.2԰l��p�U���lP��9n�����:�*2���)�l"@�Em�9�re�1w�NJ2v�0��6�Uw�QQC�æ}wbn��A0��`�`E�z"�ps�-�5���n��L�����2�ɁgW���__��T�9��|���c0v������ F�m����n7.fT#<�: Z�"S�Q��XlxVHYEB     400     120ܰ�z�
Z�f��
�7Pc���Uk�HL1�xp�
�g�Z���wr�	���V��l���x����`���E����P3�@�iPsS3aA�@�����)D{p׌H��E=k�"���S�&�U��K�g��v�zS�7��S�E~��A{(�irw�E��8H[�i�H�-z��@���DG�'�Ac�xw��n6r��i�}EK ��ӥ�A�P[s
��t��_���xT3��담S��Ь����)����i��.�6��Ѵ�t��֙'MiX]��4�ʋ�pBZ��pXlxVHYEB     400     140$�$)CH�Vpޫ��t���ө����^�Ù�	�u;8p��������Y���fei�F�j e����)��^�^��:aJ���d2��r���(�<����Sk!����c�dn���Y<Nm���ny�*��i������{?�sk1�c�\*�9֏�]����!԰a=�a8��<�{j��Či�iO4�u������ ����;�`Qb_�mڟ�Ln�lO��0ɱ�L��M�$�7�i�*3U�.��(@����`��\l+e��1�;9�V"=I^�v"Ν��zv�� �\��-��s�U����u
���Y�@^XlxVHYEB     400     140b��/^rV�"���~/���z���=5a���`&!�ƘS�Ҝ X\��F� �+u��Ę���F66�<���Z������T�ېE0��X��2�������:�����[H{��ʨ��q�t3S��*�0BX�.[��A�����8lfq䎞`Р��2ј8�\�t��l0��`��i�ES�l��J_N�g�wj���:���5i��t&tC9�)��˃��b��_b�5����,Hт���I��Hav9L�1!��;�����TjC�����<�B�~�2[�Dش�;6�oR�dZo&�4������9��������?XlxVHYEB     400      e0q�A��?�ͤW<s(��`!M<�^|�2��T�
��&�a=%y�̄�yk�dx`M6�.�M酞V��S�]��!
��Q�����\3j�(Z!���u}�R�-~1��H=o(V�*�1�/��$|��@eV������Qt�4����^�S��}R�9�/ ؟�N\��>� �������+m�l���n���9���:���Ȣ�]rڒ1���j^�A�`�XlxVHYEB     400     140����v ���%���mo��.I�>07�r���z��M�^�x��9U|���=�go��g(���]��K��Z�w8В�V���g��p�6�ySC^	�Ƕ��2��t6���vثX�7��us�}�������ߥ������Q��=���lB��6K�[�����i�T�6j��n|b�� �?RD�Ѫ�w,��� � ��(�رi�]I3��ߞ�`qsh�*��W��QɌ��s��8�R�\D]'�Ϲr╞�Kk�s~"���}d�x�UTv�Z�]I���oD�����"�-}���y8���`�I�nj�XlxVHYEB     400      e0��>8ְ�eQ�F2�|ܬtlY�����j�]ͧ����b�9���Fx���D)����?��Q��L�Wg��8Q-U���{�Q�/O���E[8���,?qH7��k��?5�)�<z1�
�	�A��:̰fS�fU
�x�}�4`�J>z5,�p��R�6Wt6t"�ڥHT�@���Z��ʐ�����d�����9kr�� �5E�����5؂nǱ#��x�����XlxVHYEB     400     190�Ci�1vXe���8Cf2�Sg<�� [�8�ܨ�Oh��#/h��Ջ�
�)T�9�̀�ya{�7+�s0��
���L�[k���7ؐ/G�a�1z�]����X����~����mŮƿ2-װ��������T~� =@	�Ք�C��MkT_��E
��q�d	��+�'��魓v6��{x��~��=z�r~�/��]l�Ǘ�ML�sD��e���2>>`v��J"��"}(N伎��;etw���Q�7�� U�Ix�}��)�/���3ף��1�T����O����f��bvME��>����D���h/j%�����rp�9�����'$�?����?&�Y�=<��[��P�W��HU�I�PJd���dj�G\ ���������`�د��R�A��XlxVHYEB     400      f0��JpVQ�务;mp��<3@����y��a&䥷~��_��[ԃ�m��fF�[�>�)��8Ad�'{P�}���{��\1���2�i�@�X�q����,�KZ��h�7��;�C84b*�5����l�±V��+����v6r��l����������'�}��$���7�\�Q���Ȭ@��H�Y�@#��@MTRs�3(��K�K�v&L,�8|�u��T�2�?rl-�XlxVHYEB     400     120o������������ ��E=�;��<mr���CE^a H�')Gv@�߳��ٳ��_+w˯g���l�����&���f�<���*�7�΂���+��p�������	-�S����[���fy0;�CCb�~��Z��z�����Bc�ςc�@�Bw�J�@��hNXn�q��J5{c�*8���ʇ�c>�Q��C�s�4?t��6�2�	�%$����Z�H��t�h8�)
�_��������M�����_���������H��k+Է>v� �[{r�{D1���XlxVHYEB     400      d0�>g�.v
UV����l�q���z���s� �`G��!+�m�Tç�.4��̰�E.<�R�+��b>K֭��AR����2f_j4����e�O� +s\�״�����	�B<RIP���5��G��P��ci�.J��+L�� �f���ܼ����O��{_��1���s���r����^�<�o۳��_���V��ˈ�XlxVHYEB     400     1504�Gj��e��D굊5C��Rv���GIy��+�'�EV䭑Y��uy.;n`� L{��F5Y"_Qe�����R����A*�NB}&�bp:��>[��`|eIT��̵�Q�^dH/��I�(7%�|�Κ�������z�4������s�5n�EƁ���w*/PAv������ܤ�{T-�(���nN�y� d�������U	�O߂>���;o��[K�0�l�:�랢����s����|�^]Ð�ש}��#���v"�9�w�Q3�@����4�:��ר�@I�7!�g�/&�1�6%>yp6ҡC~��R^laXlxVHYEB     400     180�ԫ�@�ż�����;s�G/�����\�k�iJ����Vt��yzͮN�lz��N��������ܱ����Mj�����E8Of|�����Wvd?� 70j ��^�ly^,����I�6f��x��\�<���_������iv�K�Q�ؒ)�|;n�9�^�~�&�m@$�31fi~=8��繿bdh���05%Lzܖ�f��  ��j~��/�@x^����S�-k�*-���N>hܮ=fw�$#�h�M
P�Ea ���k�=�X�ƱQ �`fAA�I�5����Y �k���I�1f;}ڒ}��Y7p��Ѵ�v%7�N>H�Y`O�O�m������#9}�}|����hڮ�$��P(�E�t.,^��c��M�����XlxVHYEB     400     120�=e_>����-m����f�ݍP��Xr���Zf]�x|X|"
��f!����i~
BAEmix"R�,yv��D6�bW�����teo�(�b�G��de'#�?���ի��t�ȗ3,�Ȓ���`��tp��$#i@�,��������r.m�ȣ��E�V���a�G�x�u*W���f*g�@�D8���N��D�i?㾏���1~���Iz*�ߋ�:YF���1 ��>O'�EX�*����%C�i�zy֢�z�&��!ko�J��m��.>�g�J-XlxVHYEB     400     180M�(휶g�=�#�J�\IY�� ���beO�A�4�k9��r��Jޝ�X�2�He�L=��]"܋�<�<\�24)�2�C0U��8����QB@��[�E�
��ZZ� F=!����i>[��lhBI��roG��G�_3d��s���;C���ٞ)��-ld8�<:W�3�3
䡁\�d�QQ�*�s��r�W�eK�a#�,X��N��^���$���������:>ϬVٓ
2�s|z�W�!�-��9b �<y�r防��,@e�i�6�)t��^�r�4�څ�DJ�N�?��5G�GȂ�X	D��~d+Ek6� Y ���ޣ8n&b��a|�K��zEę��I2�jVS��w��z�D�sT5�4'��x��8!�(���XlxVHYEB     400     120��m�Gҁ�T�{�=I�J���z���q��h,�� �����Eg��e�Ó��.�Ŭ�7�iA����z�������bF�-աȟ�h�UdgӶ?�(\��En	#*@�e�Y^(�>���h1rL�rX����3J�}r������'�:3��:g�$�ۇ��`�?��Z���|Ѫ���&�O{n���}8�z�x/G�,���C��X�������E���#�w�#��Oԥ�#~�^��'��d��h����[[lrk$�zU �?�&�Ė\!T�XlxVHYEB     400      f0�8�$9ߵ�P���AL�]�I���&�F�0����`LFg�J�1����	P�C�H����̄`<�AX|�]��`��K��
j��.6d78��'�
��~���!=�F���WIB��M>�LJ%N�Y}=�!��J��>:���G�{zk�8�M�1��f��4�Xm~�:��6�9�� e/�����ۭj�O�>\
:#NK��}�NVr2���\3)J|o� �CZ�NUXlxVHYEB     400     130z@�&�2y!��r�E����<��8{�̽��ؿ������N�5�:��Xܞ�<֐�E%"�H���p<)<c�(77m��=K��QA��g�#�I�x�����|?��)3�Yټ�YԎ8ώ�X$�2/#�dn�ׁ	M ��\i��侊�zd�,E��g�P�nu����,�ߟ�Z&婼V��*�l)Q����
�*�@��/齏�N����_����y��%�,��-*�{��ye��H1�m;� �K JvEX�:�9�?�i;kI��x�<H��֑���c<;f�ʵQr��lXlxVHYEB     400     140�aU)˔��\4}'�c�Jt�����{K{%��^z�5�ȢB���X���ݘ� ,P:��HB���ؤ��ǃ��6��A���ˍ��'�z�{8��د< #3����9[03�9Jqq�ܓ���%��v�$�BF�G�9��L�D$<��?ȳ��[D|�g���@E�M�$o�W���}�o!@��h��m�7���v�j����y�)�z3�c���M���W)� ��LB�*�@Ԧ���N��z�@z���S���(:ͻg��&� �9�GP<�ea���Ѽ��t�x2�`6��3��Qz�zSd�P��"XlxVHYEB     400     140���E���\��<q.����[��)#�u/t�׬���>2�e���L�^�í�kS��j���q���e�����7�ㅧJ؈Y�ݨ�S��!�`��vc+�፠mpU���^�}8�F�$��p����}X д1;F��%�M�3�
5tf�{�Zh`dzm�ޅ�&~��_ف�N0�5J��(���=d�Q���	����cSw�]=�n��׻�ꉆoAc�E�ܐ���]I�s���ŇF������=liYdi>���{uB��0\Ȍ������/�>j����a�J�	��fT�E�v��U,��7-q+��p�<XlxVHYEB     400      f0��v�Q���`�w��Tf���y�0�T�J#ற���W��Z/vGGh�׽-����d�]�%��`�� C�\`|R�a��>�5��Tv&�t�S���#����2����̅Q�b,mޘ�y�����E欉� �#�I&R?���Ņ�A$}��R��P#��E	��uzc� `>��l��m.ŝV��V�?Z�i�'��29)Z��-��sIj���pOH�j�9,�n/@���.���fbwXlxVHYEB     400     1401��m���%��{�0p,9�Iae
2�dڎ�e�|�T��
��ץ��ݖM��@H"z�!��<~=�N��%�5(�HH3~��`�&	�:���M�o8���@�����/���>[��Go�Np� b�]S7��b�v�AK�k�nn���!\��X�ȡ�4!,P�Hc�c��M�t�h�^n}yl���P�U���m�7�Q�~�S��7B��}{�<c8ϭ�,�A[��t���[>>J��
�Y��`h���\:�����;�;$�yWт�$���lෝ�8k�${k�I�k���d�`��u�9ψ�}��XlxVHYEB     400     120jf�4�c�3�4@Vk�e�E�������.qD��a��v1�DW��Ōs��y��I�7�z�쏸�����e.��*y��v#�DmK�m0:[�����cglU5�q���a�ƹ�F�Y�Ͷ�6�̈́=Ɇ����@�B�F�{���\t� �
$�5W׵���Z�qg���\�ǔ����>�|�_�$���C'�s(�!�^�Z ��FQ4�*eS���e���a0Iz��*1N��3Z3X��L���~���zs��b����\�}�/UK�1F���_������'�ZXlxVHYEB     400     120�Cl9q��n���*�_
oZQ� �/��p�^�a��KJ�s��:�wV3��ZQ�!�#�De��/���4�S*α��=�CPY;q�Hwρ��T�ByT��/,����&W��U�Y�����=�L�4�������ԭsH�Ne�$iRo	M���%�g"]�hA��C���26�p�#�G]�i7�c�$-�doo�q��ח��>��|e�Ҁ"�JC�A��WD��[g�V���|��V����ݠ��&��e:�=�������ˬ��-��2B��o%�_���XlxVHYEB     400     110lYL�c�"�[�C5����"�a�?^�[��}�U&�/�������U�Zq��]Lb����ћ�]T,��W!3���Gu[]��ϻ�]'��ޥ�|���^�'���N�&S�ǒ\7*�->=�@��Z�|��qr���at��	����R�S�c#���j��[-f�iϲ�>�c��2���Jo�	U��J1]tA�C$Hޛ��1]��	A|�������)�~w+��Gh��I��qI��u�<4�U7����n}�Ϯ~È��`W�t��XlxVHYEB     400     160Qk���=Ox��¹��J㠰����#H�z���#��E�����FC����^��~�$)W�P�D���ߕ�S��Q7��O������g�o ���2�R��%��(��󩭂ɭ��R���}_��e�jH�a���W��Ce�6?��LW�C���|axb��d��1�+[��}�\��Pܔ����B��ȡH1����.	b@�P��=[7bb���N��Κ�LL���;���3<���L�GR�|x�^-!x��{��89�wf�@^^V#<X��p��,"`�9��0��e�w�Q�,��Pa:�72񪗒wiBr�o�R՜�Ō�K&Rw�XlxVHYEB     400     130�SB��U�ޔ�k>ly߬J���Z+��?�Y�����(Xb�X{��n�7hzdb-M
�'��3ާ<� (���PR,$?��� ���O�f��oQ��	.�����n)�\�r�%�5���Ýi��(`I�F�v�� ��2��1?��zN 4�FA'᪄Ki���v-5����aOl#6�@�FH��௶&��H�-��]Ek7k�p�B�U��ru�l��K��P}_�	N����z�8��-��,��iT2d)�0���|j��F��\��-Ov5u�8�?�z*�W��U���XlxVHYEB     400      c0��� ��}��k���xi<�7= .#�=_�f�^��®*]τ�"�/vt����Gn��	���.񂲇��@�|j����_�)��J�_D��~z�9���'g�i�c�)�w^��ؒ�[�ݪ�υ\w�-��"y5��)`W~Q�M�?m��&�����= ��Z#"<�'�<;�V�z$G1RA�����XlxVHYEB     400     140M-��ٹ�h��j�Mak] ;��U}���ʩ#�f��H�$�u�����_s��:r ��+fp����W�e�?|KJh^�:���N6i��x1p�#$���v��BT�8��=���g�GCY�c!p"=J�F�sk<��iV��Uf#ħ�������*wM��2�ǣHv˺�x\cp�q�g�k6�E���	� ��t������/�Lr�����b����h��Gv��9|OF�Y;2���&�"^�rA���~.��[��)"�:	�7���dH6j9d�5EwWגFo/Y4���F�<Y��`�V�=ů3���zXlxVHYEB     338     100���R�Oם5^�:�ϮiS�ئ��$�}ﰷ:	��&�w���8��-^��Ԉ��a���^�Q�:&��e�n��q�|$.敫�D��{|�O�-a3�;D��=�uP�"��0���R?��aѣ�����_��LT�}����.Κ̼����E�3��n�2s�b��}��~"�w6O�L�|w3UN]*Y��{�7��&b��t�S|NN���F1��r^/A�<� O�C�j��l|�����Y��uޢT�kv