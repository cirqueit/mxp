`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qLWc5SxmRlKkU+kNIFpgRwDHD6kvqgqqb8xonn1hFRoXG4Cayt6hQ0LlZkqI1t6y6v+adi9YaziB
zKR+Z5vUV9q19yIN9581gLjmd9JqlTrkvKv0DjfoJc1JiKDH2ZQgOXGfKW6iwsPG2DGteAjm+QZh
nmtO07FLu2LPRv5O1UnZ05j16qwh/3NdHP7AsI2PBLuas0CtstgcnR5Va76P2FG+Gqo/nt4CazF4
H/hKZLpVt7QaIyvshDQcbVI+stLktgLqLEDnRSPt8MzdQIRZUMosiaty7ua/YAr3uf0ptSnPnkqM
9rb2n2TS4ZNJQMGe86EI8dVEZ9xPFwZYHEq1tA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12016)
`protect data_block
mBKRaEfR9Cp8NazrgB4sidhuLN00OsDNrz362fux1ezUFx06RweJYF9yckJH/rS7OY6GJMOSJzi6
s0gr6dq+6OoKsl7CZaB3O2DH00hedL9yLRMu48jPS2kENgjhGlEwQVpJS6YRwIMp9VmJWJ1l9h94
UFx0N1b0JQWDEEJFeDn9R1KtsSbCJUPKEJw58jDkZ/VYmHdJ8TeeiwM7WW4zbgPBpUJ/URptAAU7
uO5k9R1K975zW6rRC6wQb7JqRMv0KQws9OjX5UVlnWyc0a0CCOzt6OzykvS784LGH78cObI+038B
KRrfNOA1uukf7Ax00DURMAzgQzwZGxDjD9pK+9cbFwm86zij8qHHu85zFlWRnAtpGzFuvef++OZW
HG0HfZqT7BaJAwr/VkjWFH3sm7VwUQ8Z1VFHKLxusG0CQ8L5WrysVxnrBYlmGr9QXPaBIBPho1SL
f244Qu+8nL0AS6N0DD/IyPptX728APesdu72loSiujDYNGpSFpDazRoB29puo4lTGBNbFkOrpAGC
0nbGcwYMY8wU25szgvcTGGGVy6uQI6gZVy8/wD5MoaKRJc1Wl/kiXO/3vXpUHcSx4LUz9TGTYNQl
BVdtxTaTODKNf3K+bCmH5Eg5QQUuWrFykzV8oftxbZCR1kAiNeZCMYyb1EpWPQi4PhBv6uK/zIsC
E6af6hZ2r80JlCzWeh9vgcb9fAjlGbRvANYDiGuQu2NZaTUPZQgAIa7Eerww2wyq/aLhWtEhuTgN
2GuJJSUQaAO24fBrLYFCX8rfqbjWq2+u/jwhDqQKIkjONRkGo14IXHej57qPdIZA8FPkfarDE9Kr
Dqu22y0HwRFMvok8xJmjpLKF2cO5enqDVC618KwHmg757i/frGCH/3LrqNjFoiVWa5PIpMJKx5wf
6n9jfO4iKVPMNhCS+swaLH0LuFL6sqSR65AT1C7+mDnbQC/MggsDr8zxG14eJgE8v8+efxcZiL6f
l5udSN8weJ9FU8gOXTMNouRn5tv7XMcEmZm5prgub50S10dlwR6SMaSL9gyB05tAtzfvlBdZWWg7
fGeTQTWdl4J9LTMfr6EUkAABIEwZIXnC1n4wpFTQ4Q3d0ZsMQr52Y7SjGyviG13PoNuiKSg/9FjP
yhAxvK8MsVLxckfztSSxO/E+7Faq4ArKX1GaTjqphFKX3g/F7TH0crmm5CF72S/Oat3W/fcTdnS+
ulvDlb9mCh4KdbaybMgSHIsFuu388JIpBp6kccSu8Uor5p6Xop2AVTYeJ/3XxGKR1G97zfXE91Fa
Bbgh7vNzrHStYoCCo4QWAqpP0FU76x1GZv+ThSDmGAod49llz8a0tfmm8AXIs9WKJNcSWwX3th1p
4+bwGbIXtEUHiy6kQ7pZkyBWtvBMhe8WUBqXMnb/0q9syyfcRJvld24PJZx2yhpuYXScL8RGxyeQ
MI/ZVk9h6egouoHU99GCKNIwoB1lhB3uo6r3k97I6LtIylRP8Sac3DDLj20sQ/eRkiPPReNVvSdW
Wb/wf37h/Nf66+tEA3h6t//70dlEiolOa5ZQJtNpjYv7CY8wft6NZKgEmXifY7NWJbegwRgcPc88
3RaP6rSyOluO6xkRl58TV/oaUHFI4KwNjVIfd6xc5T288WtrZEud0Ar+Ei6BdXzvTar92HmwEWrN
dFBGcFukKt83CvbUp4sgaoO+G+V2oNwN1aKYOIekK+955wRHy4ZUj/7LyEI/SdJDM5PQyli/FiNc
0Ydk+4Etw5EKjoMgq22NAHaLwYcQopFaJJmD/q3ztv47+mt6PFGKBNHFk6SeA91+2z/mTivQ6bNK
58ZHhhuaCBk5daisCvJQvUFj+nvdyVUILZQyaKpvgFoT0IpnyLc/B4UgN2StPuA9VW3CJQoCugYX
+lMFWI1Ld7QePm/krWAEB4+6cLDNpmZqLXCejf/9oXjbL6/W9/Bk9iX8fIqXA4ob66FxbuTwDUkt
dlMGzLf8eU4+C6tNsVr3plJOAD1ayd+l0KjonspIKb+j/tfMaaAjKfETpV6MSilkClGSx/gZlpsp
ZkannfGUZFjt/Pc+ClegaMg3F8hERJElgH0JEPmuqgckeGgiYoJ08QzztjPGEyXP0djaE2GZ+Hof
Jrq4Mlac5ZFrEDr/zjql2R5phOg5PI+5XgJuxyrY4qg54gPmNOAle4DWZu37G+GUyO8VNoBSNLCg
85eGNFGASdmgaqlLVXbFMXm1CQSIJAnohjcE55dXf8ihT8hn73wCOAEVVi2DVTjzbwurUlLk10WU
pLoePffnV1B+T5Y+M/a3PkmhvT+6uLRjLFd1kiKcR1UsczHIFyZ78dkq2t5cQuBqv9ijp/y0c6t2
b8XqRxcoWCTrJeHbtTPrlfI3fDMeS94Ue5xF2YHucAfse9spydigEvoXbKkdgZfySt4Aczb4dX3I
NYP/REen5HXW955Tl8/etZ7UczrSk+xpqfMsKYpCnvJD/QFbgOP8ELkOHe9MTYP+5HkljFxYZuAi
IlBK7kEWNOsSmx8RgdyE7NX7/lIkptd9KbgtCX2EVJ5mVoJRVxS4diYao3A5ZmjNLaOX3aKblTq/
v2HLbYhVWdYiW8Byjl4aouCCOf1WdXEfLtqRTuZoGOM8d1PiCr3KniUwakcJ9PcFvJu1BztUOFsb
G07VpPdG0gl/yIMU9nK/1QUN2NtgHa7Jsmlss3xDNATUh5wo/ay46ZzmnBICU+ZabbBRJ7zZod+u
ZhgYXycCqEdPoXhpIvFbvHRH5o4nR2prRmXO/+N5qN4kgBawAZiPAhS70Y3CZAgeWAmyD2H+KrAR
EbNa+6s/ZSvWeWc2L57VE9oAPP3ROJUaMvI7ervKmOzNM+kBr5AY/ri95b5sv4snFgiv9g/6NTjl
NMS3Q0Sl5/kV0UrN2PSv7BBGipi2Kh8bDFvjtVn4rTNjHby0JwWt+x/5YqbuoZZleZ16PhaPspld
twCDbhOY4ZDnbsQ091yKBW0CgdO75vI22ywlcQ7kZZfdeoA3ivoYWDOfkTJw/i+7A8DC3uvhMrMk
8g7xa8jdawKtTZCshrpN1AG7YQAn+q1HyOudJyjmXBJUMH4HO5bdHQO0PW+MwzZW6AvC2pb0HAf4
0t/TrutYEUZ7EnsjwwjpqUFWhAoGkUbWtsmqyA7UQWlbMUaYXAvzfEeVRKmFbHyrgLF9ODJ2JV/K
GjTs4AidSFuy+ZuHX9+bCuc5+M325DQlvEIh0utFCtCCsCRAs0I9Y0gJudWhz7gtwd7KS/GCvACy
SBFEq1OhfGG2KhO26+Py5mesp52IS6686A4R7jmEi69dRQOTjyzHf4CeGS0Y5/H/UTzBHsIyfXuY
813PuV5EEWPXIL2LQaK9jA/U/HBDAtWTHWM9Fv878p1WLkmY9I794cjk7hwXKFchwKzY7yk76qYw
BzHJ18H8TB36eyllsvbdXB5KdCTlHf+HLa3m3uXeOIqZXMsnGymmj3d0uJPvkNH29so9e+JRQlaK
GjCXm1l29It/hhRRJrsZUvlJa5cy9n6+rfY5fnL2MEgVHcxQGMiHm+L+GpcPosmrHYyVaogLlw6O
bAwvBIlH7LR4aQ9s5XalJmljYwVvM+C40qZ08x1lw/FkR0RG5c+TztUe2iFdeSwG9eIdZ27rKFij
oCFaceOqindOTurJz/5n0224sRbe427fkazJ1FEV2vu4pBRbeT7POOThl6POh0jzZqybSsCFShvy
mF+oAtQCdMbb2eZ5rNN74JzNVyD7IxeIPfFjnUgB5tCSwQdRNtUWy0b927FaYa4m1Xn9kwvaoYbd
MY89+ZGzIpZxH4126g4xChlKj059qUFkO8snx2cVvCcfzorYCIqAu8WnbHpL9rFqnxvC1FGSUlAi
44fgOx+QFzEPg19+hRslvuDrJ+QkVHLtj06Eh+oLgwEGF0AeoVqCLQtOBJdLxVhaLNG0CifQao6f
dqnjWUG3mUxecOYqmsdTh/3xYDqcUcU5T3CPEWls8vMZpkIF83zyC+xGIC0oPzuwPsU3xcTRvHxC
EIyF+Y+F6nN9EehJ3LuG3p+e/NXmPx4spKvVBkhSfEz47lNJzmezBo0LbFqUzFE16MY0eQSP43xg
BoPNjNrhz2MyZIt+42llTtBdjdaQUh+XXofFThbIW2bsMhyvNH9egEjgBaFAMOY9fS3OECGYBbcC
CdPDsN4JsUDm+A3BTrxlz2agum1+5MZXXZZKG9MRUMROanWw2PMrnL82LQts0gPa0qG6XG1hv8bu
4ZL7EFLS0a3Uuw5q2OY6dOcJXjL0CiOb5cyp67UrAi59iOV33jOUGB+ZVoU+UaVlNiVbREqD2KCp
1JZfV+/yqD8yu7peQKhhXXU1Fwl7K9MIk/BOEODFTXeMikJUDArYMcxJZGBy6NjQRWlMPTOspoyT
N9ApBDy9BaIEO8vAYW/TYPU0S6mxIMVig4eiU9ucFfP/8wb4nCiRMEpffTnz73EAupdEKXFV0Oqk
npEP/oUDnqI1GwI5YT24FkhiTC9CtmEeP+w7yKPUXn48hNhYNo6hDGlX/9kpcHJ2P9KBaQbb1EU3
jsS9++WJeEkTky6D2p+M0VMObWcsS2Ke7yN7GyOd3wm6YgHSV5vAb2y8X1WRf0kKNqRtZJOK/0uj
ViFbUEKti2DTDofvMr9TojCoT9wWJex5xeDezACKbWgYFc49ajwNal4dZJAtzxGNFd7Hwv29Juap
B+FfKT8fqytM0NpyQn7Xgs/zCuXubmKnR9oriQmoefSTVAgnKQ0PQFNSzMN0p0GRmglU3IY5ysy4
vh3RgB7fyVIR5sb8vtMUalS560AkCMGGbUD9uZ54t+bdCOntk93H4ZxJAoOF7kcUI7GWZVS74J94
WogFv8l6TN6MjP6nWNHINTo5KromdTo30WaeywneYpB8HVe32MRwR8hPwxtOaan1mWclbtlFJUzr
xMZ4C5BG/lj4BqQGDOpt8rOhMQr8GyRdU/gDGPXHHcLzFX+eJEYz8xW/rGsgxH7Uq8cEcb4FR3Wx
5q9zelgOERzcOp9RJ3YRMISjbXTgpHEsyM2EB/quHrno4SawhFOBLqo9OObZBisv2vSM7qmNUvdc
pPWahw6oDcCsETCbNakr1w5erKP4OvLCPNPeu0e+Aq+wsc4gjYTO4+KPrARbachISCIM1jQ2+EQb
NJEsaRxtkiT86ZEBRYaR4ufKaWqXp/ers3g/pNOjrr53z/U9auoHHti897fqr7za6pZJb1R2iTSl
mBbInNwRl1GgyiuxmQuCoT3gZTEuW2yKLPBEfoEU5LZabczBdeQgnBntbhiFQxEIXv1F107jX27X
2pKPM/5Z+ipIv3vqe+bYXWpHPVguzSIAapjtNvUHaBv9fuJtAyfiPW9Btt50xWGfMDLsNRGExzAI
p9n6GWNgo4A+RJ2ZBDUrD1VDMDMcm6UR5w5LO3owhnqelXshrqwWl8oa5Fp7zpKD1B7ED2B+SJmv
1jQauybG1SHQUb7G3J8/gatKXnd3qRwO5mF9WdNd5n6mgMnpmesU7KFD+NBrF9XHWE9OT2STv+cE
pJljZUqRKkaBv/LBIVmGGEiKURPBxYNPHFvvtzavpNT19zKndi2qoCBUcUxYUIDmRKvx+IAHDCju
gtkoCifQ6IyaMijMSOuKwEGt9wVm7JHUPgL5B9EOsC4FLpaI1GANgl73Dlvf2j4sQEiZ+hTT8YB+
6jQYQwNpl6AmWx2hsFX1lP/cpAfRtE0lllTMIWaAI5UOtanL0OLC6XeONJFhhZMLndKRsYkI34ct
d3x4tAA08ZRXiZodo2dOpZd8txJ77+lrvMyR5ZMN+eaEaLA1mJxbgP319cpjUK1tgCRC/VhknDFv
TdbmItAmt88lasyrwKp5hZoQS66Ix8sURS0Bm4EaEkOde7ndpd7P83C7U7LAH45zqEnC/IonmWTf
d1RP37MgddJ/41/owOlQAYcQuxu3g1IWbj+idtC5e30OtmRz9tLBjkElwgP0+BygGt4ve3wBiTkU
50jvJo3EJAIo6iqw9Z2rXmOWE1eICsp3QWd4h6wPn/Z/FQyA6sz65MUUiCMNr49TZpPBwbdKXQ9V
VY0i+DbopLI/fMQZkT4bNkTH8zL4arblJELBrNqc2+uTKD9035/nrRLTzHD9DXmCmLa6Rc3dgbw9
dkeWKlvoGh45QJ7UPcRYIWj7Wx3oc93hAMwQQ2cWRx6EvkrKgru2n4mhM9Bm5ppPbDN6M0AY8xXG
V4BwotczRemryS60pnQOOu4pjDfV4Z7QpmV+mMh+cCtS88NCjIF2xnytcBff/5XSw7JIumqxC8CX
BefuJaNHHh0TYo4oVIRMHL2yT+NrvV8ohYxDFsVT/T4aHz984GhZ6W9PKrtmZ7m4daUt1Pfvxez8
pZ1PL/pEY/dchtp4utAYI+3dmRtBQxNg5PUaXVfj1L8PCOOAxy8O7wntKy5WsRxzfzL7fwKr7FgB
vxYT45a/hfFJxNhy19olCb//d7KcOpSPW1U/i4s1obH0wf/gPfpgvsT6tMk+O5X7Difu2utXb2/0
1nT+ulytAWeS7cui5/6FOjh4vD0uMLK/LFgSVOI3ItXQ7fM/+7KXIPPi3mF8fKp/3BXgnNL/6tP3
gOB893rtbO1VG/mTVndiBBoCgWWuJg4TCQgF8gucuieaxkj1SuKZ3HMbfxuSSjGH+73L/lhXMU7R
KpqgZ7zj5ijrbICZeSsTkEBlQ5LQfgAPhRsgBr4DfFe56Z9erUXBK1eoYYamUeIwJEFvq0blKQbW
3duWDmELW6C/82HjoJDKiIysBD/fFEC+K+DOHxz6Bvy8eoQbPnY4c9OEmEQFzIzQWHUDpeGvMlmG
H6iYC26D7aG5PiKyPrIk49cHE5k1ex6jM/FcFWjqrneVdaVGBAlHtQZwejan9BVXdVnQkF3Db8FV
N3SJe4kaIlzrJgmEmVG5qMr2uBHvT07o3ngbSIWh3Lshi/PcIfybQ3/sXgxZYtyOU2F5brMETvCV
yJmPyURvxcCtDdZtMQgxpvlPiKxz2mQY2ZCyweY7apGBHxq6yfGpb88y2h7Zl1HaI/FjrPMNbGkX
cWL4Rmwa3zbuPzHqkWmBDwyjWvRINISygAd0XXshZumAL9miETaZvwvSjemrNeW/K1c/UfIjxmxr
VliR6p64Pt8v3dVmGYL9NgRZ466dbNpMa5awsPsUlT2ttwN6yGaAEVN3FhskuWf26EmJ3dBVsHgV
/Lye6dME6jMMkfyEFV+05OJf4PPnXER8y2GgFlfX8q+eKtMAMEM+mSulMkw0+8kTOVOtEHBHMPcD
8FGk7CDD2DkGhPtmPeTjnqjTU34tP6bs1YdIiUEQyoKP5SvBtziuVCP8ajuktax0CiryzDuO+0kj
2xOTxfU36NOVSXVn/xBrNfJNW8TASmSRLvzQYBpbfLa/dCfhxXygNthJ3Vujp77I39mnqJ7fO/ch
FSm3Jln5jYItxtMnzoR/pFOyNF05fpl2qljzkiSBv8YHSSFU6oe+k+SkZUERKnwIaR0O99PRSyR0
IwWlTsUIlbN7aG9D3Uwzoaeje3s+H5CBttWR4LhV+ah5HEg3+j9M0l7BQ7GfeO3Df6nEadU+pYfu
LSZLHjxErNijlzMtJB7ioTPr6IyRzyItAWVg3IJmBu9c3kFrM8i6a/CaKpOusxPbYS9pxa2pMlPt
Zh0OuvIh4vWnv4tL23n7uZR04E1+y1U6RUXKtdeKCd7oW+78VkdEfg23FCQdcebmH+67B6HsqLjp
7ZHcKi+ax62kFp4prSHwUJAW1ed3ARS3M9UX1g1+kreztvZ+87Y4nil99EWkD/hF+Jo6Kf08u480
1i8ACvRy/gbNJ6BpmrDTGjBUftpNTP3irj1w5OOG+UMoC4kNhJxsKxcSQ6swFZQu1zT9CQAbeobO
2D39DKMXZhBOwJefgZpw1g/yywsZMl9keYRbvNHkAxBOsyqQPx+GcyssilhIgitXYqN6vUbHHCdb
bG+vjSzODCXxf3ydH6uYLfUa43bSb4MSzWfROSBkDFHyMPaqL54J1kcI/mLHnHuC2PBp+/2r0aK5
u2lmh7XsBG/LwbeiCrDA8atR4M+muNpaJL/vwWzoLnfqwxLzZKuHNskmkMnvGzPMJgjCf6PinV0E
2U1H94+0eYsPcHZnLY+jRaN1efyOIU2aBRJYH81S0imHXMGS7+o5CbPPfggA9cgy0kwjwN4T4XbX
WHkgESikaD6vLS4v8OPLpFBoyE/JwVd40NqKk5vJd7xIp3VFDcPKT63/wdHudAwF3sS55esf7ABR
4paHKoC5bWg6ruCiJqyV8/gDTvAzhbVCrY2HJiFvOVwAU2zD6vsuZ2dDFli8QCMFLzbyw5OJ+ugL
qkO+35DflmflOTaZ4Xhicdegi8o5+L117PqrTvybTvr2wtiBxoX21yMQ201jicTvEfaqnGdyCx1R
pcwLzvyG96tCoqz6E5ervF6fIe8f7nqQo1XP3VI2b9RHcfskRT/3JA4vhDYuHFCN99tdNdJwvP+V
xdAD7cmHs/qGzGsbZbR5ZIfIeNeYXgJ9GV+dLPT0jDW2u55Vys8hp3pxMYOl7OtDG6vIz8Zf5r/t
d3AuAmpcFo7foqx1kfdJj9E3o829O1zjkkwf/eW7/OFhjaAecEqPGDfpX9GMy9LegnV0I/dmq2VH
3RLi5fI+ytafeo0jIKeTi+w0ePBPLhX65e2+68Qaex8mtRjY5o2gTT0gwdsAexM7uQaqZ9+wFmbk
lQf0Rd/02Q/ngSWdG5/opw7DT+fW7d4N8KBgGjrXP3A95auFZdl5ir3npFdFgR9OQEubICIl3mKN
ijSuJZyjyozXOdz3Bq12e1EKj2nc0UaxFzFp29rp1JcFD63qsetBf9oX8w1XQ9npaTB1mGe7xMoZ
fwDJ6X3Lawro0GOqTGVdbiXDhEVAPUll3ExfHeJp5rILpROAw2flIUbbcOy9JZqABENQN622mdJL
i50BvhNEx7pJnlgnWGWFxNXFqjMvHFK2+71CT2k9iIjsswoy8cwYW/3JEnB6Rl0uSMhigP/g6N7G
Z6D0nDBtFmrGXjCtPu24XGC8kYdnTDtjTgCSy2IPcfTtQk2LzSvhXIlU2/KcLWKZ3HA+i7WVoKcE
qR2uQjT/BXgT3JJ67Pee2s6rpHAIdC7RhhhyO82yPNqGIYDMkLzYCMnmW11tNCoqxMFFfbPqPlX8
D2OvGYlAx+3ZJYJzpSEiJum5YtFhSa1IlU8WryS8/JPEAn6ArW2YZvQL04HhWpRbNiob5e/x/tpB
K1rOkA43ortKDlsatg9COqgKzRehNVHzWYE/10FKDMHkmcROWW+74A96goFGcU/MQIijklo6N3rN
ud4xPsCornwH9q5/5arcgGjQeMz4waNHk71H/7a+7MLJ+nA+0heRjH/gA3EZ9OCtR55fms9eggZq
eRDcSkhLop2iIHU6USQm+5YavPZ6Yk4KoluAgvv2yYD0cTxQrfjpuj5LgmLJ/Sx6gjNQVMpr740T
GhQF8gXyJVacdoQBF8DWrus/BmbiXcj4YFcD2x2uAPNPvdnEoctoVn6pSNxTQpbFTUcUlM8oSWwp
S9i9aUC2yThZPXLOSeOjXbaiQ/zDNTKKZqO69SQXyIGiXmTgSx/S8azjjVPNGHmuy+RMjnhsMvF9
Rkgr4ZPbZ6A8oYp3WYPFG/skqNEOeMvKFFJNikI8hBozxB9/HrXf9W0h6hZBPhUwzq0z8DXXHgIw
9UxKMwy2y2Po1cbHZSKRNmWlv0WpguTzoEJYEj6iISv3rJZxKizsRwBg7VRQMx+dDnWLRmFFKrYw
lg7pzuRcqvYOkqHvnItjuY2mm/gCbB1tIzp7mYbYfA0Tye44Wb0IPlvv1TzMbfpahJRMo500r8Tj
VVNZxLoU9az0zxkwNy3ey/nQsbxjz8Yf53APAtWn3jCh9Fp8b+ncbiv1peEuNmRTbhuGal4q70oG
kBD3gG1VEUU1TQ/EAh1mGjWEMC0rXTWNy4FgFdyoA5QkWWgTIHXklwuEr0VxN76+ccAqFQbNCQ/p
u4nuOpugpyUan4qK6c6GlKXCtQYpFfYaTviT7M5+l1nvGUX5IH+R4IgtTpKao4YzYQR8DuDz2Qi7
FZpYsYyVMrAo6mpJQeO9NwCfySf6Ey1O7W1gtUCv/lPkEM6SjGlvdTSKRz2ic5EBhgTSj8rTdvt2
rKCP0CXFmp1IT72fKrjxR46wVrGU5ZdmLSmXy5ULuFnHjIjinDuiR53Dgs0qzSQ1EnlsUdsyhcg1
ESryjem9+9LGbraKyK1881lX1DlSxTiqxd6r5LXhbPSB3ZEq4ZoYinobTTH6KjmvzX3I1f2aAenr
FB1u+nO05yjOUiFe7QIqTOTB7A0BJm5E7LCBESEmwbKrwcs8enmMA9z2cm2+f2TV42QVPoeGhfJj
zXdXmdLojryfE5llOPtLYj4EYoggLWLsj4kSNPlsaANThKuQ76DBKqpe+TwwmNGSO8tai+6Wb9Qc
wsq12UTjBLBhAYHDM//MoRmExTjqDzO9RSTYMbm9rllZUnDU7VVkNNgvCqsBDJ107Wl8VTBuIuEd
coM+CiguUvlC9964Vh2HxyEPuveJfZQlD3oF7LwDsiMra/SBsVIlI9S07aMC15TQhPrNRahBCFSV
BKNva6trXa/hlC2qZpDGFkwhI5wa9J7xscGb7J8jerfHAY/QIl7NwhLv0KgNH4MrXEFSW/c3QoiU
r2iouD3CehaLIqO181Kx7BZYGkj4ZEwnew4zIRykMNsEzvMZQ/99OQzj+i03Bw65zbL3a4RtZ7Be
CN+fnoEZRFyJBXR8OYmfWK0Ja5Ha3d0LieH7sB9ObWY2FnOt4FyB1xYbQm/+jMiOP9E50fVeI34r
xdXZLsqOBPhLZbl01eQUpo9nR+Nh4A9643EFknJ8dK5wvqQ2pE7mKWlhEs2133mt6Vh4e/Pic12q
Dzktj5iJJAjXLkZR078B7YFjWxWLmcHQCqpDZU1TSxr05QBFHhxcs5YQiiiHke5dmDmuPbgxm1/9
vv01zwcHTX4muOhYWxMTtSxEnzYhWYedtxwYS9PEF7MkZpzi1PboW+W9u++vXtF3+QyX5orQQHAF
QGAhel63p+eH9FjAGTSv1eih55r6AcafTI/VEdbB6MGCS+9M/jRD1thQCTSWGMiZbrZK63/iQdw/
jyGFFxxyJ0lISdcv7neOArvTt0kg9IdLokuWtVk6qOgwYaPezBzruoyJGbU6C80hUIKLw6BmLHVS
T7P4PXQ8yTAVR+iKW2QZ7yIPe3ZuFWf7aJaLL5T9Sf0RJOYAVY3syM397JRp+B3uBJrj+teY/KRE
1XBIwURc9YK1d/bUX5Ar4KVSiaPArQm0nnC+tCLKDBoyY+8R1xm0MPCUzozlV6Lf6UhzpG6pr+Ee
xBlyHgtfEQoKS0NM0BW4nOvMFmr1itY/kyqkuOY/MZwh8ARtNZNyROrHbMLjnGgIgpF8oAK7iOzc
JnoVS1c/O/GEey9luPxvwPJ6oKIH25nLyVEHZ2R6yW3YxF/xLxD3wLX/AlOxNVb4x4GWzi4p7DMj
kDc6g8Sz4J391DWz4YTGDYp2Q3jxUx/UL7IFtTyzQx/oQP7jq0jd+ItaYezRcrTCCcgg76az2UfN
C802g3Sd+EoyRhx3pDrJeSlrEyLkfTibvYf/Kvfcr9Y5JEo+tfIXN1E6zhyRbbxuK2HBL4xfB2V2
+/vgJT7jHsk9HYS4phLJqALrpMwYtxqpZwjadNHoaGnt5DyYljrh0ICk6RtYN4kmdFxEBJtmPkvM
8lOjvAF4e3zRKbElyF3TgreD++NaSNnpNXlNXKsdT2rKG1uSCFxPb1AbSXP6vJx8xO8DCljWbacb
SDsVs39GQuk4wJsTygH1f2vavq8hkTDgJvgdkoL4aGK1/gih7Sp/ddEIw6z1SYtAHYj6emW4toRI
SjpJ+N5KtTjSuhJy2qwwayXkveUOtpbRinT08KgeZ/aIrEQ09A7fv4HjUpPX8Hx4TW7+NE+TccMA
Ty4ROxD8EluM4sgkDiBivXEx3gHzOGrNzucSMqQ1QoUWC2OuQbXAc+eHr9WKwem2ZBdOuFsGVZtl
PFKw7QTdJh8ucIWfni4i0Z6mcCN/EZFPINyZoMNhCnWHY5zIZPWqgLaVuCRTRQmlIQqekT07lCGC
lOZ2uf8YN0UnPYCSPFnbBul+2ODBKP0uE+4xDEejaPtjMk3Tw29dIT1sdzgcaHnOmON85ufJhQQ8
ymrCvXXx43ubOzPNbq19Um0u61He/5PNcISNDDzniGKvqDwqez2tKXv0rAhTWdWJQFyeHi0okB3w
NcMAW0Q1Qb1ELFHDrMGwtiLsKJR7jk06AVaQmLNR68yOzuJqvPo4Ko/8mU1H5IZEqLBpPxO/V7V8
grDlLX4s+2VXeF03K6MXZkePQVj0igmRdhyfENom+7M7n+Hf777kQgJa90gznu8xg46KFGnpK2An
M1KT+QhKdXTOZIqM9cgIWxm3a2gW9l5xbcV5b073iZ4BZ6uQ1/3j0Ml/GMHbDnx9D5oqnD9eFDcB
eIaU6gjsDhy8baOQ9aKC2OID2ypuBdbuF1chIIXixY/CUlM0sQZkPAm7/m2bw2Xjeiyp9x9jBpw2
H3xTnvU6YosIsiiVEueFhM+tVbSFppDb1WtBlwYDiRy2hWIEFXdJLBSmU5nzlwb71qwouS7/gMP8
TCfBSuzeUEuIi4OT1bOAZfbrNbX9RuemQVsAigTH/3zjDuKCUqZzdtt26le/yfH4MWdX1e9GYV2L
p0YwNzzHY20RVwLN9PgUxVQfr+5iK+LkGVOkdxnmFlvs2tAVCm4Elbb5pbHXyruKHXwH23Jk0xNN
w2GyZmowAW0yyVhT0aM0C9P8RZs7Z8voAadojCefjDUqMFoWApP0TX2IMYJApGlR5PtmPvdOPnbr
4DWTbFqf6nWqOMuzMB5gJWI8EszBLLf9EQ4kAj+iqGxndF0FGPIaEjcfQA5fRR5jGzHqwbmAXYzq
UBv2iYMsepB/aCBc9g5Y0I9VZOl5VvuwlX1gVkkT4ljLGkHE4dpFTQDqAeTsiciYVlxvl9DbvuJa
HlZvsLv5XkD/o6LS5EDNzzLjOGLR6ECAdemyglDk2E+MY1dGFm3Hb0DFR/ZSaUzr953cTfQ+Y0+/
LN7Ax6ttd56zk1VK7Ow46hINpJ774QIgTCXvUHvwgnHqWOM6Ne6x65iYZvClDFHz45dmlicgZtfh
GYzlN/ICNv1/CDvWJqSqhC/thaPSJ2hLAtjqq3nZpNMtVoPQZ/gLAuJwLOsdJSei9frnEa2xA9Li
ZPbBLoPZqnyHk2Zu8fhoknIeXLy9SIVdE82mSB/F0XYJC9D24q2GcH1fsK9tOsHikvJ1sdOFEHWJ
MeXVNwZzBx+gW+/kcvdZms0NLgo0f7/HXh2KBqxvWu5DXqDP3b/Zbh3jXc32NhbZ/6yzneWMt+uQ
hlzLIIfaGfb5/XgcFoKtD3uH+oYFz3hrmHHCUCdhgHYYWMTxafivKjUcITTtcjngI3jPmWkYtJUW
eHXa/izcR7TME6NmJf3Q9v2Pa8NcGLshFRjq4RNq6Nq+0dChwwPO1DDl+KgBLvEZ1ym7lkGJwtrm
xzBLWF1LVKY0/B4SQBuJdAuHEE07dfPslVlnqwswcP0dpqy3/AKO24r3ei0hNoVkPvpoJQQ5uNdW
t++Ga6yHW/0Q95JPPJ/1Qmd2ojQBqCeE6mNakbwuGD8kUPw1FPa5614I267b/JEXcJwxSaYBYqbl
fZk9bBq1ZT1oyIDJ9M34gJSnLZQeMpzbj+XRXqi3yxCdeTe9539p87SLtvwfcNpohBnBkY3cIK4N
BFydBjUSI816eESwKMJZA+naZdJRF5hZehL34ub3OpEGslBAf7Hj0xv/UevQByqwbRaJRSGaCr8m
WZG37UOZnsnDa+EXkq/KMLo1yGlivmQ+BfDDx/DVcxykzlB1duS+WtYzGbKNj+EGWI4eaFIV3dG7
jABtQF7WRI1qQ4ok8GIOozNl0EiJLDalQ/bCbdmlFZ88S0A/x7Xw6Kzo6p55wdX8WihdMvK3yboG
4549WU1vGV5ynRePSojlbuVs4+9jq7Z/Xyb3Fq+NEwiPXoPd5MxgpBw9umRjKiVX5LuiuIEM+LJW
l3qJUmzL5LYiYbHnQzhKNeZi191ScwW0Yj67iVFm/u8g2sSOk/c0X0PuwPS5gmFBRqAjIOIHmB+Z
araI36W6OMB6SO/biiKG/y6QfY6B8ZBzkAExspJ7OQ4sLEA7CAdg7BGAiHoqMpl11Hz95XMCh/CJ
FC5ehB/w0s/sTKtA66r3qurT7cOUiTCJQeKYHHKy6JIxLoohdzjyQQNqGa9IaXQX2l/tKdR9tCVO
LyB8NRKmkE7QNwii9QQ3FRavrrOPhlqLNUpqCt7PAZGK23Yu191J9Qem5fO/atclw68dbxSpTHan
ajKO/uaI+a7fEGnPzKKpBiihW4QLMWz3us3mfvjx3cAERiPbMuCsWZICJ0TFYQyrl5ST03h3c+YP
IadzJIp8VHLKR7hbNSOR9bVqO0l9g8WuRgS8gbyIfF7J+aC935mVR30OJ3FeXS+9yUGRXE27EXJN
CY0nQsEzrRc7REdDvAvmDz3ThQ8hnLz2aGPufeN7pGv32O9s02Ogg61P+XhxnRebDCZ08MYg36aI
UZySAz6GpWGU7tW61MGJGvNgDGL6hHbg2S4/2UonwIeiVy/kFW6YqKwJTpIR/7HIKS5GlzHevJFR
0rSQ3hM+xhPS6OrRVFwHMIqASY7wv8ysBjKz7hQWWdFMZboiniV51fyQ/mJ3hianBMx/zWG1Xw1S
PHW6H3A82SsuGvF3fnnjqSrUsdgvbcpX5hYeaVaXcYXLF5XFR2wvMHqQgX5ouZClXBAPo6vbF87T
Hp5YOkbKgy9PWnTK1rD89oUjqY9X3bMl6CF7CSud6ggDmTsAIrXoAbO6wZ2fmx6/ByP2ZXz5HZvr
4cPQTDYiJR4n7DUXC5eRZQwV7vq01WgxlyhaLBksnSYdT05q8/t/VgwPBljcgkddfxVwWN2bFiNa
dLA34WPS+BBVRCf8Ks3K+Fdkan9NQU23g27OBeKDoa3xzTm6oEXLG2EWWlyZsoiqZKWkA7nIaQy7
tlyF3km2XuhKORknaS5fuDMqHfYXLF0vx++gVEW6FcTD1AqltgXwBb20OsKLKcablugdCtYVz09Y
YbROq7/J6/sEductSjSFbYyfmdgpNBTtfDO3xfIRT1fGglbc7dG+yYDyjOiKzehV2IvV9cF+FFux
T2nU5OnhxwI2sGXxC107Rn7tKeKz3I91KWjmtu6H+74bPKb+WN6AzDS1eLqj3ADYCZAGblkxcj6M
dpiTewaC1j8TIt3Gg8Gxa7hibiu5aYzm81hm7AGZjmdOxtGb4b8z/Q4YgdeTZKRhUWl9nnti3LXA
hl+2YAHD0U0CZwVvp0ddbtTp49aixuE1XCjVciKsefNGG01KoBDiMsVc3N0DBBd7TN/ydWD6dPnI
ULoioxhmJ97ltrFIzmM7yfazoqzzBZB5Y2oaovctMwiIAxF0Ss4KOqaj+E9iut1VL1wG+i6rj3LR
CN37dZYh4wgZVooIRM9ef3d1cKkGfEs1D4HsQ2urlQGA/X508Su3eCR489iuF7OVITVf1X5Ceipj
xiVILrMedjjBVSOuTeq0rwxVgZ6QDRfxja01OAUpS+Pz19W22G0QjopchnuNZr+6cSKVEU/nGNxM
Dq5ZzaDwM3GMyWWkGZYp+li1s+8Kuu4hPLPAXPJrcbbaRsH7bnVIqRMC1KqYEZTH9NHNWXoDv35Y
NS3ktEnmQ3gRtt/+rakzDONACHilwREIG6TlKSJ8NKPo5GHbu/QgOh89KXb0OIvnzUa67hK7eGhL
prpQrgeeygOi0MbpuvFnsKhLMPs63tPQcQyha3Zsdc/9oNlgqaOp4odC9QrFmBmseP40U4f7ITZ1
rEy7sL7Z4DsEYulboi7UDOk0IZGRs5Fu/B6bkpfZGaI5ghrUSmmfwN9Mtv1hJw==
`protect end_protected
