XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~��ʧ�d ���L;�p'�Z��(v������}"3W��ul��b�},+O�k����yl�SnX�h����n�P|��R���|��$E�;��M������n���
 ��p�p+���E�
�J4-j�G�T`�U@w�rÁ��c��wIX#+�7���vJ�>7���`�2�U�����''σV �"VӀ���^���'�L���Vc�H�99� j`���*Z�f�-M)rWi2���Xd��~�e�\�M��q�<$���x��ƻKG���ēg����9�L�(�5���H\S�����20���q��8��!9m85ꕴL^ �ӧh�VҮ��|�IT��,��3!A�ϻ�e(��QW��
ײeU����>a������e���-d��P�+(}jj�K�?F�Gͻ�k���>\�u�Q�-�9��������E��uQ�s�f]@i%G���|mI���Q��v>OʲX���@�}`B�����nq2`r@�u��"��|�	E�1#AX���v"��0>�����'[�/W��!�I���o�a�^`c�ϸ�a����>�ب7S�@�!�_eG�ޱ@��ӡ����^L:[�	�_p8ۇ3�>����
Ť�8��<Ϯoʻwڋ�UCu�[�n�c��ᷳf��lTKͭ�x�=����0	��N/����Sb�����E�怗0�FR�[�^Ԅ+Ўv@��Te��`Lf�x4N�z�*��cQV���m���Sx����XlxVHYEB     400     1d0I��
��c��Jw�'�;uˀ����ԺK�%t�M΅��ΒIku������52jZ��N��)��FAy�KMj�\Q�`���N-�N�<�>Q�o-eā�����%��9n�/���Ӛ�
�_�sy1(����Y�I����=�J;V͓��oӬX��A��]-d�7�bX��L�&|�����u���z^��e9j��||tU��,�Ŏ�W;ܳo^��Y(_��)�}�ʡ�t�������pl��J&O�6Y�u����`��c��8����΃;��~����5��v6&t#M�[�W��(�V�F ���b��ypހمqbx��U��e�v�?J)~c��-z�si���ą���?_��RC��9��$-�M٩��_�٧��;�؅+����&g]��K�x�A�
�(�3w�u�\$���dGO�����8��n�\��w:-(������XlxVHYEB     400     140a��kb	@�rB��3��g����9��4Qƨ�ğ��Àpw�B��v�]jf��ǽ����V:?�����>��w�_7q���WI���Ӿ-@{����ջ �E�#�О;b�{&u�|�9܇Ũ%(�n7���%�>��)�e9R�գ��O��'�P�螐��Bw�>H��ݞo����A`�GG��M�}�0K�BV�򚌀P�]��ܐ7����iL�x{Jo���|�ٜY�����-����+����B
麰���]�����6y�p5H.���B�{�g.H&��h��N�`��0��xO��R���?�'��b��XlxVHYEB     400     170�fT��-��=A��.��G��Q�IA�~_�!Gǂ���T�>��/9�bl�ۈ���ѤQ��U�o��O\�]!��7�h�y�Y�V�tTɶɟ1RA�3�.����AP�ě��=Z"Ba��D�Tc�ԋ��{#-��2(m3)��F�+w]�L� �L���W�c��@ ����Ң`�����KH���h��q�f�D����&���I��	_jn	����s[��TL�+(�J R�aΉ7�*U��aw�%t��T�iO��r�� Ji�V����拖��03(ZiYQUMw-qJ�lXp�/ƢVo=��O>�eD"|O$:���*���Ѡ#|�h�o�C)���J��p ɉ^n��+w�XlxVHYEB     400     140Q����B�)���Q�yP\"@V�o���)��*�Z,���Gv��9/o����{>ǗP���`9\8o�#�&C"�7�(}��BT E�?�8�ޛu�>��sZ����8��07�l��B�-Q�AN�R��#�������S�ø.j9��!w��9[u�ӛ+u ���'�j�MOduK�Dꂢ���<�����L3��e�O9;�rW߹���� 
�9~]\��sp�54�6��=�<���?�U���o>M)��}�	�D;$ʠa�̏�8+��m���a��o��,[��Rr/Mg�m$2]q���րXlxVHYEB     400     110�Moe��L��#���|�~�� ML���.�������A�K6w*OV{Hj`R��,W��6[�H�w8�Ռ�<�=#{7Ė�����9Ov���I��G+�})�3K�|/�YжP��L8,�S�P�����y`��{���^��"=E���6�y�(cf�������y���l��L���`0� �*k�PT7��䯮��]eujBe�K�4��d)ϐ۳ٱ'��O��J�W5��ɺ��6��&���X�i���d�M�q`U}uXlxVHYEB     400     120J�퉱0پ���y��F�5?�X;�w~�͡�C�uV�H!����QAmEO�W��گ�����u�t�=��r�:����K�Ho1�?��6�!����H���X��p�k��י��J�=yFm�Ь��D-�H��"}Uf�� ts��G\�Hթ�j��M�|�9~���?X���ObP��6���(Cx���va��4#���%�8��#ʛ�ىc��׼GN*����NQ!�h�`^�P|��i���F	d��kSG[�	Pwt�M.\["�#t�e{H�9��\9��;�XlxVHYEB     400     140F*��}�Ą�#��t>��0L�Ч�kN�杋��S}R��Bz�*��KDf����Ryc���Px�R������= ��˰h|�$�(�<��i��~o��/��?N&B�8�Z��K�ג	6��8#����D�i�tZ���!{&�!)�sDr �mF�xg/T������ݞ��7�i��@��09v��{߶����73-���x��ѐ�X�V:���r�>�+#��"Μї�)�1����;6qG�[���YY�uQN��ga�J���"�_���e��1�h���,NZ+S��O��Q����݂���E\�<�X�/Y���K�XlxVHYEB     400     150��[�ls�,�7��]B@a���]�"}���1L�E]o�K�fs�SjJ\_+��/&��Z�6ds�L�͢��u���Fj��-���>6��y�Ǝ��7�^����J���-NlF��s1��Ս: #WPg�a	��uf�J՛�����֌�Z����y��Jj��E� G�~a0R��^�Lm�az�9ć��MI�j�`E����Qޖ����ۼ��Ò�cz��O��z�u�@�w�l��G9_W'���MqM�{���x�Yk����Ik����`�|3ܷ����NH�m�T�EL�����Up��҃�9"��r���Fw�?��B�L3�XlxVHYEB     400     140'������X��M=�Df�0"�Y�������sԣ� ?���v�1��'��e�ڪ��kh�%�Aye�8�WJ�5ce�����0��?�_Õ������b�xefW@V_�"n������ aU=�X�5���g����by�x�J��$��ܮ���{����E��Kqf�h��.��S^�oSm�+ע�.֗;j׽��"	K�?n
KG�/�2u�ؔ���hT�/����8�� Ԟ[�	'�j��|�z�u
�+����H?��r��ULE }q��:��12_W�����U�ph~c2�8W�8���Χ�i��XlxVHYEB     400     100\7�F��j�_���ݖo	 ������i�n���H��}�Wb����S�>kwӤ�+�{�\d/p��>/��؅�x��8�x5M��V2�]D��3�ɱ�b~m.�����R�j�g0ge2�����>�F�T]���T��Nio!�e��?�3� ��κ�z;%+��;@6����|ƛDt�xh�t�S<��ۛIg���}�2�i��]]�gZw��+4�1��2�<"W��%�rg_FAX�����OV��#XlxVHYEB     400      e0�tv��#�����K���j���6J: �R�@�+��Č���B��ƈܪ��S�"�+v�=��Ӣ4�nD�4��W~wO���OY���6�6������4���Uw�m��K�1vt��Ĩ��eވ�/<�H�̬�6��'����S��#f�T����f�+����D��N�w�.0l��&O�F�HfZ����������B���Mߥ��»9ͷ<J�%��XlxVHYEB     400      e0�bN>_jV����ZZ\xgQ�DV^�F��=$!�Ϋ��יmA�3Ƣv�8e��<f@� ���K�cr*��cqA�_�+�r��ɱR��}����
l1��r�|����q��>��5��j�S:x�&�������g)�k�z�b7�׏�s�$"��d�Aٜ��Wׁ��U�-�c�:e�r!)��D��k����;��lH��Z�����S�r�T��UփXlxVHYEB     400      e0v﹕?�q��,~���Lz���^r�z$XN��T��_��}kW���x�i��<Ŋ�1=��xkH��,�*t���yg}��\�p�o���߀�q�F׆�i�w�N��W��/փ�@���)�G����������!��{%���y2�����0WI����9�W5m�5���qP�Ͱ����m .=����9����%͉��h��{BQq+����V�!XlxVHYEB     400      e0y1�c�Udˏ_�N��8�ZPـ���ٙc�l`��H����6�GO��Bg2%���8� ���]�����`�������@�xZtu��[�[$���W1^�]�20<��ge�,�Kʵ�>�C[�$Y	�Jc�6����G
e|ͻ��b�n&�|���%|���1ؘ�-���R�#��!��;��@�zt-+�VG����{ec�
�W�^}�#����H�RW�q��XlxVHYEB     400      e0�����a�4��U��Z�J��u��+��r�>�8��ٟ���*�2����%+���Ma:e���\ó��>0)$��O�m�cR�xZ�ە���Q$�ByVCK��Z1v�Y�{�Z5���ǜG\��u]pxP�F� �:|0(�r�.��~��u1s9b �H��n�6=�#/��P�t9��Eb�"�螺�q� T�W�ҟٽP�4��D� XlxVHYEB     400      e0㘦��8yRa���
%*���;w�7t$��dDL�[�yE��e�-�G5de'~!��x���̎1��f�6�7��N�0�ⅎg�����"�C�U&�X�)~ϒ,�b3�(-�l������*m�,�.����� �p7����I"����'%DVDЋ��b�����VZ5��Tp:���-=� =���5�P�7��)?�"cVd�t@�w�~�,-r�B����XlxVHYEB     400     1c07�\:��ʶ	�(�##��]G-\�(��$���Lׅ���&���IQⱒ���׺<t�?�hb� M�G��Y&`��T�Ͳ�gCj9�����A#/�эK�z��L�4�p�~<�0f��s�'�YmS�sշ�e�T��a�7���ӟ%��>�@4K�@7��qu���ڌ���4y�&9g0�O^܂G������DBb7��)���xV��;�7�䷑\܏%51������̾����/O(�!� �6�Tz���'��(��&3�>�#v?�?��Z@�����8OZt��xp��ܗO���M�1 Aܢ�k�U�"��#�4�/X.�ɵ�'���Y��L�Op��P����%k���s��@&äCE��'V"f��0[T��K�b"P�i;I�����XHT{�i��z�����lu�e��"���C&ۯ-L��y7ZwX��cXlxVHYEB     400     130N�ԅ��h�\I{���_U��)�z�N!EhK%�+�ES��0o�;����yt^���0,(�ी��MA6��!r��-(�[����g��s��l�3���6jùc�Z�^���}w��k�id#�1��)��7�Y����p�ɓ���w��{Wfk�ٙ�x!���R��u�b������ �����&��.�|�����~;�
i��)4\��>�^L�,�.�3��qoT6�5�&;+�s�)��		hG�t��#�J�@�b��K��k��G��D��OAS/j^�A^?�e,4j���S��XlxVHYEB     400     1001='���<�U��^��9��������*H[�7ZNw.nXX����@c��Id��@5����C�d�[;�\�6@�N^�����b�H�:�>uё�I��op���@i7�h_�[0$t�-�z �
<=%o�-s�бk�W�R#���-��3�~��&$�\An�.�f߈)��3f́�v��8�񞧭ζ��5\�/{*Rkn�����	3��Lc��}.���ǖ���Ci�?��;�PjK+XlxVHYEB     400      f0S��K����x�pF�������榙�:n垵�\a��x޷h�g�����43�_	�������.�`}L���?�����}&A��Q�������o����i?C���W_���������B����yv�W$�z�cZ+;N�#݈���;��3�W���Z�1ш7�����g������͐cr|�lZǬ�mi�Iq�-I"qF@l�0�����Yc�c  �SAǒ�WK��Z^XlxVHYEB     400     140�Y-���!�G]�l/����n@�d����o(}O��vH���LP�M2�n�ج��b��a���TiH3����w�U�*e�*u�kp=W9>�Q�$���#N�1��B�\�l1�YL
�9?�C
��Z�SǤ'Kߘ���N�=5���{J�U�|��x��^���RȻQ�m�x�>�4���{R\ޮv�,L;}�(bڍ��6�W�t$f�7�� C5�@B��)_}���i�	��J�/p�S��2�$&6"Z��|3�EB}a]�� �~pqq8����aK0���LF�6��d�J��Y��0y"�/��/XlxVHYEB     400     150��q�C��q0X������_���1-��O�&�%���k��y�0y)�K��x����Iz�����l����6^��V���i�l�7Q�/Z⼡�����*=�<5��N�[�Ă�?8���o���Qb[U�HiZ
�+��\�!�A���vg��(2T��A���^����\sH�$����f�C
�s��?^ [��C���wΞ�՝v��GA���*X�og�R�1/�{�+M��L�&ߎr<r)�k A�MF �H�|#���j=D��r���e}�:�h&N�r�7*�6�l��_�d��Ǟ/��}Հ�.4<��������KXlxVHYEB     400     170�_�$�m�y`"A ����qPT�ty���HQ
��<� �[�5�V(�!�-�뀩y�������^�q:��HS0D�J�}$�u�4��a�~���һ&���>�$��%������̍G1uE�]$�/n����S�������ǚ&���B4�;�wh��j`����i�y�I^��Z�`�9�_��޴	4G*�^���wF�4��#��w{,���;}P}ƚ.���[s�^o�:8�qnB��F�P�1��,��V��;D�����dr�w�F��)��4S�˃K5��d�z�5�:g�t�{.�Vf��ͥnǯ+�5{R����<l�����Sr�N>t��k��XlxVHYEB     400     160��f��[oQ�WU��r��h3>b�Zс)I�,s$:�Ό_�U���(u#4�Sk�Z5^���$���yxH�A��:��4bLg�����e@y�kإTK��}$�5ze�X�"������4=�ɶֳ�OAd\��D1\=����>vQ�%"����6���4��$P�%��w$I1�?��z�}4:�g����ȅ_=9�R܊`���E�3�d���a��4�̛FV��U����ύO��o���\�rĦ%��]1��s�py��'�O�`%���.��[Eں�'���k��h`�K�Փ�
�*���b�2L)w�#�I���C"nXG��	���.�lݕ=���6)�XlxVHYEB     400     180�C���4,��"e�֟>f�^xX2mA�x�2��ݽ0ӛo�U7��-��K�����Հ%����n��4�N��ҫ��m�ƇO<�牸�U�$����9v\N~ÜK\�ACO�e}���š/�YG;�w�H��i�}( ��$���TvJ/�L�Q��ź��������o�� Ι=�H�f�[c�F��S&�%�8	Uo�m?J�co������"��fF���Sa�Kvuʛtϑ� �9���K�5���n�}�c����<��ﶽ<̟��Of��{-�q;e}h��N-Z�V��6�_\M�7�O9>���+b)�~��6���[���v���FPAM!���O_!�vP���|�����FXlxVHYEB     400     100�P�Aعa�ߨ����g���2��p�!��I��4��&��MV��;��e���Tv���r�3�!�/�K$�'QF���kDq�� >�zE���=p�&�͵B"qC[Q��Y5E)�4�i���l���y�������쏥<�� ��h���j�N+�w�t��#�'�� 9��6�0�4:�J��
#o���D���Z;b����o� Lq��hO ��}�ϴ"G5,Y��eab�@�Y.�:��k.�.��f[���?XlxVHYEB     400     160�`Oh�k"/X�ff���m����e�W�Rz��/Y���Ry-Y��<'B� >~�&��"d�g�w��u$N]���]��O-�	��d�Of/�M&2�EPMbj��#��^�Ыc�9�Ҳ�d��as�-z�/�	:N/.Qs���+e����t �"��h[���F고p����+�sk�*  e6��@�����mr7�j�5�|{8�����\j!�N��JU������J%�i��z��pۑ�w�p�E�@�w4pq�ϓ1�1����ڎ�8E�,1�ܜ\��PcH&�?%�=��1k�� @��Qرv�.�.�w�a�4��^g@v(5��W����&�p�B-fD�	XlxVHYEB     400     160�����E%�O��]��+�d�B��V|mbWz��J�u��Jb|���Ư��w1I�-�L�9,q���]\�i���$��]��i��`�����d !�Vja�܇a�`���E���������)������i��D�b�c�خ֢^f�;m�SG_�ɲ��/^]�h����f���u@cCSe���<��[�s>���xG�`���0H�ouW���B ��{(�@-����y�(|SF!n�~��m���i�ع���������$��+ٲ㆟3���]w�e��.)�(�7;IkO"M;�4P�=��}qf����CIh�E����pV�F*���Í^�M-/G��bXlxVHYEB     400     140��!������p˫�����N��r��B�L�\�pģ�s�Z�Lm��P%� ����P�'�!�G�GO���>����ܦM征\S�݅4�솵-A��]�vKZY{
K �,Ղh�S����0�V��,jB�:Hp�)z��<����
�ON��0�!\��p�פu��с����j�&1��w���.��ʑ5}.2ũ(�9J��O�[0�D��g�| (�����' �"z��(��KUˇ�D��xp��v�`�@�k�#.FX�{��!+���*Z}�S�����˓�d�>� L�J���G��XlxVHYEB     400     180O/����6�Uݡ~�����`� �*�~���C`�{(L�A����w��E��lf@u@�ݝW5��h�����DH��*9��@k1%? ��[E��u��Hl�3�6�l0
³�5�.Hi�~qЄ�}�*dz���.�"{���7���|E?<�+v�s�P�$�kqT�!�����f��z�F��tA��O��6U�o'�`Y �N�Jn�h�|b/�m��`�<8*I�T6a�I���8Nm}��k@�\�!x�����֒LWڀ�����C�h6?�N�i��	Q�؏&����#������ �����g�{�C0�7���&'8ʫ��ܛ_�z��:/*=�,�=�pU���&���v��be?|	��t�W��V-3�rXlxVHYEB     400     140�9�*�EQ����/�B��:1����f`�JZX�y%1���	K��]Li��3��R�'*lϴ�#3J��
x�����X�3��e�0���zd3�(�'=Xi�,4�Y��5́T;g��5���u,�v~�hR���Q�A?�,3z�ӲJ6)��H��f���'8_n�Vَ�֖o�yǾ�%xx�/Z�!����\Xq*g�SY��t��%,�S���S���"3/��Y9Tp�S4�/��¯QBG��ĥIMLK0cv�.��&��jܱDכw[��	 N��p��Ӗvs��+R��~|��
������*���&3�XlxVHYEB     400     140xzB�M,Z���pw�1[m��WE�^�i�I��zO��o�Z-ٝ�<p�3�ܫ6����f�%�8B �\]�WC�OG��¢�jT�\$C�g/���'̝al̢yVC�����d��&1S%�~�u��,q�!,Bm�
�-x�7��n�c��x ���i�u�9h���g��8����2j+&�*V��w%`�ݑ[1\y}��,�?����!��::LT�?z�y�&Q�I}����[OS�a^���e3O*�^����i��^�TW:��Z�&+B`yș0�?b�4?�Հ��>oԀ�2���IUv��q�fƘ����V8��@R��XlxVHYEB     400     1308U�6R1��:���X���\�`滎N��o�9�3�'��y��Q�nK8���důUY��Vk*��dB��ǽ�=H�}}��~�Ko*�?پ]����$J.����@' ����T_e��f��g��#��T2쇍(mn����8Z��I'w��.�P�]�">�~gw�p���/���{�[����9bO�L8�O�Ǌ	{C#����-]N�B��'���D�B�-��Kc���x�F���{kZ���l[d�<sb�����!��p�3�&��`J�)@H-8��� �0Ӷ^����*����{7=:��ZXlxVHYEB     400     170��"�����5�@_P������Qq0��I~��sP�q������-��&=YV˥�Z��|Gos9�pj4�$&G���ˍ�m��Y*k��"U_N�Ȉ�84����Bپ��քO�s��Z�hyǾ�J�c6dI�k���88m;�9�p�/*f5{&m=�8�=�m��P�.�J����auX����@�h������v�u4�-� Ό%��t<��Ke��*F^�@���.��8��E��}�(�sE�t�3�`8�A�%���}y��Q�7��KuJ@c4�.lF9,��̫�)*S4#R����f䝜�����ރvҿ�{Df����]^�L�4-� $G �`j>T�d2�45o���]XlxVHYEB     400     170o�7�Vw�?�yP����~��0F�����S�ѓZ'_.��_�љE��v�$���}"_B	J=D5�3�v��E��@Gm�u	N������c0��R�QݟOjk9���	s_K�<�ԠL��� ���
'��KxBK��J�(z��,c7\���.�l:��8d6|�w�`'���>nF����iN�_��-��  j�K����%n��^2vۮ����1�Y�W(��s�6D���>�t,���Z�|��cީ�:԰�9�3:Ы�3 �/����H�����.��4V	{�vbH�YQMP�?ucr����/avx�J%ɓ/��祴�۳ٍ�;��
q�PD��ͬԐK�{�}*���k���Ž^��7�XlxVHYEB     400     190/�z����F���c�<:����~2�s�� ��$v�l�<D�0��c�aMB���d��#詐�������R�kGՇ�ѽ(_��4: 03���)c�\~���{�+��W��/t��8-~^v-�XΗ�"�@�2��A\��}9��h	�o�>���|� �v1�,[L�q��b�i)����I?��o�R��|���[LK�}������\���J`��^5!�#0�h�}��nï.~��)�*���ق��s��5��κ?<� B�a�1 ��lV���3;�p�+��T4+	ףrm{]�}��M	m�*�M�BjS,j��X���3��p�M�� �#m�t�z5w��uϔu�t���V�<>J|���e�,����q���8�k�XlxVHYEB     400     150�H���)���H.��Y��Ռ?�����fk(�t7��$�����j��8��,�gxCn�٤�/����^�v>��c�hn#�*�<�A��$qǘRE�M�|��s�g��9�\{)�5�U�8���X��q����L�`���]�R�a�|�R�>��MCE�����+3�9��<�1�6�Cn�p �Q�SZe�cC�k�d讋訾6�ؙꄶ��s�2�I��N �/�<�]�Y���0�E_r�ƪ�4���X)�L2L�ד�:7�8�:b{���ZW�ՙo��?�?��!��ȳ�`|m��z�p|��Z�%N8V�V]��6�?��f����XlxVHYEB     400     150�1�7	�@�O�G��;�n�'Vs�����C{��.��*6(%JN^U��`��<�nB�걻ZßZ�&o[����c>a��}gH�E]q��A������D-I��O�M7�4Q�S���P$|�ܻ$�+f�`�1vGK�m/t�a�b��{r&��%H h �|�%����xnLT���/����Ў8^3�����c����iv.�fƙ��i	�"H�{�����ņFO��^y ����E�y�X6�|
�2Ź������e:�G��[���J�%��N2���-v$�~/���`gF�Y��_�"�f|�i�D\�Ma�#��Og!��XlxVHYEB     400     160�d��#3E2ub$�c���ʩ<`��܊���q�k؄L�u�^�XB�A���\�Ձ����zC�~��c��3�Ǝpt@qFd����(���F~��^��r�=�g ��}��^x��66��/�3�Q��@A��P֏P3�����(o�2�&�$I}p��~[[<*��vϴj�c&'Ѭ?Q��ܒ�b�<�~�Id�o�/G��7#'�4�{	�~},Dt�#Q��T ����g�i_�'&���-��e��M�nٸX���9��Y�xWd�����IpMlV��e��T��d��8��ƞ+�T�DJ*�x������L!��(�A��b�����$E�XlxVHYEB     400     140H@�)��&�7���G}�H�GZ�\�7�8:��$Q�c���A����[0x�{s ���+��
^�&� �ɲ~\���^d��B�rh�W��&<��1�0����-����y����X����<|c�p��R������`ٳ�O�«J^����D��{>ƃ�P������]�cS J���w|%��o��X:�\��nr�in\�����7IS�^yOW#x.�1�l�dMJ6�o��>=�R�H��z�2ˤ����x����*��Ȏ`[D����$n��b��%/W;5;�uP��6sY1�9D�CE�y+�XlxVHYEB     400     170({���1Ίqx����,�O��=��:�j��Fٚ
/���a���b�C�?]#+w� twZTg����F��ܵR��Z��[���_��|�� ��m>��*?|��	}�9J�~b�}�B�(�r�Ҏ#��9T}�ϓnN�Q:�B���/#D�(�,b�Y&5��k��[�h�?�i7�2�p��u����@�X����"��
,i�vM�#�Z�	��ep�O
�i�<I�4:�|�2�B����-Z9B���*#���Xr���CGUjn"ʉ*�L���_�TpoC�DZ�y@	M��g(�Q���PH�Cs��������R�'�t�<�:�]G������x%��'�W�|����a� �F�A��XlxVHYEB     400     150�F������,T*4�)d)H��3
Ęt3]�֯�,Os��J O�o�q��,��ԽŚ��>V֥��{-e��������~<O���X�f�*��!��ЏO6�x�i�O$� ���.�s_
P>؂��&2�7Z�%�dvڀ��'�1g���[�9��H{�G��}��m���[K#u\��?z�7t\^co�v�г��}�Ӷ|	�r*L�y_��7����I+e�����ιᤂ�CC� �9��>_7��tƍ��W�_h���]�zЍ�5P�C�g�&��!,�8���{�@��鄜�_��|o���29dv^׺���>���X�z;<P}�B+��XlxVHYEB     400     110B�D��/䱐G�ŷ�t�s��>ƶ�e�"E5a�_{�ݾ�mJ�YuJYփ�#�R��W��2��1�G6��ٕ�"bS����ز�'�)�M�_)�y�hG�-fG��Í"��,c�Y��CTe�uf]�hq��T�ĥ��::��
(�	�G�nH�cFtP��$z�
���U�'\����Z|z���g^�3r��8��(P1�c����k%�q��x�"=��"�܃)f$A����e|�k�i��c<>�z4a-��:$a!���2�rXlxVHYEB     400     150Ĺ^r����ӕ���32b�S�I�Fb��Ӝ��ÙA4/*��5�I�D75��D]N	��"&-����'��	T���0�йf��AL�񆙋i���SƘ���$�~|��!e��>�OطP���ժV^��lχ�nx {A�G�
�	����Z)V�:��t�dk|���`
��Mޓ�*P�u��CP�!)������X&��A[9ؕa�G�.o�4J�Z؎��)jt��*��ӗ�M��GNV�](��M��̸��ݎ��Gd���w��¡�\�ȁ(~����{�Cv���VB6}nL��o��0qݟ��,����oa_]Ruyr�r���yXlxVHYEB     400     1a0��`�/&�zo9.�w��mW�3� �3�>s8�5	^��	m�>
��z[2�g��F���=�Z�'nL��K������%m�~�<�� �l+үz��Ѭ��t1���ш~�L�Y������aoz�4м����&�_Ol-C/��������o)n����}߱CdK�]�����{�t���=*�rƛ7�L)���&�jQ��*K;��a_���,0V;�r��E��r��kp5��ҘƏ~2C���qi��Kď��6�p;8l�Z�>�� 9БvZ���A�%�KQ`^���H`=Z鑳��F�7E˪� ��s�-[.�f#�|��4f-�4g��������R�[��e�Vf�]߁�n�h>M�ڠ�#gC����w1�Э���m�Bw�ǈþ#�o<�.�)�XlxVHYEB     400     130���"���u��L���k�d�F���7!�͒�ʁӭ� F�=`BQSǕ�?�+Ҳ
HWZ'[~��b0�1���n�lxN�)�AE�C<��_� �F���:v��뷣���@,ѓ�%t�p�i=��[ծ�G�E�n�����v�|Y�\���'�=�k]n�'�`��<A�{�k�*��������sH{�8CiVwO+��B�ñ�l$�� ^���S�u�n#����R.�':�Ύ7<��>�e/����X�1�b1�z�?[ZQ���(���X\_�L	��W�밻��*����vXlxVHYEB     400     120�8�)�Y0:_�+!.�Le��w���Ѥ�Kc�n��3�-:x�V�T�:�ڢi�S�^�`�ѵ��m�!����+<�t�.g[=kU���U�U��c̺4�T�(��X�p+�< �K;~�z\5A�l!���_�g���O�L�`Ot:�{� 6%�-��f�,1�2����b �UJ#+�Q'���soL����zr�J*�uv��Ꜩ4d�!�	����z�^�����,��<�#+�d$W��>r0;vE�P>�mS�� �o(Aɮ��8idjZ��TZ��@-��<){XlxVHYEB     400     170����f�r�c�FADZ/��y�z��_��!�0$v��b��?ӊ��U%�w{u�2����\���E�`�xG[�v���F�MOC�{�H�j6�m:��)Q���>��^Jw��jÅ۠K�Z��a����ӽ�� MQ���:��B��_h]�Mb Q���z]�9�3�����Bk"�� 6�Qɘ�1�;��K/�kf�C%�U�*{	�V��f��5��4�'`_3ә�^�mZ�4����2�CQ�<�ޢ�zb��M'�<��t0�?���F�ݓ"W�4�������·F�,�I;�B���Zpq�rj���p�3%p���?g�V�j}8ډ�|(c�� ���|̊rwT�����d���Fe���!W�z�V�ji� V9�yXlxVHYEB     400     160� �k�'2��KԵ�\�"������j�psҽ�.�<�/F���HD�Ê��$?�\p�QGL��A�@ˆ^}�"�,*S�L�E��{Й����%$p����'��,���YUo��p�|��9f���C�ƌG͒�9MuaP�.�.��.��`�N��,�|k��/e�� ��{�A�xZA��\��2g��~�@~6&����"6���F�ơduB���Q�ܕ�?[�V�E|X>XP��kҒ�D��@��T^�ț�����5��pp�%�%�=Z"�5k2c�����?/(��@f6��Cɉ��D�D)R�$ln.�jyy���oZ].�͋��I��<��O�!d^�XlxVHYEB     206      e0�e��`6�с2�Z@�Cծ�}U~��j+�7e��� ���0;C��Z�s�5}�[SB�i��IB�aDAl�䮉Z�IB_�`�I[K���/��PPmP���A�>(L7P�y��q���A_�mrT2�?Ed��!��e20�=�{�<�{�ж���H��SH]F
�G-V)L�<��@7t"J�}��?�IY6)БMۆ���ў�R
��I�f��#mdF��Mgo��� 