XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����}�e�$�Bo������D���O9*(����4�7����y����&����4�J��Zq�9��Y�` %�ì.�9z%8f9�f����p9���2�:h�T5L:U1]iQp:D���y]o�0�{��dpRJՁ��"�󤲹1,7����h�n�E�ƣy�Cv�}�{B|�);R�E���$���w��_d]/-�ۡ��Q�ŧ�*�&-|l9����a'6:�p)ۯ�����p�u������2��������nz����n><{#��&��-��o��Q������<��6"%X���T1�2�`�츗-���j�m���?|���]��*Rڜ�2�= ]����� _�G˩ai�rɡ^��;�B6�;�,lѦ}>}����;�$�1?ƭn�:�B��/�p��Щx�� �ïnX1�}������Y�M�3t�Q%���p��D����I�(yQ�҅(��fOa�W�c�Y,0�N�1d"��~��dOC��-��vT!�+��l��o�ȁ�<e��8���S���Cz���t��o:X�i���%�|�Y*K4<�N��hC�	$���lY�L���h��}�$�|C��<��k��wx:W �H�&�8������ҤhR�G/��ғx�����*a�K(���<���S[��
\l"�>��u�n썵$�M����)��s7'�(�O��އDZ���#��2<��k�/!&E��ܨ̝ǀ����R���<fe1hGH�XlxVHYEB     400     1e0�P��Z� ��Ȁ�^]��Q?�!�C�jS`�L��$��a$8�5�ꅹ3�y�k�����0��Y��g��d�Y�>5���b�N�h��{s�X��8�.�Z��B�L1��|A(�m!n
Q~�����4SI�����7������hn�f�J>G�u=���L��?mz|B��A��< �anr�u���j�D������
"����D-���G iֵ��R:�С���>\]:|�m��V�\?<Y)"V��һ� ��?mc6.����Je�>f�9�)��+o�)���\,mɅma��}�h�*����y�Av�B�tX����^�GSC7�I
b�'>�ll�{�7�i�Cy�o�K�-^����6�`�90k]��P����O��Rg�����o���U��du��o���t��u;��R�L��b	Q~�oܼBV��d�!�k����kz�z��Q�w��~1�ؙ�B�%�=C@��XlxVHYEB     400     1a0w9D85��9�*9���aU��G:�7!��O�S�"��10�;�2��8m�	�Q���E�n�ؤ�,U��p�λ�6G����0G.G�L�
T�:݊`�ɵ�'��=3���p%�s�B���
�Pc��SP��8�D�R:�N %#8�zX��ݍ7�oT����[�z�	�6{������IN?t�˭dMF����9��T�2sN���l���.�0�T�q��`N{;���A9�JHq(^!m��0�E��L�0e+	m��_<��@ 뵾������/�)�V�^5A����k��`>�jHa�U��V8 ;d��I�x��.����R�8{ָ� �o��|��0�Z��o#~��A%
��h�/k]����e6�U�ܮ�~�t#}Pfb�G���9�<�f��g��XlxVHYEB     400     130�ND���(�p%e��. c|�����$�5�[���@���RD�d�\�����V��dN��C�����.�1�=)����I@���L��{��h�<>��r3VѼ���E�XB
���*8�����5[���~Z�ߕ>@���>��"Y*b�!#���i.��Cg?��Ў��\z����Z�R��������л�C�_�����w��SZW$�5䬎Q�+M�؛8MP�-��g�����ꌊ���]�%$�����o{?�T"��誝vU��׊�A+wXW�W�_�xa��a݊~�XlxVHYEB     400     150 �t����=Ƒ�"��oB�/��	3g��6gyH�R�U_�$RU��s"��;�j�*]p���8���:��H#+ٹ�_2M9�g)�n{l�^	�~*��3$C}^������ a�7�ܥ�;>c|_���9/KU�V�qB�n�G��V�	ϐu7N�D��&@lp�ާwH��J
X]b�4j��#-8v! �ܧb�n�Rf�=7�\B��L��#�xX �.���9�͜�v�)z��2�ڹs�G�+⥰��xw�u��Ŀn��;(#���,N�G�Ԟ�:�ծD q�����Jz���~/[e��;<G�����m��KT^
�]Sr_G�XlxVHYEB     400     1a0��e���(�f�����(������:�����M��"#��iv�C^���|6"��S=S�X���О�Wβ���l��Ps�,2B1��:�m�^�����w��lA�Kq��F���2�՝R�NK4���\�.�[�d��~���zS��R�ȏ��ZP9�"����Hn0���U�"�X��{���d���q"\�(�ٯ�(D7�9T`�E1*O$>���qZ�d�卋����c�R��l��뫤����)$�qy0�KA���5ɋ͢�D7�j(Ko���xN���S][R���]��&���Lx��5c�_��r���hRK��mm�����BJ��D�����Eɳ��(c�j�P�I�G���B֑���|'�2W�/�x&�X���9����k��#����LުbI=�� XlxVHYEB     400     180[ӵ+���KU�'���Ƶ��u�F�Lccv&Kz��՟���Ӻ5ѐ�ϵ��#�s��*�"u;�9HK�r�nD�h� @{�*�h����������V`a����œc �A�`���*n{P�i%H���Fj�c�!�Ҩ7,�O��愆�;��f���'��E;�R�܍&�6|BaJ;g%��Q-�[7�q7B ��E�*�P(�h�&/�����B͡��󋥔Z�^8�&���*.���C+�1���Y���7,��f��w��@�T䅥2�F�Rq�:iI3Ij��	�X���f���o'��c�cF@dJc����ӱ��'��d�#�D�8�o�h�?���z�]������ &sN�hX�h�_�Qyr��;WXlxVHYEB     3a0     170��O���$K�;�=W�#`Qt �f,�����5�H^�#E�Y}���9��t�=�`��ԢYfC|Z�%G��Hk�js�1ڢ�7��fi31ku��3���f��/ⷿw�rv�:RIq�(H����S~��p�����(��u�t�t{�1V�#��R)�r�M��K�$��]��rJ���T>�o>|7������u��yX��:�1��>p^��v�����:r�>w��f�S��[�*�v�ub�f�uX����[;��U��Hhڶ#��b�$mhf��.�B)ģ���Hwc&l�#k7�^e'ov�\_�c��ܒ�M�+���b������)�as�BQѺ���N�K�}�fca�g�