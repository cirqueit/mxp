��/  ����W83|�yx����C`�sO0��b�D�u����4���3[L�8�V���{ٹ���#7[8x�C9���U� ѱ,��A�ׄ�n-�H��pN��qw|�0X���ږ�sdX�*
���p-��S�����E]֟�3���4DO�l�����<VF��B�k��o�*D������b
/�G�d�}fW:GW�h6��$6^W���z�`W��Y0d#�G'8�y����	��{~�W�C�������^��z����O�:*4�$3��vƧ9=���Vù���n����atu���V,Mr���Ͼ���ӡ�[ȁ.d�0�JV}$�����MS���I4��9w1� ��U��ՌMԤ�Z�F��øǼ�bЬ� ~J񮅴�ў��v�z�o����G����)W�SOw��\���,u��W���'w�+i`��:�)������|<��cZ�=<{b��N� !��~@��]?�R!��Y��l9���.|-�6Ng��`е_����.o@�axA46Ӧ�Ҏy,�um:�>�m<e�h��ʎ���g����Toy\!J����f�."	8�
���wd�13A�+��.��$gd��5�����0v�Y�n�y�Iw���B.m�WcTJY�h	��5Q)+��?79��Ⱥ��s Ė���0k��7�":
�6%�.T���F��"6�G���ÚN	&Ԁ�b��Pۋ2Y23))��e�Z��.	�?ʗ���,��=A�=0�jlfF�!	�,U�������~	�iY�#~�Y��h��ױ�h���; ����:9��9��Љ��y$$��1Q�c�\iSn���S�7�(dRm�Ҡ_��'���^Bv��Q�s����vn3n�ɹfI���YY����$b�P�c��0ׇ=��NW!�!�Ĉ,����ڵUb�ۺ���J��h�E��9���u���=:�wqG��F$��|�a�^��� ��T�,��<��?:�]�J��� d˙�`%�,���۱�0هsLM(:9����>zM	���*��j/DFntO~/��Q<�$dkT����bP�Ϯ��'2�&�E��W�&��LAz�2��1���u���I|�L1ac���eB�yW�?�6�83�����{A�����6�]�<�������D�J�m�R��qy��+�`�5m�G��2ѵ��qu��6ŧ��M*����c��^��[�>�2�"��E�0,ҹ����)��]~U��	��<x�!/��&݇���@��Q�u��
�7�5��ϱ��sتS�f,J[��	���S��OM��S�+��:ڀ��m��PB�QA� ���|u��@��;��P�=ywp�r��L)��Pe�~�>~!�`�8崁�s,9,涆|XɒQE�1�c�nrs`RT����c���lb�+6
D��1nԑ�7ӷ-ESNĲت��i���	�!��[��=�&����5��w�k�tĆ%���z\��}��>fo���u�����_�)K/��ϱ�s�[̚�{��0vy�%{|�� R�u���q'�^4�����x��3��l���5�z\���� ������w�t��ْ��&A%Ƚ�;#��I;S޴��S�_U>�ұW��b��
�B�"���1M�6z�B��>p���!�V����P05U�~�h�^(0QXI7�|��0=�ȚoA/����%٥���P�{�ߣh�G��A�}�HLm/z)J��un&(m�N����X��S�#��]�[Ǝ�}��?������t��{ P���!uR��r���:�L�����f������	u�*a�8�5�U��!C�7N��kG~e��qI\Zﹱn�\dPO�Q�8��C��6����3~r��\����'���ĝ�DY�Y8�C��NMo��W�N�ȋ}L+bX��oc��桤(�ȹ��Ժ��HR���	�b.�I�*e�:[B7t�=����ބ�ŹtT�|lQ́���N�)4N���q�ud���Mx�|��x�s�����z�EΜ��
��9�o�Ka��Y�RD���KX1%�4����J���jY��IC�|5,T|�Y��	���������wZ�Bt��|�m��A��VU��e�U�|N���o�'�C�!lI5�6U���>O�so���i޿K��9/�t�\�Ai.��>DK��ɕτ9�/��
��qG	<-Oy��i���T �&LS���J��]�p��fV
����]���y�Qb��ɰ&B���%҅�ŝG��������hў����{� J�>[y�j<�!�7�p�B΄��|j@��ĵŝ�Ʌ(�,Hm�W�m�p���>���Up�?���Hƍ`n���tLC�H&���7��q�dP,��kS.���^����a]�ՑW|�8_%�T�k�2|F���Fkv�����.��ݚ@��/n��6��j@I�r��ӑ<Pjo\��Dy?Z�R���07	��d��FU�PR�jr_�)�Ow�z٢�Z�Z荊v���n��=Ƞ�4g�8P�n.]�ػ�Œ��E@����y�	��SsF3Q���T*BS6T��R�m1�����e*G�T�D�"��L�Ib������;�7G�"�X�K�5�ω)�d����� ���4.�{�>x���)�IO��ZFv&(�����������i6�S���%��I,1G�����������-�?XC�%����n���tZlI">���S;~��uc���N�ˍ}���$�"5��iֽ�1���eI'{q�Y��K��)>�%��a�t��d���K�*��g�e�?�<�;�n�h��"�~�� X����5�v�=p�.Ћ�[Vd#�9CVPfᛆ�zT���TLW�����1g�$�zzV�����_�b�fJ��f9^��Ô�����N�	-c���%��F�E��!��>_�򀯈*�34%�, �z�M���ß^�+�	p�/	+?�G��o�1o`�Su�9�?�aF��H4^!��jk8���T��
�^�gLr�[��'�ݲ�T&Dky���W�W�忣��y�N���8� ������������J0�[^��w�vꅓn����t�%w��k��,VУִ��_��x��ܭ��ῶF�D�ꍨ@J��|"Bb,��l� d��J씸�XN	 ����\?�k������.O5i��
&OBF1��~x_��V����L`�0b�լs��w�V��i��w�w�}�#[!kg���;Ҝ���U�1�C���&M�w��Hd��Py��:�Ag�����-uG��qf<u���Λܟ����*dg��{X�9݂�BІ���ۣt��0��P��L���'��3*�pK��$���!����\�Ihg�h�\n��0�n"��5S���Ni��q6}�͕*i5z
/-]k�w^(�V�n���:�	~��$��+/M��8Q������jS;�v�����N��N�!9X.C���Ʉ8[���(w�gc���=`be"���&!�q�Ri�9%=oD,D���/��/9J
���9��[2��^�Py-wN�+��pO�o
CY���h���#2���N�v􆢸�T�smB�5����d
��3c��~Tu%pwQ��{�ݹtn�"�h �W��/Px�#��PP�[��� ��Ĉ���V�P�0�9Ğ6����s�@�e�Z0��ml3^u`?n���,�iz��\.!nZ>�ʻBU�F�.��E������L��j�ԃ9z"A�Q�,��<>>��2�D��^<'�Lʒ0gG�>>���;�XK@D�B�`q�W�����B���Ji4��A���3�N�lX�C�QJ5!1`��~��a���g������o/ꕺ0>f1���U�m\:�M������t(0�,r�|�Jwt�u� �m��S�ۏf�b:�i����m����lCI� �ȃ[��Fd�yNc�>�*_<��WXǛ�>�-g6$f0D��:�H�Cx��S�XgCM�O�R)��z�����HQ?
�Z
Qx�*��f�g���H'�#��-. ���jx3����?��8*P �TŇ�z*��:|0\�˴ˣ��-UdD�;���z�[��_Jv<�a��p��j���ݨ.!(�$p�G��d��a��-���MC�bw&q;rA�s�4�DͺC��!��Z����MI(br�K��JVY5)[휹�?� �Uv����pk�Q�-T\��i���s�m^1��ҧ���)�&�u�]����}�$�d���w��eZ�[,���V�'E��K@���G_8����i¿h*�t`�*�^B��s&f�U����M��c�UB[�b^|��+1<�N��G`0"y�߳(?<�.2��	�H��$<�OQ>mwě�xun�&$�A���?ZG�poE��C�EA��y�w�I�+��r��(�b�b�q��2!q����J^��l[�	��)4��2M�=窰�O��)j��=�r��YL��#��W� ���'4��a�I�I�	lׯ]� K#��R�5�gڴ�"��q;I����<Bp<6W5���?01j��c�4����I��dfD���K8ٔY[�PY_c����!�}�a���2*�����>F���~.��؈J=����+5�Hb�ԋ���C�7N��e)�#C�4?��i2�������|�X�������ԫ��%S�)�(�<"
��E��r�BlMnK��p��Lݭ��a��3��v�]/�����t��c��Ï��5V�J�[E������}��hB�g�2��p�E���@��tlT%\ZʐY<�#���l�O?E��G�7���(������ҥ�$L�+���<:�ٔ��3!��%�a�	.m����URI~�\JsI�Vw�^E�1�QǊ/��ǫL(A�,�}&���D7h?=�4�6X��:j�E��2xN�9Ik0��	C>�֫�<w!�)v1�c�����k��{Up*�O'�̨�hbXozjK�Q��9]d��w��S>='��P��<;?t;P&gf̀��T��{��u��P�<5��ms�)�lIˉ�"�~��]�ff�sFT�_��g�̛�? X��Ӎ��OhB&���X��~A}l��x��t�݆0n�m��=�>P��N�����	�wA��`�xJ��vJ��B���˰����ˢ��xC��Ȥ�|EZg�ŧ���n[�P�o�jp�뜳��9�� I-��8�&,���e8��~[���������.���ꪝ�I2��]uZ;j#�Z��Q_.6[��{�����Q,oU/�ǃ�v�G� �Z� UAz]-˯����>s��EW<�gh���>.6����XF�Z9bWa�D���kr���H�늶�m�8����̈́��iBiůyY�!����l�R���X�/���w������$��C�e�L���+_g|��,y� 4'ن8��V��?���lnD�g@`ř�� ���-hb:a*�Gm��/=瀅HJb��P�LCm�G�RQ����@�+#ϹH��I_��p�y���w�������1_)�M���� �4v��E��T����%)X��b�fH��lZ��ȹ�Jt��ac���ʵ�<D =ٟo��-�S��S�gpC��c�/���������ǲ�Q��5� X*c:������1�m�2���6Iwh���z�e՘^�s�V�x�WѾn�%9�k#؇��?�>m�-�ȳ%/�( ;��n+��t�Rq�{�y�e����L��\!���w���-R�a�g��j ���?P�&��>`p0k�/��T7�|�KA�u+,�6�����!t�F���5;���ܮPu�G���vv|P��5���ׅL_�W�g�Um��$�Q��f��O-d<2b2���/D"� �1���A1�*((`��u��X�ȩنH︸�׆�X	�|�Hs�`䦽ǂp4��D!�l�a�!/��9	�����<��i|{�Wb�[�goF�K�U�j��	��z�t@_U��^F��C�ݎ����S=ڃ��-��e��d.r��jTmV���ǻ����O줂�������1�:z_.�0���'�6��m)������� x�ؓe��j���TՂ����S��Tj��z�"�)�zwH|r�B����\~R��|TZ��"J%m�h054�b�k<_cA�#�w�S�W��4�(��;���$��n5C��1/Ggy<�rV4��(����59.S�*�8O������:����P�n+([�h��"�`g����'"�(C
�0��	���}���4�$����Ā!�9\n(����~W���?}��
g*tz����A@3W����Y�'_֟ �\�=]�fj��h/�(~��df����E���g���f�֋�l�o���6$!c��$�HH[���a�@���)�n$Im���9|���������(�͆~���X�V1�h��[!c��=�7$35�3��3�2ܛ:ﵝ�X7�Gz�>ƭ􉹼�9-o!�N���xbd~raݼ�"l�㲤 ����hԠw:����K[���ӝ1�1b�	`�ş�0��ǀGc��o�^D�w��qB'��A)�m��5w��;�90��M�=��n(�܇�њ��[&%�m<���,��(�OC2-Kf�}�;��$$D�+rֈд�N^�4���%15���\��!����"Q�ݜ��r]˯1Dm�0 '��=Ak��ȑ�>��:\I�q��V�^�6��k-ZV�?��ȶ����yry����̬M���[��k�?�o��=t�Q�|Sv�d�p����`#�!�Y� ���u7g�%�ʵܓ{x��+�l`�1�z��7r��:�6�v'�(X�nb0�#g!=���X�P4����w'8��(h�oK�mlFǧ�R�:�Jo�|=���8�S��A�Q�8bn��=��Z�8�ˎ�/-�1=�)X��S�t�NE,� �8	�����a���*�^K8*��m�/	�Uā@��>���k�e��?��Y�$���
X�,E�'�.���9�a⍮*��`�;i�[�&)�A���fXN*D�OG*����\J����(Sб\�/���m���89�ß��F.��c�PS[�v�F�i�e�+W�UCؾ��5/U.���PxM��#���	&��q�`���//���,H�:�?��*���ǅ��Űi1-��-h����=��.�pѥ�V�'�۵����~Es��?ئ�}ڞf�b��TNO��M�;�ͳB�,�Т}Q��y�^��$S��A�����#wTy����J�S�>4�u�o��-L4�f�tk�4��n���T͝*�۵3`��,�����b�# �ԣi��0)(:�C�D;�i,�'�9�N��n+1pX ���H���A�TC��o0�g�,-�D����#G���'�� ��4�G��d�o�I����ӵ�� �5����8j���	�U*��ˀh[���jz?����Z�@n�+���SʣvSã�Y���#V|���t�7r�EH�\Cl�忳'x�jJ�T]��`�|E�.e�k(�5�o���H)	�]����XF��n��;��ҧ�-f��;m�"���v�W����ƽ��́
������_Ó���2��F�Vl�u;��%MR�u�@��z�p-��z�)3�d>��G[��3@�'}ؖ܏���݄�骑-�����RI	�(}܁�������N�@�䒮-�b��jp랢>8X�< �������?L�Q�g�D��(n�L����~���#*�'e:�'J0�3u0B\��PA���QBMe�4ae�n��wׯ��w!Y]ӭ�A��X���Y�k�y��*��R��[�j�/�L���_"z��u|�����2�?�!&�F�o35ϋ��?w�Dd�O��k�:5�Z���?tTX�E�G����QX��#��H��m��f�ǳM�RCٌ6�f����D��y��l��۝�N�����d%k`��f_	X�*�Q����#����L�0�]b/"P�S����q�X�<�g,�cY�,�H���kG�0T)����-�[�NkH��КMj���)�A��<�K.g�_w;��n,(JzwXN�K�Z���؝"�3ֲ5㳒,��5������j����H�N�D�b���/���dN�T�����b��4�����������R9������g���D���GW�f=��D�i�њ��[�N@p�������-�C��I�y��30b�tM�̯�@!*p��m���D~c�����M,aďz��9��r����/�� l�6���L���+��r2?A������Қ�,p��y-.��k-���|y����w��69Hp�¸�k�@d�}]�t�%p_��2�qߏV��%*N������K�@6�m������$��B�����|�
"��5=x��M^'!�g�O>��b,<��{`�܌�]���N�53	U��":	��X)���l �wT���$��b�Z,����b'/<W͹�[�����s�Ged0�ψ���p�d�>������ ]��/D���FF��ïitI�#��v�t���b�4>q�Mc��;��.�|��ϭ�	%G�^=S��L=�t�h�x�`��a�o6[����y��r1���0�D�-o�^�������:�6ɬ��Y�dԾe9#O	 ���(*�'�����Pǆ�o��}�X����MPΉɆ�؞�*&4gAu	��~�8�ѡ?�f�m�����/��͸�W�x�/�&~��5T7<-Ejkϖ��&��*%Y�L3>���HӗW�+[�A�I�uV�Qի���F�Gzz�>?u�}A[���-����ҠS]k����1\��z�FZҦO��\�Ne�����hI��[8-ɗ=�J߂�fx�H�qߠ�������1}>�=ҸP��_�,�a��[6bMaDr�G2��X�=r}6�.S�&2��?ʩ�s=rx.e��|$�xq�y�o�K�x,maH���H˗s��b�H!�9��������1�Xt�8�ʑЮ�ЫR�U�&�-�n��&��o�8i݂��U�>�Ej
g Iq��(�O��L�D��d����ث���J-6�8�+�f�#h
fKXP�\uӚ����3�>� �i�R�v L�$�ju�D|q;����b�u�Q/���i��x��]�b*	�
c�e�m;O�<�f��wp��RD~���Kb���kS�n{��u)��/)m]���B*�hq�<%sc��-��v��]M��e�*�N� r���"�e�Di�tg8C4r�'F���j�%7l5XJ�~�u��zl�c����o~�+�-�+Q ����hs*���X��B��K���/)	�m�('z��PX^Y�f��uy��.k)�e����
��.v�|���5V������%���S��,K��Vׯ�=������ކ�}	�x��4
6�����;�e.#�W�:�f4V�i++\����X?m��>%%!�\T�.�=۬o��� �\�Bی�{���L_�]�$o���?�9�G �w�@�(1�G�>��(y{���	N�/Ax^?�azS��|4ޣK����1��
R&�JI�=7��=N˻
���ȹK<#�קC�Ǟ�'&i����jO�g�X��|%� �� ����5�T�j����5 _|�ڐm��<<TOX���)@vX2
���I4R�!��ľ0A��G6��'��Q�hG�~��+�.��M��ơ�8����T�tBUF�H�a��$��>#���Q`��&è�΀�� ����D�j�KF�m�*��%�dByГ�϶Yl��й�c�~�m�ldlg+Z�~�^�=����-����WNN"� 1O.G��8�
��(��ZL���G��>��3i�6?��W������v�
��i��� ���a��;0>%N�[�an9im����B���RQT�|�y�^%�- �#升|���N�A��c� �AL��n�!��乕���b[n�Y}��0�z� �p@��@	�濦�L�P_L;��$�L_ZU��+W%`קZ���0��/#���@�~='�Nvr��}P#Z7��:�miA���J"/`���LV��avRFa�k6��� ?0�$e@�(s����~����	�!��aܒ#�D��7������}�)K]�P��+ �QԆ>=�.��0���6�~�a�]y��H�<�H�;�:J��6xMO"���Fh����ĩ�1�ʅ�?�˦���"���p��ȉ r}s]h�qpQ��R��i@���(N(��	�^�_�Ɍn��Y�w����0G�0DW�	!	��uW(�t&vߵ�(*K��' Ւ��?N��j�䐍����:���+�`o��e�u���K�z8�@�$f�R���j_��%7���k|����e��'+˷�d<���r���^�U��� Bᕝ�Ƭ{ :�F�Ү\�sGļ�&7�|��O�O���_���O�S��D@5r�1Pj�o��*ay�A�Xt�~6`�eճ�U�ܪn�"C���L���3|%�v��öBk呍-��`���5���Ҳ���u�M�H�jI�T�"a��-\q>��4vcT�a�Ó~b�Z�|5�.���=q���N�|rj�{[�%����nC�1�|�x����Cb�Q��z&
)�������\�M�_�r��<*�og$��}�A�j�H�O��{Dd]ʄ%?d����	SC�C�B7�����N�w!W�V����¸$<`clJ-��n"�bM�LV,-���a`����dE�v�[l��,-;P�F,/��%�p�V���s4�a
;\��'�<C�p�o3�-�,�6�!�mAJ�c����*Pb:�:<08಼vm[�O������K�J��j��no�Y��o�.���)�Oi��,�Nް�oL��*JӞYkYꛊ����g��ĭEV=�d��;��3��aP�ϥ�����Mw	WYA�]oM�lK����a ��_n�i�X��h_2�b1h�����Vi���ȩ��(X�u:��4���
�;�n��ϔ���@���#����S@G�"%<#���+���z[Y�t�h���ʼL��Y�G�9}v���[�_Ƣ�%��:@� (&��nt��E���g�Q�}6��@N���O��{sG�	O����O��0#���y�R�(r�'�=�	{�����p��eɉ���V�W���o�u�q��zj;�?�>�U���v�O�x�,�0�Kb��Rjw{B��-]��ˍ5&��|(ۓ����)\�0��Ll�*�.�.�}�/�� ��-u`�-��40�^?�����[[�iМ�=�s�g�8�"�~���O��ؼQ�tI��w{jך����h<�k�h�9-�<8����<�B�$��l���H�̿ڗ�����&���RQ�16k�o~��#�Q?��R�^���������,�t�����,�o8׷#��_�t� ���u�F��rQev� �Nr�1o�N�?��XC�n\��^�9�$�?�9r�-�M
+Z��ԭ�5�d  ��?����R���bɤ巯Vd�zo�rN��N�u^��qa�ſ(����Yy*
I��f���,o<�(�7U-��}�s��������RS�U	�
��wT�u@r���e�i	�r���SI���B����$vR�!*��Q߫�3r�z'�m��Ͳ�<��)Q5+���5*���dU]���\rz��?�෪�:)��Z7#�U��z�\:�b1�v�;#�V��,U�C�E��@���7�U��hUٶ	׻��˰l*=Z�}��~��j��Gj���2mm�'����۱,7��1�`=�.���4)�n���Ю	)��:�Q� ���N����q��8&�?g}s)HLM�I.��v	*]0@m,��X�	�%�i�i�IDiO^�u��l�0*{Qe^P���Hn�C�2�E�T�y��ߙo}ț��2ڀ8Փ�f�B?��/_�In�E?
{����C�1��^��k㢾b�W`qe~�&q�_̴�G��yo��4���V����hy������b�B+���C��Ȳ��~�v��T綽t����1�;:�\s�SiB�$ewg˯>g�c�jC�����ǇE���Я�0�H����08����_�XT�����'�6�������ɛkP���W��cΪn���t'&�Lꖓ�^p����6�"����Tg�K��k]
�
���V�J@4��s�Y���V3o:M�2��"�ޘ�e_/W�(����4���ʮ>ط��U��&#ܕk݁��SIt�s>��%s�g��m@��5qN�
��݋��.w��w�I��(�ݖ��C��&Xd�/k�RH0�U�6]
�}Þv��b���}@��a��Jm�p6tP�J��s1_�W ��L�2p��/�$�M�vpK�)$mjP���:J�"����~gګ�Έ`
&L�	��;��S��V�a5;)����\Y܀L��h!྇�}ӽ�Q�����S���M8��-�G��k�%9����pJAtYA>F���&?��z�,?�G)�?+hukP
��GkO�=�荆i.�	Ԩv�+r�N��Z+F�a����WR�ο�D��P��;�?0a�I�A����sU�e��������N��P7��|����U��\��-U	�-E,���[욻�kI�kC�9�ۿ ������C�	Ҕ�v���aPe.%i���Jo5�M���}�4�����	��F�RK�t�,h=��s%���x�6�P@���5�=ڳ+n�Q	(mIѨCJ���N~]j���n���"m��:��ԑ�@^�@G?WmxK���x�&/s9ת�������r)�V@"��L�~g0Mԧ��Wh�e�/�f��������z�Ǟ`"n7���yR@�%�־���]�3�@.pؔ���]�ֈ����m��Y��.��|��.O&f���x����b�B�K^L�:�nLj�E���k���e�ϱ���zX��\�1�ƾ�b!���H�A`O�P�h)�l�"�r�FB���ׯ-�Ǖ�[ߤ
Ԟ�c�7;�����4G���{��᫷2�Mdi~��)��{����?&���3,;Ď#V��/�<��յ>C�֦�4脁dT*�Q@�di
Q�,	���,yS�
`K��
_6��Qo;���E�6����;v�a������W� �XO-Ȣ�L��S�W�l	0~F,��Է�IN��s�o�%b�Y��WF���.�t�Yx��,|o�nD!S�ҝr,껺��:B�8��MD��$`�A�[�O��ދ�|�iy�Z`b�9�U�ޢ�Ha�l̈́�S�O������"@�R�ٷ�i��=�8��+!�Kт�s�ߋ���ٝ�|Ƞ�Rk��E���c�⹂|Phrd
�����)���`�ڡY��	@�߼��,�(��]����6��{M��g0#��������^`p">�k)�=s<�^!){Z��{	��O���R��:������ի랛����F���d���5?�.2;���ё8�i1R�ؗ��mؘ��䛚�y+���v�����e'�\�~��GS�8/�c
�UXu	�8t�$�"8A�ސ7��$��,,H���/E�����[�
�P ��&��֣۩J �A�KC���qi�4a4;��@�~ذO;�(&� T�$�Y��a��΂Ц~>�J��)�k:t��-wFnC�3^i
F2�:�^�#�Y��N�Om��7�d��{�Ӭ�&0-i)��p��+l����U@�$�3f�V&A�s��ɡm3�-��4�3�(�e��J^�mQ.*"���Ȃ�w��Q��s�9/�(�c�|)���o��Ɨ4�E��4]W������'�!I�W<� .]���mME2����������*DV�o�V�{o�7�Nȋ����
d٭�d�%��<����@jU2�сV�2D�7�E�KD�\w~����`�{��Y@���o|�[���Xqጠ�[o��TU|c�cCe��&:����sF�����Mi�C՛�0��+����S����M�y`�VI徥S��|n��w1����d�ݟ,X�=�����< ���:���or��[��L�X�	� 1j�����u;+�እ�9�� �mQ6��/�f�n��-I�Q��N�JȪ~ �Uh�~5�q��	�J����j��@�������,���ܴ
��Í+M@��~w|^���D����t���u�����ZDjFg�F�_��`:8q��:�F	��"B��12ez�QFd��ľ�R�;*�O�P�넄��b��W��40�ݨK�|K���ԆiE�_θ� '97:�R]I��W?6ʀ&��C\O:5d�іQ�v��a��W�i/5�&a%��Z�T{<Z��+����Z���_Y�oZ��}���hϸ���)H���&��C0)�Y��ɖ愓�\Y_.G�w��7�
YG�E����RSQ�[:���v� �25K *t��L��RH�JFχx����-;P��+�Y�%���8�w���z]���#��E�d���`�-�M��I��k��' ��|*��S^hz�C��Ж����[`�$�+�j]���ܣ֍�.Q�1�)rn��a���	+��4_�C���L)���]��ϔ��j���=���ʃZ�q$��	�p��
IG xg���DhP�2S'B�
ss�\0%���a�L�����G�}�`��������R�f[�Q5����;���$�T�o��"����@���@1Pfs��/�sۆQי�R�2����u���u�
�m�M��d��jj�Y	m5�(S���pW5�[�l�t�z���$_&�x��IN�?︥�����G������	��h�ӿ YB��~��l7���/!HP�R,la��xN�O�Xm���n7�y�4d��}V����H>��Hi�"g��:���ԍ�%PQ����>>/|�5����ksL��4���tcA�s�/`�k\q:bM����^��
S+�3i�&�`�t�XǄ�c��!�G�3د��K3�$��/��4�9�X��4���� i$�b;�& ��r7��|�E!���A{�����̪)��x(���7[����o��uw�Mg{Hi�,w��D��ɨo=��q!��Nh�8bs��%*
�b*�ɭ�4����[N�A�Iؖ���7o���Zj��7g��K�/��Q�N�gZ+E�"�@Tk#A��\�ng��r��������e��'�.�b,��c��&JZ�hvRw�Lf�+C��]52!t�S���2�w�b�SI���q�:k`8q�/��^/0a=$tfF���ډ����.�����P�Ju��aJ��ve�0H�o�G�$,ր��`w/2Ei�h�@�fʒ���
/φ&C�������/����5���� ������iQ��w�@+B��Ma��3�iz�[3"��S�vC(i�n'�8����C)>"f+ם�n.4+J�� e A�n��/�!���a˵dX�|�+ԩո�`G�T|���r�4��7�.�SYG�����@��3�l�|=�W�
��~ĕ��e�3��X�T�G��Z�\I�xg��n����հ�я������
�}у�e�{A㩏�Rs}ή�*�����!��(��Pg�%AZ�k��J�/�8�
������ꯎ���&�J��S���:���������Ḻ,{����*���b�.��^2��]�Cf���p�,��<�Ab���v$I����o	0�)��������j'H���=q�Y����p�`�!��R��ܰ����+��D��cs&���lS�J����Mڑ�D�#cr����b�d+��E��Z$GD�m�zZ�2�t������m(��At��RON�
sMy"_���v˹� )��:�f�����8��G�C����h.�Y�U�=�*�WX������Vm��5tj 葑
B���0*�v�i|�@���ǜx6ȁ��I�jk3Q�yP@d��y�Ah��J������%���v����E��[��I�N�@2���2<fQӁ�� �����v;���H��[j��/��f���~��gy�L7 v�)e�+#���dT&KMZ�������:�a3�)�b�uZ�b\DAGϏ(>�-�x�B�(51O��.Y��=�FZmmuI7�����(B00A�7��<p�8��'�)[��\�ra:y-��]�����n] {Rd�- ʧ�wL�Œ�o��&�Ӑ�8r=/����,>��`�L���)Hg�M�:c����ψ�sǃ��|���ԋr�C��t�OM���a<#�"*.�������?���}f�N|���a*�+�a�}*�*D�6b ���>�R']a�Bu�d�3���hdפ����@"��S	�@3};� |jcO�rُ����+�zZ��������5B��K��˘�ڷR$*͸Xvc��]t)&��M�1��o?i���!3�7�U�$B����<g���Ɇh�=E9ZF�����6������CX�B��"����������v�L�{_�Ǉ��i D�k?��a0gχ������bu���-/�@Mu�����/�hA�v���ee����"�,w��1����lE�0�]l�𤘽F����#�~Fd�)Pΐ�E��4�j*ц��J���sܖP��o�iʇS��;\�Es'Z��=��O��㼖��I�?���6z�A(����YE��4e�ߍ����0%��jN�%�:��>�U'w�����c�S�J�	B�`�
����
{�ɔ�+���{%���B1�:� $;����7��?G..H�M�G#�*|�XnJ�_*���R�v}c�~�ÿ~
4�f�?����)}�,�}ع�	�R�Z��.`;l8�IH�.�3dx/~����g2N(U L�����*xy�Ur�k�)�IV�i����9ø�@�	�DHW!�PE�k�nZ?+�
�mАF�a������qe�����M�}����?TL�	۲`�:	���;z]Z3�2+G �ȇkCp�#i�?B����?������`c6�>�����,��z��p�h���q�X��5�O��}Q`�Xsksv�9���A/�)����3:�5�֦�@{Ƚ!Π^��t�;\���k+����9z�~�n� p(_8�2�
%�l5Xb�3%<���'Ԯ<�?�${�nd|
�4\���u���|�]�ڝ4Jq�i�����{�[�96Z�ãL�tb��`�ر*���ߦ�s��Y'$�YC��;���P)�1w|�����)��S��Ow	�mD07�{���f�}0�-�!���a)�m�A�қ�]�;K3`�io*ǩ2K�e���?�C�;�ץdfr8گ�O8�d鿱V�����
��JYk#a�ww�û�������$��=����nLw>�~_x�N&�cm�GO����q���2�q�,���+�]S;w����4�:}ɷ�J'v�m<]F��d5ֹ���y)�d%�׾IMX���15ow�/�b���/14��XlG��\�%��4睥 9F���w������J|`j��Ņa�*r�#��<Z�:�^|�JS�0�/C�y��-�����,�����M��g�w���8C��j @h��ؒ�,�,�F�W�r��%	��	�C;���N�x��tc�{����H����T��%�n7G�E�
��(5�9P�T�e���B�A?�r*G@�<��1h]�Vf�	���,,��k���͉�T b�T)��Q,���tv�����]X�S�Y�>Z�����m�������N��o��	?R���L  �g�bA��IL�Q�E�ez񞴗'�4w���#L�����nx�����	�w�<��g�Ҡ�'��R����R�P��d���D�o�
79l���).@�C�L[�t�I�14\�/1�oF3[�o����#E�sT����}�X����+rg���=S�ɽȻy�����%�#F=�rzփ��9g���3��c��.�F��~Lv��N,�2q>%��N�r���4PrO����2B��ҋk���G��y����h�F��y�H{qd��l�!Ь(�J�s�����I<L��7��Wl�b�~2�:i��.Uʚ<������tR�����-����s�C����RD�ٰ� �fqx��c�����R#E5�ol>*������j���d�S���H��F7ּp�zaww��r*���|��z��G�� �/F��c�=���P��h�����_@����\�|��^D8�1g�Ϡϗ��S{ĕ%��?a��e�&#?V���X����/=��Y���E�!�7~m7��5��6�����dE.G3��Jg��T����~%C*=2��]�yaO ���"ө�Va��7h� pd����"�=A�u��.�L�$^6�����{���J`4d�D[	j�GB2�Lqr�r�2.������.��r)���X�X�b�$W�3y�#ـ�d%��m�BXgB`��&��[)�#��9j12@���������X�a�G#���` `�����v>iB���o2�(�v4��~�m~\��gA��S�*���1�����i
�f��J�s\(Bm
7{<<���όg���J(Z5o�?˷�u��s�f�1:�>�a2�v�0Z��E<� �v���@"��YmR�����Z�97�;E�� �{-���=�NV�<9�'�e+"G��n��sG���jh��Tq�+���0��:�<'�)\!>f��W���k!/��� ���+��T���:C2���~�%�{��CF�ZWu�I���7�ڔ���/z�	蜇��!�k�/ ��Ǩ��Ɗ-�����Zڧ�0:�U�r�h�j�4T%��ɳ�a�CK�ͼ�r�֧���!�?[�4��f��C��-�U��*agcW����u%�u��I#�ˆ�y=�#�i��^�����K�#���<+��.J�����e�cYp�]�;`�И�6��r���S��\�g
��녬 Q�)�~{?\c�tb��l����O��?�h�<g%j��`$|[�1l�@C�\�g�s��Y��pޥ�gi�z���+Ž�-kb$�̆��S�����t�ڀK����uU�b���E��Sv�� ����}��;���+�{+���9M)���[؅R��ƕ���;��)��K���er|�������~jȺ�A����7��y ��8�zK�,�n~^�=>�����>�P.���X�҆5!��(���ۊ4\����s�U��L}@Fc����mCU��P>�x��slDk���<͐�Il�^��e3t���[z�H�:뉇��?��O<�g�)|9�90Ք���{oK��k��kA =�=n�na��T��1��01>5�n�]�^'e2?�jQ��=bpųQ󊩈�3�s?�Ҳ��0Ը�m����~ �,�e�W:�W>j���\�����Xb�n�l���|ˑqw��(/;��NRӞ#��)��t����#S-�>g<�p�ȷ����KU$�W��{ú�n���h7���Fk��v��I}	�s`����=�߸ �^\"
��	Y��5=ZX�5�=[ZkѰR�Cθ�!$"�!X:�	$���)Z�2�1���	V��"�?3�S*ijp ��rTxѻr�_h<{4}�oE }Qq�>��7�}"�I�V�6��L�Y���N�8;O,��3B-KH��v�{6�w+H�t�HN]�&�"g���1���F�A��u�����[�R�)Sv��D�F�����YG>�԰��Xu%�6���G������C�g43��|�	P+���;n�n	���9>�Z����^�7C�]�
H{�S:�6(q��U4�21y��7�z���gD(�G��U�k>
~�o�]��a������,�;aB�y���um]�@���K��}�Z��7��&��/���� �W
���"��qW&�u����E�,�K�/N�〈H�m�����|���=�]�ۊvFGi�0*�bD����zi�1�h�Y?7��S�#�#��Ԇ1>���V�"�� �ѬS���{��6�]C�x��	`,�gk�~G؜SGs�p(e�����K�2S��W�Ka=pg?*F�_4�F&�0j�%$7�2-e�
���0�0���p1`�nm��JM�X�
=0o�֕xwkc-��jz�C(����Z���4o��nL� �U�T7�|ܸy�h�,��.^��z;:[�d�
L뮕R�#��u�7�Yz�o��(Ă�/�2f��H����K$,�F��R���FV�ݟ�r�wy���wUM���Ї׊?I�p�{��=h��n`���O�[^��8~B*�ۀP�C�s3P���Wr�l�����/�O �by2*������xְ��ǯ�[���:ץ�d|)���j�arFiq�8��
�b�'�;����@Gs�E����N����֍NB=VꞖ6��o�+>I��(V>S��B�-�t��Ӯ���ѷ!��y�� -=8���6Y'T��ܹ�C~������~n�n.Rx�o��S���&�8�Co$P	y�Q��d~c��Tk���}=�'0֫�A�X�^�-~R�OLgz���?q�ViH�)�8�z&t�P0���A���ʾ}9�IنU
*)�s�8]���g��b&4j�x�q}M�ETͿ+0�!\E��q%���5�F��87X��'M�D��6Б)�F{1iS��� H��r�bl�{q�J��?/pw�H�&�E������2вR�CN2��<�d�!�.�g/U�Έ��H�%ҭA��H�����t��E%/:�Q����ZO�E&�W$�!;r�jC�ݭ�#H��LO��gS��B���5�r�ץ"A��O�1��srbY�i@��~,��\n�|H�ҷ �[ft���N��#��8BP�#��;o.E�p��<�����X��%?��-��ч(�Dx� 2�z&h�a��P^=�d,��DqUn��cr;����:�0��1�[�y b��-�L;�aVD쀘W�9I�1>_�}���k�-J�@�U��^�����22cv��
�1Ə$B�9R|�쥌`]�7$���yQ_���!;6 �޽W��󲎚�*����(�5�чWp8x�6�zP��H��`�G��@�7��w/�#��?jr<a���W���u���$�$'qY�@�᪟u3��E�}���<�	�i�����Ә'CN���4�)�$�	�W��0s��6(�.��BtJ/ĔU	��~I����y��'��rw�^�Tt�"Kl�^h��Wp4ᵹP���T��ۗk,�����Z��Km/�eY-�5�"��Y�/�c�Ā�@�k�"���B� �O��PF�H�/�@53��4,�d���B%}��U�|:7j,�q��G.��0��Av���\�bB�kus<�nt�Ck|��!f]��?�g��z�^7"�dR�#;p��J� !���Ĵ�7�d���	�N*m� a�"��d��O��1 ��5B��>-���L�f�j1.������z0t ��" ZMFH:�9��R���3���u�k3��O0�wF�e)~��7�?��S=L�4U}�VdZ�Ov/�8�&{%y�1��"O�߅!:ܟ;���8o%]s��c�	&�ϬPWfڧq-LA�Yw��i؆L3K0�YWhq��M�jԽW��~Պ��ґ�J!#7f���d�����c���(�� p����U��y1��	���;�Yf�A�Ƕ��u����YˋȿIŨ�tcnjPQdA�Q�E��U {�P�.�#�c]��o�X�:ޛ��@1wD����Y�p���o��(Yo/v��i�\�1�I��eM/��R$�uN%q��a*�uRO���On��=��)�y�g�=�gt��:7k&n;�C�z!-d�t`Ȑ+���ͺ����oluZN92C>��a��K�ɷ� а,j]�/]�a�
�kꠇ+��9�ZK�r�:͹X�d������QDQ|I$.���)�p�'�e���� <�TL��tBa-A0�vҠ�L-g.�Ro������{E�'F�+��P}�����o�;=�m�O�ua�P�2)�M���ɣ��٤���5A���pϜ�ge���]]�tVdn&~�azx(�n�����-�G��yr](署X[�m�C���( v�7�ᾺI!���~� ��*L�+���t���LxӢd��i�
�ޗ���!9�}	�#��f��/,SY+ز�N�@*ݼ�y���6�JlQg���ͫB�4�0,�kS)~�񖄩�&���A6G���n����z�s�_���qm��i\\?�-�;m�}.�Y��C���*ʐ¥<������t���VEtq�i�u�S��MmL}��Τܖ1W���jm���-![R't�q>�xͶ�(3]��VB��~
h��|��L��&�pC�y��yP��!� ��4mv<��Xղu�7�@� ,�@(^Ç�q��)������os����l+yG�-��N<�z��9#�"��w�sɺX����a�"�^�XǇ�� ��S�V@b4�qN�PK�%�x_��y�� }�, ���,�C�"%���'�����o�Y7��No^x)H�g���O]k����G���s���ۤ�e��
��:s�|�e�������s�˯���
J�:������i�z9t�/�{����O���N#�d��k�[L]I\���NZ�J�tcS+����HRL'����	�T������#>@������S�ɯZ�~Aը\Vp�qob�$�տ�&[�� j(�M�eU�o)K��> X:40����-8Gض�}[�a\���$	��PjK��&��݈�pY;����K��M�\a�"����,F���Nu;�*��y$=��27�+}�&n>��?g=�^Kܖ1.A���I󫞏�sV�����a*��\��dC�۶BÒ2MZ��P�^i�L�����$}u[��	*�a���d��Vw�B/��W}6�o �<��FN�r�dVu���E'��.��ŠP��1�@t��Ѣd5�p�C��[g�����=�s���)C��5?f�1�BN��ʟ��|J6`y�s3��~�91��~}G��M�Ŵ�;���"R�N$�uo(��h���iqq�fV!�9�u)�p�Z��'+0P�6?-S���\Aӫח�z/��v����ϠyQX.��j��u@����=����#)q썄Y����<�� s����5��4����ztb6��.6?��dTMP(UN�IuV�bQl��7�^��gJ�{�,��ğb�	�s_T�]��b
 Π�M|4��lu5�8_�ς��@��B����m=[�ĕڅ��h��2�6"u<�v�>1�+��Bhw�<ˀ�
�n�(a��Uz&����o���R�Z觓!�N���
�Q�׍�n1B$����2��0�3p�C_#��X������K޳�͏��3�\M��-�*O��^C���Bd���2M$�_$��e����+�8�ܞ�*.;.����s�%�:��zp�	pz��0�3L��	�Bc�ͺ��-��ʖ�$�]汣����"�	sl	߲��bT�g��f�԰�\�7��L�6�>#u����¢[�w��]�Jy1��_$I�:��b���YY_C-���$��)F	��8�,��.��S�;���ME��sK��|}���`��9��f|��>�gZ�������ᩦphc{�x��s�?����:��JF
=�{�k�?�7樍C$7/����������h�u�̚3z�K�\�!X��B�[k��]g�u���w�O���
�7�ՏH;й[�^O�P�)����DۦRh#p��w D�hD���]��8Tw(��e'P��3�%��".?��3
�b������F�8��-�*r�H�]��Y�I��r��+���FJd��ޫ)y�,
������$$��:��O>چʪ�t�K�p�mlYȺ13���4��o��I��lr�t�pM���\Q*�"P��хu]�.�`W�e���-���ɾc$0��$t.`�'���X3�����*����EHJ�|�Y��%��Q�y�[�5W���S��ahW�p�5�ܭ�E�S*�� �����p&����}v��=�������fq�?�.��>��a;:��B!�-~�-��R���z��Ć{��5Wf8�ⲯ^t�ˁ��,��5���:<9��\�Q/�w��g Pm�S2��҉x���?���}�'T�5v�S)�{�O�w������ Q�q�s(5f�Ƭ��ź	<�����%bk��K�.�P�C��
��ӹ;��c������>K��.p-�?E��%j5X�:��P}[�M}1X?t��;sfh��\`hKw���E�ķ�5�F3��q �`��Ĭ���.�|�A��j���+�Q���� Cdv��h��q�)��D��G�	�:+3��	-���l!�Q�%��s3	.ͯ���pmD����2�A������`��Lj�y�D�Ȉdo3���Z���3���[����*�ޔ�3�u|�g?�l��X�o�"kn$���8����m4l�~��-/�8��m�l4�����7�Р#���`i�vIN()^���B�@r�E���~gxL	D�.jܪ�S.4�0�BC�..�CY�r�Y̲����<r�6�JCk��$�G\�y�G�-�Hh�v��L��L5���ĳ��R�Sl�հ�+rp�� �T�=�;�!5�t��q5q�)�R��)��+�]�@��I�ə�=ij=GbApj������ ЙRp� �c���5�S}�(xo��b���RI�쬺�0�%4��A9��K���)ɇ��
��N�x�_D <C��'��<!��;U��7/�]�yS��^Bj{u��_������Gf)���%����#̟۸@�m��V����V�>/M&�d�2 �,|�c��nن���-����5���軞J{+���|Aj^�mA��#���N���.��v��� ��Ԋ����}n�ˆ�������W�y}p�����C�J�����C���ݼZ������<5� `�d���Vd��&��lW�T�$�#T��f�|�~W�p{ޟߋڰ+}�g��~��F-ex���F�_��v�Iހ��@�cèΐ�I�yj�ݼf��D��,Hy� <��B�=S��Yj�P@Lmn�p�i���Gw�!;ϡ�� �n.T��]���{C��-��"	Ƅzq��Id 9�֓��i*H�GC�k#N��I�_E�o�mR*C�&�� %��;�A�,����)zm��QV��	M���ȅU{bo��k/��sK_�Ⱦ�ӎ]�÷�J&��jˌ�S�\ᇄ�����������^�	׽ʌv@7��NpEp�������9Ѷ�U��伪����H�F���uͣc�NeU��m����d�
5#$�&H�,�س^z\��j!�� 
^z^`��!a��;M�h����DD��wN<[N�y����6��c]l7M�{]옛�%�3г�d�c@��ߍiҘ-9�S9�h)h�PjWi���7��y�#�_V�^�����I-��hs�}h3���� �*�F�A�tʎ_+#/�H���f����w�#�˖��e��H�Dy�k�{��5O�hן��
�lw'z����d���xM��g������tB&B��+5�jx�9�_c��?7�b�oN��iʃ{w��ғ���,�A�͗�ۣ>>໖���M�H�Q1�q��c:�	�Zt�r٨C��0%Zm��M(�����L�i�q '�TR�S��T�9�Yg��H�/A���*��~,���'����M��'^�F<:T�ת���l]i֦��8����������X?�EUZW��d㢂��apY�7$������<����~��"��W�yE�.U������x����M�3���.�r�9����_�یȸ�3�
7Ы̃���J��nB��)��m)���zQ�V�EX�����H�ռ,/,���a�{x������0�Ϧ��zBL�"Y|��@��Gda�)���E��j���~F����#��E�����$	��Wa׊��u��2x�!�Ԫ������F�L��;gUh�PSB�SX���I� � ^�;=0�VmQ�|﯑�Q�6�z�XOT&���TMk3���-��	:s��7��|b��wV���S�Ђ���2��O�A����İ?_�G��	̇���b�H���\&l8�/lV6��;Ob�q���xބ& *�s0���tQrvЌ|m���7��YǗ�`�7!��Z7QB��=ƅ�j���ԝ_��&��Fbx�_e�>�f��D� <�����s����@�z�^�_e6��FbG7u����(b����C
�^���*�s"e.	)����ЊL9���W֛en�^��[��\Y�������Q�!��4,���R� ���s����E/V��c'mlB�9E}�"oy�L*>�Ə�S�q�p#��_�(YE:��
��i���3�VھJS�nO`-$� ��ƲL�sK=0��Gӏ�,�(R
oݘI�4e���Cu:�ܒp�3c\g	��e�j�H�(��k<W��O݊�؃Z0$��_l˱��9	�$?�N5ڌ�́���UxF��h�����>V��8��G=@	6n W�>�&S���Yv�Z��q���0qT�w;�%�sf�)��ܟ_���0p4?Xt�t�<�SzHS�y\8p��ı�q�k�	_����(��1V@���7q���(���m�a?��T��f{�n�:}�����zt�����b�ʡ���4-F�,�h�	fݵ���eQ�|?A���ެ�'o�k��Z���?��ЖQ��G�q��b�BU���"v���O*�a��b5i��"���.㫲C���^9Ǝ4����z���t ��O�9�fr��J|��9�;�Dp�Q&&�`̑�ʀ�/�pZ�6	Z�ۮeqS)L6cj�$��S(�[�U�B�
 �w�{��ҧ��I��,=}��3�4��6f$���wcW�	�1�ۤ�������OUA]�A�^�JeF�a�!��g'C�5��I��*Q�@}N�M�'C�;��R�S~��$_/2�^���=ϟ'�X��F�7�����|=|U���G����H��ܥ�!�֞����q(�&���o����Ow�=P9�M�m �8ۂm?�Z�"(�_�.�$1o��Y����B��cbzmm���y��:��
ze�!RN�'��Gy�$:zx`M1����	���ŚD�����uoC����n$��Ё��.f_�e��y_Hxׂ���d[���GGП�������jiJ�!V��t�*+���m�Մ��8���a�����k�ڬ��?F����!���u҄;���r�ClG�WK�{���ġ����5��p���QͿ`]��ub=�g_|ч�~���Lc�5�����d�F���pqG)��EI{ѥ�����qJb��B��2��I��=�h�[2,ּ�I�s'��b����J�ܩT6���Ru�auI,F��Y��o+W4111J\�42K5�ga{�,g��<K83�i]�^��EZ�t�*g\�!.4t�g���n�X
����~��'�>��aV(���T��q#�C~+joD0�Fxb����*���*;��I��:[4��r��ar��[k�t��=3f�oz��,�=�C�_S���|�2Aߠ��6����#ɬ�(�PNp����"�J
BBc���[��ɠ��F���r�K�1�~��&�
�h�A��N��*�m2�A���v�m��]fīs��ͤ+"��vT�mt���{�86ׅ�fq�~x3R�������8��@2�:`�$[T2d]m��*}80-L���c���qq<-�����l��fn8T!��35E"9��DU�O�����I#�x��3�?���O��b���)����S�I�z��D�V�ϼ�UgG��hwI���EpJ XH�n��X~����օ�.������- ���p�G��"���X�$�����󨢸h-J2џ�@N�~ʨu^��n��@�^�C�(���X�D���m&h��@�_���a4��帖bJN�߅��k��hx�PˁbV�w�Z�;�m��8��/H^�)�H����u��Gpri.�,�Um��O8M��jS5�@��i�O$��Fs�����&'OV?H��$Ĳ���.�ּ�%Ԫ����-���s����������P̾�T����ty�28,�O�m�śX{)u�L��j�� ��P�X'l׺��د^�moC:�!����#���i���"m;x{d­��d�D�^FXyO~֤����4.�@�ѱy��F��Bsݝ;�S6�5<��\��/p<T@D�ͩ�k��^��4΅a�>�{���@��Z��~"k5�k$�Q�Y] �C��#׵x�������Ӥ�Dg�)ˮ�yD��q�o'����:Z�KZ��cJz�!���eW��8Q3{d�6����f���zi5$������|`�~*9��x����[f-��ٙ��F����.����h��UtLl��� �KQ�݄o��LlJ��a���F,m�
n��Kz,𤅃G��k&̙o�$��N��[���	�-;�_�m���J�6�ʢ��>j�3��v�B!BlqRu8�Xr�f�I���7��ҁ!��0f��B8ߐ�S�# �
��1��{4�X���L����\�8/��z`2a#9��_���i��P����yR���G��U��|���v7�qK��x,�""<s��K�}u4�O��Vf����1������S�󎹁�s6ʠ.��Z��Cև��n�S����w�5'a�35R�F�%W:d�����4;��B�R	���z��*�Z[ԭ�wjcɨ�r�
���AX��brQ��U����T,޵�O����?��-�v�3�e7���c:�(�}@M��������;V6�
�C�.���:�U���i�^�=����5�ۼ5��+m���_�z��@��OoM@H$��NG��UWB�C�Ee�Cr�	����I����js�G���_��6�G�tLL���cO�*&��(iX|T��U��%G��_pqZ�il�.ӕ<=/$wX��� ^6H���B?�"-�p4~�SiV�����'��s��+5Ly��, �
�:�I�Di:#VH�y���)�sb��of��yuE�7~֌-���X�k��W
�yH��[�o��O�d����]ʡ��O`��~#5[��Ӳ?yHe!9��T�0�c�'젲���
rGqYE��?�nN2z=�_z
��(*�.���+ǀ.�)��eU�����R�i��pG �����Nyz{[�ףp r�0�&�YX�+#}Q���6�������C�aca������ex%�=�yJ>i*�����TKQmO��c1F?�S�*��o���7��7��b��O��a�aQ.T2̰�*����(A��xo�0������Gv���6���U���T�hX5���������wN$��\��J4��&��=���34�(��~�Mv�o�]Yd8 �q&�pĒ^���Z��0�J��$#�;9��S��P�zd��#�w�ׁ�؉���C��aKBS֦�Q��8���X�y+���a�T
q�x�9�	ш��"u�$j�m!�Q�sȴ�S@�g��v�Ճz!�K�O�P�9���䰁����?[�#���<���W�'N�,��*@���kG^$ƾ~p��F�r�{�QϤ z���z]�������4�G|=gd���R5S5��)_���HH��0¼��f:�K	�{�Ѩ-G'4-�^
�e��P��O��oP�����g^>���7W��7c�wnX�{ʫ]ܕuzX���)�_Α�{�M}�؛O
Ҧ(|��	�Wp ���WhB�dE'���H��\!�ӄ@�XI����yb˻��T�ąw�,g��^�����^�7l��Yr�Y��(O�����Uj�7��r�S���k�֑�P��w2J������渔�U����<��Lxǭ���())Q�(�{2�)uԝc�����Q|�����}^�"�BTԦ�� �]ڝh���\S'���+�ɴ�}��&4��H� S=/E�wT�តI]�_�%&�&~~��5�/�
�ǿG�Ö7�L��Kɠ���?��J�Vs`^Je{�9Z��Mh�wƙ$��1m��cDV�`��0Y�72m�o�Eu������kY��2_��!Y,k��<=FJ(�6C�<�;�;�ue�m1z#�B�[�\Ks�9����~�V{:Tn�Uڀ�����S��	�O�J߱��E�V��SsF�R��uG���R�3f��a]�r� ����:R��&�+-�F E0,�n�����&�Y����0j�ؑ��:�� �L����:�a*%��,kV�o.4�۩j�������v���$X�tc,S�V|j}���TĊ�p`�|q��ݻK��umZ
|�)�|�^Ϯ�q��ٸ���{��⾅)��riMRs�݆�æ]�DDɩH9[{���8&�L��d��ꐦ��*<}��X9hA�k�t�(�N�Tm)�7�,m9iK�	����������K!�s��f���2�z��k�X�o���_]�?�{��U�O����`��$�	�b�#��M2�pō1��5��rݵ�k�9[��X��)#���C�7�>��L�~�##�a��!-��آ.�)ч���&�_���F��n�.qI���:��hF��v*��t��;�2�~|$?��C���[nH�dc��0-����gKRRy������lO�n�b���3�@J�R`גx�jQK�g`�Yx�� :�Ȯf9����o!y����Aj��ce�_��J
Ռ.�9��3넔`rB�4C�H�b�[P��ȸ@�N.�o������P�����pe�	��cQa�Q���%C����`����	}���,%1�Y[��H��W�[��%$u���	͉R�����#�A\��%����Nc��7=�a��?T��`���1��X+��7m��p�������p%�Yf��Ie����XS<��������3�mq���rT�6Dew�J�����|�X��X�5�(����l�}�h��{ ��o�e֡\eIp��n-7�K��-H_ظ
,��EqhK�|x�Xb�(�ō�K���uڢ2�1!�]5�҂��Y5;+�@�Y�R�bTNjf�'W~o����:E+uc���imQ�H.5��R��8����3P �a��_�*i�!߲��S`� e���9������k����FKFZ�&ȹ�׮]%W�P��
�#�{���)z|���F^�͈�� ]m��(xI/U'��R�E�������#�u��u]��:���:��R<WBQ|�)�O�,�/��Ā��h�D�h��n֊����{�]e�����N��� 
ZP�Q*�]��Y�вX&49(�Ȍ��w�6��G�f�o�k�`�ܞ6R>]�c�N=4��R~��h����ӳY��Kܓ��*���f��f�ӗ�Y\�;��Fa��qF��{��\��vƪ9����� �뇧��|��e�K{���O�V^�\�f:�EQ2;�ό���p�C����5ҷX�@d�~O�dsy�JqG78.fS[$o�[%�A eh�+[�u@���*�Y�����o�7�7$��g����ko�]�R
��m���s���f�p3	�-���X��)Vqe0������ss˫T�ݬZ���C�ҹ@[l�È?]q8�>B�ݾK�����jw��8�+X�ȵ_���W���eF�����Ia�� 8�(�9i5�Fh�v@h�nͯ���؝g!ԜH�
�f��� Y��#����")������0f�QZ'���[�|��t�oBN�_R��;E��Zڏ�T<�5�Ԑ(����j���T��s�b���ѷ��&�ߒ̎8����a0]��rq�!��퀽wM��(C����m�6g#T'���mh�ס�����b~��$���8����w��7��z�����6�>�&�@��f豳��L�m0,-�uk�N�q�z�q*�1�[�ץń4M	~w1��@Z��>SV�*݅Ό�+ �}u�v�>�٫X�̵�j��t���%G����i��������ɺÖ�b��F��QCu�U����R�-P����>QL�]�ʃ44�]�"�!!8L0�.|�v�U+
aV�{�p<�}�n_a��x��U9f�aTl}R�S72c���i�wR����A�˞.MR��K+-ʳ�N�IWq�_�g����g�IE�V?[(��/����g��a?�l��Y�K���M���<'���g�	���������+�3��������C�c���~oS���X�c�䉥�;�����T'��s�!V�8g�Y\t��p�g�N|�.�g57������N\�|���~��O�>�f̜��b�V�{`�])u��2��¹�*�,5�����3����Id�����	S�Fm7nY9
C~����x�%���u�W�D�.i��$���b?��ۨ�C��ʥ��������"4H�_yWA[��W(!�����)�#g�M��~U����z�~������ڴ%1���5Y#���-uA@���_\k�76�	K\���I�xC9�N߼Җk����J��ŇS@x�=�����cu՘26��| ���y���#b;��m�XQY& fpp�nD5�	޿Q8*�N�a$4"�{P��F��@�.<��T��J�ƿl?�p�[�4r����f1"�)�,����2����Z
o�J�,�%4�(<�q�vh��W��v7����̃��R��"���7����rO�)�uݱ'q ��R8亻1���ǎ5�i�|�H��Ž+)ɯ��>�� ��t�G����]SF��#y��Q?؅P�k5?�>&Su��g��#@�*f(D<��HZ��A�����8}�5"� dC(�2�0��$��������9���"j,(tNY`��z�l�oa�@d�=��4R�{�0U1��'Ҿ��Gcߝ��D���2�r6%�6ń�mc:�Ղ�8ȡ��ijj�(MTX�?=ΐDl6g`'���K5qYCh`�W��Bw$�m�olȅ�DYE�����HiU2J#��3��&��g}�����'�^I�14�9]���oBZG�ˋM�}�:&B�4e�o����{����q��f$rA]�`�|��檷�#�[_Q����I�~ٍ�l�X�M,�V��)��Ї	z�3��l���E�u��79m�lV�7-� m����J3���{=�[N��4��'> m��ooT)�����{�7�]�{$�Ga+�_��ȹ6�� �˃�}tݯ����qZ�,�EoLocqݹ�V�E�f�&5�H�0�m�{�dk��?d��,D��}KB��o��$ULZvf9H���ԇk�=%���1q\+��j�5�M�o��]!��}��{<��U������wo㉰�QZ�:5NV��~CU`��E�&���M�K.��R����Ps|ϴ���Y�;5gG�����PC(�"`�9g�!U$3��E������V�H�(�)�v�c�9�b\a$�3���E�i~7�`���V��ǭ�p}�0:����y��D���U75�:���.���Z75t�
\��CӦm�K�E�nb7�E�,�����'�g�r��ż�5��]�g��	��W���gm�$q�R�S�D����z���[. �y�]����l��b�?�����~P۩�rV�%�ζ X^�x��2c�����8Ѐ)�M�B��̔g$��~�^���ֻ���h�NI4>�u���h��]Ȉ�����m(�̹��G{r܀�rE2��\�S:|��'�-Q����P޿9!W��,dL�BY�(�.0qR��y���`�����v���Z�t"���&���H`EE���;�,�V����~+�O?�B�}��9�(��|r����P�sS��dxǻ8���C+8��VԵ|��r{W9�V5����PJ���aUy�b�|�Ma�?~���u֔�a[�#����tl��=r�1�c�)�ك���Z}�`�X,���X���?�Qc�Յ�~�h5�|�W�Ó��a� �ȓ�xMM�DϞ�M{ZB��{Ti��`�|Y4�T!�2\pW3Y�b�����E�>(gI�J��i�_Q����3Ǒ���`�]߀o�9w)�M ���JΞ��ߝ�����c\"^5�:���1L�--y���\D�Cz}e�Sɽ�:���L�����2e����r	"�f���
�yZD7�)�tz+��4\xݙ$����[��g�Q��9��N���Ж��p[�2k���Q��A!�i��Op�<|6�#�qA�TF�|̝\�5���PM���J��7~�_�Wd���e�־��оVH�rx�w/[*M!A��fA��̣���I!� eY��w��fA����dC�U��U7$H��fG����؎�APy�;��؀�)L���L[�}(��CX��쮓pPa9�l�*���)7eʠ�g��M�IQ�zRY8f�r�E<�u����'C��#l�?/��R���=p���F���ޙ�]��$����jj� �M]A�����3#����hZ�(�Ըx�:�k7����֜��O�B*E=D�ՒiՋE���5c���`�!FB�̍(Qp غ���`��U�Cr�@4���zJ2�i�BV��-[.f��Om�dd�x2������Hd̗D���j��Ƈ=��8bd�IZ���-q H?�o��vY��{i���[�n-��7B|����o4/"Q$)�]U�k���h���?�N���W`a��Y_� �6X��@�J5��^�í^��� ^�+��/��$D�[�R���{)����F0yЍ_��%���~������*"��e%X4�wC��Z��W���Ĕ�y	�	�|������(��U��@3h/�ҧ\�mǗ��Uz����A�hYI�-�����Ȋ@��O����K�%��ϖ<Q��ID,�2g��)�Сc�����P2IQ`���m��qYU�K��.�jqChB����� ��w$Ȍ?g�v�m�ƙ�`�KH��ĞTa��H�e�1���ƥ!T��W˭���4"/�4pK��.����T�?������-��XT��oI@�"?P��r]._�i�)��"�?J0�\���19+��[��z�ǉZ�q�?a�e�`�5�M�l�N��rgg�Kv���u�	��[�W[Ʀ���췪Ӌ�Z�3&��*��|&pN�p�,"ce-?/��N�h�l©�1���w9��xS~���h,E�;O^)�s�5j��9R
��ȕ���c"�b��dE���M�4x��}o��cWqK_��d����]�����x���fa F(��ٝ��#�V��WD��KuV�8�h�tjj��LV&��80��L�en �[��r��E���S�l���uA�$�!����
��[7�0��4����:
�AA�� C�&�p�<)���F�� �+uO��!�%}�*�h{�@��g`�0Z��+eQ�OO�?��{��mD~�=ci$~4��1܏Vh܆Fo�~�@׏x�H
�i]Cw�wY���Bs�яR�Z��[{(�QX���Q��K�x�#з�2Rf={��yq�`�0AĽ�0M�#�2p�*<�GF�h(��P֘b�f��)�͈�X��Nǋ���O�g�����`k<yJ����[��T���<��?�gGȱ�JH�7o0�G��A-2�9�,��9J���ϟ�2��]�爳�E�/L��.���^��I��D�	y=�"�J��3�<C�O:hK��]�t��A��JJT���땟+�x�����o�)&���O��hQ��Onj�N��*��p*�-�ju��H7����\\�a��^���"�-�N��%p3$.�9SUa,�b?��P׵�Z�U-w�8G���E��X��9%�7����D+��͌��Q���)q�T�_�B�A5���J��Y	~:Ɖ�#_����󛃈m�#�ݍh�U�W�W���6�!֧�\Q����P+3�|����_$^��&����ߔ^�9�C8�5\���U�ن���e�9�������ze��>���W��#駱I/�#��)�� o1]�S]Q�[�i�~1���0\�/R�6�_�|j�:�����k"��:���P,�*��a,fr`���u$�$N�U ����X�r<�xUŽ��2G�:�!���x�ӗ9pj �M!k�F��3$��S,:�2;G��U�1��Ԁ��GuWޒp+aN���Y��ણT����E�,ՖwCi���9�, ���d�a<G5Cgz�`K;����|-��*7�!
�~[X+��K�M�1�o���bb�?׶�B�V5�d߳K�g\dz�"�pbWp~�=�goAw&�����|�H �r��}ʍbe�\��<]�^�2 E�G��s��Ycn��4@>��.����SJ|���S��(��'�?��cL����>G�y��W;��]�e�p[�l��h4Ŋv���޹H,c��L��S��.���[�T���˗6�L�%/��������jJ�&`�[��r��yZ�J��̼����F��(�{����}ᱻk��N�V,	���?��~�2�s��aLHٍ��.7���kۖ��[��Ub�3v�[s�g���|�<��=�	�K~>�r�	�0m�����6k�^��>z�x�d�9 �=vt>��q��^J�k�$��1XM�ⱸ��j���Ei26��2)�AQ���G}GQH�,���>�<��ײ���_{Vԩڼ6����p���3����Z's!x���I28�{$v�����M�7yc���1�5�c`�����:��)o������zE�D<	LC�ak��f������R���l���Xz��wA�\a��ߵ�	��]�?�EE+��-�I�,<Qgl`Z�*;��.�W{vULi@�m#p3��EQ4p��9��n���>��ʕA[s�xu1���,�ɨ��|*/������a�@��#kY{�H�\P��,�5��w��ߛ�]���4{��e�x��[4CS�X4�ț�;|��zK����߂ӷ�0Q`�W��}-�G�ŗK�Ƿ�G/܇�6��.�I��R�<�b��K|�.E�v׊f!WC�I�� �����ӏf���o���Ρؒhb<
5�[��q�`	�����'5 ��/�r���
�O'�CH�L�)�/,7=
Vkt@*���ˉ^**����,�_���U��3���Z��"\/�&����&p�QA3��X9t��K4�������Qk1;�aU���J�����B��Q]�qe�pP��Koʉ��Ld�CX��}�oG �u�j��g;�1*d�g3D5�	h�_�{�ݍ��uӃ8#H�D�+Rn�c�X��!��.����
�ٓ��&�.F��E64K����?l�B.	���g+7��7�}��fA����:���\'^�<��L����#�(La�d�*���x��s��N��6�tk�?�p��[��HrK���ډ�e�������c6��Ks(2����M5q��Y���!��+_�.+���Xe%��$Z¿�r�3i��r�B3͌��Bb\�C�9��Q�|˷�D��)!���=�~:-��t�͓_�C��wq�eG<��&1�FB�z+�;u�*�Œ�^6�i��7�Ԥ��+9��>�n������2��ҽ���&g3_�I]�`�2��� '>�D�К�3#�^�s\2Vd�M��K���7·���O�9a�!��'�v��-K��Ŋ
\�ȗ`��-�VMH�R,b�"e�`U�t���ֆ�b�K�6��*�<�HO��1d�ט�D��n�E�CǠ'��"� ����*m�u��C�\�ZH]68\�e��?����[v�k�S�!���h��:�`5�6�a��'���`�ƗA�J�d���g�B���#�Fi�6e�,}��ْJ�/íZ�v5��~[�D�xY��?6hgM���T=�iKT[)+�{�Ds��hpW�؊�Wwd ��Z��@�>#ST}k��%�g��	H���ضj����!X�NΟj-�@���Kf��.t�;�|ҁ����<������ ��[�]�7l�M|�P7ǩ�SB�}���1g?�����Xg��"J&5NWr1�����W��sk{fO���5�����^aQm�Ce��E9[Z�7��X���.'�U�t�d�|7`�Gr�n�2R&��!���>�F~t�6O]�<�#	��`��Ze�bXѤM�V`8��$ٚ��47E�E��h�[�,��� �?ZZ(lN��p]��?�s�Tl�4
�5bn�yj�=��ކ�F���10!D�i^lú���9X��O}#c��=����䙱?���8��W*�Vȫ�L�����Ozit\A��8����1�s�g���,���3�HN�a!/?�Kl�;]Ǧ	~W�2���)2�3���Eδ��fPG#'n�����U\Y4�3陾���jȤ8���ѳ}59X�8QUd�CG��f%]@�jq�j-����H;�M�N�����-�I���Ģ��c���9'p�]Ӄ���"� �x�!mPˑ����i���#��UB߿����� �2���ld+���Ĺ�R��͑^@~F�G�W`q^q`�4���@bPgf��P�{ �Ac��/Q��/\Q�'ǈ~���u��"������x�`ٯ��в�(n���;'�C�z�q�sR�c��%:п��T�� �s2��n��d{u�R�=����<��Π\fAmY��<w˾��J�g��oZ��x]��k��uQ��f
�j&f�\$�q[�~� ��}X���y��z�CE4B�c����ƽԺq���=�ϲq'k�)t�{bŎ~;�4�ȑI��-c�
h:�^�T�H�@�y��Kx�n���$���ܒ�����8�	�!��C�^�hHm�d$7�]g�s��})�%��@N`��hD�j��y�y������2�5��4���B�~�U
��F��Bu酗jwp9�bBR�H�S�ĥ�m)C$�R�E��m[>��Q��Rgگ���s�FNdz�2' a �ta0ג��J�\���K�NRK�6SZ���r��>�d6k����:6�S���Pn����T�S����VR��/2f[��
r �A��Ax��|�uQs'�l��7ez�>���D�A��aw��V�R���KO��5�ݽ|�Tͻ�Ԛ��͏<3��ҪԲ�Ϗ;�4�
��+�X���v�0�{ހp��ݞlAX'� w"���׶z;���4%�Ū����N�4o�a$���u�s�-��7P�jT,��ϨP`[���&i��@�)���V>��^�h+�|�T _��Z}����ο���V?��C�Ͳ��r�r|�T(<�[X��N�$����jh�Q������D�t#]�  ��XI�R�ԁ�)�t�:Ą�:��n���˭zL�~��뫏Z�;������|[asv�W���� ǻ*�F�2^�X��5�3h�3q��%�~���܀K*��5�MA��)7y?O���nK�u��
Y�@i̷�rCb�Q�{V�"�{[Z!�|�ש(b�묈F���\��1�T��ĭ����ڹ���]�]\��c��ʏ�_#H�N/˅�m��8cfT��`kQ���i~��H�rh��XGFYi�^����p�O4�5���YM֎����
� &E}��~�4>/�[�s_��%]?唭K7�-d�$T�.ea��v ��B��_�n�::�=�R���Jw>�~�)�����P)���$$����=7���Ut	R�l;&�{��~��ϴ���7x'vk��CK!1C�D��.����<����2'7� ��l�~�A�@O��xz�EGCB\���`Ȫv����#��nK*�SN�<R���?UO����lv) w�1�N�춈��҅�+;��O�۔��7T��6  �ɴ�]�km �"����3����@��d��
�S�3������+͚D�Si�$O���Nd��4��n�	��3W����+���c���5��'�b�9&O/��ȇ��LǾ���-����D�O*/,���,������a�a�NP"�􈵎�|����+�Dǫ������T5�Ǭ�C���'`ssmQY�l�QjD&�{K�^�Y�/Z��`d
�����ZѣA��d��S���7��_�b�]�X4YA�q�$�F���q0K�!t��9�^� 2�_���4�yݡ����ZИ֌��a��0�\�ʹD�I�	Ip�\A���y=��E�FWAR~SZ����ߪG�:�3�u�E[-K
E�,��3�t�[0�SF*
q,vU&T1�����m�[Lm��c�?�W�ҝy�_0��������?Y�|����#A��c#�o����� �����0%�DA5�U�iD��>�/�T�7b���h�O�!].42������}�@��:%H5Ѭ������ ���]���/�����m�AIV}6�I���:�/>%��[n!�y�н�\�V�o� ?GwZ��ܙ���
��t�K.�\���u<�a�3�CK&3iT�{��]	��=�\���1OҪ���U���g���H�7��_��j�q́;�4����*�y]sMi`"tVX����~��`R|�H�cz\C�H�N���_�d��5Aɟ������{,��do�Ѡ�Z\�4^+(b?��8�'H �Y��8���>3�A}6%�Vv�L�]�J�]��Qgs��*�=7fx�<pj:��|�Ҍe�r�{잵o4B�S��J��ȟ��Ԇ�u��-��.իK�)������zg�UW�h�\`۩�C�_����4��C�D��̔��'�-z2�M�[?���01��/W�3}������
0�%Nհ<��%ΰ���L��1���v�F7Q�>��F��A*3��$I�4��l"��Ñu��(��v>?�ac�Kܠ�+զ��U����g`6�:Ī�����_	�(���`vLB�X=��S0��ݷ��_�cv��^��~S�TL �o�M}$Tr�D��2a�C���g@�_ B0�߲"�J��S��E���)պv}O���>�z$!�d�1����@�(�	[�|f��݌�Ws����f����N)��R����0���,�=
\�����`b��4� $8���8D� ��8<����>��#"dcX�UvY�خ=D&0JB�_�;�%��O�#��y��UW��=�(t��)���O�I�Q�e��S/��Bw�4�LL�6�Xi3ڈ��|��及�� c��C0e>Ԓ�i�u�Ј�OįB[��(�X��yp"�'��J��)�e����x���TC0x)���ρ�R��?i�|�?� �4ͣ2��#]��'%��b	��P��xc>V*u�HNnt��W��(z�z��$!/�Y���䴖A�w��QyeC���+2�
��H���Xx^�IϿ�Q���+�{EW�o�B�MA �k�`5��\�_�D0�x�X������h_�/p������Q��=�	�Y�И�e�^�N��{��������/�'89�%|!)��v�� ��	��R�bb�lY`���u�"_}b,Ck������0�Y��n�&�H�Y���C�X�΍k�&Hq�G&g�Z�D���h���e#yP�n�[ֿ���:�������'�<������i�ӹ����˝Pٺ)�����S8�i\F�tz��dlEr�r��Åb�%赘ߩFt??��]�������ͩs\�軸n�i�Ud�Xny?��M:�-�\��Q.�BK����v�#���5�f׌HK��a����J��q�OC<ѷ�$"�&E�� l�&���k�)2pk ᵩ��G��A��6-\ #魩�����(�Kw�:�H�����@���M��kظ�tk�7=�gaj_NXҎ-7%�bR�2�>!Ru��Y�v9�����?�4�sߵZ'K÷��=�+��2���7i�J�c� x�ޢM�3T+d��2u;�s*��uX���8�:K��EʝY�� �JR�����2�[�r�,�Ȃ��C��	��F���Ԗ�X��(�Ɛ�HY�M��^�
��o3^�k�歎�"NY���G�2�������ukʅƹ��oP���P)]u����c1����GQ����٭F3���4>{CR*У~}�C���Ù�8�p��~Zn�׽0g����V*��׀p����*�!SP9��^o�L|��"�?�� �����bx�D7X�����X�NdS��k����m0X���ܾlyA@|/�:�����ČB��,����HI��T	���"k�ƥ}E*j��ƋSY�aS�Ȯ<�J��YU\�A��][��bo�6ǲnLw�P��ȫ�s3�b0m�#�2��P��~�n!s)"�,��'l���D�x��N��g<�6���}T���8 ���D�R�!"�g��[�D&~��o��D�ʈ�c ��n���p>��"sm���@� �y9i��U�1pa�K��ݎ,��­j)�8��0��q�e'.%+7%ݶ;���"@�/~QW�*���XZwGR3ӷ �9��А��R�k����$_!fq�� ��Y���<&)9g�p
��q/��y�\��VS��V_��O��L�I���/��,gMzpnb���r}�Ќ�� ����70�J�8M�d���܊o�h��|~�btg9nxx��������eN�b������}Wm�0tj,�+*���Qn�V:���ׯR[�*���\�	���ߪ�7�l����I��:�*:����*�H�]w�0�����sɽo�m�Byk��l��߁��xvd��8v�!��R��	���ڷh�H�u�SA�&q��?��NX��!0��T�qݼ�7�Mr���o޳?J{��˝#�ET;*�cb�HV�A���.��f�'
uf������`A
خ67%��Z���º�'��/-#�3Lo?�����;Ӻ��_T(��e1M\Tґw)�rӆ�1;�s�F1o��z�$؂uxM�
�H�����N���?	E�cko�W�Q$�h��.�D��&O�KC�+<�����x�-�A=>,�z3�ixc-62B�|��ﻮ
ZHҟg�wS��Z�!�T��ySV��(�͎29���g"��ѡ��	5t�_DX������T�:��9�	0`�u�D��v��
��#�P����?��s�ɟrlb`k@豇bgsY9��|���X�y���g���׈����uf�Q1z��!��p/m��zySC63����AIo�\L�A�j	��@J�#w?T	Ф�5$���#;��2	Y��	A�"Ơ@��;61���ר��+TC��6>#�e��38�b�=a���0Ot�7� �S<�ȥ�1�'3N%Ed���p_��9�6b?��N)�'	�ʬ�%-?�N=,X�T�z��w��+��f�Cn��H��`=�}gŴ�э����
m6&T�mC`�>�#@��7H�A��Ugқ2{ii�
�g�����%���,�||�!��
H���~a��@I�4g@�oѫ&V .]
��WA(�l'���Zhl����G�z����_�i׺�͎*6�ָ;�I��m��p^���O��q21j\��S�sR�f}���{٥F/���V��Ng���� �0�Z�c�g��>CpZ���2�	|�a�u��pTl���r�QKk�<�[�Rӡ#j�M 4}@�!Q��F�0�})��0\qOt-����NG<ɍ�X6೺��ֻ�^R����@r4L�%���n��C�Onq���R�˂zV5�S��q�f��c�Y1Xcv����P�e'�%oi8��I>d{\�$��I蟉kxp��gE�ӄ ����ޞmZ�4w��6�W���ñn)�Z
ǍF�_��j���*y�"����J;rU,MSO��ͯ?-���I�:!��)8a�/\r�(�5�'��$1�5!�L�$
���t8	���3�R�;hQn�f&����~n������Qt6��/��+ئ���%Yk-Ǽ��ύ��bQ*�8����\Vn�h�:yR���Wqb�6�KL"���^O��C��p}���mH���5�5����U�P��]2��� �nk�Y��G��<gd�pf�����T���+�t���c�\��o�M�����BX����D���Sf��"�K�T��p1��q�6y~�Ĉ���Q^7��&�A�X����]$O��هq��V4Td.���$��`{⍗��\��Fq��6���J����c�Z~��V�i���2���6���)�$���d^Mn`��u��v���tkm/�AM���#��yk��P`r�2oc�c�Zo�=u�]s`E�HG�{|Z�_6wjT�iH��7��;J�7.�+��4ܶ�;)'�Y"[єu�X� ��E���xm{�.ꛢ��5p�i�X,��}E7���xu��y��ol�շ�6������
�#�%�����1�7�����: `V�Lt�ee�8�Wlc�l��G�o�,�B�*��_cP�G^�	�CV/w��ˇ½�KT`H�G&K��%g���	
�W�Y���\C�=�9>Q�K����$��w�ȬU:2��E�Zf0#	�:����(�eb[Z=�㺺��F���2��S?yѝ����S����B�m}�ѢWx��	�S?�C�,	�{��G�#�*�;v�^�3ٰo��:�
��i�M�xN+r����9i&���ؗ�~,�F�P=:$�2-J��+�exG���8�������<7���1�l�jGO2m�<cx/����ݏ��L��Y(}���;&
k���gpb��"7�>�aX��� �I�+��~����ŉZ�
3���c�F�]��}�X��
�y�9%.mEd&��J�4�ba!����n�'a��x���fX�JJ>��0�V��k|�4ͼ`# 8��zI��zФG<��t�����Pּ.@t��7�>uF\m5Y4i��|gm�L�9�}s@3qp��%�y�y�k~�QW���~jI���|rNJ/cz�ŕ� �`CSk��Dv���p��H�=��ʏ���<��@ .�d�fYf�1m� h�pZ�t�|/V^y`�[��p{5�q��[�<�9�sc)�	zÞ��6�zmˮ&[��\�lZڬ��=�9]�U�?�L�+��h�Pb��\ 6�\I�˻�'�2ό��@鋢��|帷6��v�&Dc�"!w3���nU�ӊ�%��(��5�m#5��p�/YnA����[ Zd�B�i��}�聁�gŋ�3f��3R
/���	���v}FY��.�d	���nw:�>+�Sؒ4^fnuq�wDe	_u�S�������8Z�P�0�m1lM�%��$��Ҍ����`&梩[�
�#�K ~ʯŷ����y��2�����U�x4�QM��J��7�)Um_1BSCyp��Ô�f<K��'�F���w�څ�)��7j���\��f]v�M�g�%[����q�!��ʛ�S�ǈZ㑔��s�[�w7�O�g=��W2��{�v��Mxr���c]�mT���T��K�[a�pt�
29��Q?��O$�=(�ܾ�B �#����Ж뚜{�=2��Q�ѡ����Fl���'�2~�Ze�j�μ{Ά�2�����P0~`=#��(�ue�����M��9�`��Ǻ�TH-r���"ǅ�8͏��>ŸF�� �f(��%#SM�x���6��.�*���#r��j�-.`l� �1Z�P��>�L#5�P���h-�A�N��
h�u�r	�� cl@��s��1������'aظoȽh�W�\�?��Y'�G]����Ǿ����λc۶ڬb�*%��<����jq�8xn���1��DT����ER2�M�QvB��t�ɇm�=�O�����ނ)d?��@`,�de�m3�Nx��F[@��4��}�%:�THf<-��
6c�5�h��{����4с���(�q����T�i�\d2��b?��CG�_�T�hj�=��)�h�ǒϟ�RR惡/ma��>�@�ҕ���x�u<�:J�t%xr�?�>�b摐�'_�t�+͚s���~!$t(��	����hޭ�5�Q��D�Cs79M�Q3R]��3-��%��yU�a�q���_f/nefr������pf��U�ml�|F	凁BJ�@\pk�䕥�����+����	��lQڧI��{��4��ˬ}u)��i�^��2פ����2���gz8���߫H��x��Lx��C���b�4I(�<�r&2Tf�ش�v!oA�F5C$J����WE����=�)��CʼJ�H�ѩ��ߒ�
�hH��rx^5T�l6���
�P#��R�h�3 ���� �gQ�3d^�>"+ҹ+e���A���\�g�Ō�m�VB�<���ܰ��X^���Gt�|2��`�@f6
��H�����w0ԝ����/�vǴ��u��}Л��+�����m&��{��"���WO4EF-���ES	"������Zã�� b���x� �;��WN��q�|w�A��0�C�qˣz�#���E��"����g��t{��tB�EI[Mo�F��Ax((ݛ~�:�J>h�\Ӏ��d����<NXY��ڑdJ��z0�VM��3ժ� ��D8��-ñ�����(�c�*�|0�	�7a����"_��u~\�O��\�)���f��v*��7��,%1��:������F��Z9��+�,���
�=x钘p:��K*�� �cJ���Dx�Ϫ/�t}���4beJ9	_5�ZQ�����;كcH��!�9K:���u{we�ߕjѽW�Y�&s������q�����`��e�-�8�X��g��)�2Ԥ�Z�,��y��c�]�`W�Ӓ�[;.�P�ah1��?�S����Շ�O�b���<��L�����P�x�xD�W�KQ�bffi���(�G���@Ai�c,���4��3K�����6	�T����[w�^8�*�Rf��*W)��sgiD�_�-�wO�$�?MǬ�Ri'<OU���
�yu�ϊ�`�	%��GY���J5�c#���X�Dp1r��r����r��=�촶�� Sz�]�|e?�R(^bH�G�RKjt�;�-[i��
�X���&A����0�Q��c�q �v��;��z�_�+n�ʠ�/����o���ٿ�x�0?�&��j��qM�74z �^�$��uK[A���}@6�)�P�rS5n+u��U0 �/�;��w�H�E�,M��;�� ^�D��橈���5����)KD<�-(�K�(�hI���飄eoz�2�lN��푆Uv+N#}Q[��ΗAt�_ґ\�����!7��I�7u	��ati�t/|/9�(�d��٢×#�q�/��kY�k�U�m�;��U�d�ӛ��數\�O$̇��Ppa�X����1é��:$(A`[�F!�,�^��Qi�f	�M-��	1v�/:�mқO;�
�x<�x�q	2�s����;���NU���{S��C��u��9柋��0�� t���ơ�u��)���&ٗ�|�c�Q4���lP�b��بFQ/%Db*,���:��1aR��+�U/�'��O���׸@�����3� ߅��E���Qd��*�
����~6�,퉊q43�[>޲]8�SjirGz�\܎�����r���o����EFXuOt�����б4�ɥ]%�
K�O�b8���\ZŎ�T����m��Wգ- J4�ִ=��cD��=�����=�U>Jj���|'�(,�3m���B)1�=��0���P����s�������37㊆��a��E�U�Wx=\+�-�ٝ�s7G��(��M?�S���䬜�BPyT!������I�Ġ�&��]а��d֠Fbǌ�k`� ~7��Xfl�&��I'f��ʆ>�p�5B�ó�n~<�C�NBB[�MB���B��6��P�{���B��oڮ݀$�^��εC�I+�2M+��#�x��4��*:���p�`��fNؖ���W�fL�.Nf-���h׮�L�E;A�z��S��A�q���FT��=�hUv
� F�q޺xeܻ�"9wBm�A�Y�Alf[d�x�n/?R������2���߇������y[�x�Z�|:�$�g)S�v�ݙ�<�%
���j�h�*��ѿ&�K_��qQ��+=�� J\"���Cw�T��O��	�	�6�U��n�'r�jf� ���t�<_�/���`��/r_Ytl!�~؋L����uK<�c����p���*�}�_c	�#�d�*�f�3NO<#N�k������d)W�����/�X���a�Z�n���3w���UG��I�۴�((>̖8M9)�VM͊X�a_��Q2��J�1�%!HG���~�V��x7c�2v�Y왵�����S>�x�'�[�4�6*�K175�1��Z�[P����$Jm_x��b�&�20.:F��1�2�TF��r ���ݘb����6��?1���	y�2����QG���Ls�l�DreE.������(v�p/X=��NW��Z�K<h�ɛ��&����%vm2�����Ʒ:�8��^�!��K�5�B����ʅ��
E�!o�ЛN�
�MHs�X0mc��i� <.r��p��L�@~:�Fke��
��E7��)�A�3�G_�,�̻I���X`��Y���*�$��]v�&F;�]��~>6����`bǕ���o��T}+��on�KK8�s��u��w4b@���HK,Y详�����z��7׉���I_�֫�$�_q?��R%�(�us$n��|>�o�N�g�?t�_*ܨ�z>U*�.�ߠA.$�I�pM�z�[���Iy��Ne������~�*O0�Q��>�HB�.F3�����$Sw��ڕҶ���@@D�>�c|B�N��^G���ˇ[�b���`�����Y��/��;��s�<v�@�����{U�'ޖ�TT�o9�,�O��s��B�h������p=�����>�,�Q]L�KZJ���6Q'SXwގ��m�[�@�aWn���Q�>�b}+b�1_S�.9�����'�����<����O_�'#�]�B>p�FY0/o�d\}�N��20��}Ė��7�N2��ف"�՗{�&�Jʈ���p���%��1}P;��X�hFL��'�{v0cXː��;n������������/d6��&��e�����S�访��7LV�'�G�b���s(��BȘ���ϧ�&*�w�l �0�	�J-�ӻ�4�We���d$� O3�w<�zYK;���N�d����o�$|�Ea�a�69�z�2\�I+x7(�l*s/���z�����A���� 2�G�0�(D��'WF��-q��݋�M\MJ'n���C�j���8��_��������I5炆H�|�S��@}�+<�?����aR�FJ�oݺ��N���|
����ϓ�SX�cgAߦ���S�������9MDO@W�/C�;���w�W����
�Y��ׄt����칿Ѫb�Mcc<�t�qR,�i�̊6�����ܰ��� �]����z�[��ú �I�Fz�.�<ı�����i\�|f�k�n�|��� ��d��&���`�_y�2[B]���kM��rK{�S
���a����پȶ@SR�Jr�,*�BE��}�xgJz*>����'B���B]��a�v��>�f�[s�!�j���(���{7�md#�x�1
�x���y�����S.C���T,L ��,?�j������5i�%�*��(��k��z�ch�Y>��F#v���n��̗� �����s�	?��.\�"<x�ԯo�Q&A�M�9�r���>��죘P��r�l���ò�K��Q��0�*>����6�;-?%����%H=e'Ke�Uֲ�Y;D62��pcDK�'kՉѳ������b8�S)$+�d�`g$.6�M�<0i��S�iD<�0���vΏ�;������v�'$C_�g���{��'x���%1ub���)�"p��W��6P$$�J2}��e#<�3p�����3F��.�}����+���3�j�V���Z��>�U[-CJ
�ѿ�����2^�-b���ل�.Cx<t���A(�+���4�{$��O�c�S&�sČ�?�Q�0��@�BQ�Mx]�ES��eկͼ�=z�G�Y ��!�ˡ���m��4�6\��x�2��'����xD/��g�ħ�m�����Ρ�rH[��]�J [�x9Y,XY����1�ۙ��_G��֕4�4���=����-e[2���x��
!}��J�<���=��l�6犹u)�gjnV��Q�D��p�B��:�O�&���щ�5���<���v��,�dh�Е�y4(��,s��UMiV�^�$��{��zK˹�r�rD��B��o�Ltd�K'�Rx���c�i��tpS	������ �s9��h�e[��dE��[xlfq�&92�7+Ro�\#O~9�o������Fn��i
k�]�,n� Y���5K��!%ԅ��Ơ�X� -�T&y}q��!mK�܋`����3ܗ&W�D��{f<����ʻƈ�>#�ə��q��F�˲�m����[b�����G.�ȫ��/^���J�+j	uk}�ˣu���9T%,\�����،��~P���G0��;� M$P���)�He��c}L�q�ܖ����:`�H(]Ql8��F�o�([+5E�0J��z���G��&MU�=y>�+��mdO9�p$@�k�\�\����}�(��d��IFw=��t�MK�eȿ�p�l��gĝ���A;ȓ����]��֝S�Z���*\�-�|-��9
3�Y53��a�I����8��'@�O�����=��?��ѡ4�k&�L�H`�fa/��̟굌?���]r���"�Ŕ�E�{'����䦬�q��S��%y���:?��� ��	�	&����F(`U���ucm�?��5[`�2��4B��̫~o�
�G�K�0�!BM+b.˟��!���<�ل���t�'#^��w������&F��cʯ�^���0y��FN�9��v�S���V7�#jxņQ����i�[��)�����s�o������7B��x�9���[@^�����)Лx��P�d�Jmm�c�ك�EN�{�z�y�LSu��<�}�aы}�i�n��*���ꭊX���yco��?.Y�\8�vc�]�f�)�H�L7��#�1/Rq3 UT�ăe������5��6
��	Ԓ�vE��25����l\lQ{A�K���Ų�V[r��`���~g�Dj؏�m�.�'3�f1~�{l���n�5��T��L��K8q��,+��@�8�>?i�Z]d�-��z�0L����˙D��{��1�};S�3�@N�j��ͺ%o�-�V�*��������9�+�P����O��*y��6��eb۝ش�Pgjkio8>`�hm���夡�����?��렽�F�žBbmD����^�C��w��d�����0�4eNK�� ~<��ע��~ԃ�e����4��sF͗�/�F.��B'��2te[�ľ\�|���%�*wr�c������n�J��)�&6z�4+~Y�s/Q�G��0HGʫ���M�9A��wZS��<��r�k���|+/�=����0�i�n�h���o��0�@����t�Bpe�?�	��px�}��K<��_z	���=T0�8�gk˙����lnƄ�f!�B��PX�d�;����k;G����jo��(�Ӡ��5"�ؒ2ݺy�8`��)o�7@T��*�;��? w�D�a8l�<R�Tb�a�_��I��߻gb`-�6���ĂC�� ݜ����$�O�wt�Y]�/&_z{1�8�CI`��	�䖽j��|f��cT#vC�b���~�p>���O����d�1�Z�(�y[ @pO��!*�j�v~��#�څCЋS�`�r ΔD�����.�e-wo�=���`鳸�+Ѥ6������`K��kYDT�\c���o�AlV��J۳NAzG���B�ٔhz- Kw��wvyR�J�[8y���L�Ld��2+�ؿ��h�W7����M��
���H��9��mH�n����:Q2�Kg�m�շ���Z���ng�th��+M��x��c�Ds=д������(i[G�5*���WD�5�K��.jʴ��QΏU��-�4�v�!�X��BI�y��)wE����G�dROS�k7 ~h_vG�yvѻ��\�_<s���'�jq���\0�yP���_㣭���ľ�[r�@��ŕ6���>�@��4M�V�"?�zl&��b�h��1�?�0M
Hm�?9�S���[x=\i4�9����*��t����6��I�A���v� >��p�(��|��O��ٚ�N)��u�l��l3֢��Gb&ЦF"��iߚ��|�s�q�ɺܙ��[��)�9����K�Z����3Y���q[�[��u��k ��`�kg�k��H�]�5�/� h��IZ?��/��>Ջ]��j�5��;�D3������k��*]J�E~\�N���շWj�*�6]&�J���4j�����4���cv!�f'�Z���'ް"@����-[_��̃<Z
�{[��hS�(�<O��S��3Bi���؝�q�U��_|�T�M��m��S�����Q�B�lK\�vۤ�:�f��ε$��&�Xh 뽁�I�!�l� ���d<���kA}G��R��4�̡�(�e��OTۅ�\y9�v�T@���{��@��2�~Ŷ��ϚҮ������Se���<J�v-����N��'�zHJ�����>����[Pu��ż��|���,�Ӳn_�S){{nW�z�lS���V�R�PnJ�:-$)�(�jG3����G%�� �k�1�S�m��Ykb0m��RJu�?o�r�F�����	�p&�g�%���H�ő�����i�r���
#/Mk�Ms|�u3H0�?)���u�U������([���~v����n㏕�ȉ�!�(+G��3��j8��@(���U��g��طA���׷��B�Ve�ާ>	��c,`+�@(L���|����x\;u�k��yLWC�ݗ���M�丛9t����Q�S����m�yt-E��1v�=��(��U�H\����821U�FD�&{Oce���0�va��}��WS��UJ��7����4�Po�	�n��Sښ_�<D���g�Ae{ڭ͌���e�O�}���D3��������L�3T�2�� �#1��#�5ڍ�:��+��������6���q@��g��*�K ~t9S�ӻ].��@$�͍)���]�+��o �p�Z+磛��r����9�*��\�+�IPG��	�%,���e�c6�d�a�F�gѭ�j��)�/ V�_���\���;�4���D�a��T��V��'*"��3�naX�W�@>cZ��mL�q�(�׉XUhq40�`��*U���ie�!z+qQ�ȹ����|B���$�o@gB�׾�7��w���Z
��u�r@R���V���˰��?�\2��<��ؤ=��'��8��D�B����.�a�bB��/��R�9n���Q�_�,� K����;O��5��d�]�}/�C�i���nIWＶ��2�"pϧ�.$%BR��L�A�5=8�c�$�%��ӆjʪ��nIzvw^"���G��/L�\x�eIh��7fpk��I�V��rJ_!�� ]ґM���N������9|�h���<I�6�h�HT�'r]g&��`,&�aK�\���U{�)�5cP��O�{��O D!.x[J�_�lr��=��q	��	�� s��{byC��FFV!��������p{�H��xTC��,h��`��M%g����Q5��Q��nJV���=�'Jw�l������^���Tb�'�Ս��4w��ζ�3�h���B`��z,���'�rw����'X��_���4��n��0S�����Ɵ��� �p�c�#����6+h2�Ɩ>�
薬IH 8HBj
7kHd��l_�4gSb��/ډI����~jQ�X��� 	�5��O֬��q򰰐m� K6st]YH#� ��\��D=l*�L���9�i�T��������%h����$r�c����HkZy�:�(��Ը�Q;�:�
�K�&Nc���o�^J`�����;YC�/�xh�p�� ����_���`�A�9�B�xHV���ò����\d�Lv��@�Oo:5��kձ�qΥFԍ�K���N�X������M=���/��ߒa)J5>����6�j0�)�c����!�|h���~;��>�mpO���:�@O
�<�\$��d�qlwb�O_�^��:���w`�_��h���ƍŲ���\x� ���6c>f�#a2oa���coҸ�9�c5�Qy���V_��#�p��(���"�����K���9c�(ɭ�iA/��Ye	U��-Y�(��j��U�F��������9�7N��������.���Q��ة|�`Ctzr �~�Fte8���B�<�Q_@�����#�� X�5 ���9b�u��^���>���0g���%ǬZ]�Jί�pe�H�3�E�me8�@"��A�v��F��Q�gN(�6�s�4,�n�o�ٞ@'��Z"�3N� �����1ٱ��$X�j�/3o�2�:vR[Ҷ���%�*�E�\aj,�������˼u{���I�\ &�	T�=3�ٝ�(�@4��%U�b1^}�VI6��KA�3UU�cL���{R��:ƱGx�������h�h��
��=�3��þ1�4�gN�ȩ)���g��d�s��{�si����6�n�}%����Lf�)56d�<H42��k���>��K^6�����cq�!(jN�;[w���{�z����?�m.�oVMV��8�2�p�MA���C���f���-���� IR��"<>���J��ǃ���<r�M�9f1��i�O� 䜲���ti��a�tw�*I�j暘����@�P�r�{x����(�<���� ��Ȧ�a�%�J��jt8���u˯O�)�,2IJ`��ǉX!��) %�U�>��;�#����b�h�z�5�����-��3�t�\��}$���ݛ5�h��=�8q4�	\gL����z���M��iA��
{��DFF(� ��`��P9
����7q�O�;=	,�;4�8�D�䫶q�p�A�e���Vd���՗��و�J��\�Sj#I��Ά���cl_F]�c�*�&'(�Dm��A�����p� �rˌ<mw�����p�(�e���2{"�`�U�n0�@��KJ��rr��eqwx%���� 1r��VR&y�6ff�<@� ^�cЊ�F�E���U�E*�'����-��'Lգ7�e�~�F]&��<B��h�:�� *i>.�W�(���g�'A�s\V�<����>ŀ��h��jʚ�Lm����6Bʮ�W��*��2�^���W��k��pd��{Й��L�ҍ�@��F ��U�ԗ��K6%\�� �(��.�U[����+�F%�<ž@齢P��3�p��v}����7�e
�vYdy�Cl@�c��		�eYDײ���"E1�]K@=6�Y`�.	Wa��7������Ct눲���i�%̬�����XmAp��L���/_htny{Ƶ3�x���E�f�	C7�����A��~I�-���ĆC��	6��M�!D,|NO�=C�WE#4T�}�c��<Eٜ�����&��	����M����������/����#�0c��܌]&Ï>2dz�h�ݠ�V�J݅O��U(�cV5:/�OP��P_H8X<m�����V,��z���
��e�V}&glvcu�kv��ﳃi��t�r��_�6��j#k�4��(\�d���o�ĉj�'���W�b'�0<FM��Z�k~������%|_b���h['�����l(�����%_q�.��`3���,���t�I�>8��¼�h�DHKlki��3-	�;U����ǲ�Cix�����g&�`�+Lν���y1Z=ǥ�<� YT�2�+�S3���r�l�L[�#�X���OSY@��!$x�qO/�+"ԶLn��6]�ߏ�jM.������f6]g�Y�ʴ���O$C�ō�Ǡ��YǍQ�߻�Y��������"�p���8�?�:F��&���s��2�h���7Q�(�'��4
&T׾��w۱�A �h6�S����z}MU�LWDπ��<v�M�,�E�.B���ɥ���7ya�$v)o\��'N'�6{;!ܲa�F�ޢ����n�5Z��4�N1֛�C1p�`Ύ���;#S?S1A�+#J��9(Im~V�I�Փl�`/+@���e6n=����~�ڑ�`�2Q�T�}�E������l��;���c�]+/�� ��d�NLߑ���?�OH����;�-c[m�N[�Q�^Ƽ�/Z�7���0J�L?V�ێB���	�t4>�r:nqpW�����Ήo%�ɺ&,b��_���^I���"<&U�v�i��Mp=4p9V��o>�<��R�lp�?��k
|�S���ǈ�&��9���d�SU��2ڪ�G��j�Rg����*;�{mp�3�<x!��L*�R�a��b&�OF^�ֽ'F�ղKY�ֶ��|�o$�9+��f=H{�$�D+�!m�ۜø/p[�RV²�� �lM[X��s��x��l���z�[�p�[&�օV�{�g��ۀ5���m�=��ʈl�e�C'����ʹ��5��1��d�����h*9Q��Ix�)�Y�QV_�=K�t(��@�1A@x~�Q;{��3�p��>�w>�W�~���!ڧש\v��>�&�[S_�y�i��$̡^�9*X>�s�ux���F_�s��$H�?8��n��Y����8v�K��s�Jţ�����O6�L\�j���~���N-���(�)�F�vЊ;R[L�3��1��j+�������b��  �FG��w�0������d4QH��$�C�WgL�ڶ֚�v?v0;r�#�X����$F�,�Rχ�S�-�7F��Vh�ܺ��O�eP��+;��5dw��� TF���F��p�õ6QSe���ݮ�E�����f|�`����-�t������`��Ѹ���*L�j�0�:�+6&\�~ՎѪ8,r�7��;�}M֐B
���\ԧ��4���}�M2��(�{{6�w���m��4MT��X�$ް�\�H�)du:C�"���d�O��SԳ�
�����yѯ^�c��^d��5oq���)�FYʤ�8b!z�q�A��q�nb�f�!�[3���,|�{�AY�^�Ȅ�:K�K�cW,���22��d�
'h�t��a�|d��nT��\�F ��A:�F�j��g�M3������$�����ش��(gdb�(�
M+�U..��ש��ߣܷ*�E�r�c��q����<�3����SA�kk)0���4"E	���Z��ҩ���^�d��&��)�.'q":w�w��}MGA^���-�hs&�<��}M<ķ�Ha$Br$��Osr��ģ�p�˃�� \��p�k%��n7�������=n�����$�����_q��(9o���*'�^��8ve������xcʆ��]��lǣl>��X�9�4�Y��b栍�D�X�S���Q����:K�W��j����}����{�؎PB�,�Z8��*�f���D��~�XC���Co��m5�ѷD�hN��L��� ��(Ww<h�do� ����f)*d���ä��k�[l�U�{]��큔�O\�osU?��6!8Ѳ��Ӏ����X�fv�K����I��L�t�]J����́����t�P0�i稑W��m�[��g��_�f,��ɦ��I��9��`$�͊@,��_A�n�m��L�j�u��_�믇���-��|#���V�{�u�0���:QW��ޞ�j�;Wc��G�̙$!�r9�~�x��z��p��?X���
0�TK�r۩��;�PܪkG�u��>̈B�0<����P�)��N���F{3�J�+��G�m�t{ٰ2�I�h欰08n���n�B-��8z}r_�@�-���3T�e^4���A�d���d��ᅾ�e%���ɵZ����OIS^��wI�r�����������f��9��Ȉ��gX� &�|PGS�_���La����PM|_����x�AJ>��#����z�lđ�uG�GZ���fB��("�7.�b��H�ٳ�0@�bR����l��5��ݭ�2C7�&����HNx:u��������!{��q����Qc9���e s�[�O���
 /�k]���Zk?'�K��˃.It��G
�X�'w=��<s�F-����@���G+���"n"x-x���it]3�Qp���%��\?�>дM���u[$"0�ń��E�U�f�a�`��_��_Z���j�_�?fo��al0�BM>�m�6��j �s��B��r���E��+�c"	6|�dB��~�V���>7}C�h?f���W��j�c��ZBB�È����Q�0�z~��' �-
�l�P��AF�Q�;�|�Q��:�D��+0��8���ّ5�DrW=������!���=-ew��l ?��M<u�� '��-�9 ��+��Ww���SM�!��A,��O���(�{TFPf�p+�Y��\'��<�4��t>�2�O��^�7���2SD9�kvÙi��b���}�  ���ƀ����D���&|pK�ۄ�U1q�{3<D�`N��q-�
\�K�g��@�����>�U��a�ĕ0���8uoD��$7x[�n�����J�I�r�^6�< ���D5�k��v�ͽ.Fq����ՆG0�R+98�K)A�5�m�&<�Е���Do_l����,��Kc��Pv2����O|�6���TZ�/�qXk;_Z�����$��r[Y�!��>Z�>Nt�������}ƫA�06��7�ZSP	O�0%�aRч�Wh��]�Bl~(��x=�O����lu�9
�����Jj���nia�̙�l�����-"���<�:�C[��x��|��(�8��A3єT����y�c��-�݋�E�����m�=˘�*� ��|�M��0�\�i�`=#�����P�Z*GXq���"���Va0G|J��cH�R��0p�2��L��`*�/
����h�U�0i�F�&�������ST7���,�KNv*��}�h+l�\ɏ����!������"�yrg����'�M�
��Yȕ�0�$�xqC#��L�l����^�e��πh�8�ߦ��Z��q���������r��?[h�ٴ�b�,��a� (!�"�]��A�0mO��J���g���ȁ)1���Z1R����܂�D����.P݄�,��L_׃��X���1���p5��z���0Q�V8{v"�%`�4����s:<��x�4x�t�i?�j��k�,~��R�������H���I*�lj$����k)��V´5�'J|�*�G?��F���4*!��ܚ�^%���&�*p<�D�ͪ��D*�S���Ӑ{�+k������@<5�Ѱ
f5�HQ'��M9��F^L�N۠�K�b�݁(&��/~��~��/Q���8�H ��ˠ�����|*u�\8�T߈4�}x���oS���Ir@�;7����E���X)-�?��?����|��Fa��9[���CC�#Q|���{�>G\��3SE���qC��m���E��%��\&(BȠ��=�ٖ�>m�y(�,}��b,�6���(Cz-_vy���3����{�auf�([q~����ך�1�������N��c�� �>�kp�^�fu��a�->j�Vg@.��޺��(��S5E7&z�����I�nv�De�g��?�����0�@K3�@�7#{����j�g�a�q�j�]�X\"��WL�������F�C����,�3_�J��0�P�������t�A��Cz9-�?Xyf���#�?���T 
��J^��}�G�� F�����j�FS���}
�\��+�C���ŀ}.��Jlh�����U��~����'�d��ӃFl�2&�`M���s�=�[���L�bq@0ޥ�pq�{j�㉳^��m�T��Q�(G"���U�`�BX[���l @�S�r��ĿCLSU��1 ���Ol�ߤ��(w�մ���+F�����Ʀ��Cǂ�"|��\
����:l���u�cs������V'���ǱT��M�a[�������m'$5�u�9��sS-���S=� ԆI�*-�Vv��#�"���f��g�)��1}HsZw��z�l3l����͗�W3R!qe��eTM�K�Q�D<��;V����*aq�ŏP�X��z�����ԅk��*�W�]��]��ue"݅�b7�:׋<��,I�p��E��\u%*�h3������c�5A�ָ���S��
�W؋���έ<!��V�k\j.��Gf�gsI�3��4��w1{��ࢩ��Am�S��R��� �"D��H�%¦wڢ��r:�A!HY?��u���o��o|�2 ��2x�mb�g`ap�.�p ����g="5�^����p��Z�C)�#'��"՚kc���E�]D��n$w����Ð���Gm�_V��Rh�&,����3?MVއ�+9�.�>�G#ٗr�43ƍw�� ��8@U��fl���4/%~���Kl덈�|FS��-�]r�.�-%Ҷ�8x9!z���w�;���l�y��� jY�s��r0�U1��aDjY;�V�ON�w
m#�;g�نK�5���o�Zgw����?k^�`��11L�>�IS���ƅu�/����4�]�CQ!���Je�\�K�����~^�?�,o���,�`���	|N=�:$�)j���.�Eq91[f��)��X�Ҡ�� ]/[3����U�Y�
�IU�\}�2��=��{8�	3:��wC��1h���{r�����I��
=����Ѥ�k������+��;w"����	��2�?�|��L�M��J���R�UYw�E�`�l=�h����	����작���ɋ��j�>t�2ƿ
sĵt�H�W�2��a^���Oy�I�V׊szO�哸�l�hP)�|���IG��dN��(�q�b���b�A�|�&���+�d��9e��7�vq	����!�~Ur��]Ht�Nv ����3�ڙE�O�U�Ɩ}/��(�)5��ǡ6]�L����<A�w�lAi��DW�9J&�~Ũ�������J���PMQ#A�<�KP��,5���W�<1���Mз����F��of��a+H ��f����?,|+Ƅ��|i=�m}p�o�6�W��~�6����������2�k�JT���ﮬR�=z��b:ک�y�����No��n<�U��������<�����h��8��Q���WEKj��˵'1�(�:uBw:��x�}HG�^�&%���ݳ�KΤ�%�e!R�B��9���m$�M�ΕJ&o�����>��I���VW]K�![�)��zN���Z���B�Ovp8�]�ƫ
Lfm��? ����hD�o��V��؛L�)x�B��'x�m�:�����6v.�Ԯ�0�g��[�)�55z ��D��4N�������k����(PQ��F��R��b�F�@�����Fq�X�����p6N�f� ��A)�kZk�<���g%(	'�͵R�nVŽ@<�^RUV ���>aF}B>�I`N�n����d�����c
���)��Ф�8�w_d<!.�U�3t3����C5bя�m�c�[?�a&��O=��v�+�kJkEĿ�`/8b��u���M�2��ݟ�9���0䠐F��L{���I1�\��������ؚ�$%�Ͷ7-�z&��󃺏���ޅ��SI��-m6=����'���z�
��r�)�:c;1��T�#;��߽��X:;�L�����p!u{�q5d���w:@���8qfv��	bM���p�!�D��s��y/�#k-��ӄj�@/�J��U擙Y·� ��N�e��^�b���ܴ@a�Fcm���5�Y��c��������GZ5�ژ�Pʑu7���ziBK����~�}�� �%��|��
��)������Y�sX����5�3��<�c��G�ߛҼ�U`K}�۪�:��������P3uUAE�Xl�2�H2�� �m�0���P��O�0��dG�� ���`;�GB}�����
#3F�ة/�g�1Vt�	�����Ѥ�tO�A$
�@g���	^�z���$�2i%+g�#�	�f3�l��^�?.T�	Ŧ����E�j��<�9[Y�aj��bT�g<������{��E"���%�o���q�{������\`x��A�˽��%��Ar�f�'m���,C����?�F���/ޜ�f��+W�p�Q��\dMq�Qöp$�D(!e����9�qY3�� ���r"�8�ي&�G)?񫙸Ē�����w�}Oz��{'x(�T���.~�� ���1	^X���m����	��ʊM���\����I�3n{�r-)���P�4�n=��}���{	U�ڏ���b����d�Ê��繠f�_�jqXx��c'��w?�
쟝��;3h�IJ1��w!�>{��Cb�$��ӁQ=iJ��Q*��ʿ ���1�ƣ4�ٖ{��R�P]�:�ޝ�̚�#��mm�������P��,1�Ic�izOR�!-w{��Rtg��ĺ�P�}>1薀y�!�H�vq��GFTtEN�D�|��M�!E�2�A�����~i��(��q7�/���_7�db-���S���=tT��D^$�itI4�I~��������ˏQw���ri �ǝ=��*s	�uC�zP��{]��(<��3�,��6֟����V�a\�/SGUخ�]�,ܬY����^��a8&��x�T]�u�Ё�.��_,}��#��E��?4�*Ns��HzG�ӛ�%~
b��W1x8�3'�4������5*�o�Z�Mħ�c��Xlc��Z��i�؇q�4�Q��тM	~)�� d�*��>�ڞ�����<SjQ���Q���<r�t�4u0�$�z晧;�M�q��Y�4��/b� }��j���Щi����6��y|5�k�˩�6��fi���z;C��=Yl�ၳ!+��Q0�~��l��r�8_ܼ���Km?E�ݭ�W:rvk��#$���Լ�MA��э���������Qo5����J�[�bL����_DZG>�;���M/�&����)�(�ˌ �l��$6��]H%�0�F0����Q��=��q��F�"k$=���|��\P7�Q�u� ���➊��t L�g�w�x������㌊?��Aj�QE���/����=N�X�=��U?wpvH�S��&?�4�&��0����(��S�S��E���m��o��|�i�W�!���4и�g�9ʫ���O���/�JZ����<�r(Q�'gh��RRC���+T6&�KP>y.���]�'�-C��r�%
'c���9�6��kE��t�	�~��;�?L��������E2g��X�LJjӘ}�����C�]ďO�G�F��|�q���Ƈ��A��6�Iib%���К�������w�[0��HGou7ь�i��g��Vt��-Nx#���s� 99n�Fm�b�VR~���I��Ob�o]y���(�D[eĲ	gP ��J�{�M���D7�0�0/��J�q�F�d�T[���+�є��%8�0
��6Jѐ��ߦ�}]C;'�w�o�bȹ�J�-^9�ң�h=�=9��^|�l�K><��O���*>F�h���9�%P5�M���c�*�����5��\S&J��a�6�bL�Ы?�OԨX�t3	����"�C���I����2�*���EY���_˲����W��3آq���v3������Av�P���*���׋o����V&�E�p��/%�MJK}��5���"���
z5��+�OM���%Z�{�����Ec�gQ�Put֜�uti�I����6�L��ĩ�j|VB.ѴF2�Y�@ғ3��f����b�p,/���<"�G'5��K�=��l���x�shTW**8dd�bT����u�NEsj����
�8����(���+���x!�t$J͑�cz	= E�k=(
ӄИ�wu��@g���!@�2�vw�Dx��cF�	h����WT�ĸ�>*p��Ɲf�IA;h��n��b+�:I���3��Xa��E1�Tyue�K�sW�,������b��c���rIځtw�762�̒�=�2�p�;�kF��;����1;��7G�ߞR`�@,�KG^�G�[�fj��m�N����C��#u`�,��F,0!˩���BA�����F�l!٘�Q���:���j�{&>�z���y+}rG<3�;�("h%���ۆ��yc0��0Fӌ��<��ќ5u�����pv6* Rg`$8�x�Ҷ�jr�7�3���\��Ǹݫ���E�r{��Ԫ�9�,g=t�m_QmҹZ:_��C�����4c��б���1oQ
��V��=ҫ�����I�u���h�p���6��\U��2��V�:+�#��0�����h� �{�ig�����L��7$ʼ��kV�����nHGU���mA,�@��5���"����2��VW�D��)L4s�]�O�������͜��ɵ����U�w�d>p��[	��T������m¬\)@��BW�9mA��ɔ�k1A2�ˬx�(AJ�ٓ�^`��M�gP�X�xa.��i4�6�6��Y���D�.�J�=m�~^�*�%X4�*�8��
��4�O��F����ͅx�I����B�5ۻ�Ɲ��E��=h[�$�pa�$w>I��[(o�M�@;�*OyLi���P.��%v���� ���.��UN��M�)�,7F��p[���/&QpdY7мҢ�jq�ܬ��APr;�������h3��G�*���RS��A�B��п��JXJ����=9,��^fw����*U*E�[��:o����*�-΁K�I�a����6*CB����w�~�d]�X�Fb܌�"���	c�5~Myކ0K=�yv1�� �e[�>@ʓ%�p��P1o;���T�J� �3�)�����nn�'��|4\��d�vq�1�Ӿn�}��t>}�V�P�!�I��ۣRs���������O�CV���O���o��q���C�ui}3��K��ݔR>�Ƃ��> �t��Օ�gvjVP�r2�@o�E~�{x�U����c�k��$q��gb4~�hmh�����Lk�F���������S�#�'�Zy�<!��w��D0�SU3���e^�IGm��[�G��K���y��4蘼�3�X���,��u.��]���W�Y?6D���+�_JX
�f�Ӿ��ฆ���1���}����I�K���۽tr�4h����=��^�mnt	B/'�I�����	O�G��ϓh.]^�|I����
@��42((e��rF6��Yrc[�q�摒s5*�ݍ��6�,���MO@ę�m|t�g�~�j�/��i{���p��t�B�~x?��o��f��w?8���ع��9���&P�<��݆-�.�3Kr�%��=)�P�Ò�~����k�מ5�i�P�/%�--܋<xS�,�2B��JN�]8����*�ݗ~|�'���,�ǖ4/�A��p�1�hD35M��<c�`8D�MP��O}�����Xổ�(%+�Z�:{i��ǡ|t[A}���f�D�霃��7�QL������ߠ�ԫ����y�@x�E|����o��:��J�� ��@�dx��ݰNjќ�V�ܗ�s�Gz~��dD��1��1	��:IG���܃��F�y|nǜ�7��O�Z8��=�n��^�������&����r�$���U��`�q�,?��h1М��<�>/�Jo�w����lKH�Q�����z�x��<4�@#��f��IYa�Ӂ��x�lz�Y���N�,��A���E��!(�m����Y�z��MD^��q����
2C�2Fk�mK�L�G�G����_�